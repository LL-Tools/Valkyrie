

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944;

  OR2_X1 U11018 ( .A1(n14559), .A2(n19908), .ZN(n11230) );
  AOI211_X1 U11019 ( .C1(n15383), .C2(n15404), .A(n15409), .B(n15382), .ZN(
        n15402) );
  OAI22_X1 U11020 ( .A1(n13966), .A2(n9942), .B1(n14882), .B2(n9940), .ZN(
        n13992) );
  AND2_X1 U11021 ( .A1(n14766), .A2(n14767), .ZN(n15316) );
  NOR2_X2 U11022 ( .A1(n18519), .A2(n18532), .ZN(n17939) );
  AND2_X1 U11023 ( .A1(n11735), .A2(n9699), .ZN(n9995) );
  BUF_X2 U11024 ( .A(n15856), .Z(n9581) );
  NAND2_X1 U11025 ( .A1(n13156), .A2(n15505), .ZN(n14823) );
  INV_X2 U11026 ( .A(n18896), .ZN(n18915) );
  AND2_X1 U11027 ( .A1(n13512), .A2(n9702), .ZN(n13710) );
  NAND2_X1 U11028 ( .A1(n11112), .A2(n11111), .ZN(n11113) );
  INV_X1 U11029 ( .A(n18094), .ZN(n17185) );
  NAND2_X1 U11030 ( .A1(n13151), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13152) );
  NAND2_X1 U11031 ( .A1(n17694), .A2(n17695), .ZN(n17693) );
  NOR2_X1 U11032 ( .A1(n11518), .A2(n11496), .ZN(n19360) );
  INV_X1 U11033 ( .A(n15592), .ZN(n9608) );
  XNOR2_X1 U11034 ( .A(n10365), .B(n10364), .ZN(n10462) );
  NAND2_X1 U11035 ( .A1(n10325), .A2(n10324), .ZN(n10454) );
  INV_X1 U11036 ( .A(n16815), .ZN(n16965) );
  AND2_X1 U11037 ( .A1(n11529), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12140) );
  AND2_X1 U11038 ( .A1(n9601), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12169) );
  INV_X1 U11039 ( .A(n17065), .ZN(n15641) );
  NAND2_X1 U11040 ( .A1(n9988), .A2(n9990), .ZN(n11464) );
  CLKBUF_X3 U11041 ( .A(n12475), .Z(n17036) );
  CLKBUF_X2 U11043 ( .A(n11999), .Z(n12014) );
  NAND2_X1 U11044 ( .A1(n11448), .A2(n12748), .ZN(n13350) );
  INV_X1 U11045 ( .A(n15592), .ZN(n17053) );
  CLKBUF_X2 U11046 ( .A(n12470), .Z(n17061) );
  INV_X1 U11047 ( .A(n16815), .ZN(n17062) );
  NOR3_X1 U11048 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18672), .A3(
        n18522), .ZN(n12475) );
  AND2_X1 U11049 ( .A1(n10222), .A2(n20132), .ZN(n11063) );
  BUF_X2 U11050 ( .A(n12474), .Z(n9579) );
  NAND2_X1 U11051 ( .A1(n18690), .A2(n16736), .ZN(n16773) );
  INV_X1 U11052 ( .A(n11927), .ZN(n11916) );
  OR2_X2 U11053 ( .A1(n10206), .A2(n10205), .ZN(n10222) );
  CLKBUF_X2 U11055 ( .A(n11424), .Z(n13139) );
  INV_X1 U11056 ( .A(n11424), .ZN(n12798) );
  INV_X1 U11057 ( .A(n11737), .ZN(n11440) );
  NAND2_X1 U11058 ( .A1(n10086), .A2(n10085), .ZN(n20122) );
  NAND4_X2 U11059 ( .A1(n10168), .A2(n10167), .A3(n10166), .A4(n10165), .ZN(
        n10229) );
  AND2_X1 U11060 ( .A1(n13118), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11408) );
  AND2_X1 U11061 ( .A1(n13118), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9606) );
  NAND4_X1 U11062 ( .A1(n10046), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10161) );
  CLKBUF_X1 U11063 ( .A(n20092), .Z(n9574) );
  NOR2_X1 U11064 ( .A1(n20091), .A2(n20090), .ZN(n20092) );
  CLKBUF_X1 U11065 ( .A(n20141), .Z(n9575) );
  NOR2_X1 U11066 ( .A1(n20090), .A2(n20089), .ZN(n20141) );
  NAND2_X2 U11068 ( .A1(n13461), .A2(n13460), .ZN(n13456) );
  NOR2_X2 U11069 ( .A1(n13036), .A2(n13157), .ZN(n13156) );
  AND2_X2 U11070 ( .A1(n13511), .A2(n13510), .ZN(n13512) );
  NAND2_X1 U11071 ( .A1(n9970), .A2(n9851), .ZN(n9576) );
  NOR2_X4 U11072 ( .A1(n17217), .A2(n17738), .ZN(n17598) );
  NAND2_X2 U11073 ( .A1(n17939), .A2(n18529), .ZN(n17956) );
  BUF_X2 U11074 ( .A(n11505), .Z(n14847) );
  NAND2_X1 U11075 ( .A1(n11505), .A2(n13057), .ZN(n11514) );
  OR2_X1 U11076 ( .A1(n11505), .A2(n11501), .ZN(n19327) );
  OR3_X2 U11077 ( .A1(n11505), .A2(n13057), .A3(n11510), .ZN(n11665) );
  NAND2_X1 U11078 ( .A1(n11505), .A2(n14861), .ZN(n11511) );
  OR3_X2 U11079 ( .A1(n11505), .A2(n13057), .A3(n11512), .ZN(n19247) );
  INV_X1 U11080 ( .A(n10840), .ZN(n11039) );
  INV_X1 U11081 ( .A(n10154), .ZN(n10308) );
  OAI21_X1 U11082 ( .B1(n13647), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10280), 
        .ZN(n10301) );
  NAND2_X1 U11083 ( .A1(n18682), .A2(n18672), .ZN(n12426) );
  AOI21_X1 U11084 ( .B1(n10454), .B2(n10453), .A(n10329), .ZN(n10444) );
  CLKBUF_X2 U11085 ( .A(n11528), .Z(n9588) );
  NAND2_X2 U11086 ( .A1(n11379), .A2(n11378), .ZN(n11737) );
  NAND4_X1 U11087 ( .A1(n11423), .A2(n13139), .A3(n11440), .A4(n19157), .ZN(
        n12049) );
  AND2_X1 U11088 ( .A1(n9588), .A2(n11530), .ZN(n13703) );
  AND2_X1 U11089 ( .A1(n11409), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11602) );
  NAND2_X1 U11090 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n16736), .ZN(
        n12425) );
  INV_X1 U11091 ( .A(n14089), .ZN(n13105) );
  INV_X1 U11092 ( .A(n10509), .ZN(n11057) );
  CLKBUF_X2 U11094 ( .A(n15017), .Z(n9610) );
  NAND2_X1 U11095 ( .A1(n15421), .A2(n9835), .ZN(n15085) );
  NAND2_X1 U11097 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18522) );
  NAND3_X1 U11098 ( .A1(n11156), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14419), .ZN(n14402) );
  XNOR2_X1 U11100 ( .A(n11082), .B(n11083), .ZN(n13151) );
  NAND2_X1 U11101 ( .A1(n10387), .A2(n10386), .ZN(n13503) );
  AND2_X1 U11103 ( .A1(n15315), .A2(n9713), .ZN(n14886) );
  AOI22_X1 U11104 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14710), .B1(n15022), 
        .B2(n18737), .ZN(n14711) );
  NAND2_X1 U11105 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18517) );
  INV_X1 U11106 ( .A(n11320), .ZN(n14087) );
  NOR2_X1 U11107 ( .A1(n11160), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14373) );
  NOR2_X1 U11108 ( .A1(n12598), .A2(n12597), .ZN(n18062) );
  INV_X1 U11109 ( .A(n19955), .ZN(n15810) );
  INV_X1 U11110 ( .A(n19993), .ZN(n19981) );
  AOI211_X1 U11111 ( .C1(n15889), .C2(n14399), .A(n14398), .B(n14397), .ZN(
        n14400) );
  OR2_X1 U11112 ( .A1(n12757), .A2(n11420), .ZN(n16168) );
  INV_X2 U11113 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9751) );
  INV_X2 U11114 ( .A(n10161), .ZN(n10700) );
  INV_X2 U11115 ( .A(n10161), .ZN(n9621) );
  INV_X1 U11116 ( .A(n15892), .ZN(n15856) );
  AND2_X1 U11117 ( .A1(n10209), .A2(n10210), .ZN(n9577) );
  NAND2_X1 U11118 ( .A1(n11703), .A2(n11702), .ZN(n15215) );
  NAND2_X2 U11119 ( .A1(n11138), .A2(n9983), .ZN(n14514) );
  NAND2_X2 U11120 ( .A1(n13749), .A2(n11136), .ZN(n11138) );
  INV_X1 U11121 ( .A(n12438), .ZN(n9578) );
  NOR2_X1 U11122 ( .A1(n12425), .A2(n12429), .ZN(n12474) );
  NAND2_X2 U11124 ( .A1(n11348), .A2(n11347), .ZN(n11424) );
  AND2_X2 U11125 ( .A1(n11920), .A2(n11416), .ZN(n11448) );
  NAND2_X2 U11126 ( .A1(n11482), .A2(n11481), .ZN(n11942) );
  OAI21_X2 U11127 ( .B1(n14802), .B2(n12300), .A(n15404), .ZN(n15182) );
  NOR2_X4 U11128 ( .A1(n12425), .A2(n12431), .ZN(n15615) );
  AND2_X4 U11129 ( .A1(n19890), .A2(n19883), .ZN(n12079) );
  AND2_X2 U11131 ( .A1(n12967), .A2(n12996), .ZN(n10160) );
  XNOR2_X2 U11132 ( .A(n11943), .B(n11942), .ZN(n11940) );
  NAND2_X2 U11134 ( .A1(n9783), .A2(n9781), .ZN(n11927) );
  AOI211_X2 U11135 ( .C1(n14561), .C2(n20075), .A(n14554), .B(n14566), .ZN(
        n14552) );
  XNOR2_X2 U11136 ( .A(n17237), .B(n12509), .ZN(n12523) );
  AND2_X1 U11137 ( .A1(n10064), .A2(n10060), .ZN(n9583) );
  AND2_X1 U11138 ( .A1(n10064), .A2(n10060), .ZN(n10197) );
  OAI21_X2 U11139 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18710), .A(n16393), 
        .ZN(n17735) );
  AND2_X1 U11140 ( .A1(n9956), .A2(n9953), .ZN(n11160) );
  AOI211_X1 U11141 ( .C1(n15391), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15390), .B(n15389), .ZN(n15392) );
  OR2_X1 U11142 ( .A1(n12329), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12330) );
  CLKBUF_X1 U11143 ( .A(n14120), .Z(n14132) );
  NOR2_X2 U11144 ( .A1(n15063), .A2(n15231), .ZN(n12329) );
  NOR3_X1 U11145 ( .A1(n15085), .A2(n15062), .A3(n15276), .ZN(n12313) );
  CLKBUF_X1 U11146 ( .A(n14248), .Z(n14249) );
  NAND2_X2 U11147 ( .A1(n15215), .A2(n15216), .ZN(n11736) );
  AND2_X1 U11148 ( .A1(n13736), .A2(n13735), .ZN(n13737) );
  OAI21_X1 U11149 ( .B1(n20027), .B2(n9973), .A(n15911), .ZN(n9972) );
  NAND2_X1 U11150 ( .A1(n14976), .A2(n9746), .ZN(n14958) );
  OR2_X1 U11151 ( .A1(n15856), .A2(n14540), .ZN(n14492) );
  NAND2_X1 U11152 ( .A1(n9905), .A2(n9904), .ZN(n17515) );
  AND2_X1 U11153 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16850), .ZN(n16855) );
  NOR2_X1 U11154 ( .A1(n16518), .A2(n16868), .ZN(n16850) );
  BUF_X2 U11155 ( .A(n12898), .Z(n13057) );
  NAND2_X2 U11156 ( .A1(n11483), .A2(n11484), .ZN(n11490) );
  NAND2_X1 U11157 ( .A1(n12751), .A2(n9616), .ZN(n12359) );
  NAND2_X1 U11158 ( .A1(n12840), .A2(n10169), .ZN(n12914) );
  NAND2_X1 U11159 ( .A1(n9616), .A2(n9584), .ZN(n12970) );
  INV_X2 U11160 ( .A(n12686), .ZN(n18089) );
  AND2_X1 U11161 ( .A1(n9584), .A2(n10222), .ZN(n13630) );
  INV_X1 U11162 ( .A(n18716), .ZN(n16410) );
  INV_X2 U11163 ( .A(n10209), .ZN(n10233) );
  BUF_X1 U11164 ( .A(n10212), .Z(n20127) );
  INV_X2 U11165 ( .A(n20122), .ZN(n9841) );
  INV_X1 U11166 ( .A(n13368), .ZN(n11895) );
  NOR2_X1 U11167 ( .A1(n16175), .A2(n14723), .ZN(n14722) );
  CLKBUF_X2 U11168 ( .A(n10576), .Z(n11034) );
  NOR2_X1 U11169 ( .A1(n9862), .A2(n9861), .ZN(n9860) );
  AND3_X1 U11170 ( .A1(n10183), .A2(n10185), .A3(n10186), .ZN(n9858) );
  CLKBUF_X1 U11172 ( .A(n10260), .Z(n10978) );
  CLKBUF_X2 U11173 ( .A(n10197), .Z(n11033) );
  AND2_X1 U11174 ( .A1(n12967), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9622) );
  AND2_X1 U11175 ( .A1(n10046), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10061) );
  AND2_X1 U11176 ( .A1(n13118), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9605) );
  AND2_X2 U11177 ( .A1(n11531), .A2(n13343), .ZN(n11523) );
  AND2_X2 U11178 ( .A1(n11531), .A2(n13343), .ZN(n9607) );
  INV_X2 U11179 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13343) );
  INV_X2 U11180 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9875) );
  OR2_X1 U11181 ( .A1(n14381), .A2(n15892), .ZN(n9856) );
  AOI211_X1 U11182 ( .C1(n15889), .C2(n14417), .A(n14416), .B(n14415), .ZN(
        n14418) );
  AOI21_X1 U11183 ( .B1(n15051), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n9764), .ZN(n15041) );
  NOR2_X1 U11184 ( .A1(n12315), .A2(n12329), .ZN(n15034) );
  XNOR2_X1 U11185 ( .A(n12356), .B(n12355), .ZN(n14379) );
  OAI21_X1 U11186 ( .B1(n15160), .B2(n15161), .A(n15109), .ZN(n15146) );
  NAND2_X1 U11187 ( .A1(n9722), .A2(n15105), .ZN(n15160) );
  AND2_X1 U11188 ( .A1(n15496), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15461) );
  OAI21_X1 U11189 ( .B1(n13966), .B2(n13965), .A(n13990), .ZN(n9939) );
  NAND2_X1 U11190 ( .A1(n15097), .A2(n15096), .ZN(n15098) );
  NOR2_X1 U11191 ( .A1(n15515), .A2(n11755), .ZN(n15496) );
  NAND2_X1 U11192 ( .A1(n11837), .A2(n15310), .ZN(n15097) );
  NAND2_X1 U11193 ( .A1(n15419), .A2(n15416), .ZN(n15183) );
  AND2_X1 U11194 ( .A1(n9723), .A2(n15194), .ZN(n15419) );
  XNOR2_X1 U11195 ( .A(n15021), .B(n15020), .ZN(n16101) );
  NAND2_X1 U11196 ( .A1(n12304), .A2(n12303), .ZN(n16186) );
  OR2_X1 U11197 ( .A1(n12026), .A2(n14873), .ZN(n16053) );
  OR2_X1 U11198 ( .A1(n14704), .A2(n14707), .ZN(n15255) );
  NOR4_X1 U11199 ( .A1(n14547), .A2(n14546), .A3(n14545), .A4(n14544), .ZN(
        n14548) );
  NAND3_X1 U11200 ( .A1(n12296), .A2(n9829), .A3(n9828), .ZN(n15206) );
  NAND2_X1 U11201 ( .A1(n12342), .A2(n15228), .ZN(n16023) );
  OR2_X1 U11202 ( .A1(n13885), .A2(n13884), .ZN(n10017) );
  OR2_X1 U11203 ( .A1(n12338), .A2(n12264), .ZN(n14935) );
  NAND2_X1 U11204 ( .A1(n17400), .A2(n12554), .ZN(n12555) );
  NAND2_X1 U11205 ( .A1(n11664), .A2(n11663), .ZN(n13587) );
  OAI21_X1 U11206 ( .B1(n9995), .B2(n9627), .A(n11766), .ZN(n9730) );
  NOR2_X1 U11207 ( .A1(n15313), .A2(n15312), .ZN(n15315) );
  INV_X1 U11208 ( .A(n14476), .ZN(n11152) );
  AND2_X1 U11209 ( .A1(n10029), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9830) );
  AND2_X1 U11210 ( .A1(n14941), .A2(n14940), .ZN(n12262) );
  AND2_X1 U11211 ( .A1(n14941), .A2(n9748), .ZN(n12338) );
  NAND2_X1 U11212 ( .A1(n12004), .A2(n12003), .ZN(n15313) );
  OR2_X1 U11213 ( .A1(n14614), .A2(n14611), .ZN(n14531) );
  INV_X1 U11214 ( .A(n15125), .ZN(n12004) );
  OR2_X1 U11215 ( .A1(n15123), .A2(n15124), .ZN(n15125) );
  NAND2_X1 U11216 ( .A1(n11733), .A2(n18880), .ZN(n11734) );
  NAND2_X1 U11217 ( .A1(n13497), .A2(n12280), .ZN(n13565) );
  OR2_X1 U11218 ( .A1(n12306), .A2(n12300), .ZN(n12305) );
  OR2_X1 U11219 ( .A1(n13564), .A2(n13597), .ZN(n9826) );
  NAND2_X1 U11220 ( .A1(n9769), .A2(n14845), .ZN(n13483) );
  AND2_X1 U11221 ( .A1(n14926), .A2(n15154), .ZN(n15152) );
  AND2_X2 U11222 ( .A1(n11062), .A2(n11065), .ZN(n15892) );
  NOR2_X2 U11223 ( .A1(n13422), .A2(n13421), .ZN(n13511) );
  CLKBUF_X1 U11224 ( .A(n14766), .Z(n15340) );
  AND2_X1 U11225 ( .A1(n14527), .A2(n14526), .ZN(n14674) );
  AND2_X1 U11226 ( .A1(n10434), .A2(n10433), .ZN(n11098) );
  OAI211_X1 U11227 ( .C1(n10476), .C2(n12996), .A(n10475), .B(n10474), .ZN(
        n13455) );
  AND2_X1 U11228 ( .A1(n10424), .A2(n10502), .ZN(n11105) );
  CLKBUF_X1 U11229 ( .A(n11088), .Z(n11089) );
  INV_X1 U11230 ( .A(n16846), .ZN(n16849) );
  AND2_X1 U11231 ( .A1(n11692), .A2(n11691), .ZN(n11693) );
  CLKBUF_X1 U11232 ( .A(n13612), .Z(n13695) );
  INV_X1 U11233 ( .A(n15425), .ZN(n9795) );
  AND2_X1 U11234 ( .A1(n11730), .A2(n11729), .ZN(n12298) );
  OR2_X1 U11235 ( .A1(n13514), .A2(n13515), .ZN(n15425) );
  NOR2_X1 U11236 ( .A1(n13721), .A2(n13722), .ZN(n14681) );
  NOR2_X1 U11237 ( .A1(n9757), .A2(n11516), .ZN(n9756) );
  AND2_X1 U11238 ( .A1(n13503), .A2(n9838), .ZN(n9999) );
  AND2_X1 U11239 ( .A1(n10447), .A2(n10330), .ZN(n10463) );
  AND4_X1 U11240 ( .A1(n11547), .A2(n11546), .A3(n11545), .A4(n11544), .ZN(
        n11558) );
  NOR2_X1 U11241 ( .A1(n14268), .A2(n11293), .ZN(n14269) );
  AOI22_X1 U11242 ( .A1(n19211), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n19111), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11520) );
  OR2_X1 U11243 ( .A1(n12956), .A2(n12957), .ZN(n12958) );
  INV_X1 U11244 ( .A(n17582), .ZN(n17566) );
  OR2_X1 U11245 ( .A1(n11511), .A2(n11513), .ZN(n19419) );
  INV_X1 U11246 ( .A(n19564), .ZN(n19556) );
  AND2_X1 U11247 ( .A1(n11519), .A2(n18929), .ZN(n19211) );
  OR2_X1 U11248 ( .A1(n11511), .A2(n9670), .ZN(n19487) );
  OR2_X1 U11249 ( .A1(n11511), .A2(n11512), .ZN(n19521) );
  CLKBUF_X2 U11250 ( .A(n12980), .Z(n9603) );
  NAND2_X1 U11251 ( .A1(n11077), .A2(n10302), .ZN(n10330) );
  NAND2_X1 U11252 ( .A1(n17647), .A2(n12539), .ZN(n12540) );
  AND2_X1 U11253 ( .A1(n13013), .A2(n13012), .ZN(n13034) );
  AND2_X1 U11254 ( .A1(n12904), .A2(n12903), .ZN(n12905) );
  OR2_X1 U11255 ( .A1(n11514), .A2(n11510), .ZN(n19591) );
  OR2_X1 U11256 ( .A1(n11514), .A2(n11512), .ZN(n19684) );
  NAND2_X1 U11257 ( .A1(n11495), .A2(n13347), .ZN(n11518) );
  NOR2_X1 U11258 ( .A1(n16552), .A2(n16897), .ZN(n16909) );
  INV_X1 U11259 ( .A(n13057), .ZN(n14861) );
  NAND2_X1 U11260 ( .A1(n13598), .A2(n12113), .ZN(n13000) );
  NAND2_X1 U11261 ( .A1(n12728), .A2(n16410), .ZN(n17738) );
  INV_X1 U11262 ( .A(n18929), .ZN(n13355) );
  NAND2_X1 U11263 ( .A1(n12797), .A2(n12796), .ZN(n12901) );
  AND2_X1 U11264 ( .A1(n9903), .A2(n9902), .ZN(n17668) );
  NAND2_X1 U11265 ( .A1(n10369), .A2(n10368), .ZN(n20251) );
  NOR2_X1 U11266 ( .A1(n9737), .A2(n9735), .ZN(n9734) );
  OAI21_X1 U11267 ( .B1(n17693), .B2(n9901), .A(n9899), .ZN(n9903) );
  OR2_X1 U11268 ( .A1(n10336), .A2(n12996), .ZN(n10369) );
  INV_X2 U11269 ( .A(n18988), .ZN(n18983) );
  NAND2_X1 U11270 ( .A1(n11472), .A2(n11473), .ZN(n11475) );
  AND2_X1 U11271 ( .A1(n11753), .A2(n9697), .ZN(n11757) );
  AND2_X1 U11272 ( .A1(n11181), .A2(n11180), .ZN(n11191) );
  NOR2_X2 U11273 ( .A1(n11742), .A2(n11739), .ZN(n11753) );
  INV_X1 U11274 ( .A(n9731), .ZN(n12098) );
  NOR3_X2 U11275 ( .A1(n18716), .A2(n18062), .A3(n15761), .ZN(n17099) );
  OR2_X1 U11276 ( .A1(n11699), .A2(n11698), .ZN(n11742) );
  NOR2_X2 U11277 ( .A1(n15689), .A2(n12535), .ZN(n17608) );
  AOI21_X1 U11278 ( .B1(n11477), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n10038), .ZN(n11457) );
  AND2_X1 U11279 ( .A1(n11637), .A2(n11631), .ZN(n11696) );
  NAND2_X1 U11280 ( .A1(n9609), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11427) );
  AND4_X1 U11281 ( .A1(n11454), .A2(n11453), .A3(n13390), .A4(n11452), .ZN(
        n11458) );
  AND2_X1 U11282 ( .A1(n12811), .A2(n12812), .ZN(n12810) );
  NAND2_X1 U11283 ( .A1(n16392), .A2(n9774), .ZN(n15650) );
  NAND2_X1 U11284 ( .A1(n12367), .A2(n10435), .ZN(n13014) );
  BUF_X4 U11285 ( .A(n11477), .Z(n15019) );
  NOR2_X1 U11286 ( .A1(n11639), .A2(n11638), .ZN(n11637) );
  NAND2_X1 U11287 ( .A1(n17715), .A2(n12524), .ZN(n12527) );
  NAND2_X1 U11288 ( .A1(n11218), .A2(n10236), .ZN(n14692) );
  NAND2_X1 U11289 ( .A1(n12083), .A2(n12082), .ZN(n12811) );
  CLKBUF_X1 U11290 ( .A(n11248), .Z(n14090) );
  INV_X2 U11291 ( .A(n11169), .ZN(n11200) );
  NAND2_X1 U11292 ( .A1(n9807), .A2(n11903), .ZN(n11888) );
  NAND2_X1 U11293 ( .A1(n10281), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11169) );
  CLKBUF_X1 U11294 ( .A(n11999), .Z(n15014) );
  AND3_X2 U11295 ( .A1(n11418), .A2(n11417), .A3(n11914), .ZN(n13389) );
  AND2_X1 U11296 ( .A1(n9616), .A2(n10224), .ZN(n13252) );
  AND2_X1 U11297 ( .A1(n10370), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11215) );
  NAND2_X1 U11298 ( .A1(n11883), .A2(n11430), .ZN(n12069) );
  INV_X1 U11299 ( .A(n18072), .ZN(n12685) );
  INV_X1 U11300 ( .A(n18081), .ZN(n15557) );
  NAND2_X2 U11301 ( .A1(n10224), .A2(n10222), .ZN(n14089) );
  AND2_X1 U11302 ( .A1(n11434), .A2(n11433), .ZN(n11437) );
  INV_X2 U11303 ( .A(n16343), .ZN(n16347) );
  CLKBUF_X1 U11304 ( .A(n10210), .Z(n20132) );
  NAND2_X1 U11305 ( .A1(n10210), .A2(n10213), .ZN(n10218) );
  AND3_X1 U11306 ( .A1(n11430), .A2(n11446), .A3(n19131), .ZN(n9779) );
  AND2_X2 U11307 ( .A1(n10222), .A2(n20122), .ZN(n11320) );
  NAND2_X2 U11308 ( .A1(n9841), .A2(n10224), .ZN(n11312) );
  INV_X1 U11309 ( .A(n11422), .ZN(n11446) );
  NOR2_X1 U11310 ( .A1(n11422), .A2(n11420), .ZN(n11421) );
  AOI211_X1 U11311 ( .C1(n16813), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n12481), .B(n12480), .ZN(n12482) );
  CLKBUF_X1 U11312 ( .A(n11934), .Z(n9602) );
  CLKBUF_X3 U11313 ( .A(n11440), .Z(n12321) );
  NOR2_X2 U11314 ( .A1(n12587), .A2(n12586), .ZN(n18716) );
  INV_X1 U11315 ( .A(n10224), .ZN(n9584) );
  AND3_X1 U11316 ( .A1(n10058), .A2(n10057), .A3(n10042), .ZN(n10027) );
  NAND4_X1 U11317 ( .A1(n10145), .A2(n10144), .A3(n10143), .A4(n10142), .ZN(
        n10212) );
  AND4_X1 U11318 ( .A1(n10130), .A2(n10129), .A3(n10128), .A4(n10127), .ZN(
        n10145) );
  AND4_X1 U11319 ( .A1(n10159), .A2(n10158), .A3(n10157), .A4(n10156), .ZN(
        n10166) );
  AND4_X1 U11320 ( .A1(n10149), .A2(n10148), .A3(n10147), .A4(n10146), .ZN(
        n10168) );
  AND4_X1 U11321 ( .A1(n10175), .A2(n10174), .A3(n10173), .A4(n10172), .ZN(
        n10187) );
  AND4_X1 U11322 ( .A1(n10080), .A2(n10079), .A3(n10078), .A4(n10077), .ZN(
        n10086) );
  INV_X2 U11323 ( .A(U214), .ZN(n16340) );
  OAI22_X1 U11324 ( .A1(n10260), .A2(n10726), .B1(n10999), .B2(n10900), .ZN(
        n10047) );
  AND4_X1 U11325 ( .A1(n10134), .A2(n10133), .A3(n10132), .A4(n10131), .ZN(
        n10144) );
  AND4_X1 U11326 ( .A1(n10153), .A2(n10152), .A3(n10151), .A4(n10150), .ZN(
        n10167) );
  AND4_X1 U11327 ( .A1(n10117), .A2(n10116), .A3(n10115), .A4(n10114), .ZN(
        n10118) );
  AND4_X1 U11328 ( .A1(n10084), .A2(n10083), .A3(n10082), .A4(n10081), .ZN(
        n10085) );
  AND4_X1 U11329 ( .A1(n10138), .A2(n10137), .A3(n10136), .A4(n10135), .ZN(
        n10143) );
  AND3_X1 U11330 ( .A1(n10181), .A2(n10180), .A3(n10179), .ZN(n10186) );
  NAND2_X2 U11331 ( .A1(n18658), .A2(n18591), .ZN(n18638) );
  AND3_X1 U11332 ( .A1(n11326), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11325), .ZN(n11329) );
  OR2_X1 U11333 ( .A1(n10260), .A2(n10125), .ZN(n10128) );
  BUF_X2 U11334 ( .A(n10126), .Z(n10999) );
  AOI21_X1 U11335 ( .B1(n18534), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12566), .ZN(n12572) );
  INV_X2 U11336 ( .A(n16381), .ZN(U215) );
  INV_X1 U11337 ( .A(n12427), .ZN(n15614) );
  CLKBUF_X2 U11338 ( .A(n12497), .Z(n15627) );
  CLKBUF_X1 U11339 ( .A(n10516), .Z(n10840) );
  INV_X1 U11340 ( .A(n10262), .ZN(n10154) );
  INV_X2 U11341 ( .A(n10882), .ZN(n9586) );
  INV_X1 U11342 ( .A(n10858), .ZN(n10952) );
  INV_X2 U11343 ( .A(n13853), .ZN(n9601) );
  BUF_X2 U11344 ( .A(n10267), .Z(n11012) );
  NAND2_X2 U11345 ( .A1(n12981), .A2(n10049), .ZN(n10262) );
  NAND2_X1 U11346 ( .A1(n10064), .A2(n10061), .ZN(n10260) );
  AND2_X2 U11347 ( .A1(n10064), .A2(n10063), .ZN(n10858) );
  AND2_X2 U11348 ( .A1(n13446), .A2(n10063), .ZN(n10849) );
  INV_X1 U11349 ( .A(n9623), .ZN(n9587) );
  AND2_X2 U11350 ( .A1(n10064), .A2(n10065), .ZN(n10601) );
  INV_X2 U11351 ( .A(n16383), .ZN(n16385) );
  OR2_X1 U11352 ( .A1(n18517), .A2(n12429), .ZN(n10015) );
  AND2_X2 U11353 ( .A1(n12968), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12967) );
  NAND2_X1 U11354 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18690), .ZN(
        n12428) );
  NAND2_X1 U11355 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18682), .ZN(
        n12429) );
  NAND2_X1 U11356 ( .A1(n12981), .A2(n10050), .ZN(n10087) );
  AND2_X2 U11357 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11531) );
  NOR2_X1 U11358 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13348) );
  AND2_X1 U11359 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13494) );
  INV_X1 U11360 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10873) );
  INV_X1 U11361 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10830) );
  NAND2_X1 U11362 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12430) );
  INV_X1 U11363 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10046) );
  NOR2_X2 U11364 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10065) );
  INV_X1 U11365 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18534) );
  AND2_X1 U11366 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10063) );
  OR2_X1 U11367 ( .A1(n10257), .A2(n10240), .ZN(n9589) );
  NAND2_X1 U11368 ( .A1(n12326), .A2(n12325), .ZN(n15003) );
  NAND2_X1 U11369 ( .A1(n9801), .A2(n9804), .ZN(n12326) );
  NAND2_X1 U11370 ( .A1(n9576), .A2(n11121), .ZN(n9590) );
  NAND2_X1 U11371 ( .A1(n13718), .A2(n11121), .ZN(n11123) );
  BUF_X1 U11372 ( .A(n20213), .Z(n9591) );
  XNOR2_X1 U11373 ( .A(n10332), .B(n9847), .ZN(n20213) );
  NOR3_X2 U11374 ( .A1(n16638), .A2(n17075), .A3(n15559), .ZN(n17020) );
  NOR4_X4 U11375 ( .A1(n16730), .A2(n16749), .A3(n17102), .A4(n17086), .ZN(
        n17089) );
  AND2_X4 U11376 ( .A1(n9771), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11477) );
  NAND2_X1 U11377 ( .A1(n11123), .A2(n9595), .ZN(n9592) );
  AND2_X2 U11378 ( .A1(n9592), .A2(n9593), .ZN(n13749) );
  OR2_X1 U11379 ( .A1(n9594), .A2(n15903), .ZN(n9593) );
  INV_X1 U11380 ( .A(n15902), .ZN(n9594) );
  AND2_X1 U11381 ( .A1(n11122), .A2(n15902), .ZN(n9595) );
  NAND2_X1 U11382 ( .A1(n10211), .A2(n9577), .ZN(n10215) );
  AND2_X2 U11383 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12968) );
  CLKBUF_X1 U11384 ( .A(n13151), .Z(n9596) );
  AND3_X1 U11385 ( .A1(n10071), .A2(n10070), .A3(n10069), .ZN(n10072) );
  OR2_X2 U11386 ( .A1(n10258), .A2(n20213), .ZN(n10335) );
  NOR2_X2 U11387 ( .A1(n11233), .A2(n12970), .ZN(n12367) );
  CLKBUF_X1 U11388 ( .A(n10231), .Z(n12961) );
  INV_X1 U11389 ( .A(n12961), .ZN(n11218) );
  CLKBUF_X1 U11390 ( .A(n13749), .Z(n9597) );
  NOR2_X2 U11391 ( .A1(n10477), .A2(n13534), .ZN(n13537) );
  OR2_X2 U11392 ( .A1(n14120), .A2(n10012), .ZN(n14108) );
  CLKBUF_X1 U11393 ( .A(n13586), .Z(n9598) );
  BUF_X1 U11394 ( .A(n15451), .Z(n9599) );
  INV_X1 U11395 ( .A(n11498), .ZN(n9600) );
  XNOR2_X1 U11396 ( .A(n11701), .B(n13600), .ZN(n13586) );
  AND2_X1 U11397 ( .A1(n19119), .A2(n13368), .ZN(n14757) );
  NAND2_X1 U11398 ( .A1(n13368), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11422) );
  NAND2_X1 U11399 ( .A1(n13368), .A2(n11521), .ZN(n11934) );
  NAND3_X2 U11400 ( .A1(n11459), .A2(n11419), .A3(n11448), .ZN(n9771) );
  AND2_X2 U11401 ( .A1(n10463), .A2(n10462), .ZN(n10430) );
  AND2_X2 U11402 ( .A1(n9771), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9609) );
  NAND2_X2 U11403 ( .A1(n13001), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11082) );
  OAI21_X2 U11404 ( .B1(n11070), .B2(n9982), .A(n11074), .ZN(n13001) );
  OAI211_X1 U11405 ( .C1(n9761), .C2(n11489), .A(n9760), .B(n9758), .ZN(n12898) );
  NAND2_X1 U11406 ( .A1(n11489), .A2(n11492), .ZN(n18929) );
  AND2_X2 U11407 ( .A1(n11439), .A2(n11438), .ZN(n11455) );
  INV_X1 U11408 ( .A(n10160), .ZN(n9604) );
  NAND2_X1 U11409 ( .A1(n11391), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11392) );
  NAND2_X2 U11410 ( .A1(n12798), .A2(n11737), .ZN(n11442) );
  INV_X1 U11411 ( .A(n9726), .ZN(n13679) );
  AND2_X1 U11412 ( .A1(n10257), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10332) );
  OR2_X2 U11413 ( .A1(n10220), .A2(n13018), .ZN(n10257) );
  NAND2_X4 U11414 ( .A1(n9728), .A2(n9727), .ZN(n13675) );
  NAND2_X2 U11415 ( .A1(n14514), .A2(n11139), .ZN(n14474) );
  AND2_X2 U11416 ( .A1(n10227), .A2(n10219), .ZN(n12751) );
  NAND2_X4 U11417 ( .A1(n11393), .A2(n11392), .ZN(n13368) );
  INV_X1 U11418 ( .A(n15017), .ZN(n9611) );
  INV_X1 U11419 ( .A(n15017), .ZN(n9612) );
  INV_X1 U11420 ( .A(n15017), .ZN(n9613) );
  NAND2_X1 U11422 ( .A1(n13389), .A2(n11421), .ZN(n15017) );
  NAND3_X2 U11423 ( .A1(n10124), .A2(n10123), .A3(n10045), .ZN(n10209) );
  AND2_X1 U11424 ( .A1(n12967), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10268) );
  AND2_X2 U11425 ( .A1(n12967), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9623) );
  NOR2_X1 U11426 ( .A1(n12649), .A2(n12648), .ZN(n9615) );
  INV_X1 U11427 ( .A(n10222), .ZN(n9616) );
  INV_X1 U11428 ( .A(n10262), .ZN(n9617) );
  NAND2_X1 U11429 ( .A1(n12981), .A2(n10050), .ZN(n9618) );
  INV_X2 U11430 ( .A(n15059), .ZN(n9803) );
  AND3_X1 U11431 ( .A1(n10211), .A2(n10233), .A3(n9840), .ZN(n12840) );
  AND2_X2 U11432 ( .A1(n9768), .A2(n9803), .ZN(n9802) );
  NAND2_X2 U11433 ( .A1(n12030), .A2(n12805), .ZN(n11459) );
  XNOR2_X2 U11434 ( .A(n11086), .B(n20071), .ZN(n13467) );
  NAND2_X2 U11435 ( .A1(n13152), .A2(n11085), .ZN(n11086) );
  AOI21_X1 U11436 ( .B1(n11467), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11476), .ZN(n11943) );
  NAND2_X2 U11437 ( .A1(n11455), .A2(n11447), .ZN(n11467) );
  AND3_X4 U11439 ( .A1(n9751), .A2(n9800), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11409) );
  NAND2_X2 U11440 ( .A1(n11900), .A2(n11934), .ZN(n12038) );
  OAI21_X2 U11441 ( .B1(n12288), .B2(n11814), .A(n18893), .ZN(n11701) );
  NAND3_X2 U11442 ( .A1(n11427), .A2(n11425), .A3(n11426), .ZN(n9989) );
  OR2_X4 U11443 ( .A1(n14847), .A2(n11503), .ZN(n19389) );
  AND2_X1 U11444 ( .A1(n11523), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11611) );
  NOR2_X4 U11445 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13332) );
  OAI21_X2 U11446 ( .B1(n15079), .B2(n15081), .A(n15080), .ZN(n15059) );
  NAND2_X2 U11447 ( .A1(n15098), .A2(n11840), .ZN(n15079) );
  OAI211_X2 U11448 ( .C1(n15003), .C2(n15002), .A(n15001), .B(n15000), .ZN(
        n15009) );
  AND2_X2 U11449 ( .A1(n13736), .A2(n10005), .ZN(n13769) );
  NOR2_X4 U11450 ( .A1(n13656), .A2(n13744), .ZN(n13736) );
  OAI21_X2 U11451 ( .B1(n15192), .B2(n11830), .A(n11829), .ZN(n15308) );
  OAI21_X2 U11452 ( .B1(n15451), .B2(n15454), .A(n15452), .ZN(n15192) );
  AND2_X2 U11453 ( .A1(n14182), .A2(n10001), .ZN(n14131) );
  NOR2_X4 U11454 ( .A1(n14248), .A2(n14250), .ZN(n14182) );
  CLKBUF_X1 U11455 ( .A(n10511), .Z(n9620) );
  AND3_X4 U11456 ( .A1(n9751), .A2(n13343), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11349) );
  OR2_X1 U11457 ( .A1(n11414), .A2(n11737), .ZN(n11402) );
  NOR2_X1 U11458 ( .A1(n12680), .A2(n12679), .ZN(n12566) );
  OAI22_X1 U11459 ( .A1(n18682), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n20885), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12571) );
  NAND2_X1 U11460 ( .A1(n13083), .A2(n13082), .ZN(n13142) );
  NAND2_X1 U11461 ( .A1(n9738), .A2(n13240), .ZN(n9737) );
  OAI21_X1 U11462 ( .B1(n12044), .B2(n12037), .A(n19884), .ZN(n11438) );
  INV_X1 U11463 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9800) );
  INV_X1 U11464 ( .A(n9742), .ZN(n9741) );
  OAI21_X1 U11465 ( .B1(n12999), .B2(n12116), .A(n13037), .ZN(n9742) );
  NAND2_X1 U11466 ( .A1(n10232), .A2(n12961), .ZN(n10253) );
  INV_X1 U11467 ( .A(n10245), .ZN(n10232) );
  NOR2_X1 U11468 ( .A1(n9876), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10048) );
  CLKBUF_X1 U11469 ( .A(n10316), .Z(n11032) );
  INV_X1 U11470 ( .A(n10423), .ZN(n10422) );
  NOR2_X1 U11471 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12996), .ZN(
        n10049) );
  NOR2_X1 U11472 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10050) );
  AND2_X1 U11473 ( .A1(n13468), .A2(n20054), .ZN(n9963) );
  INV_X1 U11474 ( .A(n11087), .ZN(n9965) );
  AND2_X1 U11475 ( .A1(n11087), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9966) );
  INV_X1 U11476 ( .A(n12966), .ZN(n13028) );
  OAI21_X1 U11477 ( .B1(n20772), .B2(n16008), .A(n13448), .ZN(n20096) );
  INV_X1 U11478 ( .A(n15739), .ZN(n13448) );
  NAND2_X1 U11479 ( .A1(n11424), .A2(n13675), .ZN(n9726) );
  INV_X1 U11480 ( .A(n13674), .ZN(n9944) );
  NAND2_X1 U11481 ( .A1(n9823), .A2(n11475), .ZN(n9822) );
  INV_X1 U11482 ( .A(n11474), .ZN(n9823) );
  AND2_X1 U11483 ( .A1(n12249), .A2(n12248), .ZN(n14985) );
  OR2_X1 U11484 ( .A1(n14791), .A2(n11791), .ZN(n15105) );
  AND2_X1 U11485 ( .A1(n9666), .A2(n15486), .ZN(n9992) );
  NAND2_X1 U11486 ( .A1(n9750), .A2(n13432), .ZN(n9749) );
  INV_X1 U11487 ( .A(n14824), .ZN(n9750) );
  INV_X1 U11488 ( .A(n12112), .ZN(n12232) );
  NAND2_X1 U11489 ( .A1(n11475), .A2(n11474), .ZN(n9761) );
  NAND2_X1 U11490 ( .A1(n12078), .A2(n19119), .ZN(n12112) );
  AND2_X1 U11491 ( .A1(n12077), .A2(n19883), .ZN(n12078) );
  CLKBUF_X1 U11492 ( .A(n12030), .Z(n12031) );
  NAND2_X1 U11493 ( .A1(n12795), .A2(n19883), .ZN(n13081) );
  NAND2_X1 U11494 ( .A1(n9987), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9986) );
  NAND2_X1 U11495 ( .A1(n9985), .A2(n11530), .ZN(n9984) );
  NAND2_X1 U11496 ( .A1(n11871), .A2(n11870), .ZN(n11910) );
  NAND2_X1 U11497 ( .A1(n9784), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9783) );
  NAND2_X1 U11498 ( .A1(n9782), .A2(n11530), .ZN(n9781) );
  NAND2_X1 U11499 ( .A1(n11372), .A2(n13115), .ZN(n11379) );
  NAND2_X1 U11500 ( .A1(n11377), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11378) );
  AND2_X1 U11501 ( .A1(n12035), .A2(n13675), .ZN(n11914) );
  NAND2_X1 U11502 ( .A1(n18533), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12679) );
  INV_X1 U11503 ( .A(n12689), .ZN(n9774) );
  AOI21_X1 U11504 ( .B1(n12572), .B2(n12571), .A(n12570), .ZN(n12684) );
  OR2_X1 U11505 ( .A1(n10012), .A2(n12413), .ZN(n10011) );
  OR3_X1 U11506 ( .A1(n14128), .A2(n9873), .A3(n9872), .ZN(n9871) );
  INV_X1 U11507 ( .A(n12414), .ZN(n9872) );
  NAND2_X1 U11508 ( .A1(n13469), .A2(n11087), .ZN(n11096) );
  INV_X1 U11509 ( .A(n10212), .ZN(n13016) );
  NAND2_X1 U11510 ( .A1(n11213), .A2(n11212), .ZN(n11217) );
  INV_X1 U11511 ( .A(n12366), .ZN(n11214) );
  NAND2_X1 U11512 ( .A1(n11386), .A2(n13115), .ZN(n11393) );
  NAND2_X1 U11513 ( .A1(n11753), .A2(n12077), .ZN(n11854) );
  INV_X1 U11514 ( .A(n16236), .ZN(n12850) );
  AND2_X1 U11515 ( .A1(n18737), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13076) );
  AND4_X1 U11516 ( .A1(n11610), .A2(n11609), .A3(n11608), .A4(n11607), .ZN(
        n11616) );
  AND4_X1 U11517 ( .A1(n11601), .A2(n11600), .A3(n11599), .A4(n11598), .ZN(
        n11618) );
  NAND2_X1 U11518 ( .A1(n15146), .A2(n15147), .ZN(n15136) );
  NAND2_X1 U11519 ( .A1(n9736), .A2(n9734), .ZN(n13598) );
  NAND2_X1 U11520 ( .A1(n13599), .A2(n9732), .ZN(n9735) );
  INV_X1 U11521 ( .A(n13412), .ZN(n9732) );
  INV_X1 U11522 ( .A(n19695), .ZN(n19452) );
  OR2_X1 U11523 ( .A1(n16723), .A2(n16482), .ZN(n9910) );
  OR2_X1 U11524 ( .A1(n18729), .A2(n18062), .ZN(n16412) );
  OAI21_X1 U11525 ( .B1(n18523), .B2(n9778), .A(n15658), .ZN(n15762) );
  AND2_X1 U11526 ( .A1(n17307), .A2(n16410), .ZN(n9778) );
  NAND2_X1 U11527 ( .A1(n17920), .A2(n17608), .ZN(n9906) );
  AOI21_X1 U11528 ( .B1(n11196), .B2(n11195), .A(n11194), .ZN(n11205) );
  CLKBUF_X1 U11529 ( .A(n10601), .Z(n11044) );
  AND2_X1 U11530 ( .A1(n10404), .A2(n10403), .ZN(n10431) );
  NOR2_X1 U11531 ( .A1(n9981), .A2(n15892), .ZN(n9980) );
  AND2_X1 U11532 ( .A1(n14470), .A2(n9718), .ZN(n9981) );
  AND2_X1 U11533 ( .A1(n10494), .A2(n10493), .ZN(n10503) );
  OR2_X1 U11534 ( .A1(n10279), .A2(n10278), .ZN(n11076) );
  OR2_X1 U11535 ( .A1(n10361), .A2(n10360), .ZN(n11066) );
  NOR2_X1 U11536 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20088), .ZN(
        n11208) );
  OAI21_X1 U11537 ( .B1(n10252), .B2(n10228), .A(n10223), .ZN(n10238) );
  AND2_X1 U11538 ( .A1(n12947), .A2(n10226), .ZN(n10239) );
  NOR2_X1 U11539 ( .A1(n9876), .A2(n10259), .ZN(n9850) );
  NOR2_X1 U11540 ( .A1(n10059), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10060) );
  OAI21_X1 U11541 ( .B1(n11888), .B2(n12321), .A(n9806), .ZN(n11638) );
  NAND2_X1 U11542 ( .A1(n12321), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n9806) );
  NAND2_X1 U11543 ( .A1(n11539), .A2(n19119), .ZN(n9752) );
  OR2_X1 U11544 ( .A1(n11592), .A2(n11591), .ZN(n12094) );
  NOR2_X1 U11545 ( .A1(n18089), .A2(n17111), .ZN(n12687) );
  NOR2_X1 U11546 ( .A1(n9841), .A2(n10210), .ZN(n9840) );
  NAND2_X1 U11547 ( .A1(n14109), .A2(n10013), .ZN(n10012) );
  INV_X1 U11548 ( .A(n14121), .ZN(n10013) );
  OR2_X1 U11549 ( .A1(n14692), .A2(n10259), .ZN(n11023) );
  INV_X1 U11550 ( .A(n14261), .ZN(n10762) );
  NOR2_X1 U11551 ( .A1(n13550), .A2(n13659), .ZN(n9996) );
  INV_X1 U11552 ( .A(n13549), .ZN(n9997) );
  NAND2_X1 U11553 ( .A1(n10233), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10653) );
  AND2_X1 U11554 ( .A1(n10032), .A2(n9979), .ZN(n9978) );
  NOR2_X1 U11555 ( .A1(n9980), .A2(n9582), .ZN(n9976) );
  INV_X1 U11556 ( .A(n9980), .ZN(n9979) );
  INV_X1 U11557 ( .A(n14252), .ZN(n9886) );
  AND2_X1 U11558 ( .A1(n14256), .A2(n14262), .ZN(n9887) );
  INV_X1 U11559 ( .A(n11317), .ZN(n9866) );
  INV_X1 U11560 ( .A(n11310), .ZN(n11299) );
  NAND2_X1 U11561 ( .A1(n14087), .A2(n13105), .ZN(n11310) );
  INV_X1 U11562 ( .A(n13474), .ZN(n11247) );
  OR2_X1 U11563 ( .A1(n12914), .A2(n14089), .ZN(n12357) );
  NAND2_X1 U11564 ( .A1(n13107), .A2(n11241), .ZN(n13474) );
  NOR2_X1 U11565 ( .A1(n20127), .A2(n10259), .ZN(n11064) );
  OR2_X1 U11566 ( .A1(n10260), .A2(n10684), .ZN(n10173) );
  OR2_X1 U11567 ( .A1(n10126), .A2(n10113), .ZN(n10117) );
  NAND2_X1 U11568 ( .A1(n9603), .A2(n10259), .ZN(n10387) );
  AND3_X1 U11569 ( .A1(n12941), .A2(n11231), .A3(n11221), .ZN(n12918) );
  INV_X1 U11570 ( .A(n13434), .ZN(n15708) );
  NOR2_X1 U11571 ( .A1(n11859), .A2(n11858), .ZN(n12320) );
  NAND2_X1 U11572 ( .A1(n11785), .A2(n9644), .ZN(n11834) );
  NOR2_X1 U11573 ( .A1(n9812), .A2(n11777), .ZN(n9811) );
  INV_X1 U11574 ( .A(n11784), .ZN(n9812) );
  NAND2_X1 U11575 ( .A1(n11785), .A2(n11784), .ZN(n11807) );
  NOR2_X1 U11576 ( .A1(n9815), .A2(n11796), .ZN(n9814) );
  INV_X1 U11577 ( .A(n11770), .ZN(n9815) );
  NAND2_X1 U11578 ( .A1(n11757), .A2(n13425), .ZN(n11768) );
  INV_X1 U11579 ( .A(n12108), .ZN(n11697) );
  AND2_X1 U11580 ( .A1(n13401), .A2(n16183), .ZN(n9787) );
  AND2_X2 U11581 ( .A1(n11529), .A2(n11530), .ZN(n13876) );
  INV_X1 U11582 ( .A(n13958), .ZN(n13987) );
  AND2_X1 U11583 ( .A1(n14940), .A2(n12263), .ZN(n9748) );
  AND4_X1 U11584 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n11617) );
  NOR2_X1 U11585 ( .A1(n11855), .A2(n15070), .ZN(n11856) );
  INV_X1 U11586 ( .A(n14894), .ZN(n9788) );
  AND2_X1 U11587 ( .A1(n13697), .A2(n9703), .ZN(n14766) );
  INV_X1 U11588 ( .A(n15341), .ZN(n9744) );
  INV_X1 U11589 ( .A(n15182), .ZN(n9721) );
  NOR2_X1 U11590 ( .A1(n15424), .A2(n9797), .ZN(n9796) );
  INV_X1 U11591 ( .A(n13579), .ZN(n9797) );
  INV_X1 U11592 ( .A(n15471), .ZN(n9763) );
  NAND2_X1 U11593 ( .A1(n12287), .A2(n12286), .ZN(n12289) );
  INV_X1 U11594 ( .A(n11471), .ZN(n11472) );
  AND2_X1 U11595 ( .A1(n11531), .A2(n11532), .ZN(n13828) );
  AND2_X1 U11596 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11532) );
  OAI21_X1 U11597 ( .B1(n12934), .B2(n12933), .A(n9672), .ZN(n9731) );
  NAND2_X1 U11598 ( .A1(n12900), .A2(n12899), .ZN(n13072) );
  NAND2_X1 U11599 ( .A1(n12898), .A2(n13076), .ZN(n12900) );
  NOR2_X1 U11600 ( .A1(n11518), .A2(n13057), .ZN(n11519) );
  NOR2_X1 U11601 ( .A1(n12426), .A2(n12425), .ZN(n12470) );
  NOR2_X1 U11602 ( .A1(n12426), .A2(n16773), .ZN(n12497) );
  AND3_X1 U11603 ( .A1(n17633), .A2(n9634), .A3(n9925), .ZN(n16424) );
  NOR2_X1 U11604 ( .A1(n17596), .A2(n9926), .ZN(n9925) );
  NAND2_X1 U11605 ( .A1(n10031), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9926) );
  INV_X1 U11606 ( .A(n9900), .ZN(n9899) );
  OAI21_X1 U11607 ( .B1(n12532), .B2(n9901), .A(n17988), .ZN(n9900) );
  NOR2_X1 U11608 ( .A1(n17233), .A2(n12526), .ZN(n12530) );
  NAND2_X1 U11609 ( .A1(n17535), .A2(n17521), .ZN(n12545) );
  NAND2_X1 U11610 ( .A1(n12507), .A2(n12702), .ZN(n12535) );
  NAND2_X1 U11611 ( .A1(n12534), .A2(n17666), .ZN(n12537) );
  NAND2_X1 U11612 ( .A1(n15650), .A2(n15649), .ZN(n16407) );
  NOR2_X1 U11613 ( .A1(n15555), .A2(n15554), .ZN(n15656) );
  OR3_X1 U11614 ( .A1(n20766), .A2(n13619), .A3(n13618), .ZN(n14217) );
  AND2_X1 U11615 ( .A1(n9687), .A2(n10002), .ZN(n10001) );
  INV_X1 U11616 ( .A(n14148), .ZN(n10002) );
  NAND2_X1 U11617 ( .A1(n14193), .A2(n9641), .ZN(n10008) );
  NOR2_X1 U11618 ( .A1(n10650), .A2(n14211), .ZN(n10655) );
  OR2_X1 U11619 ( .A1(n13008), .A2(n19901), .ZN(n12790) );
  NOR2_X1 U11620 ( .A1(n11158), .A2(n9955), .ZN(n9954) );
  INV_X1 U11621 ( .A(n14571), .ZN(n9955) );
  AND2_X1 U11622 ( .A1(n9631), .A2(n14402), .ZN(n14382) );
  NAND2_X1 U11623 ( .A1(n20028), .A2(n20027), .ZN(n20026) );
  INV_X1 U11624 ( .A(n9966), .ZN(n9960) );
  NAND2_X1 U11625 ( .A1(n9962), .A2(n9964), .ZN(n9961) );
  NAND2_X1 U11626 ( .A1(n13469), .A2(n9966), .ZN(n9957) );
  NOR2_X1 U11627 ( .A1(n20093), .A2(n13503), .ZN(n20343) );
  AND2_X1 U11628 ( .A1(n20565), .A2(n20101), .ZN(n20433) );
  NOR2_X1 U11629 ( .A1(n13479), .A2(n20095), .ZN(n20504) );
  INV_X1 U11630 ( .A(n20480), .ZN(n20342) );
  NAND2_X1 U11631 ( .A1(n10259), .A2(n20096), .ZN(n20257) );
  AND2_X1 U11632 ( .A1(n12031), .A2(n12032), .ZN(n13378) );
  NAND2_X1 U11633 ( .A1(n14737), .A2(n9638), .ZN(n14740) );
  NAND2_X1 U11634 ( .A1(n11854), .A2(n11790), .ZN(n11785) );
  NAND2_X1 U11635 ( .A1(n11767), .A2(n9814), .ZN(n11799) );
  NAND2_X1 U11636 ( .A1(n11753), .A2(n9817), .ZN(n11756) );
  NAND2_X1 U11637 ( .A1(n14878), .A2(n14013), .ZN(n9934) );
  NOR2_X1 U11638 ( .A1(n13144), .A2(n9937), .ZN(n9936) );
  INV_X1 U11639 ( .A(n13140), .ZN(n9937) );
  AND2_X1 U11640 ( .A1(n9637), .A2(n9747), .ZN(n9746) );
  INV_X1 U11641 ( .A(n14955), .ZN(n9747) );
  NAND2_X1 U11642 ( .A1(n9948), .A2(n9947), .ZN(n9946) );
  INV_X1 U11643 ( .A(n16103), .ZN(n9947) );
  AND2_X1 U11644 ( .A1(n9688), .A2(n13513), .ZN(n9945) );
  INV_X1 U11645 ( .A(n12049), .ZN(n12829) );
  NAND2_X1 U11646 ( .A1(n11359), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9727) );
  NAND2_X1 U11647 ( .A1(n11354), .A2(n11530), .ZN(n9728) );
  NAND2_X1 U11648 ( .A1(n14737), .A2(n9889), .ZN(n15044) );
  AND2_X1 U11649 ( .A1(n9638), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9889) );
  NAND2_X1 U11650 ( .A1(n14737), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14738) );
  NAND2_X1 U11651 ( .A1(n14732), .A2(n9645), .ZN(n14736) );
  NAND2_X1 U11652 ( .A1(n14732), .A2(n9636), .ZN(n14713) );
  AND2_X1 U11653 ( .A1(n14732), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14734) );
  OR3_X1 U11654 ( .A1(n12306), .A2(n12300), .A3(n16199), .ZN(n12307) );
  NAND2_X1 U11655 ( .A1(n11941), .A2(n11940), .ZN(n9792) );
  NAND2_X1 U11656 ( .A1(n9792), .A2(n9791), .ZN(n13572) );
  AND2_X1 U11657 ( .A1(n11945), .A2(n11950), .ZN(n9791) );
  INV_X1 U11658 ( .A(n13569), .ZN(n11950) );
  OR3_X1 U11659 ( .A1(n12323), .A2(n12300), .A3(n15232), .ZN(n15001) );
  AND2_X1 U11660 ( .A1(n15105), .A2(n11792), .ZN(n15167) );
  AND2_X1 U11661 ( .A1(n15417), .A2(n15181), .ZN(n15103) );
  AND3_X1 U11662 ( .A1(n12195), .A2(n12194), .A3(n12193), .ZN(n14808) );
  OR2_X1 U11663 ( .A1(n14823), .A2(n9749), .ZN(n14809) );
  INV_X1 U11664 ( .A(n15502), .ZN(n9993) );
  AND3_X1 U11665 ( .A1(n12164), .A2(n12163), .A3(n12162), .ZN(n14824) );
  INV_X1 U11666 ( .A(n12289), .ZN(n12292) );
  NAND2_X1 U11667 ( .A1(n11731), .A2(n12232), .ZN(n12113) );
  NAND2_X1 U11668 ( .A1(n13564), .A2(n13597), .ZN(n9827) );
  AND3_X1 U11669 ( .A1(n12107), .A2(n12106), .A3(n12105), .ZN(n13412) );
  AND2_X1 U11670 ( .A1(n11933), .A2(n12850), .ZN(n12316) );
  OR2_X1 U11671 ( .A1(n12389), .A2(n11932), .ZN(n11933) );
  NAND2_X1 U11672 ( .A1(n18945), .A2(n13076), .ZN(n12797) );
  NOR2_X1 U11673 ( .A1(n12048), .A2(n12047), .ZN(n13354) );
  AND2_X1 U11674 ( .A1(n11414), .A2(n11927), .ZN(n11415) );
  AND2_X1 U11675 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19519) );
  AND2_X1 U11676 ( .A1(n19281), .A2(n19851), .ZN(n19690) );
  NAND2_X1 U11677 ( .A1(n12397), .A2(n12396), .ZN(n19695) );
  NAND2_X1 U11678 ( .A1(n12395), .A2(n12394), .ZN(n12396) );
  NAND2_X1 U11679 ( .A1(n12393), .A2(n12392), .ZN(n12397) );
  AOI21_X1 U11680 ( .B1(n12684), .B2(n12682), .A(n12681), .ZN(n18498) );
  NOR2_X1 U11681 ( .A1(n16441), .A2(n16738), .ZN(n16434) );
  OAI21_X1 U11682 ( .B1(n15656), .B2(n15558), .A(n18711), .ZN(n15761) );
  NOR3_X1 U11683 ( .A1(n15557), .A2(n17185), .A3(n15556), .ZN(n15558) );
  NOR2_X1 U11684 ( .A1(n17366), .A2(n9919), .ZN(n12694) );
  NAND2_X1 U11685 ( .A1(n9921), .A2(n9920), .ZN(n9919) );
  INV_X1 U11686 ( .A(n9922), .ZN(n9921) );
  AND2_X1 U11687 ( .A1(n17447), .A2(n9648), .ZN(n17368) );
  NOR2_X1 U11688 ( .A1(n17511), .A2(n17512), .ZN(n17487) );
  NOR2_X1 U11689 ( .A1(n12540), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12541) );
  NAND2_X1 U11690 ( .A1(n17668), .A2(n17667), .ZN(n17666) );
  NOR2_X1 U11691 ( .A1(n12437), .A2(n12436), .ZN(n15689) );
  NAND2_X2 U11692 ( .A1(n12540), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17920) );
  NOR2_X1 U11693 ( .A1(n15657), .A2(n18520), .ZN(n18523) );
  INV_X1 U11694 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18563) );
  NAND2_X1 U11695 ( .A1(n12930), .A2(n12791), .ZN(n20766) );
  INV_X1 U11696 ( .A(n14290), .ZN(n19999) );
  AND2_X1 U11697 ( .A1(n11236), .A2(n13012), .ZN(n20003) );
  INV_X1 U11698 ( .A(n19999), .ZN(n14297) );
  AND2_X2 U11699 ( .A1(n12371), .A2(n13012), .ZN(n14365) );
  OAI21_X1 U11700 ( .B1(n13008), .B2(n12913), .A(n12370), .ZN(n12371) );
  AND2_X1 U11701 ( .A1(n13238), .A2(n20011), .ZN(n20009) );
  XNOR2_X1 U11702 ( .A(n12352), .B(n12351), .ZN(n14086) );
  XNOR2_X1 U11703 ( .A(n11321), .B(n14088), .ZN(n14550) );
  CLKBUF_X1 U11704 ( .A(n13647), .Z(n13648) );
  NAND2_X1 U11705 ( .A1(n10344), .A2(n9845), .ZN(n10347) );
  NAND2_X1 U11706 ( .A1(n20218), .A2(n20342), .ZN(n20260) );
  NOR2_X1 U11707 ( .A1(n12802), .A2(n16236), .ZN(n19878) );
  INV_X1 U11708 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19883) );
  NAND2_X1 U11709 ( .A1(n12389), .A2(n12388), .ZN(n12757) );
  INV_X1 U11710 ( .A(n19861), .ZN(n19413) );
  XNOR2_X1 U11711 ( .A(n15010), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15238) );
  NAND2_X1 U11712 ( .A1(n12398), .A2(n19094), .ZN(n12408) );
  NAND2_X1 U11713 ( .A1(n15010), .A2(n12330), .ZN(n12391) );
  AND2_X1 U11714 ( .A1(n19100), .A2(n12762), .ZN(n19089) );
  INV_X1 U11715 ( .A(n19102), .ZN(n19094) );
  INV_X1 U11716 ( .A(n19091), .ZN(n16169) );
  OAI21_X1 U11717 ( .B1(n16023), .B2(n16204), .A(n12345), .ZN(n12346) );
  NOR2_X1 U11718 ( .A1(n12344), .A2(n12404), .ZN(n12345) );
  XNOR2_X1 U11719 ( .A(n9724), .B(n15111), .ZN(n15339) );
  NAND2_X1 U11720 ( .A1(n9725), .A2(n15120), .ZN(n9724) );
  NAND2_X1 U11721 ( .A1(n15122), .A2(n15119), .ZN(n9725) );
  INV_X1 U11722 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19865) );
  INV_X1 U11723 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19857) );
  INV_X1 U11724 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20880) );
  INV_X1 U11725 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19842) );
  NAND2_X1 U11726 ( .A1(n18711), .A2(n18498), .ZN(n17305) );
  XNOR2_X1 U11727 ( .A(n16434), .B(n9914), .ZN(n9913) );
  INV_X1 U11728 ( .A(n16435), .ZN(n9914) );
  NAND2_X1 U11729 ( .A1(n16582), .A2(n9918), .ZN(n16536) );
  NAND2_X1 U11730 ( .A1(n16723), .A2(n17443), .ZN(n9918) );
  NAND2_X1 U11731 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16782), .ZN(n16774) );
  AND2_X1 U11732 ( .A1(n18094), .A2(n16909), .ZN(n16894) );
  INV_X1 U11733 ( .A(n17117), .ZN(n17113) );
  NOR2_X1 U11734 ( .A1(n17365), .A2(n17186), .ZN(n17181) );
  AND2_X1 U11735 ( .A1(n17244), .A2(n9776), .ZN(n17224) );
  NOR2_X1 U11736 ( .A1(n17106), .A2(n9777), .ZN(n9776) );
  NAND2_X1 U11737 ( .A1(n15763), .A2(n17244), .ZN(n17239) );
  INV_X1 U11738 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18675) );
  INV_X1 U11739 ( .A(n10431), .ZN(n9838) );
  AND2_X1 U11740 ( .A1(n11167), .A2(n11166), .ZN(n11179) );
  AND2_X1 U11741 ( .A1(n10243), .A2(n10246), .ZN(n10226) );
  AND3_X1 U11742 ( .A1(n11509), .A2(n11499), .A3(n11500), .ZN(n9754) );
  NOR2_X1 U11743 ( .A1(n11517), .A2(n11494), .ZN(n9755) );
  INV_X1 U11744 ( .A(n19111), .ZN(n11553) );
  INV_X1 U11745 ( .A(n11215), .ZN(n11171) );
  OR2_X1 U11746 ( .A1(n10402), .A2(n10401), .ZN(n11106) );
  NAND2_X1 U11747 ( .A1(n9967), .A2(n10241), .ZN(n10305) );
  NAND2_X1 U11748 ( .A1(n9969), .A2(n9968), .ZN(n9967) );
  NOR2_X1 U11749 ( .A1(n9875), .A2(n10259), .ZN(n9968) );
  AND4_X1 U11750 ( .A1(n10251), .A2(n10250), .A3(n10246), .A4(n10249), .ZN(
        n10255) );
  NAND2_X1 U11751 ( .A1(n11200), .A2(n11063), .ZN(n11211) );
  INV_X1 U11752 ( .A(n10198), .ZN(n10954) );
  AOI22_X1 U11753 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10516), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10130) );
  OR2_X1 U11754 ( .A1(n10126), .A2(n10975), .ZN(n10091) );
  AOI22_X1 U11755 ( .A1(n10273), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10198), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10100) );
  INV_X1 U11756 ( .A(n10260), .ZN(n10511) );
  OR2_X1 U11757 ( .A1(n10385), .A2(n10384), .ZN(n11107) );
  NAND2_X1 U11758 ( .A1(n9680), .A2(n11854), .ZN(n11851) );
  AND2_X1 U11759 ( .A1(n11916), .A2(n11521), .ZN(n11430) );
  AND2_X1 U11760 ( .A1(n11921), .A2(n13675), .ZN(n11443) );
  NAND2_X1 U11761 ( .A1(n11423), .A2(n11737), .ZN(n11432) );
  INV_X1 U11762 ( .A(n15615), .ZN(n16815) );
  NOR2_X1 U11763 ( .A1(n17226), .A2(n12508), .ZN(n12507) );
  NOR2_X1 U11764 ( .A1(n17734), .A2(n12509), .ZN(n12710) );
  INV_X1 U11765 ( .A(n10210), .ZN(n11078) );
  NOR2_X1 U11766 ( .A1(n14170), .A2(n10004), .ZN(n10003) );
  INV_X1 U11767 ( .A(n14183), .ZN(n10004) );
  INV_X1 U11768 ( .A(n14260), .ZN(n10000) );
  INV_X1 U11769 ( .A(n14275), .ZN(n10009) );
  INV_X1 U11770 ( .A(n14286), .ZN(n10677) );
  INV_X1 U11771 ( .A(n13770), .ZN(n10010) );
  AND3_X1 U11772 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A3(n10471), .ZN(n10495) );
  INV_X1 U11773 ( .A(n10653), .ZN(n10669) );
  NAND2_X1 U11774 ( .A1(n14110), .A2(n9874), .ZN(n9873) );
  INV_X1 U11775 ( .A(n14139), .ZN(n9874) );
  NAND2_X1 U11776 ( .A1(n11144), .A2(n10032), .ZN(n9853) );
  NAND2_X1 U11777 ( .A1(n11148), .A2(n15892), .ZN(n9854) );
  INV_X1 U11778 ( .A(n13740), .ZN(n9870) );
  OR2_X1 U11779 ( .A1(n10492), .A2(n10491), .ZN(n11126) );
  NAND2_X1 U11780 ( .A1(n11255), .A2(n9880), .ZN(n9879) );
  INV_X1 U11781 ( .A(n13557), .ZN(n9880) );
  AND3_X1 U11782 ( .A1(n10299), .A2(n10298), .A3(n10297), .ZN(n10302) );
  INV_X1 U11783 ( .A(n11128), .ZN(n11133) );
  NAND2_X1 U11784 ( .A1(n10463), .A2(n10462), .ZN(n10470) );
  XNOR2_X1 U11785 ( .A(n10470), .B(n13503), .ZN(n11088) );
  NAND2_X1 U11786 ( .A1(n11210), .A2(n11209), .ZN(n12366) );
  OR2_X1 U11787 ( .A1(n11207), .A2(n11206), .ZN(n11210) );
  OR2_X1 U11788 ( .A1(n11211), .A2(n12366), .ZN(n11212) );
  NAND2_X1 U11789 ( .A1(n9849), .A2(n9848), .ZN(n9847) );
  AOI21_X1 U11790 ( .B1(n10240), .B2(n9850), .A(n10256), .ZN(n9848) );
  NAND2_X1 U11791 ( .A1(n10257), .A2(n9850), .ZN(n9849) );
  OAI211_X1 U11792 ( .C1(n10176), .C2(n10952), .A(n10184), .B(n10177), .ZN(
        n9862) );
  NAND2_X1 U11793 ( .A1(n10182), .A2(n10178), .ZN(n9861) );
  NOR2_X1 U11794 ( .A1(n10068), .A2(n10067), .ZN(n10069) );
  INV_X1 U11795 ( .A(n11070), .ZN(n20095) );
  INV_X1 U11796 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20505) );
  NAND2_X1 U11797 ( .A1(n12094), .A2(n9808), .ZN(n9807) );
  NOR2_X1 U11798 ( .A1(n15075), .A2(n9891), .ZN(n9890) );
  NOR2_X1 U11799 ( .A1(n9818), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n9817) );
  INV_X1 U11800 ( .A(n11740), .ZN(n9818) );
  NAND2_X1 U11801 ( .A1(n12823), .A2(n12798), .ZN(n13958) );
  INV_X1 U11802 ( .A(n14884), .ZN(n9941) );
  NOR2_X1 U11803 ( .A1(n9950), .A2(n9949), .ZN(n9948) );
  INV_X1 U11804 ( .A(n14915), .ZN(n9949) );
  NAND2_X1 U11805 ( .A1(n9951), .A2(n16106), .ZN(n9950) );
  INV_X1 U11806 ( .A(n14923), .ZN(n9951) );
  OR2_X1 U11807 ( .A1(n12761), .A2(n12112), .ZN(n12083) );
  NOR2_X1 U11808 ( .A1(n18831), .A2(n9895), .ZN(n9894) );
  INV_X1 U11809 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n9895) );
  NOR2_X1 U11810 ( .A1(n19099), .A2(n9898), .ZN(n9897) );
  INV_X1 U11811 ( .A(n14719), .ZN(n9896) );
  INV_X1 U11812 ( .A(n12094), .ZN(n12274) );
  INV_X1 U11813 ( .A(n11851), .ZN(n15006) );
  AND2_X1 U11814 ( .A1(n14706), .A2(n14872), .ZN(n9799) );
  NOR2_X1 U11815 ( .A1(n14902), .A2(n9790), .ZN(n9789) );
  INV_X1 U11816 ( .A(n14910), .ZN(n9790) );
  INV_X1 U11817 ( .A(n15353), .ZN(n9745) );
  INV_X1 U11818 ( .A(n15107), .ZN(n15109) );
  AND3_X1 U11819 ( .A1(n12221), .A2(n12220), .A3(n12219), .ZN(n15429) );
  AND2_X1 U11820 ( .A1(n18809), .A2(n11814), .ZN(n11825) );
  NAND2_X1 U11821 ( .A1(n12299), .A2(n12298), .ZN(n12306) );
  NOR2_X1 U11822 ( .A1(n12293), .A2(n16198), .ZN(n9831) );
  OR2_X1 U11823 ( .A1(n11690), .A2(n11689), .ZN(n12108) );
  AND3_X2 U11824 ( .A1(n11595), .A2(n11596), .A3(n12282), .ZN(n12281) );
  OR2_X1 U11825 ( .A1(n11538), .A2(n11537), .ZN(n12100) );
  INV_X1 U11826 ( .A(n11595), .ZN(n9820) );
  NAND2_X1 U11827 ( .A1(n13987), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13070) );
  NAND2_X1 U11828 ( .A1(n13987), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12902) );
  NOR2_X1 U11829 ( .A1(n12035), .A2(n13368), .ZN(n11414) );
  OAI22_X1 U11830 ( .A1(n11422), .A2(n11910), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12393) );
  INV_X1 U11831 ( .A(n12473), .ZN(n12588) );
  OR2_X1 U11832 ( .A1(n18517), .A2(n12430), .ZN(n12472) );
  NOR2_X1 U11833 ( .A1(n12429), .A2(n16773), .ZN(n12473) );
  OR2_X1 U11834 ( .A1(n12431), .A2(n16773), .ZN(n10022) );
  NOR2_X1 U11835 ( .A1(n12426), .A2(n12428), .ZN(n12515) );
  NOR2_X1 U11836 ( .A1(n9924), .A2(n17728), .ZN(n9920) );
  NAND2_X1 U11837 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9922) );
  NAND2_X1 U11838 ( .A1(n17633), .A2(n9634), .ZN(n16634) );
  OAI22_X1 U11839 ( .A1(n18690), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12680) );
  AND2_X1 U11840 ( .A1(n12573), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12575) );
  NAND2_X1 U11841 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18672), .ZN(
        n12431) );
  OR2_X1 U11842 ( .A1(n14692), .A2(n11232), .ZN(n12966) );
  OR2_X1 U11843 ( .A1(n10531), .A2(n10527), .ZN(n10565) );
  INV_X1 U11844 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19927) );
  AND2_X1 U11845 ( .A1(n11281), .A2(n11280), .ZN(n13774) );
  NOR2_X1 U11846 ( .A1(n14208), .A2(n13774), .ZN(n14282) );
  OR2_X1 U11847 ( .A1(n14366), .A2(n10207), .ZN(n12383) );
  AND2_X1 U11848 ( .A1(n13015), .A2(n12358), .ZN(n12913) );
  OR2_X1 U11849 ( .A1(n12357), .A2(n20687), .ZN(n12358) );
  INV_X1 U11850 ( .A(n20091), .ZN(n20089) );
  AND2_X1 U11851 ( .A1(n20613), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12353) );
  NOR2_X1 U11852 ( .A1(n10993), .A2(n14395), .ZN(n10994) );
  NAND2_X1 U11853 ( .A1(n10994), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13621) );
  AOI21_X1 U11854 ( .B1(n11020), .B2(n14399), .A(n10992), .ZN(n14109) );
  NAND2_X1 U11855 ( .A1(n10895), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10896) );
  OR2_X1 U11856 ( .A1(n10896), .A2(n14152), .ZN(n10922) );
  INV_X1 U11857 ( .A(n10868), .ZN(n10895) );
  OR2_X1 U11858 ( .A1(n10828), .A2(n10827), .ZN(n10868) );
  OR2_X1 U11859 ( .A1(n15776), .A2(n11055), .ZN(n10807) );
  AND2_X1 U11860 ( .A1(n10754), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10755) );
  AND2_X1 U11861 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n10755), .ZN(
        n10802) );
  OR2_X1 U11862 ( .A1(n15862), .A2(n11055), .ZN(n10760) );
  NOR2_X1 U11863 ( .A1(n10718), .A2(n10717), .ZN(n10754) );
  INV_X1 U11864 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10717) );
  CLKBUF_X1 U11865 ( .A(n14260), .Z(n14266) );
  NAND2_X1 U11866 ( .A1(n10699), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10718) );
  NOR2_X1 U11867 ( .A1(n10678), .A2(n15818), .ZN(n10699) );
  NAND2_X1 U11868 ( .A1(n10655), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10678) );
  CLKBUF_X1 U11869 ( .A(n13770), .Z(n13771) );
  NAND2_X1 U11870 ( .A1(n10594), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10650) );
  AND2_X1 U11871 ( .A1(n10006), .A2(n9696), .ZN(n10005) );
  OR2_X1 U11872 ( .A1(n9685), .A2(n10007), .ZN(n10006) );
  AND2_X1 U11873 ( .A1(n10569), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10570) );
  CLKBUF_X1 U11874 ( .A(n13656), .Z(n13657) );
  NAND2_X1 U11875 ( .A1(n10507), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10531) );
  NOR2_X1 U11876 ( .A1(n10472), .A2(n13529), .ZN(n10471) );
  AND2_X1 U11877 ( .A1(n11159), .A2(n14572), .ZN(n9952) );
  NOR3_X1 U11878 ( .A1(n9626), .A2(n14128), .A3(n9873), .ZN(n14111) );
  NOR3_X1 U11879 ( .A1(n9626), .A2(n14128), .A3(n14139), .ZN(n14127) );
  AND2_X1 U11880 ( .A1(n14269), .A2(n9885), .ZN(n14173) );
  AND2_X1 U11881 ( .A1(n9639), .A2(n9712), .ZN(n9885) );
  NAND2_X1 U11882 ( .A1(n9674), .A2(n9979), .ZN(n9977) );
  NAND2_X1 U11883 ( .A1(n14269), .A2(n9639), .ZN(n14254) );
  OR2_X1 U11884 ( .A1(n15922), .A2(n14645), .ZN(n14636) );
  NAND2_X1 U11885 ( .A1(n14269), .A2(n9887), .ZN(n14258) );
  AND2_X1 U11886 ( .A1(n14269), .A2(n14262), .ZN(n14264) );
  OR2_X1 U11887 ( .A1(n14195), .A2(n14196), .ZN(n14268) );
  AND2_X1 U11888 ( .A1(n14282), .A2(n14281), .ZN(n14284) );
  OR3_X1 U11889 ( .A1(n14294), .A2(n14207), .A3(n14206), .ZN(n14208) );
  NAND2_X1 U11890 ( .A1(n9869), .A2(n9867), .ZN(n14294) );
  NOR2_X1 U11891 ( .A1(n9693), .A2(n9868), .ZN(n9867) );
  INV_X1 U11892 ( .A(n14291), .ZN(n9868) );
  NOR2_X1 U11893 ( .A1(n15970), .A2(n9693), .ZN(n14292) );
  NAND2_X1 U11894 ( .A1(n9869), .A2(n11268), .ZN(n15972) );
  AND2_X1 U11895 ( .A1(n11137), .A2(n10023), .ZN(n9983) );
  AND2_X1 U11896 ( .A1(n11261), .A2(n11260), .ZN(n13552) );
  NOR2_X1 U11897 ( .A1(n13545), .A2(n9877), .ZN(n13688) );
  NAND2_X1 U11898 ( .A1(n9878), .A2(n13552), .ZN(n9877) );
  INV_X1 U11899 ( .A(n9879), .ZN(n9878) );
  NOR2_X1 U11900 ( .A1(n13545), .A2(n9879), .ZN(n13560) );
  OR2_X1 U11901 ( .A1(n13545), .A2(n13540), .ZN(n13558) );
  NAND2_X1 U11902 ( .A1(n13543), .A2(n13542), .ZN(n13545) );
  NAND2_X1 U11903 ( .A1(n12994), .A2(n10259), .ZN(n11227) );
  AND2_X1 U11904 ( .A1(n11247), .A2(n9863), .ZN(n13543) );
  NOR2_X1 U11905 ( .A1(n13457), .A2(n13473), .ZN(n9863) );
  NAND2_X1 U11906 ( .A1(n11247), .A2(n11246), .ZN(n9865) );
  NAND2_X1 U11907 ( .A1(n20061), .A2(n20076), .ZN(n15950) );
  NAND2_X1 U11908 ( .A1(n13034), .A2(n13028), .ZN(n20057) );
  NOR2_X1 U11909 ( .A1(n13024), .A2(n15706), .ZN(n13722) );
  NAND2_X1 U11910 ( .A1(n10464), .A2(n10470), .ZN(n13478) );
  OR2_X1 U11911 ( .A1(n10463), .A2(n10462), .ZN(n10464) );
  BUF_X1 U11912 ( .A(n10456), .Z(n13631) );
  AND3_X1 U11913 ( .A1(n12926), .A2(n12925), .A3(n12924), .ZN(n13434) );
  NOR2_X1 U11914 ( .A1(n10109), .A2(n10020), .ZN(n10124) );
  AND2_X1 U11915 ( .A1(n20097), .A2(n20096), .ZN(n20142) );
  NAND2_X1 U11916 ( .A1(n13479), .A2(n20095), .ZN(n20480) );
  INV_X1 U11917 ( .A(n20424), .ZN(n20567) );
  NOR2_X1 U11918 ( .A1(n20093), .A2(n9839), .ZN(n20539) );
  INV_X1 U11919 ( .A(n13503), .ZN(n9839) );
  NOR2_X2 U11920 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20624) );
  INV_X1 U11921 ( .A(n12914), .ZN(n10188) );
  NAND2_X1 U11922 ( .A1(n11832), .A2(n11831), .ZN(n11841) );
  INV_X1 U11923 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n9810) );
  NAND2_X1 U11924 ( .A1(n11785), .A2(n9811), .ZN(n11813) );
  AND2_X1 U11925 ( .A1(n11810), .A2(n11809), .ZN(n18780) );
  NAND2_X1 U11926 ( .A1(n11767), .A2(n9690), .ZN(n11790) );
  NAND2_X1 U11927 ( .A1(n11767), .A2(n11770), .ZN(n11797) );
  NAND2_X1 U11928 ( .A1(n11753), .A2(n11740), .ZN(n11752) );
  OR2_X1 U11929 ( .A1(n12231), .A2(n12230), .ZN(n13578) );
  OR2_X1 U11930 ( .A1(n12161), .A2(n12160), .ZN(n18969) );
  NOR2_X1 U11931 ( .A1(n9938), .A2(n13992), .ZN(n14876) );
  NOR2_X1 U11932 ( .A1(n14883), .A2(n9939), .ZN(n9938) );
  NOR2_X1 U11933 ( .A1(n14882), .A2(n14884), .ZN(n14883) );
  NAND2_X1 U11934 ( .A1(n14908), .A2(n10017), .ZN(n14900) );
  OR2_X1 U11935 ( .A1(n13709), .A2(n13708), .ZN(n13711) );
  AND2_X1 U11936 ( .A1(n12804), .A2(n12803), .ZN(n13131) );
  OAI21_X1 U11937 ( .B1(n12208), .B2(n20815), .A(n12087), .ZN(n12812) );
  AND2_X1 U11938 ( .A1(n12086), .A2(n12085), .ZN(n12087) );
  CLKBUF_X1 U11939 ( .A(n11442), .Z(n12817) );
  NOR2_X1 U11940 ( .A1(n14746), .A2(n12880), .ZN(n19063) );
  INV_X1 U11941 ( .A(n12745), .ZN(n19103) );
  OAI21_X1 U11942 ( .B1(n12744), .B2(n12743), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12745) );
  XNOR2_X1 U11943 ( .A(n14709), .B(n14708), .ZN(n15022) );
  NOR2_X1 U11944 ( .A1(n15046), .A2(n15029), .ZN(n15027) );
  NAND2_X1 U11945 ( .A1(n14705), .A2(n9798), .ZN(n15011) );
  AND2_X1 U11946 ( .A1(n9799), .A2(n12027), .ZN(n9798) );
  OR2_X1 U11947 ( .A1(n15044), .A2(n15043), .ZN(n15046) );
  AND2_X1 U11948 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n12403), .ZN(
        n14737) );
  AND2_X1 U11949 ( .A1(n14731), .A2(n12402), .ZN(n14732) );
  NOR2_X1 U11950 ( .A1(n14729), .A2(n15169), .ZN(n14731) );
  INV_X1 U11951 ( .A(n14715), .ZN(n14730) );
  NAND2_X1 U11952 ( .A1(n14730), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14729) );
  AND2_X1 U11953 ( .A1(n14722), .A2(n9893), .ZN(n14726) );
  AND2_X1 U11954 ( .A1(n9628), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9893) );
  NAND2_X1 U11955 ( .A1(n14722), .A2(n9628), .ZN(n14727) );
  INV_X1 U11956 ( .A(n13423), .ZN(n9786) );
  NAND2_X1 U11957 ( .A1(n13161), .A2(n9683), .ZN(n14830) );
  NAND2_X1 U11958 ( .A1(n14722), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14725) );
  NOR2_X1 U11959 ( .A1(n14720), .A2(n16189), .ZN(n14716) );
  AND2_X1 U11960 ( .A1(n9896), .A2(n9630), .ZN(n14721) );
  NAND2_X1 U11961 ( .A1(n9896), .A2(n9897), .ZN(n14717) );
  NOR2_X1 U11962 ( .A1(n14719), .A2(n19099), .ZN(n14718) );
  INV_X1 U11963 ( .A(n11488), .ZN(n11498) );
  NAND2_X1 U11964 ( .A1(n14941), .A2(n9715), .ZN(n15228) );
  AOI21_X1 U11965 ( .B1(n15039), .B2(n9719), .A(n9805), .ZN(n9804) );
  OAI211_X1 U11966 ( .C1(n15039), .C2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11856), .B(n9802), .ZN(n9801) );
  AND2_X1 U11967 ( .A1(n14705), .A2(n9799), .ZN(n12026) );
  NAND2_X1 U11968 ( .A1(n9768), .A2(n15069), .ZN(n9767) );
  NOR2_X1 U11969 ( .A1(n12300), .A2(n14744), .ZN(n15038) );
  XNOR2_X1 U11970 ( .A(n9766), .B(n9765), .ZN(n15051) );
  INV_X1 U11971 ( .A(n15038), .ZN(n9765) );
  NAND2_X1 U11972 ( .A1(n15315), .A2(n9789), .ZN(n14904) );
  AND2_X1 U11973 ( .A1(n9654), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9835) );
  INV_X1 U11974 ( .A(n14776), .ZN(n12003) );
  AND2_X1 U11975 ( .A1(n15358), .A2(n12311), .ZN(n15331) );
  NAND2_X1 U11976 ( .A1(n15421), .A2(n9653), .ZN(n15131) );
  NAND2_X1 U11977 ( .A1(n15152), .A2(n14919), .ZN(n15123) );
  NAND2_X1 U11978 ( .A1(n13697), .A2(n9684), .ZN(n15355) );
  NAND2_X1 U11979 ( .A1(n15104), .A2(n9720), .ZN(n9722) );
  NOR2_X1 U11980 ( .A1(n15106), .A2(n9721), .ZN(n9720) );
  AND2_X1 U11981 ( .A1(n9796), .A2(n9794), .ZN(n9793) );
  INV_X1 U11982 ( .A(n14784), .ZN(n9794) );
  NAND2_X1 U11983 ( .A1(n9795), .A2(n9796), .ZN(n14785) );
  NOR2_X1 U11984 ( .A1(n15425), .A2(n15424), .ZN(n15426) );
  NOR2_X1 U11985 ( .A1(n14823), .A2(n9694), .ZN(n13522) );
  NAND2_X1 U11986 ( .A1(n13522), .A2(n13523), .ZN(n15428) );
  OR2_X1 U11987 ( .A1(n18819), .A2(n11822), .ZN(n15193) );
  INV_X1 U11988 ( .A(n9730), .ZN(n9762) );
  NAND2_X1 U11989 ( .A1(n9994), .A2(n9992), .ZN(n15469) );
  AND2_X1 U11990 ( .A1(n12064), .A2(n15525), .ZN(n15507) );
  AND3_X1 U11991 ( .A1(n12134), .A2(n12133), .A3(n12132), .ZN(n13157) );
  CLKBUF_X1 U11992 ( .A(n13156), .Z(n15506) );
  NAND2_X1 U11993 ( .A1(n13145), .A2(n13166), .ZN(n13167) );
  NOR2_X1 U11994 ( .A1(n9737), .A2(n13412), .ZN(n9733) );
  OR2_X1 U11995 ( .A1(n16216), .A2(n12063), .ZN(n16196) );
  INV_X1 U11996 ( .A(n11464), .ZN(n9759) );
  XNOR2_X1 U11997 ( .A(n12810), .B(n12093), .ZN(n12934) );
  XNOR2_X1 U11998 ( .A(n12098), .B(n12097), .ZN(n13040) );
  XNOR2_X1 U11999 ( .A(n12901), .B(n12902), .ZN(n12827) );
  AOI21_X1 U12000 ( .B1(n18929), .B2(n13076), .A(n12825), .ZN(n12826) );
  XNOR2_X1 U12001 ( .A(n13072), .B(n13070), .ZN(n12906) );
  NOR2_X1 U12002 ( .A1(n19281), .A2(n19851), .ZN(n19414) );
  NOR2_X1 U12003 ( .A1(n19281), .A2(n19280), .ZN(n19832) );
  INV_X1 U12004 ( .A(n19832), .ZN(n19517) );
  INV_X1 U12005 ( .A(n12035), .ZN(n19131) );
  INV_X1 U12006 ( .A(n13675), .ZN(n19157) );
  NAND2_X1 U12007 ( .A1(n19695), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19158) );
  INV_X1 U12008 ( .A(n19518), .ZN(n19588) );
  INV_X1 U12009 ( .A(n19156), .ZN(n19150) );
  NOR2_X1 U12010 ( .A1(n19450), .A2(n19413), .ZN(n19625) );
  NOR2_X2 U12011 ( .A1(n19103), .A2(n19102), .ZN(n19155) );
  AND2_X1 U12012 ( .A1(n11910), .A2(n11875), .ZN(n13382) );
  NOR2_X1 U12013 ( .A1(n19757), .A2(n19491), .ZN(n13133) );
  INV_X1 U12014 ( .A(n11435), .ZN(n11418) );
  NOR2_X1 U12015 ( .A1(n18523), .A2(n16407), .ZN(n18497) );
  NOR2_X1 U12016 ( .A1(n16442), .A2(n16443), .ZN(n16441) );
  NOR2_X1 U12017 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16667), .ZN(n16647) );
  NOR2_X1 U12018 ( .A1(n17258), .A2(n17260), .ZN(n9772) );
  NAND3_X1 U12019 ( .A1(n12629), .A2(n12628), .A3(n12627), .ZN(n17111) );
  AOI211_X1 U12020 ( .C1(n17034), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n12626), .B(n12625), .ZN(n12627) );
  AOI21_X1 U12021 ( .B1(n15650), .B2(n18555), .A(n18714), .ZN(n17252) );
  NOR3_X1 U12022 ( .A1(n17366), .A2(n9922), .A3(n17728), .ZN(n16254) );
  NAND2_X1 U12023 ( .A1(n17368), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17366) );
  NOR2_X1 U12024 ( .A1(n17421), .A2(n9916), .ZN(n9915) );
  INV_X1 U12025 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n9916) );
  INV_X1 U12026 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17445) );
  NOR2_X1 U12027 ( .A1(n16420), .A2(n17445), .ZN(n17447) );
  INV_X1 U12028 ( .A(n17528), .ZN(n12691) );
  OAI21_X1 U12029 ( .B1(n17728), .B2(n17482), .A(n18204), .ZN(n17579) );
  AND3_X1 U12030 ( .A1(n17633), .A2(n9634), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17580) );
  NOR2_X1 U12031 ( .A1(n17662), .A2(n17663), .ZN(n17633) );
  NAND2_X1 U12032 ( .A1(n17693), .A2(n9669), .ZN(n9902) );
  NAND2_X1 U12033 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17686) );
  NOR2_X1 U12034 ( .A1(n18503), .A2(n18561), .ZN(n12728) );
  OR2_X1 U12035 ( .A1(n15744), .A2(n12556), .ZN(n12558) );
  INV_X1 U12036 ( .A(n12560), .ZN(n15744) );
  NAND2_X1 U12037 ( .A1(n12553), .A2(n17608), .ZN(n12554) );
  OR2_X1 U12038 ( .A1(n9907), .A2(n17639), .ZN(n16287) );
  NAND2_X1 U12039 ( .A1(n12548), .A2(n10040), .ZN(n12549) );
  NAND2_X1 U12040 ( .A1(n12545), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9905) );
  INV_X1 U12041 ( .A(n17521), .ZN(n16244) );
  NOR2_X1 U12042 ( .A1(n17639), .A2(n17920), .ZN(n17618) );
  XNOR2_X1 U12043 ( .A(n12537), .B(n12536), .ZN(n17648) );
  NAND2_X1 U12044 ( .A1(n17648), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17647) );
  XNOR2_X1 U12045 ( .A(n12527), .B(n12525), .ZN(n17705) );
  NAND2_X1 U12046 ( .A1(n12509), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12522) );
  AOI21_X1 U12047 ( .B1(n12684), .B2(n12683), .A(n15672), .ZN(n18499) );
  NOR2_X1 U12048 ( .A1(n15676), .A2(n15653), .ZN(n16288) );
  XNOR2_X1 U12049 ( .A(n17246), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17725) );
  NOR2_X1 U12050 ( .A1(n16407), .A2(n9773), .ZN(n18515) );
  AND2_X1 U12051 ( .A1(n12662), .A2(n18716), .ZN(n9773) );
  OR2_X1 U12052 ( .A1(n18517), .A2(n12431), .ZN(n10014) );
  NOR3_X1 U12053 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n18715), .ZN(n18398) );
  NOR2_X1 U12054 ( .A1(n12639), .A2(n12638), .ZN(n18072) );
  NOR2_X1 U12055 ( .A1(n12659), .A2(n12658), .ZN(n18076) );
  NOR2_X1 U12056 ( .A1(n12609), .A2(n12608), .ZN(n18081) );
  INV_X1 U12057 ( .A(n17111), .ZN(n18085) );
  INV_X1 U12058 ( .A(n18399), .ZN(n18300) );
  NOR2_X1 U12059 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18563), .ZN(n17489) );
  INV_X1 U12060 ( .A(n19103), .ZN(n19101) );
  NAND2_X1 U12061 ( .A1(n15738), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19901) );
  NOR2_X1 U12062 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20772) );
  AND2_X1 U12063 ( .A1(n14097), .A2(n14085), .ZN(n9883) );
  INV_X1 U12064 ( .A(n15838), .ZN(n19925) );
  OR2_X1 U12065 ( .A1(n13637), .A2(n13636), .ZN(n15838) );
  INV_X1 U12066 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15818) );
  INV_X1 U12067 ( .A(n19986), .ZN(n19928) );
  OR3_X1 U12068 ( .A1(n13637), .A2(n13629), .A3(n13628), .ZN(n19936) );
  INV_X1 U12069 ( .A(n19936), .ZN(n19982) );
  AND2_X1 U12070 ( .A1(n14217), .A2(n13635), .ZN(n19993) );
  INV_X1 U12071 ( .A(n19971), .ZN(n19983) );
  AND2_X1 U12072 ( .A1(n14217), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19986) );
  INV_X1 U12073 ( .A(n20003), .ZN(n14288) );
  OR2_X1 U12074 ( .A1(n12383), .A2(n20089), .ZN(n14326) );
  INV_X1 U12075 ( .A(n14323), .ZN(n14352) );
  INV_X1 U12076 ( .A(n14326), .ZN(n14354) );
  NAND2_X1 U12077 ( .A1(n14365), .A2(n12963), .ZN(n14364) );
  OR3_X1 U12078 ( .A1(n12930), .A2(n12929), .A3(n15754), .ZN(n13238) );
  INV_X2 U12079 ( .A(n20009), .ZN(n20007) );
  OR3_X1 U12080 ( .A1(n13254), .A2(n9616), .A3(n20687), .ZN(n13396) );
  XNOR2_X1 U12081 ( .A(n13622), .B(n14093), .ZN(n14377) );
  OR2_X1 U12082 ( .A1(n13621), .A2(n13620), .ZN(n13622) );
  INV_X1 U12083 ( .A(n14484), .ZN(n20025) );
  AND2_X1 U12084 ( .A1(n11061), .A2(n20624), .ZN(n20031) );
  AND2_X1 U12085 ( .A1(n14484), .A2(n11226), .ZN(n15889) );
  INV_X1 U12086 ( .A(n19908), .ZN(n20032) );
  OR2_X1 U12087 ( .A1(n12790), .A2(n15724), .ZN(n19908) );
  XNOR2_X1 U12088 ( .A(n14092), .B(n14091), .ZN(n14534) );
  XNOR2_X1 U12089 ( .A(n9855), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14568) );
  NAND2_X1 U12090 ( .A1(n9857), .A2(n9856), .ZN(n9855) );
  NAND2_X1 U12091 ( .A1(n14382), .A2(n15892), .ZN(n9857) );
  NOR3_X1 U12092 ( .A1(n20049), .A2(n13727), .A3(n13725), .ZN(n15983) );
  NAND2_X1 U12093 ( .A1(n20026), .A2(n11104), .ZN(n15912) );
  OR2_X1 U12094 ( .A1(n11227), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20065) );
  NAND2_X1 U12095 ( .A1(n9958), .A2(n9957), .ZN(n13525) );
  INV_X1 U12096 ( .A(n9961), .ZN(n9958) );
  AND2_X1 U12097 ( .A1(n13034), .A2(n13019), .ZN(n20062) );
  INV_X1 U12098 ( .A(n15950), .ZN(n20056) );
  INV_X1 U12099 ( .A(n20079), .ZN(n20048) );
  INV_X1 U12100 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20536) );
  INV_X1 U12101 ( .A(n20624), .ZN(n20622) );
  INV_X1 U12102 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20425) );
  NAND2_X1 U12104 ( .A1(n20251), .A2(n9845), .ZN(n9842) );
  NAND2_X1 U12105 ( .A1(n10346), .A2(n9844), .ZN(n9843) );
  NOR2_X1 U12106 ( .A1(n20251), .A2(n9845), .ZN(n9844) );
  NAND2_X1 U12107 ( .A1(n11089), .A2(n20093), .ZN(n20481) );
  INV_X1 U12108 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20088) );
  OAI21_X1 U12109 ( .B1(n13449), .B2(n16009), .A(n20257), .ZN(n20087) );
  OAI211_X1 U12110 ( .C1(n20108), .C2(n20613), .A(n20433), .B(n20104), .ZN(
        n20147) );
  OAI21_X1 U12111 ( .B1(n20275), .B2(n20259), .A(n20572), .ZN(n20278) );
  NAND2_X1 U12112 ( .A1(n20343), .A2(n20424), .ZN(n20372) );
  OAI211_X1 U12113 ( .C1(n20393), .C2(n20510), .A(n20433), .B(n20378), .ZN(
        n20396) );
  OAI211_X1 U12114 ( .C1(n20438), .C2(n20435), .A(n20434), .B(n20433), .ZN(
        n20470) );
  INV_X1 U12115 ( .A(n20426), .ZN(n20615) );
  INV_X1 U12116 ( .A(n20441), .ZN(n20629) );
  INV_X1 U12117 ( .A(n20449), .ZN(n20641) );
  INV_X1 U12118 ( .A(n20453), .ZN(n20647) );
  INV_X1 U12119 ( .A(n20461), .ZN(n20659) );
  NOR2_X2 U12120 ( .A1(n20619), .A2(n20567), .ZN(n20670) );
  INV_X1 U12121 ( .A(n20465), .ZN(n20665) );
  AND2_X1 U12122 ( .A1(n15734), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15738) );
  INV_X1 U12123 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20510) );
  CLKBUF_X1 U12124 ( .A(n20779), .Z(n20765) );
  OR2_X1 U12125 ( .A1(n12748), .A2(n12747), .ZN(n14746) );
  NOR2_X1 U12126 ( .A1(n11883), .A2(n11890), .ZN(n19872) );
  XNOR2_X1 U12127 ( .A(n15004), .B(n12322), .ZN(n16026) );
  OR3_X1 U12128 ( .A1(n19878), .A2(n19090), .A3(n14752), .ZN(n18873) );
  NAND2_X1 U12129 ( .A1(n11832), .A2(n9651), .ZN(n16071) );
  NAND2_X1 U12130 ( .A1(n11832), .A2(n9649), .ZN(n11842) );
  INV_X1 U12131 ( .A(n18950), .ZN(n18892) );
  INV_X1 U12132 ( .A(n18873), .ZN(n18936) );
  AND2_X1 U12133 ( .A1(n14748), .A2(n14747), .ZN(n18906) );
  XNOR2_X1 U12134 ( .A(n13137), .B(n13138), .ZN(n19450) );
  CLKBUF_X1 U12135 ( .A(n14742), .Z(n18901) );
  NOR2_X1 U12136 ( .A1(n14711), .A2(n18934), .ZN(n18949) );
  NOR2_X1 U12137 ( .A1(n9932), .A2(n14870), .ZN(n9931) );
  NAND2_X1 U12138 ( .A1(n9934), .A2(n14038), .ZN(n9933) );
  OR2_X1 U12139 ( .A1(n12205), .A2(n12204), .ZN(n13513) );
  OR2_X1 U12140 ( .A1(n12192), .A2(n12191), .ZN(n18963) );
  OR2_X1 U12141 ( .A1(n12180), .A2(n12179), .ZN(n18964) );
  OR2_X1 U12142 ( .A1(n12149), .A2(n12148), .ZN(n18970) );
  INV_X1 U12143 ( .A(n19851), .ZN(n19280) );
  AND2_X1 U12144 ( .A1(n12830), .A2(n12850), .ZN(n18988) );
  INV_X1 U12145 ( .A(n18984), .ZN(n18954) );
  NAND2_X1 U12146 ( .A1(n14976), .A2(n9637), .ZN(n14956) );
  AND2_X1 U12147 ( .A1(n14979), .A2(n13676), .ZN(n20782) );
  AND2_X1 U12148 ( .A1(n14979), .A2(n13680), .ZN(n20783) );
  NAND2_X1 U12149 ( .A1(n13141), .A2(n13140), .ZN(n13410) );
  INV_X1 U12150 ( .A(n14996), .ZN(n20791) );
  INV_X1 U12151 ( .A(n20787), .ZN(n18989) );
  NAND2_X1 U12152 ( .A1(n19049), .A2(n19880), .ZN(n19017) );
  CLKBUF_X1 U12153 ( .A(n19061), .Z(n19081) );
  INV_X1 U12154 ( .A(n19063), .ZN(n19086) );
  INV_X1 U12155 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16175) );
  INV_X1 U12156 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16189) );
  INV_X1 U12157 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19099) );
  NAND2_X1 U12158 ( .A1(n9792), .A2(n11945), .ZN(n13570) );
  INV_X1 U12159 ( .A(n16168), .ZN(n19095) );
  INV_X1 U12160 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12784) );
  INV_X1 U12161 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18930) );
  NAND2_X1 U12162 ( .A1(n12757), .A2(n12399), .ZN(n19100) );
  AND2_X1 U12163 ( .A1(n12390), .A2(n11420), .ZN(n19091) );
  NAND3_X1 U12164 ( .A1(n19837), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19695), 
        .ZN(n19102) );
  INV_X1 U12165 ( .A(n19100), .ZN(n16156) );
  AOI21_X1 U12166 ( .B1(n15238), .B2(n16192), .A(n9695), .ZN(n9780) );
  NAND2_X1 U12167 ( .A1(n15104), .A2(n15182), .ZN(n15168) );
  NOR2_X1 U12168 ( .A1(n14823), .A2(n14824), .ZN(n13433) );
  AND2_X1 U12169 ( .A1(n9994), .A2(n9666), .ZN(n15484) );
  NAND2_X1 U12170 ( .A1(n9994), .A2(n11750), .ZN(n15504) );
  NAND2_X1 U12171 ( .A1(n9740), .A2(n9743), .ZN(n13038) );
  NAND2_X1 U12172 ( .A1(n13000), .A2(n12999), .ZN(n9740) );
  OAI211_X1 U12173 ( .C1(n12295), .C2(n12293), .A(n9832), .B(n9833), .ZN(
        n15214) );
  NAND2_X1 U12174 ( .A1(n12292), .A2(n12293), .ZN(n9833) );
  OAI21_X1 U12175 ( .B1(n9825), .B2(n13565), .A(n9827), .ZN(n13592) );
  INV_X1 U12176 ( .A(n9826), .ZN(n9825) );
  NAND2_X1 U12177 ( .A1(n9663), .A2(n13490), .ZN(n13497) );
  NAND2_X1 U12178 ( .A1(n12316), .A2(n12029), .ZN(n15521) );
  NAND2_X1 U12179 ( .A1(n11486), .A2(n11485), .ZN(n11487) );
  INV_X1 U12180 ( .A(n11483), .ZN(n11486) );
  AND2_X1 U12181 ( .A1(n12316), .A2(n12072), .ZN(n16217) );
  INV_X1 U12182 ( .A(n15521), .ZN(n16218) );
  OR2_X1 U12183 ( .A1(n12901), .A2(n12800), .ZN(n19861) );
  AND2_X1 U12185 ( .A1(n13074), .A2(n12907), .ZN(n19281) );
  OR2_X1 U12186 ( .A1(n12906), .A2(n12905), .ZN(n12907) );
  OR3_X1 U12187 ( .A1(n19108), .A2(n19452), .A3(n19107), .ZN(n19163) );
  OAI21_X1 U12188 ( .B1(n19214), .B2(n19491), .A(n19218), .ZN(n19238) );
  OAI21_X1 U12189 ( .B1(n19295), .B2(n19294), .A(n19293), .ZN(n19319) );
  NAND2_X1 U12190 ( .A1(n19354), .A2(n19594), .ZN(n19353) );
  OAI21_X1 U12191 ( .B1(n19362), .B2(n19377), .A(n19695), .ZN(n19380) );
  OAI21_X1 U12192 ( .B1(n19356), .B2(n19489), .A(n19355), .ZN(n19378) );
  OAI21_X1 U12193 ( .B1(n19386), .B2(n19634), .A(n19385), .ZN(n19408) );
  OAI21_X1 U12194 ( .B1(n19444), .B2(n19418), .A(n19695), .ZN(n19447) );
  AND2_X1 U12195 ( .A1(n19383), .A2(n19690), .ZN(n19445) );
  OAI21_X1 U12196 ( .B1(n19496), .B2(n19511), .A(n19695), .ZN(n19514) );
  OAI21_X1 U12197 ( .B1(n19490), .B2(n19489), .A(n19488), .ZN(n19512) );
  NOR2_X2 U12198 ( .A1(n19518), .A2(n19517), .ZN(n19584) );
  NAND2_X1 U12199 ( .A1(n19625), .A2(n19594), .ZN(n19617) );
  INV_X1 U12200 ( .A(n19677), .ZN(n19629) );
  OAI21_X1 U12201 ( .B1(n19642), .B2(n19641), .A(n19640), .ZN(n19679) );
  NAND2_X1 U12202 ( .A1(n19588), .A2(n19594), .ZN(n19677) );
  AND2_X1 U12203 ( .A1(n19695), .A2(n19126), .ZN(n19708) );
  INV_X1 U12204 ( .A(n19748), .ZN(n19734) );
  NAND2_X1 U12205 ( .A1(n19588), .A2(n19690), .ZN(n19737) );
  INV_X1 U12206 ( .A(n19737), .ZN(n19744) );
  NAND2_X1 U12207 ( .A1(n19625), .A2(n19690), .ZN(n19748) );
  NOR2_X1 U12208 ( .A1(n19692), .A2(n19687), .ZN(n19742) );
  INV_X1 U12209 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n18737) );
  INV_X1 U12210 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19763) );
  NAND2_X1 U12211 ( .A1(n16501), .A2(n9911), .ZN(n9909) );
  NOR2_X1 U12212 ( .A1(n16493), .A2(n17419), .ZN(n16492) );
  NOR2_X1 U12213 ( .A1(n16501), .A2(n16738), .ZN(n16493) );
  NOR2_X2 U12214 ( .A1(n18554), .A2(n16412), .ZN(n16763) );
  NOR2_X1 U12215 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16529), .ZN(n16514) );
  NOR2_X1 U12216 ( .A1(n16535), .A2(n16738), .ZN(n16525) );
  NOR2_X1 U12217 ( .A1(n16536), .A2(n17483), .ZN(n16535) );
  NOR2_X1 U12218 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16589), .ZN(n16577) );
  NAND2_X1 U12219 ( .A1(n16723), .A2(n10036), .ZN(n16582) );
  INV_X1 U12220 ( .A(n16582), .ZN(n16595) );
  NOR2_X1 U12221 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16714), .ZN(n16705) );
  INV_X1 U12222 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16749) );
  INV_X1 U12223 ( .A(n16774), .ZN(n16759) );
  INV_X1 U12224 ( .A(n16768), .ZN(n16785) );
  INV_X1 U12225 ( .A(n16763), .ZN(n16781) );
  NAND2_X1 U12226 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16855), .ZN(n16846) );
  NAND2_X1 U12227 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16880), .ZN(n16868) );
  NAND3_X1 U12228 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n17089), .ZN(n17075) );
  INV_X2 U12229 ( .A(n17103), .ZN(n17097) );
  INV_X1 U12230 ( .A(n17085), .ZN(n17103) );
  NAND2_X1 U12231 ( .A1(n17126), .A2(n9655), .ZN(n17117) );
  INV_X1 U12232 ( .A(n17130), .ZN(n17126) );
  NAND2_X1 U12233 ( .A1(n17126), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n17125) );
  NOR2_X1 U12234 ( .A1(n17326), .A2(n17139), .ZN(n17134) );
  NAND2_X1 U12235 ( .A1(n17140), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17139) );
  NOR2_X1 U12236 ( .A1(n17180), .A2(n9775), .ZN(n17145) );
  NAND2_X1 U12237 ( .A1(n17145), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n17144) );
  NOR2_X1 U12238 ( .A1(n17315), .A2(n17168), .ZN(n17163) );
  INV_X1 U12239 ( .A(n17173), .ZN(n17169) );
  NAND2_X1 U12240 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17181), .ZN(n17180) );
  NOR2_X1 U12241 ( .A1(n17218), .A2(n17107), .ZN(n17108) );
  NOR2_X1 U12242 ( .A1(n12458), .A2(n12457), .ZN(n17233) );
  INV_X1 U12243 ( .A(n17248), .ZN(n17242) );
  NOR2_X2 U12244 ( .A1(n12649), .A2(n12648), .ZN(n18094) );
  OAI21_X1 U12245 ( .B1(n15762), .B2(n18561), .A(n9692), .ZN(n17244) );
  NOR2_X1 U12246 ( .A1(n15763), .A2(n17221), .ZN(n17248) );
  INV_X1 U12247 ( .A(n17239), .ZN(n17247) );
  CLKBUF_X1 U12248 ( .A(n17361), .Z(n17354) );
  OAI211_X1 U12249 ( .C1(n18716), .C2(n18717), .A(n17307), .B(n17306), .ZN(
        n17361) );
  NAND2_X1 U12250 ( .A1(n17447), .A2(n9635), .ZN(n17397) );
  NAND2_X1 U12251 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17528) );
  NOR2_X2 U12252 ( .A1(n15689), .A2(n17738), .ZN(n17615) );
  INV_X1 U12253 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17621) );
  INV_X1 U12254 ( .A(n17598), .ZN(n17646) );
  NOR2_X1 U12255 ( .A1(n12541), .A2(n9906), .ZN(n17638) );
  INV_X1 U12256 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17663) );
  NOR2_X1 U12257 ( .A1(n17686), .A2(n17700), .ZN(n17683) );
  NAND2_X1 U12258 ( .A1(n17675), .A2(n17674), .ZN(n17673) );
  NAND2_X1 U12259 ( .A1(n17693), .A2(n12532), .ZN(n17675) );
  NAND2_X1 U12260 ( .A1(n18300), .A2(n18398), .ZN(n18204) );
  INV_X1 U12261 ( .A(n17729), .ZN(n17719) );
  INV_X1 U12262 ( .A(n18204), .ZN(n18374) );
  INV_X1 U12263 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17728) );
  INV_X1 U12264 ( .A(n17739), .ZN(n17727) );
  NAND2_X1 U12265 ( .A1(n18716), .A2(n12728), .ZN(n17739) );
  INV_X1 U12266 ( .A(n9907), .ZN(n17384) );
  NOR2_X1 U12267 ( .A1(n16244), .A2(n17922), .ZN(n17870) );
  NOR2_X2 U12268 ( .A1(n15689), .A2(n18041), .ZN(n17936) );
  NAND2_X1 U12269 ( .A1(n18515), .A2(n15657), .ZN(n18532) );
  INV_X1 U12270 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18533) );
  INV_X1 U12271 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20885) );
  INV_X2 U12272 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16736) );
  AOI211_X1 U12273 ( .C1(n18711), .C2(n18538), .A(n18061), .B(n15660), .ZN(
        n18697) );
  INV_X1 U12274 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18504) );
  INV_X1 U12275 ( .A(n18717), .ZN(n18578) );
  INV_X1 U12276 ( .A(n16739), .ZN(n18569) );
  AND2_X2 U12277 ( .A1(n12381), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20091)
         );
  NAND2_X1 U12279 ( .A1(n9884), .A2(n9881), .ZN(P1_U2810) );
  OR2_X1 U12280 ( .A1(n14550), .A2(n19971), .ZN(n9884) );
  INV_X1 U12281 ( .A(n9882), .ZN(n9881) );
  OAI21_X1 U12282 ( .B1(n14086), .B2(n15810), .A(n9671), .ZN(n9882) );
  OR2_X1 U12283 ( .A1(n14550), .A2(n14298), .ZN(n11324) );
  OAI21_X1 U12284 ( .B1(n14305), .B2(n14297), .A(n12420), .ZN(P1_U2843) );
  AOI21_X1 U12285 ( .B1(n12419), .B2(n12418), .A(n12417), .ZN(n12420) );
  NOR2_X1 U12286 ( .A1(n20003), .A2(n12416), .ZN(n12417) );
  INV_X1 U12287 ( .A(n14564), .ZN(n12419) );
  NOR2_X1 U12288 ( .A1(n12410), .A2(n12409), .ZN(n12411) );
  NAND2_X1 U12289 ( .A1(n12408), .A2(n12407), .ZN(n12409) );
  OAI21_X1 U12290 ( .B1(n15339), .B2(n16168), .A(n15118), .ZN(P2_U2993) );
  INV_X1 U12291 ( .A(n16392), .ZN(n16387) );
  AOI211_X1 U12292 ( .C1(n16438), .C2(n16800), .A(n16430), .B(n16429), .ZN(
        n16431) );
  AOI21_X1 U12293 ( .B1(n9913), .B2(n16739), .A(n9912), .ZN(n16440) );
  OR2_X1 U12294 ( .A1(n16437), .A2(n16436), .ZN(n9912) );
  AND2_X1 U12295 ( .A1(n11522), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11565) );
  AND2_X1 U12296 ( .A1(n9643), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9624) );
  AND2_X4 U12297 ( .A1(n13332), .A2(n13343), .ZN(n11522) );
  AND4_X1 U12298 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n9625)
         );
  OR2_X1 U12299 ( .A1(n14157), .A2(n14145), .ZN(n9626) );
  AND2_X1 U12300 ( .A1(n11523), .A2(n11530), .ZN(n11646) );
  NAND2_X1 U12301 ( .A1(n11736), .A2(n9995), .ZN(n9994) );
  NAND2_X1 U12302 ( .A1(n14892), .A2(n9668), .ZN(n13964) );
  NAND2_X1 U12303 ( .A1(n10010), .A2(n10677), .ZN(n14274) );
  NAND2_X1 U12304 ( .A1(n14182), .A2(n14183), .ZN(n14169) );
  NAND2_X1 U12305 ( .A1(n14182), .A2(n9687), .ZN(n14147) );
  NAND2_X1 U12306 ( .A1(n13736), .A2(n9685), .ZN(n13764) );
  NAND2_X1 U12307 ( .A1(n16110), .A2(n9948), .ZN(n14913) );
  NAND2_X1 U12308 ( .A1(n9992), .A2(n9763), .ZN(n9627) );
  NOR2_X1 U12309 ( .A1(n14120), .A2(n10011), .ZN(n12352) );
  AND2_X1 U12310 ( .A1(n9894), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9628) );
  AND2_X1 U12311 ( .A1(n13407), .A2(n9708), .ZN(n9629) );
  AND2_X1 U12312 ( .A1(n9897), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9630) );
  INV_X1 U12313 ( .A(n11529), .ZN(n13854) );
  INV_X1 U12314 ( .A(n11104), .ZN(n9973) );
  AND2_X1 U12315 ( .A1(n14411), .A2(n14572), .ZN(n9631) );
  AND3_X1 U12316 ( .A1(n15237), .A2(n9780), .A3(n9676), .ZN(n9632) );
  AND2_X1 U12317 ( .A1(n9629), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n9633)
         );
  NAND2_X1 U12318 ( .A1(n9935), .A2(n13407), .ZN(n13159) );
  NAND2_X1 U12319 ( .A1(n13512), .A2(n13513), .ZN(n13671) );
  AND2_X1 U12320 ( .A1(n17593), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9634) );
  INV_X1 U12321 ( .A(n20251), .ZN(n9846) );
  OAI211_X1 U12322 ( .C1(n10346), .C2(n9846), .A(n9843), .B(n9842), .ZN(n12980) );
  INV_X1 U12323 ( .A(n16723), .ZN(n16738) );
  AND2_X1 U12324 ( .A1(n9624), .A2(n9915), .ZN(n9635) );
  AND2_X1 U12325 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9636) );
  AND2_X1 U12326 ( .A1(n9710), .A2(n14975), .ZN(n9637) );
  AND2_X1 U12327 ( .A1(n9890), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9638) );
  AND2_X1 U12328 ( .A1(n9887), .A2(n9886), .ZN(n9639) );
  AND2_X1 U12329 ( .A1(n9636), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9640) );
  AND2_X1 U12330 ( .A1(n10677), .A2(n10009), .ZN(n9641) );
  AND2_X1 U12331 ( .A1(n9811), .A2(n9810), .ZN(n9642) );
  AND2_X1 U12332 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n9643) );
  AND2_X1 U12333 ( .A1(n9642), .A2(n14917), .ZN(n9644) );
  AND2_X1 U12334 ( .A1(n9640), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9645) );
  INV_X1 U12335 ( .A(n13399), .ZN(n18978) );
  OR2_X1 U12336 ( .A1(n12131), .A2(n12130), .ZN(n13399) );
  AND2_X1 U12337 ( .A1(n9814), .A2(n9689), .ZN(n9646) );
  AND2_X1 U12338 ( .A1(n17409), .A2(n9911), .ZN(n9647) );
  AND2_X1 U12339 ( .A1(n9635), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9648) );
  NOR2_X1 U12340 ( .A1(n11865), .A2(n15071), .ZN(n15037) );
  INV_X1 U12341 ( .A(n15037), .ZN(n9805) );
  AND2_X1 U12342 ( .A1(n11831), .A2(n9714), .ZN(n9649) );
  INV_X1 U12343 ( .A(n14865), .ZN(n9932) );
  AND2_X1 U12344 ( .A1(n9649), .A2(n9809), .ZN(n9650) );
  AND2_X1 U12345 ( .A1(n9650), .A2(n16072), .ZN(n9651) );
  OR2_X1 U12346 ( .A1(n17639), .A2(n15750), .ZN(n9652) );
  AND2_X1 U12347 ( .A1(n12310), .A2(n12311), .ZN(n9653) );
  AND2_X1 U12348 ( .A1(n9653), .A2(n9836), .ZN(n9654) );
  AND2_X1 U12349 ( .A1(n9772), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n9655) );
  NAND4_X2 U12350 ( .A1(n11618), .A2(n11617), .A3(n11616), .A4(n10018), .ZN(
        n11814) );
  INV_X4 U12351 ( .A(n12472), .ZN(n16998) );
  INV_X1 U12352 ( .A(n17674), .ZN(n9901) );
  NAND2_X1 U12353 ( .A1(n9589), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10336) );
  INV_X1 U12354 ( .A(n11521), .ZN(n11420) );
  INV_X1 U12355 ( .A(n11349), .ZN(n13853) );
  NAND2_X1 U12356 ( .A1(n11736), .A2(n11735), .ZN(n15207) );
  AND2_X1 U12357 ( .A1(n10010), .A2(n9641), .ZN(n9656) );
  AND2_X1 U12358 ( .A1(n14182), .A2(n10003), .ZN(n14159) );
  NAND2_X1 U12359 ( .A1(n14976), .A2(n14975), .ZN(n14965) );
  NAND2_X1 U12360 ( .A1(n12308), .A2(n12307), .ZN(n15196) );
  AND2_X1 U12361 ( .A1(n10000), .A2(n10762), .ZN(n9657) );
  AND2_X1 U12362 ( .A1(n17126), .A2(n9772), .ZN(n9658) );
  OAI211_X1 U12363 ( .C1(n10336), .C2(n10059), .A(n10343), .B(n10342), .ZN(
        n10345) );
  AND2_X2 U12364 ( .A1(n11490), .A2(n11487), .ZN(n18945) );
  INV_X1 U12365 ( .A(n12116), .ZN(n9743) );
  AND2_X1 U12366 ( .A1(n11814), .A2(n12232), .ZN(n12116) );
  AND4_X1 U12367 ( .A1(n10101), .A2(n10044), .A3(n10100), .A4(n10099), .ZN(
        n9659) );
  OR2_X1 U12368 ( .A1(n9626), .A2(n9871), .ZN(n9660) );
  NAND2_X1 U12369 ( .A1(n11767), .A2(n9646), .ZN(n9661) );
  NAND2_X1 U12370 ( .A1(n10211), .A2(n20122), .ZN(n10221) );
  AND2_X1 U12371 ( .A1(n12546), .A2(n12544), .ZN(n9662) );
  NAND2_X1 U12372 ( .A1(n11138), .A2(n11137), .ZN(n13757) );
  AND2_X2 U12373 ( .A1(n9876), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10064) );
  AND2_X1 U12374 ( .A1(n9819), .A2(n12283), .ZN(n9663) );
  AOI21_X1 U12375 ( .B1(n11222), .B2(n11320), .A(n10225), .ZN(n10246) );
  AND4_X1 U12376 ( .A1(n11673), .A2(n11672), .A3(n11671), .A4(n11670), .ZN(
        n9664) );
  AND4_X1 U12377 ( .A1(n11712), .A2(n11711), .A3(n11710), .A4(n11709), .ZN(
        n9665) );
  NAND2_X1 U12378 ( .A1(n9841), .A2(n10211), .ZN(n10242) );
  INV_X1 U12379 ( .A(n12541), .ZN(n12542) );
  AND2_X1 U12380 ( .A1(n11750), .A2(n9993), .ZN(n9666) );
  AND2_X1 U12381 ( .A1(n11785), .A2(n9642), .ZN(n9667) );
  OR2_X1 U12382 ( .A1(n14898), .A2(n13937), .ZN(n9668) );
  AND2_X1 U12383 ( .A1(n12532), .A2(n9901), .ZN(n9669) );
  INV_X1 U12384 ( .A(n9837), .ZN(n15150) );
  NAND2_X1 U12385 ( .A1(n15421), .A2(n12310), .ZN(n9837) );
  INV_X1 U12386 ( .A(n9834), .ZN(n15090) );
  NAND2_X1 U12387 ( .A1(n15421), .A2(n9654), .ZN(n9834) );
  NAND2_X1 U12388 ( .A1(n18929), .A2(n13347), .ZN(n9670) );
  NOR2_X1 U12389 ( .A1(n14084), .A2(n9883), .ZN(n9671) );
  OR2_X1 U12390 ( .A1(n12810), .A2(n12093), .ZN(n9672) );
  AND2_X1 U12391 ( .A1(n14705), .A2(n14706), .ZN(n14704) );
  NAND2_X1 U12392 ( .A1(n10330), .A2(n9998), .ZN(n9673) );
  AND2_X1 U12393 ( .A1(n11498), .A2(n18945), .ZN(n11504) );
  INV_X1 U12394 ( .A(n11504), .ZN(n11510) );
  NAND2_X1 U12395 ( .A1(n11152), .A2(n9582), .ZN(n9674) );
  AND2_X1 U12396 ( .A1(n14886), .A2(n14887), .ZN(n14705) );
  AND2_X1 U12397 ( .A1(n12293), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9675) );
  OR2_X1 U12398 ( .A1(n16101), .A2(n15521), .ZN(n9676) );
  AND2_X1 U12399 ( .A1(n9831), .A2(n12290), .ZN(n9677) );
  AND2_X1 U12400 ( .A1(n11152), .A2(n10025), .ZN(n9678) );
  NAND2_X1 U12401 ( .A1(n11113), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9679) );
  NAND2_X1 U12402 ( .A1(n12074), .A2(n12090), .ZN(n12208) );
  INV_X1 U12403 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11530) );
  OR2_X1 U12404 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n16071), .ZN(n9680) );
  NOR2_X1 U12405 ( .A1(n14921), .A2(n14923), .ZN(n14922) );
  AND2_X1 U12406 ( .A1(n12542), .A2(n9906), .ZN(n17535) );
  INV_X1 U12407 ( .A(n9602), .ZN(n9808) );
  NAND2_X1 U12408 ( .A1(n13697), .A2(n15366), .ZN(n15352) );
  NAND2_X1 U12409 ( .A1(n17447), .A2(n9624), .ZN(n9917) );
  OR2_X1 U12410 ( .A1(n9626), .A2(n14139), .ZN(n9681) );
  INV_X1 U12411 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9876) );
  AND2_X1 U12412 ( .A1(n14722), .A2(n9894), .ZN(n9682) );
  AND2_X1 U12413 ( .A1(n9787), .A2(n14829), .ZN(n9683) );
  AND2_X1 U12414 ( .A1(n9745), .A2(n15366), .ZN(n9684) );
  NOR2_X1 U12415 ( .A1(n13770), .A2(n10008), .ZN(n14192) );
  AND2_X1 U12416 ( .A1(n13735), .A2(n10575), .ZN(n9685) );
  NAND2_X1 U12417 ( .A1(n12289), .A2(n12290), .ZN(n12295) );
  OR2_X1 U12418 ( .A1(n13550), .A2(n13549), .ZN(n13548) );
  AND2_X1 U12419 ( .A1(n11832), .A2(n9650), .ZN(n9686) );
  AND2_X1 U12420 ( .A1(n14160), .A2(n10003), .ZN(n9687) );
  NOR2_X1 U12421 ( .A1(n13612), .A2(n12239), .ZN(n13697) );
  NAND2_X1 U12422 ( .A1(n13074), .A2(n13073), .ZN(n13137) );
  NAND2_X1 U12423 ( .A1(n12542), .A2(n17920), .ZN(n17631) );
  NOR2_X1 U12424 ( .A1(n14928), .A2(n14927), .ZN(n14926) );
  NOR2_X1 U12425 ( .A1(n15428), .A2(n15429), .ZN(n13611) );
  XNOR2_X1 U12426 ( .A(n14898), .B(n13934), .ZN(n14891) );
  INV_X1 U12427 ( .A(n15060), .ZN(n9768) );
  NAND2_X1 U12428 ( .A1(n14900), .A2(n14899), .ZN(n14898) );
  NOR2_X1 U12429 ( .A1(n13672), .A2(n18958), .ZN(n9688) );
  NAND2_X1 U12430 ( .A1(n15316), .A2(n15317), .ZN(n14986) );
  OR2_X1 U12431 ( .A1(n12077), .A2(n11775), .ZN(n9689) );
  AND2_X1 U12432 ( .A1(n9646), .A2(n14788), .ZN(n9690) );
  AND2_X1 U12433 ( .A1(n9683), .A2(n9786), .ZN(n9691) );
  OR2_X1 U12434 ( .A1(n15761), .A2(n15760), .ZN(n9692) );
  INV_X1 U12435 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17551) );
  NAND2_X1 U12436 ( .A1(n11268), .A2(n9870), .ZN(n9693) );
  INV_X1 U12437 ( .A(n13473), .ZN(n11246) );
  INV_X1 U12438 ( .A(n11063), .ZN(n9982) );
  OR2_X1 U12439 ( .A1(n9749), .A2(n14808), .ZN(n9694) );
  AND3_X1 U12440 ( .A1(n10530), .A2(n10529), .A3(n10528), .ZN(n13659) );
  NAND2_X1 U12441 ( .A1(n15236), .A2(n10037), .ZN(n9695) );
  NAND2_X1 U12442 ( .A1(n15315), .A2(n14910), .ZN(n14901) );
  AND2_X1 U12443 ( .A1(n14203), .A2(n13765), .ZN(n9696) );
  AND2_X1 U12444 ( .A1(n9817), .A2(n9816), .ZN(n9697) );
  AND2_X1 U12445 ( .A1(n11320), .A2(n11242), .ZN(n9698) );
  AND2_X1 U12446 ( .A1(n16177), .A2(n16178), .ZN(n9699) );
  AND2_X1 U12447 ( .A1(n11320), .A2(n13644), .ZN(n9700) );
  AND2_X1 U12448 ( .A1(n10016), .A2(n10762), .ZN(n9701) );
  AND2_X1 U12449 ( .A1(n9945), .A2(n9944), .ZN(n9702) );
  AND2_X1 U12450 ( .A1(n9684), .A2(n9744), .ZN(n9703) );
  AND2_X1 U12451 ( .A1(n9905), .A2(n9662), .ZN(n9704) );
  INV_X1 U12452 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13053) );
  INV_X1 U12453 ( .A(n11020), .ZN(n11055) );
  INV_X1 U12454 ( .A(n14711), .ZN(n18896) );
  NAND2_X1 U12455 ( .A1(n13141), .A2(n9936), .ZN(n9935) );
  AND2_X1 U12456 ( .A1(n9935), .A2(n9629), .ZN(n13398) );
  OAI21_X1 U12457 ( .B1(n13000), .B2(n12116), .A(n9741), .ZN(n13036) );
  INV_X1 U12458 ( .A(n13041), .ZN(n9736) );
  NOR2_X1 U12459 ( .A1(n13167), .A2(n13160), .ZN(n13161) );
  OR2_X1 U12460 ( .A1(n13041), .A2(n9737), .ZN(n13242) );
  AND2_X1 U12461 ( .A1(n17447), .A2(n9643), .ZN(n9705) );
  NOR2_X1 U12462 ( .A1(n13572), .A2(n13146), .ZN(n13145) );
  AND2_X1 U12463 ( .A1(n14737), .A2(n9890), .ZN(n9706) );
  INV_X1 U12464 ( .A(n12282), .ZN(n9991) );
  OAI21_X1 U12465 ( .B1(n13478), .B2(n10653), .A(n10468), .ZN(n13459) );
  NAND2_X1 U12466 ( .A1(n13512), .A2(n9945), .ZN(n13673) );
  AND2_X1 U12467 ( .A1(n9909), .A2(n16723), .ZN(n9707) );
  NAND2_X1 U12468 ( .A1(n9736), .A2(n9733), .ZN(n9739) );
  AND2_X1 U12469 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9708) );
  INV_X1 U12470 ( .A(n13990), .ZN(n9943) );
  INV_X1 U12471 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17396) );
  INV_X1 U12472 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14768) );
  AND2_X1 U12473 ( .A1(n13161), .A2(n16183), .ZN(n9709) );
  NAND2_X1 U12474 ( .A1(n12253), .A2(n12252), .ZN(n9710) );
  AND2_X1 U12475 ( .A1(n13161), .A2(n9787), .ZN(n9711) );
  AND2_X1 U12476 ( .A1(n14171), .A2(n14184), .ZN(n9712) );
  AND2_X1 U12477 ( .A1(n9789), .A2(n9788), .ZN(n9713) );
  NAND2_X1 U12478 ( .A1(n14732), .A2(n9640), .ZN(n9888) );
  INV_X1 U12479 ( .A(n9785), .ZN(n14813) );
  NAND2_X1 U12480 ( .A1(n13161), .A2(n9691), .ZN(n9785) );
  INV_X1 U12481 ( .A(n17419), .ZN(n9911) );
  OR2_X1 U12482 ( .A1(n12077), .A2(n11838), .ZN(n9714) );
  AND2_X1 U12483 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12981) );
  AND2_X1 U12484 ( .A1(n9748), .A2(n12339), .ZN(n9715) );
  INV_X1 U12485 ( .A(n9864), .ZN(n20064) );
  OR2_X1 U12486 ( .A1(n17366), .A2(n9922), .ZN(n9716) );
  AND2_X1 U12487 ( .A1(n9865), .A2(n13457), .ZN(n9717) );
  AND2_X1 U12488 ( .A1(n11153), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9718) );
  INV_X1 U12489 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9892) );
  INV_X1 U12490 ( .A(n12312), .ZN(n9836) );
  INV_X1 U12491 ( .A(n10273), .ZN(n10833) );
  INV_X1 U12492 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n9924) );
  INV_X1 U12493 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9898) );
  INV_X1 U12494 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n9809) );
  NAND2_X1 U12495 ( .A1(n15053), .A2(n15042), .ZN(n9719) );
  INV_X1 U12496 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9891) );
  INV_X1 U12497 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n9816) );
  INV_X1 U12498 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18667) );
  INV_X1 U12499 ( .A(n20031), .ZN(n20090) );
  AOI22_X2 U12500 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n9575), .B1(DATAI_25_), 
        .B2(n9574), .ZN(n20581) );
  AOI22_X2 U12501 ( .A1(DATAI_19_), .A2(n9574), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n9575), .ZN(n20646) );
  AOI22_X2 U12502 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n9575), .B1(DATAI_20_), 
        .B2(n9574), .ZN(n20652) );
  AOI22_X2 U12503 ( .A1(DATAI_22_), .A2(n9574), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n9575), .ZN(n20664) );
  AOI22_X2 U12504 ( .A1(DATAI_31_), .A2(n9574), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n9575), .ZN(n20609) );
  AOI22_X2 U12505 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19155), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19156), .ZN(n19730) );
  NOR2_X2 U12506 ( .A1(n19101), .A2(n19102), .ZN(n19156) );
  AOI22_X2 U12507 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n9575), .B1(DATAI_21_), 
        .B2(n9574), .ZN(n20658) );
  NOR3_X2 U12508 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18564), .A3(
        n18227), .ZN(n18245) );
  AND2_X2 U12509 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13118) );
  NAND2_X1 U12510 ( .A1(n15192), .A2(n15193), .ZN(n9723) );
  NAND2_X1 U12511 ( .A1(n12294), .A2(n12300), .ZN(n11733) );
  XNOR2_X2 U12512 ( .A(n12297), .B(n12298), .ZN(n12294) );
  NAND2_X2 U12513 ( .A1(n12281), .A2(n11693), .ZN(n12297) );
  AND2_X2 U12514 ( .A1(n11519), .A2(n13355), .ZN(n19111) );
  NOR2_X2 U12515 ( .A1(n11432), .A2(n9726), .ZN(n11429) );
  XNOR2_X2 U12516 ( .A(n11941), .B(n11940), .ZN(n13077) );
  AND2_X2 U12517 ( .A1(n9822), .A2(n9729), .ZN(n11941) );
  NAND3_X1 U12518 ( .A1(n11489), .A2(n11464), .A3(n11475), .ZN(n9729) );
  NAND2_X2 U12519 ( .A1(n11488), .A2(n11490), .ZN(n11489) );
  AND2_X4 U12520 ( .A1(n13118), .A2(n9751), .ZN(n14052) );
  NOR2_X1 U12521 ( .A1(n13041), .A2(n12099), .ZN(n13241) );
  INV_X1 U12522 ( .A(n12099), .ZN(n9738) );
  INV_X1 U12523 ( .A(n9739), .ZN(n13413) );
  AND2_X2 U12524 ( .A1(n9753), .A2(n9752), .ZN(n11595) );
  NAND4_X1 U12525 ( .A1(n9755), .A2(n9756), .A3(n11539), .A4(n9754), .ZN(n9753) );
  INV_X1 U12526 ( .A(n11520), .ZN(n9757) );
  NAND3_X1 U12527 ( .A1(n9761), .A2(n11464), .A3(n11489), .ZN(n9760) );
  NAND3_X1 U12528 ( .A1(n11475), .A2(n11474), .A3(n9759), .ZN(n9758) );
  OAI21_X2 U12529 ( .B1(n11736), .B2(n9627), .A(n9762), .ZN(n15451) );
  AND2_X1 U12530 ( .A1(n9766), .A2(n15038), .ZN(n9764) );
  OAI21_X1 U12531 ( .B1(n15059), .B2(n9767), .A(n15037), .ZN(n9766) );
  NOR2_X2 U12532 ( .A1(n11511), .A2(n11510), .ZN(n19458) );
  NAND3_X1 U12533 ( .A1(n9819), .A2(n12283), .A3(n12300), .ZN(n9769) );
  OAI21_X1 U12534 ( .B1(n13483), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n13481), .ZN(n11645) );
  INV_X1 U12535 ( .A(n11477), .ZN(n12333) );
  NAND3_X1 U12536 ( .A1(n11465), .A2(n11466), .A3(n9770), .ZN(n11470) );
  NAND2_X1 U12537 ( .A1(n11477), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n9770) );
  NOR2_X1 U12538 ( .A1(n17144), .A2(n17185), .ZN(n17140) );
  NAND3_X1 U12539 ( .A1(n9625), .A2(P3_EAX_REG_21__SCAN_IN), .A3(
        P3_EAX_REG_22__SCAN_IN), .ZN(n9775) );
  NAND3_X1 U12540 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .ZN(n9777) );
  INV_X2 U12541 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18672) );
  INV_X2 U12542 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18682) );
  OAI22_X1 U12543 ( .A1(n11467), .A2(n9779), .B1(n11999), .B2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11463) );
  AND2_X2 U12544 ( .A1(n9779), .A2(n12829), .ZN(n11999) );
  NAND4_X1 U12545 ( .A1(n11407), .A2(n11404), .A3(n11405), .A4(n11406), .ZN(
        n9782) );
  NAND4_X1 U12546 ( .A1(n11413), .A2(n11410), .A3(n11412), .A4(n11411), .ZN(
        n9784) );
  NAND2_X1 U12547 ( .A1(n9795), .A2(n9793), .ZN(n14928) );
  INV_X1 U12548 ( .A(n15011), .ZN(n15013) );
  NOR2_X1 U12549 ( .A1(n15038), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11855) );
  NAND2_X1 U12550 ( .A1(n11859), .A2(n9813), .ZN(n14744) );
  NAND2_X1 U12551 ( .A1(n9680), .A2(n11853), .ZN(n9813) );
  NAND2_X1 U12552 ( .A1(n12329), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15010) );
  NAND2_X1 U12553 ( .A1(n11596), .A2(n11595), .ZN(n12283) );
  NAND2_X1 U12554 ( .A1(n9821), .A2(n9820), .ZN(n9819) );
  INV_X1 U12555 ( .A(n11596), .ZN(n9821) );
  NAND2_X1 U12556 ( .A1(n13565), .A2(n9827), .ZN(n9824) );
  NAND2_X1 U12557 ( .A1(n9824), .A2(n9826), .ZN(n12287) );
  NAND2_X1 U12558 ( .A1(n12292), .A2(n9675), .ZN(n9828) );
  AOI21_X1 U12559 ( .B1(n9677), .B2(n12289), .A(n9830), .ZN(n9829) );
  INV_X1 U12560 ( .A(n10029), .ZN(n9832) );
  NAND3_X2 U12561 ( .A1(n9659), .A2(n10103), .A3(n10102), .ZN(n10210) );
  INV_X2 U12562 ( .A(n20117), .ZN(n10211) );
  NAND2_X2 U12563 ( .A1(n10072), .A2(n10027), .ZN(n20117) );
  AND2_X2 U12564 ( .A1(n13446), .A2(n10061), .ZN(n10198) );
  AND2_X2 U12565 ( .A1(n9876), .A2(n9875), .ZN(n13446) );
  NAND2_X1 U12566 ( .A1(n10346), .A2(n10345), .ZN(n12910) );
  NAND2_X2 U12567 ( .A1(n10335), .A2(n10334), .ZN(n10346) );
  INV_X1 U12568 ( .A(n10345), .ZN(n9845) );
  OR2_X2 U12569 ( .A1(n10257), .A2(n10240), .ZN(n9969) );
  INV_X1 U12570 ( .A(n9972), .ZN(n9971) );
  NAND2_X1 U12571 ( .A1(n9970), .A2(n9851), .ZN(n13718) );
  INV_X1 U12572 ( .A(n9852), .ZN(n9851) );
  OAI21_X1 U12573 ( .B1(n9972), .B2(n11104), .A(n9679), .ZN(n9852) );
  NAND3_X1 U12574 ( .A1(n9854), .A2(n9853), .A3(n9678), .ZN(n14454) );
  NAND3_X1 U12575 ( .A1(n9854), .A2(n9853), .A3(n11152), .ZN(n14471) );
  NAND4_X4 U12576 ( .A1(n10187), .A2(n9860), .A3(n9858), .A4(n9859), .ZN(
        n10224) );
  NAND2_X1 U12577 ( .A1(n10576), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n9859) );
  NAND2_X1 U12578 ( .A1(n9865), .A2(n13475), .ZN(n9864) );
  NAND2_X1 U12579 ( .A1(n9700), .A2(n13105), .ZN(n11239) );
  NAND2_X1 U12580 ( .A1(n13105), .A2(n9698), .ZN(n11245) );
  NAND2_X1 U12581 ( .A1(n13105), .A2(n11320), .ZN(n11317) );
  NAND2_X1 U12582 ( .A1(n9866), .A2(n15845), .ZN(n11272) );
  NAND2_X1 U12583 ( .A1(n9866), .A2(n14243), .ZN(n11309) );
  NAND2_X1 U12584 ( .A1(n9866), .A2(n13779), .ZN(n11281) );
  INV_X1 U12585 ( .A(n15970), .ZN(n9869) );
  INV_X1 U12586 ( .A(n9888), .ZN(n14735) );
  NAND3_X1 U12587 ( .A1(n9896), .A2(n9630), .A3(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14720) );
  NAND2_X1 U12588 ( .A1(n12549), .A2(n17476), .ZN(n17425) );
  NAND2_X2 U12589 ( .A1(n17515), .A2(n17639), .ZN(n17476) );
  OR2_X2 U12591 ( .A1(n12468), .A2(n12467), .ZN(n17246) );
  OR2_X1 U12592 ( .A1(n12555), .A2(n17752), .ZN(n9907) );
  OR3_X1 U12593 ( .A1(n12555), .A2(n17752), .A3(n9652), .ZN(n12560) );
  NAND2_X1 U12594 ( .A1(n9908), .A2(n9910), .ZN(n16481) );
  NAND2_X1 U12595 ( .A1(n16501), .A2(n9647), .ZN(n9908) );
  INV_X1 U12596 ( .A(n9917), .ZN(n17408) );
  NOR2_X1 U12597 ( .A1(n17366), .A2(n12692), .ZN(n16257) );
  INV_X1 U12598 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9923) );
  NAND4_X1 U12599 ( .A1(n17633), .A2(n9634), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A4(n10031), .ZN(n17552) );
  NAND2_X2 U12600 ( .A1(n9929), .A2(n9927), .ZN(n11521) );
  NAND2_X1 U12601 ( .A1(n9928), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9927) );
  NAND4_X1 U12602 ( .A1(n11394), .A2(n11396), .A3(n11395), .A4(n11397), .ZN(
        n9928) );
  NAND2_X1 U12603 ( .A1(n9930), .A2(n11530), .ZN(n9929) );
  NAND4_X1 U12604 ( .A1(n11401), .A2(n11400), .A3(n11398), .A4(n11399), .ZN(
        n9930) );
  NAND2_X1 U12605 ( .A1(n9934), .A2(n9931), .ZN(n14866) );
  NAND2_X1 U12606 ( .A1(n9933), .A2(n9932), .ZN(n14933) );
  NAND2_X1 U12607 ( .A1(n9935), .A2(n9633), .ZN(n18976) );
  NAND2_X1 U12608 ( .A1(n9943), .A2(n9941), .ZN(n9940) );
  NAND2_X1 U12609 ( .A1(n9943), .A2(n13961), .ZN(n9942) );
  NOR2_X2 U12610 ( .A1(n14921), .A2(n9946), .ZN(n16102) );
  NOR2_X1 U12611 ( .A1(n14921), .A2(n9950), .ZN(n14914) );
  NAND3_X1 U12612 ( .A1(n14402), .A2(n9952), .A3(n14411), .ZN(n9953) );
  NAND2_X1 U12613 ( .A1(n14402), .A2(n14411), .ZN(n14401) );
  NAND2_X1 U12614 ( .A1(n14401), .A2(n14571), .ZN(n14381) );
  NAND2_X1 U12615 ( .A1(n14401), .A2(n9954), .ZN(n9956) );
  INV_X1 U12616 ( .A(n9956), .ZN(n14372) );
  OAI211_X2 U12617 ( .C1(n13469), .C2(n9961), .A(n9959), .B(n13524), .ZN(
        n13527) );
  NAND3_X1 U12618 ( .A1(n9960), .A2(n9964), .A3(n9962), .ZN(n9959) );
  NAND2_X1 U12619 ( .A1(n13467), .A2(n13468), .ZN(n13469) );
  NAND2_X1 U12620 ( .A1(n13467), .A2(n9963), .ZN(n9962) );
  NAND2_X1 U12621 ( .A1(n9965), .A2(n20054), .ZN(n9964) );
  NAND2_X1 U12622 ( .A1(n20028), .A2(n9971), .ZN(n9970) );
  OAI21_X1 U12623 ( .B1(n20028), .B2(n9973), .A(n9971), .ZN(n15910) );
  NAND2_X1 U12624 ( .A1(n11144), .A2(n9978), .ZN(n9974) );
  NAND2_X1 U12625 ( .A1(n11148), .A2(n9976), .ZN(n9975) );
  NAND3_X1 U12626 ( .A1(n9975), .A2(n9974), .A3(n9977), .ZN(n14447) );
  NAND2_X1 U12627 ( .A1(n14471), .A2(n14470), .ZN(n14453) );
  XNOR2_X2 U12628 ( .A(n10454), .B(n10453), .ZN(n11070) );
  NAND2_X2 U12629 ( .A1(n9986), .A2(n9984), .ZN(n12035) );
  NAND4_X1 U12630 ( .A1(n11363), .A2(n11360), .A3(n11361), .A4(n11362), .ZN(
        n9985) );
  NAND4_X1 U12631 ( .A1(n11367), .A2(n11366), .A3(n11364), .A4(n11365), .ZN(
        n9987) );
  INV_X1 U12632 ( .A(n9989), .ZN(n9988) );
  XNOR2_X2 U12633 ( .A(n9990), .B(n9989), .ZN(n11488) );
  AND2_X2 U12634 ( .A1(n11451), .A2(n11450), .ZN(n9990) );
  NAND2_X1 U12635 ( .A1(n9997), .A2(n9996), .ZN(n13656) );
  NAND3_X1 U12636 ( .A1(n10330), .A2(n9998), .A3(n10444), .ZN(n10447) );
  NAND2_X1 U12637 ( .A1(n10301), .A2(n10300), .ZN(n9998) );
  INV_X1 U12638 ( .A(n10301), .ZN(n11077) );
  NAND2_X1 U12639 ( .A1(n10430), .A2(n9999), .ZN(n10433) );
  NAND3_X1 U12640 ( .A1(n10430), .A2(n9999), .A3(n10422), .ZN(n10502) );
  NAND2_X1 U12641 ( .A1(n10000), .A2(n9701), .ZN(n14248) );
  AND2_X1 U12642 ( .A1(n13735), .A2(n10593), .ZN(n10007) );
  NOR2_X1 U12643 ( .A1(n14120), .A2(n14121), .ZN(n14107) );
  NAND2_X1 U12644 ( .A1(n12352), .A2(n12351), .ZN(n12356) );
  XNOR2_X1 U12645 ( .A(n14061), .B(n14060), .ZN(n14068) );
  NAND2_X1 U12646 ( .A1(n14866), .A2(n14043), .ZN(n14061) );
  AOI21_X1 U12647 ( .B1(n12413), .B2(n14108), .A(n12352), .ZN(n14386) );
  NOR2_X1 U12648 ( .A1(n12035), .A2(n11440), .ZN(n11380) );
  NAND2_X1 U12649 ( .A1(n12049), .A2(n19131), .ZN(n11444) );
  AND2_X1 U12650 ( .A1(n14052), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12121) );
  AND2_X1 U12651 ( .A1(n14052), .A2(n13115), .ZN(n11597) );
  NAND2_X1 U12652 ( .A1(n12798), .A2(n11423), .ZN(n11435) );
  AOI22_X1 U12653 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9605), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11375) );
  OR2_X1 U12654 ( .A1(n12827), .A2(n12826), .ZN(n12828) );
  NAND2_X1 U12655 ( .A1(n12827), .A2(n12826), .ZN(n12904) );
  AOI22_X1 U12656 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U12657 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U12658 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11376) );
  INV_X1 U12659 ( .A(n11470), .ZN(n11473) );
  NAND2_X1 U12660 ( .A1(n12918), .A2(n11222), .ZN(n15724) );
  AND2_X1 U12661 ( .A1(n11220), .A2(n11219), .ZN(n12941) );
  NAND2_X1 U12662 ( .A1(n11219), .A2(n13016), .ZN(n10245) );
  INV_X1 U12663 ( .A(n10218), .ZN(n11222) );
  NAND2_X1 U12664 ( .A1(n10447), .A2(n10446), .ZN(n13479) );
  XNOR2_X1 U12665 ( .A(n10305), .B(n10304), .ZN(n10456) );
  NAND2_X1 U12666 ( .A1(n10305), .A2(n10303), .ZN(n10258) );
  OAI22_X1 U12667 ( .A1(n10262), .A2(n10089), .B1(n10087), .B2(n10088), .ZN(
        n10090) );
  AOI21_X2 U12668 ( .B1(n14373), .B2(n15892), .A(n10035), .ZN(n14375) );
  AOI21_X1 U12669 ( .B1(n14379), .B2(n20031), .A(n14378), .ZN(n14380) );
  NAND2_X1 U12670 ( .A1(n14379), .A2(n10041), .ZN(n12387) );
  XNOR2_X1 U12671 ( .A(n12326), .B(n10033), .ZN(n15036) );
  AND2_X1 U12672 ( .A1(n10782), .A2(n10781), .ZN(n10016) );
  INV_X1 U12673 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13115) );
  AND4_X1 U12674 ( .A1(n11615), .A2(n11614), .A3(n11613), .A4(n11612), .ZN(
        n10018) );
  AND2_X1 U12675 ( .A1(n11435), .A2(n13675), .ZN(n10019) );
  AND2_X1 U12676 ( .A1(n10601), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10020) );
  AND3_X1 U12677 ( .A1(n12730), .A2(n12729), .A3(n10039), .ZN(n10021) );
  NAND2_X1 U12678 ( .A1(n17489), .A2(n17735), .ZN(n17482) );
  OR2_X1 U12679 ( .A1(n9581), .A2(n15980), .ZN(n10023) );
  NOR2_X1 U12680 ( .A1(n13377), .A2(n19883), .ZN(n10024) );
  AND2_X1 U12681 ( .A1(n15857), .A2(n14660), .ZN(n10025) );
  INV_X2 U12682 ( .A(n19897), .ZN(n19813) );
  OR2_X1 U12683 ( .A1(n17639), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10026) );
  NAND2_X1 U12684 ( .A1(n10505), .A2(n10504), .ZN(n11062) );
  NAND2_X1 U12685 ( .A1(n10188), .A2(n10224), .ZN(n12753) );
  NOR2_X1 U12686 ( .A1(n14914), .A2(n16107), .ZN(n10028) );
  AND2_X1 U12687 ( .A1(n13591), .A2(n12291), .ZN(n10029) );
  INV_X1 U12688 ( .A(n10457), .ZN(n10509) );
  NOR2_X1 U12689 ( .A1(n10229), .A2(n20613), .ZN(n10457) );
  AND2_X1 U12690 ( .A1(n11324), .A2(n11323), .ZN(n10030) );
  INV_X1 U12691 ( .A(n14645), .ZN(n11153) );
  INV_X1 U12692 ( .A(n13763), .ZN(n10575) );
  INV_X1 U12693 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14374) );
  INV_X1 U12694 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12525) );
  AND2_X1 U12695 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10031) );
  AND2_X1 U12696 ( .A1(n15865), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10032) );
  AND2_X1 U12697 ( .A1(n15000), .A2(n12325), .ZN(n10033) );
  INV_X1 U12698 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12693) );
  INV_X2 U12699 ( .A(n18725), .ZN(n18658) );
  INV_X1 U12700 ( .A(n11814), .ZN(n12300) );
  INV_X1 U12701 ( .A(n12079), .ZN(n12118) );
  OR2_X1 U12702 ( .A1(n15231), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10034) );
  OR2_X1 U12703 ( .A1(n18713), .A2(n17274), .ZN(n17276) );
  NOR2_X1 U12704 ( .A1(n11581), .A2(n11580), .ZN(n12271) );
  AND2_X1 U12705 ( .A1(n14372), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10035) );
  INV_X1 U12706 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n19757) );
  OR2_X1 U12707 ( .A1(n16588), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10036) );
  NOR2_X1 U12708 ( .A1(n12430), .A2(n16773), .ZN(n12427) );
  CLKBUF_X3 U12709 ( .A(n12497), .Z(n17052) );
  INV_X1 U12710 ( .A(n11522), .ZN(n13849) );
  AND2_X1 U12711 ( .A1(n9601), .A2(n13115), .ZN(n12170) );
  NOR2_X1 U12712 ( .A1(n15235), .A2(n15234), .ZN(n10037) );
  OR2_X1 U12713 ( .A1(n11728), .A2(n11727), .ZN(n11731) );
  INV_X2 U12714 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20613) );
  AND3_X1 U12715 ( .A1(n11456), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n12037), 
        .ZN(n10038) );
  INV_X1 U12716 ( .A(n17221), .ZN(n17213) );
  OR2_X1 U12717 ( .A1(n16278), .A2(n17739), .ZN(n10039) );
  OR3_X1 U12718 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17452), .ZN(n10040) );
  INV_X1 U12719 ( .A(n17608), .ZN(n17639) );
  AND2_X1 U12720 ( .A1(n14365), .A2(n14069), .ZN(n10041) );
  NAND2_X2 U12721 ( .A1(n14365), .A2(n12962), .ZN(n14370) );
  NAND2_X1 U12722 ( .A1(n20003), .A2(n14069), .ZN(n14298) );
  INV_X1 U12723 ( .A(n14298), .ZN(n12418) );
  INV_X1 U12724 ( .A(n12073), .ZN(n12117) );
  INV_X1 U12725 ( .A(n12117), .ZN(n15224) );
  INV_X1 U12726 ( .A(n10087), .ZN(n10516) );
  AND3_X1 U12727 ( .A1(n10056), .A2(n10055), .A3(n10054), .ZN(n10042) );
  INV_X1 U12728 ( .A(n10126), .ZN(n10316) );
  AND2_X1 U12729 ( .A1(n10106), .A2(n10105), .ZN(n10043) );
  NAND2_X1 U12730 ( .A1(n10858), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10044) );
  AND3_X1 U12731 ( .A1(n10122), .A2(n10121), .A3(n10120), .ZN(n10045) );
  INV_X1 U12732 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n10259) );
  NAND2_X1 U12733 ( .A1(n11432), .A2(n11927), .ZN(n11433) );
  INV_X1 U12734 ( .A(n13630), .ZN(n10243) );
  INV_X1 U12735 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10388) );
  INV_X1 U12736 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10479) );
  OAI22_X1 U12737 ( .A1(n13895), .A2(n19521), .B1(n19635), .B2(n12142), .ZN(
        n11542) );
  INV_X1 U12738 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10170) );
  INV_X1 U12739 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10059) );
  OR2_X1 U12740 ( .A1(n10419), .A2(n10418), .ZN(n11116) );
  AOI22_X1 U12741 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10516), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10120) );
  OR2_X1 U12742 ( .A1(n11893), .A2(n11872), .ZN(n11622) );
  NOR2_X1 U12743 ( .A1(n11381), .A2(n11380), .ZN(n11403) );
  AOI22_X1 U12744 ( .A1(n11349), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11412) );
  INV_X1 U12745 ( .A(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10684) );
  INV_X1 U12746 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11030) );
  INV_X1 U12747 ( .A(n11009), .ZN(n10392) );
  AND4_X1 U12748 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10282), .ZN(
        n10289) );
  AND2_X1 U12749 ( .A1(n19890), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12823) );
  AND2_X1 U12750 ( .A1(n11627), .A2(n11623), .ZN(n11625) );
  NAND2_X1 U12751 ( .A1(n12100), .A2(n19119), .ZN(n11539) );
  OR2_X1 U12752 ( .A1(n10260), .A2(n10155), .ZN(n10157) );
  OR4_X1 U12753 ( .A1(n10890), .A2(n10889), .A3(n10888), .A4(n10887), .ZN(
        n10916) );
  AND2_X1 U12754 ( .A1(n10421), .A2(n10420), .ZN(n10423) );
  INV_X1 U12755 ( .A(n10825), .ZN(n10826) );
  BUF_X1 U12756 ( .A(n10392), .Z(n10902) );
  INV_X2 U12757 ( .A(n10952), .ZN(n11028) );
  INV_X1 U12758 ( .A(n10503), .ZN(n10504) );
  OR2_X1 U12759 ( .A1(n10322), .A2(n10321), .ZN(n11075) );
  NAND2_X1 U12760 ( .A1(n10224), .A2(n20127), .ZN(n10370) );
  INV_X1 U12761 ( .A(n16111), .ZN(n13802) );
  OR2_X1 U12762 ( .A1(n11656), .A2(n11655), .ZN(n12282) );
  AND2_X1 U12763 ( .A1(n15759), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11868) );
  NAND2_X1 U12764 ( .A1(n15027), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14709) );
  OR2_X1 U12765 ( .A1(n12571), .A2(n12572), .ZN(n12567) );
  NAND2_X1 U12766 ( .A1(n10945), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10947) );
  NAND2_X1 U12767 ( .A1(n10826), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10828) );
  OR2_X1 U12768 ( .A1(n10296), .A2(n10295), .ZN(n11128) );
  INV_X1 U12769 ( .A(n13540), .ZN(n11255) );
  OAI211_X1 U12770 ( .C1(n11169), .C2(n10834), .A(n10327), .B(n10326), .ZN(
        n10453) );
  OR2_X1 U12771 ( .A1(n13959), .A2(n13962), .ZN(n13986) );
  OR2_X1 U12772 ( .A1(n11869), .A2(n11868), .ZN(n11871) );
  OR2_X1 U12773 ( .A1(n15695), .A2(n12300), .ZN(n11836) );
  AND2_X1 U12774 ( .A1(n12243), .A2(n12242), .ZN(n15353) );
  OR2_X1 U12775 ( .A1(n14818), .A2(n12300), .ZN(n11773) );
  INV_X1 U12776 ( .A(n12297), .ZN(n12299) );
  INV_X1 U12777 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n20820) );
  NOR2_X1 U12778 ( .A1(n12428), .A2(n12431), .ZN(n12469) );
  NAND2_X1 U12779 ( .A1(n17608), .A2(n17865), .ZN(n12544) );
  INV_X1 U12780 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12529) );
  INV_X1 U12781 ( .A(n18076), .ZN(n12672) );
  INV_X1 U12782 ( .A(n10630), .ZN(n10594) );
  INV_X1 U12783 ( .A(n15969), .ZN(n11268) );
  OR2_X1 U12784 ( .A1(n10947), .A2(n10946), .ZN(n10993) );
  OR2_X1 U12785 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13722), .ZN(
        n20076) );
  NAND2_X1 U12786 ( .A1(n11215), .A2(n11214), .ZN(n11216) );
  AND2_X1 U12787 ( .A1(n11794), .A2(n11803), .ZN(n18809) );
  OR2_X1 U12788 ( .A1(n12218), .A2(n12217), .ZN(n13577) );
  AND2_X1 U12789 ( .A1(n13675), .A2(n19883), .ZN(n12090) );
  OR2_X1 U12790 ( .A1(n11836), .A2(n15321), .ZN(n15310) );
  AND2_X1 U12791 ( .A1(n11786), .A2(n15368), .ZN(n15107) );
  INV_X1 U12792 ( .A(n16196), .ZN(n15525) );
  INV_X1 U12793 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12758) );
  AOI21_X1 U12794 ( .B1(n11912), .B2(n11911), .A(n12393), .ZN(n13377) );
  INV_X1 U12795 ( .A(n19487), .ZN(n19492) );
  AND2_X1 U12796 ( .A1(n19559), .A2(n19837), .ZN(n19554) );
  OAI22_X1 U12797 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18545), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12568), .ZN(n12574) );
  NOR2_X1 U12799 ( .A1(n12685), .A2(n12672), .ZN(n18509) );
  NOR3_X1 U12800 ( .A1(n12672), .A2(n12664), .A3(n12666), .ZN(n12673) );
  INV_X1 U12801 ( .A(n11320), .ZN(n10247) );
  INV_X1 U12802 ( .A(n12970), .ZN(n13624) );
  INV_X1 U12803 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14152) );
  AND2_X1 U12804 ( .A1(n10802), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10803) );
  INV_X1 U12805 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14211) );
  AND2_X1 U12806 ( .A1(n14377), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13635) );
  AND2_X1 U12807 ( .A1(n12923), .A2(n12369), .ZN(n12370) );
  AND2_X1 U12808 ( .A1(n14081), .A2(n11020), .ZN(n11058) );
  INV_X1 U12809 ( .A(n10922), .ZN(n10945) );
  INV_X1 U12810 ( .A(n11055), .ZN(n10780) );
  NOR2_X1 U12811 ( .A1(n10565), .A2(n19927), .ZN(n10569) );
  INV_X1 U12812 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13529) );
  NAND2_X1 U12813 ( .A1(n19908), .A2(n11223), .ZN(n14484) );
  NAND2_X1 U12815 ( .A1(n13034), .A2(n13020), .ZN(n20079) );
  NAND2_X1 U12816 ( .A1(n11217), .A2(n11216), .ZN(n13008) );
  OR2_X1 U12817 ( .A1(n11089), .A2(n20094), .ZN(n20153) );
  INV_X1 U12818 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20473) );
  NOR2_X1 U12819 ( .A1(n20258), .A2(n20257), .ZN(n20572) );
  AOI21_X1 U12820 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20536), .A(n20257), 
        .ZN(n20620) );
  NAND2_X1 U12821 ( .A1(n18737), .A2(n19757), .ZN(n13390) );
  INV_X1 U12822 ( .A(n18906), .ZN(n18941) );
  INV_X1 U12823 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15075) );
  INV_X1 U12824 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15169) );
  INV_X1 U12825 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18818) );
  INV_X1 U12826 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n15217) );
  OR2_X1 U12827 ( .A1(n15131), .A2(n15330), .ZN(n15305) );
  AND2_X1 U12828 ( .A1(n15381), .A2(n15379), .ZN(n16216) );
  OR2_X1 U12829 ( .A1(n18736), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13051) );
  INV_X1 U12830 ( .A(n19526), .ZN(n19691) );
  INV_X1 U12831 ( .A(n19697), .ZN(n19627) );
  INV_X1 U12832 ( .A(n19155), .ZN(n19148) );
  OR2_X1 U12833 ( .A1(n19450), .A2(n19861), .ZN(n19518) );
  OAI22_X1 U12834 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18504), .B1(
        n12575), .B2(n12574), .ZN(n12681) );
  NOR2_X1 U12835 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16612), .ZN(n16599) );
  NOR2_X1 U12836 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16641), .ZN(n16623) );
  NAND2_X1 U12837 ( .A1(n16275), .A2(n17598), .ZN(n12729) );
  INV_X1 U12838 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17437) );
  OR3_X1 U12839 ( .A1(n17469), .A2(n17472), .A3(n17811), .ZN(n16279) );
  NOR2_X1 U12840 ( .A1(n17920), .A2(n16244), .ZN(n17871) );
  NOR2_X1 U12841 ( .A1(n17555), .A2(n17885), .ZN(n17521) );
  INV_X1 U12842 ( .A(n17921), .ZN(n17904) );
  INV_X1 U12843 ( .A(n12538), .ZN(n12536) );
  INV_X1 U12844 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12510) );
  OR2_X1 U12845 ( .A1(n18691), .A2(n18570), .ZN(n18060) );
  AOI22_X1 U12846 ( .A1(n9580), .A2(n18494), .B1(n18499), .B2(n16288), .ZN(
        n18503) );
  NAND2_X1 U12847 ( .A1(n10803), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10825) );
  AND2_X1 U12848 ( .A1(n14217), .A2(n13623), .ZN(n19955) );
  INV_X1 U12849 ( .A(n19962), .ZN(n19973) );
  NOR2_X1 U12850 ( .A1(n14326), .A2(n16300), .ZN(n12384) );
  NOR2_X2 U12851 ( .A1(n12383), .A2(n20091), .ZN(n14355) );
  INV_X1 U12852 ( .A(n14365), .ZN(n14366) );
  INV_X1 U12853 ( .A(n19901), .ZN(n13012) );
  OR2_X1 U12854 ( .A1(n12790), .A2(n12789), .ZN(n12930) );
  INV_X1 U12855 ( .A(n13396), .ZN(n20014) );
  AOI21_X1 U12856 ( .B1(n11060), .B2(n11059), .A(n11058), .ZN(n12351) );
  NAND2_X1 U12857 ( .A1(n10570), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10630) );
  AND2_X1 U12858 ( .A1(n10495), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10507) );
  AND2_X1 U12859 ( .A1(n14531), .A2(n15982), .ZN(n14602) );
  OR2_X1 U12860 ( .A1(n14622), .A2(n14610), .ZN(n14614) );
  NOR2_X1 U12861 ( .A1(n15945), .A2(n14540), .ZN(n14661) );
  OR2_X1 U12862 ( .A1(n20075), .A2(n20059), .ZN(n15982) );
  INV_X1 U12863 ( .A(n14681), .ZN(n20061) );
  INV_X1 U12864 ( .A(n13728), .ZN(n13721) );
  NOR2_X1 U12865 ( .A1(n13008), .A2(n20510), .ZN(n15739) );
  NOR2_X1 U12866 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12994) );
  OAI22_X1 U12867 ( .A1(n20110), .A2(n20109), .B1(n20436), .B2(n20253), .ZN(
        n20146) );
  INV_X1 U12868 ( .A(n20210), .ZN(n20173) );
  OAI22_X1 U12869 ( .A1(n20183), .A2(n20182), .B1(n20436), .B2(n20312), .ZN(
        n20206) );
  INV_X1 U12870 ( .A(n20153), .ZN(n20218) );
  INV_X1 U12871 ( .A(n20260), .ZN(n20277) );
  OAI22_X1 U12872 ( .A1(n20314), .A2(n20313), .B1(n20312), .B2(n20565), .ZN(
        n20337) );
  AND2_X1 U12873 ( .A1(n13479), .A2(n11070), .ZN(n20424) );
  INV_X1 U12874 ( .A(n20366), .ZN(n20395) );
  INV_X1 U12875 ( .A(n20467), .ZN(n20428) );
  OAI22_X1 U12876 ( .A1(n20438), .A2(n20437), .B1(n20436), .B2(n20566), .ZN(
        n20469) );
  INV_X1 U12877 ( .A(n20503), .ZN(n20494) );
  OAI22_X1 U12878 ( .A1(n20514), .A2(n20513), .B1(n20512), .B2(n20565), .ZN(
        n20530) );
  AND2_X1 U12879 ( .A1(n20539), .A2(n20504), .ZN(n20560) );
  OAI211_X1 U12880 ( .C1(n20602), .C2(n20573), .A(n20572), .B(n20571), .ZN(
        n20605) );
  NOR2_X1 U12881 ( .A1(n13479), .A2(n11070), .ZN(n20535) );
  INV_X1 U12882 ( .A(n20445), .ZN(n20635) );
  INV_X1 U12883 ( .A(n20457), .ZN(n20653) );
  INV_X1 U12884 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n15734) );
  INV_X1 U12885 ( .A(n20768), .ZN(n20687) );
  INV_X1 U12886 ( .A(n20746), .ZN(n20740) );
  AOI21_X1 U12887 ( .B1(n14771), .B2(n18915), .A(n14769), .ZN(n15699) );
  NAND2_X1 U12888 ( .A1(n14750), .A2(n16015), .ZN(n18935) );
  INV_X1 U12889 ( .A(n18925), .ZN(n18937) );
  AND2_X1 U12890 ( .A1(n19063), .A2(n19630), .ZN(n18944) );
  AND2_X1 U12891 ( .A1(n14979), .A2(n13678), .ZN(n20784) );
  INV_X1 U12892 ( .A(n14979), .ZN(n20780) );
  INV_X2 U12893 ( .A(n19017), .ZN(n19047) );
  NOR2_X1 U12894 ( .A1(n19063), .A2(n19084), .ZN(n19061) );
  INV_X2 U12895 ( .A(n12897), .ZN(n19084) );
  INV_X1 U12896 ( .A(n13051), .ZN(n19090) );
  INV_X1 U12897 ( .A(n16227), .ZN(n16192) );
  NOR2_X2 U12898 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19837) );
  NAND2_X1 U12899 ( .A1(n12904), .A2(n12828), .ZN(n19851) );
  AND3_X1 U12900 ( .A1(n13132), .A2(n13131), .A3(n13130), .ZN(n13367) );
  OAI21_X1 U12901 ( .B1(n19114), .B2(n19113), .A(n19112), .ZN(n19162) );
  INV_X1 U12902 ( .A(n19189), .ZN(n19206) );
  INV_X1 U12903 ( .A(n19210), .ZN(n19239) );
  OAI21_X1 U12904 ( .B1(n19252), .B2(n19251), .A(n19250), .ZN(n19276) );
  AND2_X1 U12905 ( .A1(n19450), .A2(n19413), .ZN(n19383) );
  AND2_X1 U12906 ( .A1(n19383), .A2(n19594), .ZN(n19379) );
  AND2_X1 U12907 ( .A1(n19450), .A2(n19861), .ZN(n19354) );
  OAI21_X1 U12908 ( .B1(n19424), .B2(n19423), .A(n19422), .ZN(n19446) );
  INV_X1 U12909 ( .A(n19481), .ZN(n19483) );
  NOR2_X2 U12910 ( .A1(n19462), .A2(n19518), .ZN(n19513) );
  INV_X1 U12911 ( .A(n19544), .ZN(n19549) );
  OAI21_X1 U12912 ( .B1(n19561), .B2(n19558), .A(n19557), .ZN(n19583) );
  INV_X1 U12913 ( .A(n19617), .ZN(n19621) );
  AND2_X1 U12914 ( .A1(n19281), .A2(n19280), .ZN(n19594) );
  INV_X1 U12915 ( .A(n19645), .ZN(n19701) );
  INV_X1 U12916 ( .A(n19665), .ZN(n19725) );
  INV_X1 U12917 ( .A(n19676), .ZN(n19740) );
  NOR2_X1 U12918 ( .A1(n18737), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19752) );
  AND3_X1 U12919 ( .A1(n19763), .A2(n19818), .A3(n19768), .ZN(n19891) );
  INV_X1 U12920 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19774) );
  NOR2_X1 U12921 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n12695), .ZN(n18730) );
  AOI211_X1 U12922 ( .C1(n12577), .C2(n12576), .A(n12684), .B(n12681), .ZN(
        n18495) );
  NOR2_X1 U12923 ( .A1(n16781), .A2(n16425), .ZN(n16466) );
  NOR2_X1 U12924 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16508), .ZN(n16491) );
  NOR2_X1 U12925 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16551), .ZN(n16533) );
  NOR2_X1 U12926 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16573), .ZN(n16557) );
  NAND4_X1 U12927 ( .A1(n18048), .A2(n18729), .A3(n18569), .A4(n18559), .ZN(
        n16782) );
  NOR2_X1 U12928 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16696), .ZN(n16671) );
  NOR2_X1 U12929 ( .A1(n18497), .A2(n17305), .ZN(n18731) );
  AND2_X1 U12930 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16894), .ZN(n16880) );
  NAND2_X1 U12931 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17020), .ZN(n17005) );
  INV_X1 U12932 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17031) );
  INV_X1 U12933 ( .A(n17099), .ZN(n17102) );
  INV_X1 U12934 ( .A(n17159), .ZN(n17154) );
  NAND2_X1 U12935 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17169), .ZN(n17168) );
  INV_X1 U12936 ( .A(n15689), .ZN(n17217) );
  INV_X1 U12937 ( .A(n18528), .ZN(n15763) );
  INV_X1 U12938 ( .A(n17304), .ZN(n17274) );
  INV_X1 U12939 ( .A(n17746), .ZN(n16250) );
  NOR2_X1 U12940 ( .A1(n16279), .A2(n17454), .ZN(n17428) );
  NOR2_X1 U12941 ( .A1(n18675), .A2(n17730), .ZN(n17582) );
  INV_X1 U12942 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17596) );
  AND2_X1 U12943 ( .A1(n12726), .A2(n17640), .ZN(n17922) );
  NAND2_X1 U12944 ( .A1(n17735), .A2(n17632), .ZN(n17730) );
  INV_X1 U12945 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17573) );
  INV_X1 U12946 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17591) );
  NOR2_X2 U12947 ( .A1(n16410), .A2(n17956), .ZN(n18494) );
  NOR2_X1 U12948 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18667), .ZN(
        n18691) );
  INV_X1 U12949 ( .A(n18159), .ZN(n18150) );
  INV_X1 U12950 ( .A(n18181), .ZN(n18174) );
  INV_X1 U12951 ( .A(n18215), .ZN(n18223) );
  INV_X1 U12952 ( .A(n18266), .ZN(n18268) );
  INV_X1 U12953 ( .A(n18295), .ZN(n18288) );
  INV_X1 U12954 ( .A(n18346), .ZN(n18339) );
  INV_X1 U12955 ( .A(n18362), .ZN(n18369) );
  INV_X1 U12956 ( .A(n18396), .ZN(n18387) );
  NAND2_X1 U12957 ( .A1(n12696), .A2(n18060), .ZN(n18399) );
  INV_X1 U12958 ( .A(n18424), .ZN(n18427) );
  INV_X1 U12959 ( .A(n18564), .ZN(n18433) );
  NOR2_X1 U12960 ( .A1(n18566), .A2(n18563), .ZN(n18711) );
  INV_X1 U12961 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18591) );
  OR2_X1 U12962 ( .A1(n12790), .A2(n12753), .ZN(n13254) );
  INV_X1 U12963 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20254) );
  OR3_X1 U12964 ( .A1(n13637), .A2(n15731), .A3(n13626), .ZN(n19971) );
  NAND2_X1 U12965 ( .A1(n20003), .A2(n10229), .ZN(n14290) );
  OR2_X1 U12966 ( .A1(n14192), .A2(n14194), .ZN(n15871) );
  AND2_X1 U12967 ( .A1(n13266), .A2(n13265), .ZN(n20145) );
  AND2_X1 U12968 ( .A1(n13186), .A2(n13185), .ZN(n20114) );
  INV_X1 U12969 ( .A(n20004), .ZN(n13235) );
  INV_X1 U12970 ( .A(n20020), .ZN(n20019) );
  INV_X2 U12971 ( .A(n20021), .ZN(n13397) );
  INV_X1 U12972 ( .A(n15889), .ZN(n20036) );
  AND2_X1 U12973 ( .A1(n13731), .A2(n13724), .ZN(n20049) );
  INV_X1 U12974 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20086) );
  INV_X1 U12975 ( .A(n20062), .ZN(n20073) );
  NAND2_X1 U12976 ( .A1(n20218), .A2(n20504), .ZN(n20177) );
  NAND2_X1 U12977 ( .A1(n20218), .A2(n20535), .ZN(n20210) );
  NAND2_X1 U12978 ( .A1(n20218), .A2(n20424), .ZN(n20245) );
  NAND2_X1 U12979 ( .A1(n20343), .A2(n20504), .ZN(n20300) );
  NAND2_X1 U12980 ( .A1(n20343), .A2(n20535), .ZN(n20341) );
  NAND2_X1 U12981 ( .A1(n20343), .A2(n20342), .ZN(n20366) );
  NAND2_X1 U12982 ( .A1(n20373), .A2(n20504), .ZN(n20423) );
  OR2_X1 U12983 ( .A1(n20481), .A2(n20403), .ZN(n20467) );
  OR2_X1 U12984 ( .A1(n20481), .A2(n20567), .ZN(n20503) );
  OR2_X1 U12985 ( .A1(n20481), .A2(n20480), .ZN(n20534) );
  NAND2_X1 U12986 ( .A1(n20539), .A2(n20535), .ZN(n20608) );
  NAND2_X1 U12987 ( .A1(n20539), .A2(n20342), .ZN(n20674) );
  NOR2_X1 U12988 ( .A1(n20613), .A2(n15734), .ZN(n16008) );
  AND2_X1 U12989 ( .A1(n20777), .A2(n19906), .ZN(n20757) );
  INV_X1 U12990 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20698) );
  NOR2_X1 U12991 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20686), .ZN(n20779) );
  INV_X1 U12992 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19630) );
  NAND2_X1 U12993 ( .A1(n19878), .A2(n14758), .ZN(n18925) );
  INV_X1 U12994 ( .A(n18944), .ZN(n18911) );
  INV_X1 U12995 ( .A(n18901), .ZN(n18934) );
  NAND2_X1 U12996 ( .A1(n13675), .A2(n18988), .ZN(n18984) );
  NAND2_X1 U12997 ( .A1(n19157), .A2(n14979), .ZN(n20787) );
  AND2_X1 U12998 ( .A1(n12808), .A2(n12850), .ZN(n14979) );
  NAND2_X1 U12999 ( .A1(n14979), .A2(n12818), .ZN(n13614) );
  NAND2_X1 U13000 ( .A1(n14979), .A2(n12809), .ZN(n14996) );
  OR2_X1 U13001 ( .A1(n19049), .A2(n11422), .ZN(n19014) );
  NAND2_X1 U13002 ( .A1(n12855), .A2(n19891), .ZN(n19049) );
  OR2_X1 U13003 ( .A1(n12852), .A2(n12851), .ZN(n12897) );
  INV_X1 U13004 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18831) );
  INV_X1 U13005 ( .A(n19089), .ZN(n16166) );
  NOR2_X1 U13006 ( .A1(n12335), .A2(n12334), .ZN(n12350) );
  INV_X1 U13007 ( .A(n16217), .ZN(n16204) );
  NAND2_X1 U13008 ( .A1(n12316), .A2(n19872), .ZN(n16227) );
  INV_X1 U13009 ( .A(n15669), .ZN(n15552) );
  NAND2_X1 U13010 ( .A1(n19414), .A2(n19354), .ZN(n19189) );
  NAND2_X1 U13011 ( .A1(n19354), .A2(n19832), .ZN(n19274) );
  NAND2_X1 U13012 ( .A1(n19383), .A2(n19832), .ZN(n19317) );
  INV_X1 U13013 ( .A(n19379), .ZN(n19358) );
  NAND2_X1 U13014 ( .A1(n19690), .A2(n19354), .ZN(n19406) );
  INV_X1 U13015 ( .A(n19445), .ZN(n19441) );
  AND2_X1 U13016 ( .A1(n19456), .A2(n19455), .ZN(n19481) );
  NAND2_X1 U13017 ( .A1(n19625), .A2(n19414), .ZN(n19486) );
  NAND2_X1 U13018 ( .A1(n19625), .A2(n19832), .ZN(n19544) );
  INV_X1 U13019 ( .A(n19703), .ZN(n19646) );
  INV_X1 U13020 ( .A(n19715), .ZN(n19656) );
  INV_X1 U13021 ( .A(n19709), .ZN(n19654) );
  INV_X1 U13022 ( .A(n19609), .ZN(n19724) );
  NAND2_X1 U13023 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19752), .ZN(n16236) );
  INV_X1 U13024 ( .A(n19831), .ZN(n19758) );
  NAND2_X1 U13025 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19763), .ZN(n19897) );
  INV_X1 U13026 ( .A(n18731), .ZN(n18729) );
  INV_X1 U13027 ( .A(n12728), .ZN(n16393) );
  INV_X1 U13028 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17511) );
  INV_X1 U13029 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17007) );
  INV_X1 U13030 ( .A(n16748), .ZN(n16784) );
  NAND2_X1 U13031 ( .A1(n17099), .A2(n17185), .ZN(n17085) );
  NOR2_X1 U13032 ( .A1(n12448), .A2(n12447), .ZN(n17226) );
  INV_X1 U13033 ( .A(n17261), .ZN(n17273) );
  NAND2_X1 U13034 ( .A1(n17306), .A2(n17252), .ZN(n17304) );
  INV_X1 U13035 ( .A(n17362), .ZN(n17357) );
  INV_X1 U13036 ( .A(n17355), .ZN(n17364) );
  INV_X1 U13037 ( .A(n17599), .ZN(n17624) );
  INV_X1 U13038 ( .A(n17615), .ZN(n17642) );
  INV_X1 U13039 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17700) );
  INV_X1 U13040 ( .A(n18026), .ZN(n18049) );
  INV_X1 U13041 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17839) );
  INV_X1 U13042 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17885) );
  INV_X1 U13043 ( .A(n17936), .ZN(n17960) );
  NAND2_X1 U13044 ( .A1(n16288), .A2(n18026), .ZN(n18041) );
  AND2_X1 U13045 ( .A1(n12695), .A2(n16389), .ZN(n18710) );
  INV_X1 U13046 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18545) );
  INV_X1 U13047 ( .A(n18403), .ZN(n18442) );
  INV_X1 U13048 ( .A(n18711), .ZN(n18561) );
  INV_X1 U13049 ( .A(n18664), .ZN(n18575) );
  OAI211_X1 U13050 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18589), .B(n18652), .ZN(n18714) );
  INV_X1 U13051 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18589) );
  NAND2_X1 U13052 ( .A1(n18589), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18725) );
  NOR2_X1 U13053 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12746), .ZN(n16376)
         );
  INV_X1 U13054 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19786) );
  OAI21_X1 U13055 ( .B1(n14086), .B2(n14297), .A(n10030), .ZN(P1_U2842) );
  NAND2_X1 U13056 ( .A1(n12387), .A2(n12386), .ZN(P1_U2873) );
  INV_X1 U13057 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10726) );
  NAND2_X2 U13058 ( .A1(n10061), .A2(n10048), .ZN(n10126) );
  INV_X1 U13059 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10900) );
  INV_X1 U13060 ( .A(n10047), .ZN(n10058) );
  INV_X2 U13061 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12996) );
  NAND2_X1 U13062 ( .A1(n10160), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10057) );
  AND2_X2 U13063 ( .A1(n10048), .A2(n10065), .ZN(n10267) );
  AND2_X2 U13064 ( .A1(n10065), .A2(n12968), .ZN(n10273) );
  AOI22_X1 U13065 ( .A1(n10267), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10273), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10056) );
  NAND2_X1 U13066 ( .A1(n10268), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10055) );
  INV_X1 U13067 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10052) );
  INV_X1 U13068 ( .A(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10051) );
  OAI22_X1 U13069 ( .A1(n10262), .A2(n10052), .B1(n9618), .B2(n10051), .ZN(
        n10053) );
  INV_X1 U13070 ( .A(n10053), .ZN(n10054) );
  AOI22_X1 U13071 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10197), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10071) );
  AND2_X2 U13072 ( .A1(n10060), .A2(n13446), .ZN(n10199) );
  AOI22_X1 U13073 ( .A1(n10601), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10199), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10070) );
  AOI22_X1 U13074 ( .A1(n10198), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10849), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10062) );
  INV_X1 U13075 ( .A(n10062), .ZN(n10068) );
  AND2_X2 U13076 ( .A1(n10065), .A2(n13446), .ZN(n10200) );
  AOI22_X1 U13077 ( .A1(n10858), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10200), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10066) );
  INV_X1 U13078 ( .A(n10066), .ZN(n10067) );
  INV_X1 U13079 ( .A(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10073) );
  INV_X1 U13080 ( .A(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10927) );
  OAI22_X1 U13081 ( .A1(n10260), .A2(n10073), .B1(n10126), .B2(n10927), .ZN(
        n10076) );
  INV_X1 U13082 ( .A(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10074) );
  INV_X1 U13083 ( .A(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10925) );
  OAI22_X1 U13084 ( .A1(n9618), .A2(n10074), .B1(n10262), .B2(n10925), .ZN(
        n10075) );
  NOR2_X1 U13085 ( .A1(n10076), .A2(n10075), .ZN(n10080) );
  AOI22_X1 U13086 ( .A1(n10267), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10273), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10079) );
  NAND2_X1 U13087 ( .A1(n10160), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10078) );
  NAND2_X1 U13088 ( .A1(n9622), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10077) );
  AOI22_X1 U13089 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10197), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10084) );
  AOI22_X1 U13090 ( .A1(n10601), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10199), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10083) );
  AOI22_X1 U13091 ( .A1(n10858), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10200), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10082) );
  AOI22_X1 U13092 ( .A1(n10198), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10849), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10081) );
  INV_X1 U13093 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10089) );
  INV_X1 U13094 ( .A(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10088) );
  INV_X1 U13095 ( .A(n10090), .ZN(n10094) );
  NAND2_X1 U13096 ( .A1(n9622), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10093) );
  NAND2_X1 U13097 ( .A1(n10849), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10092) );
  INV_X1 U13098 ( .A(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10975) );
  NAND4_X1 U13099 ( .A1(n10094), .A2(n10093), .A3(n10092), .A4(n10091), .ZN(
        n10098) );
  INV_X1 U13100 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10406) );
  NAND2_X1 U13101 ( .A1(n10267), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10096) );
  NAND2_X1 U13102 ( .A1(n10601), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10095) );
  OAI211_X1 U13103 ( .C1(n9604), .C2(n10406), .A(n10096), .B(n10095), .ZN(
        n10097) );
  NOR2_X1 U13104 ( .A1(n10098), .A2(n10097), .ZN(n10103) );
  AOI22_X1 U13105 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10200), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10101) );
  NAND2_X1 U13106 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10099) );
  AOI22_X1 U13107 ( .A1(n10511), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10199), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10102) );
  INV_X1 U13108 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10104) );
  OR2_X1 U13109 ( .A1(n10260), .A2(n10104), .ZN(n10108) );
  NAND2_X1 U13110 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10107) );
  NAND2_X1 U13111 ( .A1(n10267), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10106) );
  NAND2_X1 U13112 ( .A1(n10858), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10105) );
  NAND3_X1 U13113 ( .A1(n10108), .A2(n10107), .A3(n10043), .ZN(n10109) );
  NAND2_X1 U13114 ( .A1(n10199), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10111) );
  NAND2_X1 U13115 ( .A1(n10273), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10110) );
  OAI211_X1 U13116 ( .C1(n9604), .C2(n10479), .A(n10111), .B(n10110), .ZN(
        n10112) );
  INV_X1 U13117 ( .A(n10112), .ZN(n10119) );
  INV_X1 U13118 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10113) );
  NAND2_X1 U13119 ( .A1(n10198), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10116) );
  NAND2_X1 U13120 ( .A1(n10849), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10115) );
  NAND2_X1 U13121 ( .A1(n10200), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10114) );
  AND2_X2 U13122 ( .A1(n10119), .A2(n10118), .ZN(n10123) );
  NAND2_X1 U13123 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10122) );
  NAND2_X1 U13124 ( .A1(n9622), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10121) );
  NAND2_X1 U13125 ( .A1(n10268), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10129) );
  INV_X1 U13126 ( .A(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10125) );
  NAND2_X1 U13127 ( .A1(n10316), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10127) );
  NAND2_X1 U13128 ( .A1(n10198), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10134) );
  NAND2_X1 U13129 ( .A1(n10858), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10133) );
  NAND2_X1 U13130 ( .A1(n10200), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10132) );
  NAND2_X1 U13131 ( .A1(n10849), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10131) );
  NAND2_X1 U13132 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10138) );
  NAND2_X1 U13133 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10137) );
  NAND2_X1 U13134 ( .A1(n10601), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10136) );
  NAND2_X1 U13135 ( .A1(n10199), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10135) );
  NAND2_X1 U13136 ( .A1(n10267), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10140) );
  NAND2_X1 U13137 ( .A1(n10273), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10139) );
  OAI211_X1 U13138 ( .C1(n9604), .C2(n10388), .A(n10140), .B(n10139), .ZN(
        n10141) );
  INV_X1 U13139 ( .A(n10141), .ZN(n10142) );
  NAND2_X1 U13140 ( .A1(n10601), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10149) );
  NAND2_X1 U13141 ( .A1(n10316), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10148) );
  NAND2_X1 U13142 ( .A1(n10858), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10147) );
  NAND2_X1 U13143 ( .A1(n10849), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10146) );
  NAND2_X1 U13144 ( .A1(n10198), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10153) );
  INV_X1 U13145 ( .A(n10199), .ZN(n11009) );
  NAND2_X1 U13146 ( .A1(n10199), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10152) );
  NAND2_X1 U13147 ( .A1(n10267), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10151) );
  NAND2_X1 U13148 ( .A1(n10200), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10150) );
  AOI22_X1 U13149 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10516), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10159) );
  NAND2_X1 U13150 ( .A1(n9622), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10158) );
  INV_X1 U13151 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10155) );
  NAND2_X1 U13152 ( .A1(n9583), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10156) );
  NAND2_X1 U13153 ( .A1(n10273), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10163) );
  NAND2_X1 U13154 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10162) );
  OAI211_X1 U13155 ( .C1(n9604), .C2(n11030), .A(n10163), .B(n10162), .ZN(
        n10164) );
  INV_X1 U13156 ( .A(n10164), .ZN(n10165) );
  AND2_X1 U13157 ( .A1(n13016), .A2(n10229), .ZN(n10169) );
  OAI22_X1 U13158 ( .A1(n10262), .A2(n10830), .B1(n9618), .B2(n10170), .ZN(
        n10171) );
  INV_X1 U13159 ( .A(n10171), .ZN(n10175) );
  NAND2_X1 U13160 ( .A1(n10268), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10174) );
  NAND2_X1 U13161 ( .A1(n10316), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10172) );
  INV_X1 U13162 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10176) );
  INV_X1 U13163 ( .A(n10200), .ZN(n10885) );
  NAND2_X1 U13164 ( .A1(n10200), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10178) );
  NAND2_X1 U13165 ( .A1(n10849), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10177) );
  NAND2_X1 U13166 ( .A1(n10160), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10181) );
  NAND2_X1 U13167 ( .A1(n10267), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10180) );
  NAND2_X1 U13168 ( .A1(n10273), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10179) );
  NAND2_X1 U13169 ( .A1(n10197), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10185) );
  NAND2_X1 U13170 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10184) );
  NAND2_X1 U13171 ( .A1(n10601), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10183) );
  NAND2_X1 U13172 ( .A1(n10199), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10182) );
  XNOR2_X1 U13173 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12836) );
  INV_X1 U13174 ( .A(n10242), .ZN(n10228) );
  NAND2_X1 U13175 ( .A1(n10228), .A2(n11078), .ZN(n11233) );
  INV_X1 U13176 ( .A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10706) );
  NAND2_X1 U13177 ( .A1(n10858), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10189) );
  OAI21_X1 U13178 ( .B1(n10260), .B2(n10706), .A(n10189), .ZN(n10192) );
  INV_X1 U13179 ( .A(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10190) );
  OAI22_X1 U13180 ( .A1(n10087), .A2(n10190), .B1(n10262), .B2(n10873), .ZN(
        n10191) );
  NOR2_X1 U13181 ( .A1(n10192), .A2(n10191), .ZN(n10196) );
  AOI22_X1 U13182 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10601), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10195) );
  NAND2_X1 U13183 ( .A1(n10160), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10194) );
  NAND2_X1 U13184 ( .A1(n9622), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10193) );
  NAND4_X1 U13185 ( .A1(n10196), .A2(n10195), .A3(n10194), .A4(n10193), .ZN(
        n10206) );
  AOI22_X1 U13186 ( .A1(n10316), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10273), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10204) );
  AOI22_X1 U13187 ( .A1(n10198), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9583), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U13188 ( .A1(n10199), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10267), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10202) );
  AOI22_X1 U13189 ( .A1(n10200), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10849), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10201) );
  NAND4_X1 U13190 ( .A1(n10204), .A2(n10203), .A3(n10202), .A4(n10201), .ZN(
        n10205) );
  INV_X1 U13191 ( .A(n10224), .ZN(n10223) );
  NAND2_X1 U13192 ( .A1(n10229), .A2(n10209), .ZN(n10207) );
  INV_X1 U13193 ( .A(n10207), .ZN(n10435) );
  OAI21_X1 U13194 ( .B1(n12753), .B2(n12836), .A(n13014), .ZN(n10220) );
  NAND2_X1 U13195 ( .A1(n10233), .A2(n10210), .ZN(n10231) );
  NAND2_X1 U13196 ( .A1(n10231), .A2(n20122), .ZN(n10248) );
  NAND2_X1 U13197 ( .A1(n10212), .A2(n10229), .ZN(n10235) );
  NAND2_X1 U13198 ( .A1(n10235), .A2(n10207), .ZN(n10208) );
  NAND2_X1 U13199 ( .A1(n10248), .A2(n10208), .ZN(n10217) );
  INV_X1 U13200 ( .A(n10212), .ZN(n10213) );
  NAND2_X1 U13201 ( .A1(n10218), .A2(n20117), .ZN(n10214) );
  NAND2_X1 U13202 ( .A1(n10215), .A2(n10214), .ZN(n10216) );
  NOR2_X1 U13203 ( .A1(n10217), .A2(n10216), .ZN(n10227) );
  NOR2_X1 U13204 ( .A1(n10218), .A2(n10224), .ZN(n10219) );
  NAND2_X1 U13205 ( .A1(n12359), .A2(n12357), .ZN(n13018) );
  NAND2_X1 U13206 ( .A1(n11312), .A2(n10247), .ZN(n11248) );
  NAND2_X1 U13207 ( .A1(n11248), .A2(n10221), .ZN(n12947) );
  AND2_X1 U13208 ( .A1(n20117), .A2(n10224), .ZN(n10225) );
  INV_X1 U13209 ( .A(n10227), .ZN(n10252) );
  NAND2_X1 U13210 ( .A1(n11078), .A2(n10209), .ZN(n10230) );
  AND2_X1 U13211 ( .A1(n10230), .A2(n10229), .ZN(n11219) );
  AOI21_X1 U13212 ( .B1(n11063), .B2(n10233), .A(n10223), .ZN(n10234) );
  NAND2_X1 U13213 ( .A1(n10253), .A2(n10234), .ZN(n12945) );
  INV_X1 U13214 ( .A(n10235), .ZN(n10236) );
  NAND2_X1 U13215 ( .A1(n10253), .A2(n14692), .ZN(n10237) );
  NAND4_X1 U13216 ( .A1(n10239), .A2(n10238), .A3(n12945), .A4(n10237), .ZN(
        n10240) );
  MUX2_X1 U13217 ( .A(n11227), .B(n15738), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n10241) );
  OR2_X1 U13218 ( .A1(n10242), .A2(n10209), .ZN(n13031) );
  NAND2_X1 U13219 ( .A1(n12994), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19904) );
  INV_X1 U13220 ( .A(n19904), .ZN(n10244) );
  AND3_X1 U13221 ( .A1(n13031), .A2(n10244), .A3(n10243), .ZN(n10251) );
  NAND2_X1 U13222 ( .A1(n10245), .A2(n13252), .ZN(n10250) );
  AND2_X1 U13223 ( .A1(n12970), .A2(n14087), .ZN(n12794) );
  NAND2_X1 U13224 ( .A1(n12794), .A2(n10248), .ZN(n10249) );
  NAND2_X1 U13225 ( .A1(n10252), .A2(n13624), .ZN(n12944) );
  NAND3_X1 U13226 ( .A1(n10253), .A2(n10222), .A3(n14692), .ZN(n10254) );
  NAND3_X1 U13227 ( .A1(n10255), .A2(n12944), .A3(n10254), .ZN(n10303) );
  NAND2_X1 U13228 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10339) );
  OAI21_X1 U13229 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n10339), .ZN(n20430) );
  OR2_X1 U13230 ( .A1(n15738), .A2(n20505), .ZN(n10331) );
  OAI21_X1 U13231 ( .B1(n11227), .B2(n20430), .A(n10331), .ZN(n10256) );
  NAND2_X1 U13232 ( .A1(n9591), .A2(n10258), .ZN(n20150) );
  NAND2_X1 U13233 ( .A1(n10335), .A2(n20150), .ZN(n13647) );
  INV_X1 U13234 ( .A(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10871) );
  INV_X1 U13235 ( .A(n10849), .ZN(n10882) );
  NAND2_X1 U13236 ( .A1(n9586), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10261) );
  OAI21_X1 U13237 ( .B1(n10978), .B2(n10871), .A(n10261), .ZN(n10266) );
  INV_X1 U13238 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10264) );
  INV_X1 U13239 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10263) );
  OAI22_X1 U13240 ( .A1(n10308), .A2(n10264), .B1(n11039), .B2(n10263), .ZN(
        n10265) );
  NOR2_X1 U13241 ( .A1(n10266), .A2(n10265), .ZN(n10272) );
  AOI22_X1 U13242 ( .A1(n10392), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10267), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10271) );
  INV_X2 U13243 ( .A(n9619), .ZN(n10585) );
  NAND2_X1 U13244 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10270) );
  NAND2_X1 U13245 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10269) );
  NAND4_X1 U13246 ( .A1(n10272), .A2(n10271), .A3(n10270), .A4(n10269), .ZN(
        n10279) );
  INV_X1 U13247 ( .A(n10954), .ZN(n10576) );
  AOI22_X1 U13248 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U13249 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10276) );
  AOI22_X1 U13250 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10275) );
  AOI22_X1 U13251 ( .A1(n10601), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10273), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10274) );
  NAND4_X1 U13252 ( .A1(n10277), .A2(n10276), .A3(n10275), .A4(n10274), .ZN(
        n10278) );
  NAND2_X1 U13253 ( .A1(n11064), .A2(n11076), .ZN(n10280) );
  INV_X1 U13254 ( .A(n10370), .ZN(n10281) );
  NAND2_X1 U13255 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10299) );
  NOR2_X1 U13256 ( .A1(n10224), .A2(n10259), .ZN(n10363) );
  NAND2_X1 U13257 ( .A1(n10363), .A2(n11076), .ZN(n10298) );
  NAND2_X1 U13258 ( .A1(n10154), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10285) );
  NAND2_X1 U13259 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10284) );
  NAND2_X1 U13260 ( .A1(n11011), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10283) );
  NAND2_X1 U13261 ( .A1(n10840), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10282) );
  AOI22_X1 U13262 ( .A1(n10601), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10267), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10288) );
  NAND2_X1 U13263 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10287) );
  NAND2_X1 U13264 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10286) );
  NAND4_X1 U13265 ( .A1(n10289), .A2(n10288), .A3(n10287), .A4(n10286), .ZN(
        n10296) );
  INV_X1 U13266 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11038) );
  INV_X1 U13267 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11041) );
  OAI22_X1 U13268 ( .A1(n10978), .A2(n11038), .B1(n10999), .B2(n11041), .ZN(
        n10290) );
  INV_X1 U13269 ( .A(n10290), .ZN(n10294) );
  AOI22_X1 U13270 ( .A1(n10576), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U13271 ( .A1(n9583), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n9586), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10292) );
  AOI22_X1 U13272 ( .A1(n10392), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10273), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10291) );
  NAND4_X1 U13273 ( .A1(n10294), .A2(n10293), .A3(n10292), .A4(n10291), .ZN(
        n10295) );
  NAND2_X1 U13274 ( .A1(n11064), .A2(n11133), .ZN(n10297) );
  INV_X1 U13275 ( .A(n10302), .ZN(n10300) );
  INV_X1 U13276 ( .A(n10303), .ZN(n10304) );
  NAND2_X1 U13277 ( .A1(n10456), .A2(n10259), .ZN(n10325) );
  INV_X1 U13278 ( .A(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10307) );
  NAND2_X1 U13279 ( .A1(n9586), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10306) );
  OAI21_X1 U13280 ( .B1(n10978), .B2(n10307), .A(n10306), .ZN(n10311) );
  INV_X1 U13281 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10309) );
  INV_X1 U13282 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10832) );
  OAI22_X1 U13283 ( .A1(n10309), .A2(n10308), .B1(n11039), .B2(n10832), .ZN(
        n10310) );
  NOR2_X1 U13284 ( .A1(n10311), .A2(n10310), .ZN(n10315) );
  AOI22_X1 U13285 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n10700), .B1(
        n10267), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10314) );
  NAND2_X1 U13286 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10313) );
  NAND2_X1 U13287 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10312) );
  NAND4_X1 U13288 ( .A1(n10315), .A2(n10314), .A3(n10313), .A4(n10312), .ZN(
        n10322) );
  AOI22_X1 U13289 ( .A1(n10601), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10392), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U13290 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9583), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U13291 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10273), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10318) );
  AOI22_X1 U13292 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10317) );
  NAND4_X1 U13293 ( .A1(n10320), .A2(n10319), .A3(n10318), .A4(n10317), .ZN(
        n10321) );
  XNOR2_X1 U13294 ( .A(n11133), .B(n11075), .ZN(n10323) );
  NAND2_X1 U13295 ( .A1(n10323), .A2(n11064), .ZN(n10324) );
  INV_X1 U13296 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10834) );
  AOI21_X1 U13297 ( .B1(n13016), .B2(n11128), .A(n10259), .ZN(n10327) );
  NAND2_X1 U13298 ( .A1(n10223), .A2(n11075), .ZN(n10326) );
  INV_X1 U13299 ( .A(n11064), .ZN(n10328) );
  NOR2_X1 U13300 ( .A1(n10328), .A2(n11133), .ZN(n10329) );
  INV_X1 U13301 ( .A(n10331), .ZN(n10333) );
  OAI21_X1 U13302 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n10333), .A(
        n10332), .ZN(n10334) );
  INV_X1 U13303 ( .A(n10346), .ZN(n10344) );
  INV_X1 U13304 ( .A(n15738), .ZN(n10337) );
  NAND2_X1 U13305 ( .A1(n10337), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10343) );
  INV_X1 U13306 ( .A(n11227), .ZN(n10341) );
  INV_X1 U13307 ( .A(n10339), .ZN(n10338) );
  NAND2_X1 U13308 ( .A1(n10338), .A2(n20425), .ZN(n20474) );
  NAND2_X1 U13309 ( .A1(n10339), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10340) );
  NAND2_X1 U13310 ( .A1(n20474), .A2(n10340), .ZN(n20107) );
  NAND2_X1 U13311 ( .A1(n10341), .A2(n20107), .ZN(n10342) );
  NAND2_X2 U13312 ( .A1(n10347), .A2(n12910), .ZN(n12965) );
  INV_X1 U13313 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10908) );
  OAI22_X1 U13314 ( .A1(n10978), .A2(n10900), .B1(n10999), .B2(n10908), .ZN(
        n10351) );
  INV_X1 U13315 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10349) );
  INV_X1 U13316 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10348) );
  OAI22_X1 U13317 ( .A1(n10308), .A2(n10349), .B1(n11039), .B2(n10348), .ZN(
        n10350) );
  NOR2_X1 U13318 ( .A1(n10351), .A2(n10350), .ZN(n10355) );
  INV_X2 U13319 ( .A(n10833), .ZN(n11003) );
  AOI22_X1 U13320 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10354) );
  NAND2_X1 U13321 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10353) );
  NAND2_X1 U13322 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10352) );
  NAND4_X1 U13323 ( .A1(n10355), .A2(n10354), .A3(n10353), .A4(n10352), .ZN(
        n10361) );
  AOI22_X1 U13324 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10359) );
  AOI22_X1 U13325 ( .A1(n10601), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10358) );
  INV_X2 U13326 ( .A(n10885), .ZN(n11011) );
  AOI22_X1 U13327 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U13328 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10356) );
  NAND4_X1 U13329 ( .A1(n10359), .A2(n10358), .A3(n10357), .A4(n10356), .ZN(
        n10360) );
  NAND2_X1 U13330 ( .A1(n11064), .A2(n11066), .ZN(n10362) );
  OAI21_X2 U13331 ( .B1(n12965), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10362), 
        .ZN(n10365) );
  AOI22_X1 U13332 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10363), .B2(n11066), .ZN(n10364) );
  NOR3_X1 U13333 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20425), .A3(
        n20505), .ZN(n20349) );
  NAND2_X1 U13334 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20349), .ZN(
        n20344) );
  NAND2_X1 U13335 ( .A1(n20473), .A2(n20344), .ZN(n10366) );
  NAND3_X1 U13336 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20614) );
  INV_X1 U13337 ( .A(n20614), .ZN(n20623) );
  NAND2_X1 U13338 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20623), .ZN(
        n20610) );
  NAND2_X1 U13339 ( .A1(n10366), .A2(n20610), .ZN(n20099) );
  OAI22_X1 U13340 ( .A1(n11227), .A2(n20099), .B1(n15738), .B2(n20473), .ZN(
        n10367) );
  INV_X1 U13341 ( .A(n10367), .ZN(n10368) );
  INV_X1 U13342 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10371) );
  OAI22_X1 U13343 ( .A1(n10978), .A2(n10927), .B1(n10999), .B2(n10371), .ZN(
        n10375) );
  INV_X1 U13344 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10373) );
  INV_X1 U13345 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10372) );
  OAI22_X1 U13346 ( .A1(n10308), .A2(n10373), .B1(n11039), .B2(n10372), .ZN(
        n10374) );
  NOR2_X1 U13347 ( .A1(n10375), .A2(n10374), .ZN(n10379) );
  AOI22_X1 U13348 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10378) );
  NAND2_X1 U13349 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10377) );
  NAND2_X1 U13350 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10376) );
  NAND4_X1 U13351 ( .A1(n10379), .A2(n10378), .A3(n10377), .A4(n10376), .ZN(
        n10385) );
  AOI22_X1 U13352 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10383) );
  AOI22_X1 U13353 ( .A1(n10601), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U13354 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U13355 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10380) );
  NAND4_X1 U13356 ( .A1(n10383), .A2(n10382), .A3(n10381), .A4(n10380), .ZN(
        n10384) );
  AOI22_X1 U13357 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11215), .B2(n11107), .ZN(n10386) );
  NAND2_X1 U13358 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10404) );
  INV_X1 U13359 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10949) );
  INV_X1 U13360 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10959) );
  OAI22_X1 U13361 ( .A1(n10978), .A2(n10949), .B1(n10999), .B2(n10959), .ZN(
        n10391) );
  INV_X1 U13362 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10389) );
  OAI22_X1 U13363 ( .A1(n10308), .A2(n10389), .B1(n11039), .B2(n10388), .ZN(
        n10390) );
  NOR2_X1 U13364 ( .A1(n10391), .A2(n10390), .ZN(n10396) );
  AOI22_X1 U13365 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10395) );
  NAND2_X1 U13366 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10394) );
  NAND2_X1 U13367 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10393) );
  NAND4_X1 U13368 ( .A1(n10396), .A2(n10395), .A3(n10394), .A4(n10393), .ZN(
        n10402) );
  AOI22_X1 U13369 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10400) );
  AOI22_X1 U13370 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10399) );
  AOI22_X1 U13371 ( .A1(n11011), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10398) );
  AOI22_X1 U13372 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10397) );
  NAND4_X1 U13373 ( .A1(n10400), .A2(n10399), .A3(n10398), .A4(n10397), .ZN(
        n10401) );
  NAND2_X1 U13374 ( .A1(n11215), .A2(n11106), .ZN(n10403) );
  NAND2_X1 U13375 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10421) );
  INV_X1 U13376 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10405) );
  OAI22_X1 U13377 ( .A1(n10978), .A2(n10975), .B1(n10999), .B2(n10405), .ZN(
        n10409) );
  INV_X1 U13378 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10407) );
  OAI22_X1 U13379 ( .A1(n10308), .A2(n10407), .B1(n11039), .B2(n10406), .ZN(
        n10408) );
  NOR2_X1 U13380 ( .A1(n10409), .A2(n10408), .ZN(n10413) );
  AOI22_X1 U13381 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10412) );
  NAND2_X1 U13382 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10411) );
  NAND2_X1 U13383 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10410) );
  NAND4_X1 U13384 ( .A1(n10413), .A2(n10412), .A3(n10411), .A4(n10410), .ZN(
        n10419) );
  AOI22_X1 U13385 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10417) );
  AOI22_X1 U13386 ( .A1(n10601), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10416) );
  AOI22_X1 U13387 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10415) );
  AOI22_X1 U13388 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10414) );
  NAND4_X1 U13389 ( .A1(n10417), .A2(n10416), .A3(n10415), .A4(n10414), .ZN(
        n10418) );
  NAND2_X1 U13390 ( .A1(n11215), .A2(n11116), .ZN(n10420) );
  NAND2_X1 U13391 ( .A1(n10433), .A2(n10423), .ZN(n10424) );
  INV_X1 U13392 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13289) );
  NAND2_X1 U13393 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10472) );
  INV_X1 U13394 ( .A(n10495), .ZN(n10497) );
  INV_X1 U13395 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10426) );
  NAND2_X1 U13396 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n10471), .ZN(
        n10425) );
  NAND2_X1 U13397 ( .A1(n10426), .A2(n10425), .ZN(n10427) );
  NAND2_X1 U13398 ( .A1(n10497), .A2(n10427), .ZN(n19964) );
  NOR2_X2 U13399 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11020) );
  AOI22_X1 U13400 ( .A1(n19964), .A2(n11020), .B1(n12353), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10428) );
  OAI21_X1 U13401 ( .B1(n10509), .B2(n13289), .A(n10428), .ZN(n10429) );
  AOI21_X1 U13402 ( .B1(n11105), .B2(n10669), .A(n10429), .ZN(n13536) );
  INV_X1 U13403 ( .A(n13536), .ZN(n10443) );
  NAND2_X1 U13404 ( .A1(n10430), .A2(n13503), .ZN(n10432) );
  NAND2_X1 U13405 ( .A1(n10432), .A2(n10431), .ZN(n10434) );
  NAND2_X1 U13406 ( .A1(n10435), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10476) );
  INV_X1 U13407 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13438) );
  OAI21_X1 U13408 ( .B1(n20254), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20613), .ZN(n10437) );
  NAND2_X1 U13409 ( .A1(n11057), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n10436) );
  OAI211_X1 U13410 ( .C1(n10476), .C2(n13438), .A(n10437), .B(n10436), .ZN(
        n10440) );
  XNOR2_X1 U13411 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B(n10471), .ZN(
        n20035) );
  INV_X1 U13412 ( .A(n20035), .ZN(n10438) );
  NAND2_X1 U13413 ( .A1(n10438), .A2(n10780), .ZN(n10439) );
  AND2_X1 U13414 ( .A1(n10440), .A2(n10439), .ZN(n10441) );
  AOI21_X1 U13415 ( .B1(n11098), .B2(n10669), .A(n10441), .ZN(n13533) );
  INV_X1 U13416 ( .A(n13533), .ZN(n10442) );
  NAND2_X1 U13417 ( .A1(n10443), .A2(n10442), .ZN(n10477) );
  INV_X1 U13418 ( .A(n10444), .ZN(n10445) );
  NAND2_X1 U13419 ( .A1(n9673), .A2(n10445), .ZN(n10446) );
  NAND2_X1 U13420 ( .A1(n13479), .A2(n10669), .ZN(n10452) );
  AOI22_X1 U13421 ( .A1(n11057), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20613), .ZN(n10450) );
  INV_X1 U13422 ( .A(n10476), .ZN(n10448) );
  NAND2_X1 U13423 ( .A1(n10448), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10449) );
  AND2_X1 U13424 ( .A1(n10450), .A2(n10449), .ZN(n10451) );
  NAND2_X1 U13425 ( .A1(n10452), .A2(n10451), .ZN(n13104) );
  NAND2_X1 U13426 ( .A1(n11070), .A2(n10233), .ZN(n10455) );
  NAND2_X1 U13427 ( .A1(n10455), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12956) );
  NAND2_X1 U13428 ( .A1(n10457), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n10459) );
  NAND2_X1 U13429 ( .A1(n20613), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10458) );
  OAI211_X1 U13430 ( .C1(n10476), .C2(n9875), .A(n10459), .B(n10458), .ZN(
        n10460) );
  AOI21_X1 U13431 ( .B1(n13631), .B2(n10669), .A(n10460), .ZN(n12957) );
  NAND2_X1 U13432 ( .A1(n12957), .A2(n10780), .ZN(n10461) );
  NAND2_X1 U13433 ( .A1(n12958), .A2(n10461), .ZN(n13103) );
  NAND2_X1 U13434 ( .A1(n13104), .A2(n13103), .ZN(n13463) );
  INV_X1 U13435 ( .A(n13463), .ZN(n10469) );
  XNOR2_X1 U13436 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14230) );
  AOI21_X1 U13437 ( .B1(n11020), .B2(n14230), .A(n12353), .ZN(n10466) );
  NAND2_X1 U13438 ( .A1(n11057), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n10465) );
  OAI211_X1 U13439 ( .C1(n10476), .C2(n10059), .A(n10466), .B(n10465), .ZN(
        n10467) );
  INV_X1 U13440 ( .A(n10467), .ZN(n10468) );
  NAND2_X1 U13441 ( .A1(n10469), .A2(n13459), .ZN(n13461) );
  NAND2_X1 U13442 ( .A1(n12353), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13460) );
  NAND2_X1 U13443 ( .A1(n11088), .A2(n10669), .ZN(n10475) );
  AOI21_X1 U13444 ( .B1(n13529), .B2(n10472), .A(n10471), .ZN(n19994) );
  INV_X1 U13445 ( .A(n12353), .ZN(n10572) );
  OAI22_X1 U13446 ( .A1(n19994), .A2(n11055), .B1(n10572), .B2(n13529), .ZN(
        n10473) );
  AOI21_X1 U13447 ( .B1(n11057), .B2(P1_EAX_REG_3__SCAN_IN), .A(n10473), .ZN(
        n10474) );
  NAND2_X2 U13448 ( .A1(n13456), .A2(n13455), .ZN(n13534) );
  INV_X1 U13449 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13584) );
  NAND2_X1 U13450 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10494) );
  NAND2_X1 U13451 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10478) );
  OAI21_X1 U13452 ( .B1(n10978), .B2(n10113), .A(n10478), .ZN(n10482) );
  INV_X1 U13453 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10480) );
  OAI22_X1 U13454 ( .A1(n10308), .A2(n10480), .B1(n11039), .B2(n10479), .ZN(
        n10481) );
  NOR2_X1 U13455 ( .A1(n10482), .A2(n10481), .ZN(n10486) );
  AOI22_X1 U13456 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10485) );
  NAND2_X1 U13457 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10484) );
  NAND2_X1 U13458 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10483) );
  NAND4_X1 U13459 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n10492) );
  AOI22_X1 U13460 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13461 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13462 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13463 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10487) );
  NAND4_X1 U13464 ( .A1(n10490), .A2(n10489), .A3(n10488), .A4(n10487), .ZN(
        n10491) );
  NAND2_X1 U13465 ( .A1(n11215), .A2(n11126), .ZN(n10493) );
  NAND2_X1 U13466 ( .A1(n10502), .A2(n10503), .ZN(n11114) );
  NAND2_X1 U13467 ( .A1(n11114), .A2(n10669), .ZN(n10501) );
  INV_X1 U13468 ( .A(n10507), .ZN(n10499) );
  INV_X1 U13469 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10496) );
  NAND2_X1 U13470 ( .A1(n10497), .A2(n10496), .ZN(n10498) );
  NAND2_X1 U13471 ( .A1(n10499), .A2(n10498), .ZN(n19959) );
  AOI22_X1 U13472 ( .A1(n19959), .A2(n11020), .B1(n12353), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10500) );
  OAI211_X1 U13473 ( .C1(n10509), .C2(n13584), .A(n10501), .B(n10500), .ZN(
        n13556) );
  NAND2_X1 U13474 ( .A1(n13537), .A2(n13556), .ZN(n13549) );
  INV_X1 U13475 ( .A(n10502), .ZN(n10505) );
  INV_X1 U13476 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10662) );
  OAI22_X1 U13477 ( .A1(n11169), .A2(n10662), .B1(n11171), .B2(n11133), .ZN(
        n10506) );
  XNOR2_X1 U13478 ( .A(n11062), .B(n10506), .ZN(n11124) );
  INV_X1 U13479 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13297) );
  OAI21_X1 U13480 ( .B1(n10507), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n10531), .ZN(n19947) );
  AOI22_X1 U13481 ( .A1(n19947), .A2(n10780), .B1(n12353), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10508) );
  OAI21_X1 U13482 ( .B1(n10509), .B2(n13297), .A(n10508), .ZN(n10510) );
  AOI21_X1 U13483 ( .B1(n11124), .B2(n10669), .A(n10510), .ZN(n13550) );
  AOI22_X1 U13484 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10700), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U13485 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13486 ( .A1(n10902), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13487 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10512) );
  NAND4_X1 U13488 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(
        n10526) );
  NAND2_X1 U13489 ( .A1(n10154), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10520) );
  NAND2_X1 U13490 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10519) );
  NAND2_X1 U13491 ( .A1(n11011), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10518) );
  NAND2_X1 U13492 ( .A1(n10840), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10517) );
  AND4_X1 U13493 ( .A1(n10520), .A2(n10519), .A3(n10518), .A4(n10517), .ZN(
        n10524) );
  AOI22_X1 U13494 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10523) );
  NAND2_X1 U13495 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10522) );
  NAND2_X1 U13496 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10521) );
  NAND4_X1 U13497 ( .A1(n10524), .A2(n10523), .A3(n10522), .A4(n10521), .ZN(
        n10525) );
  OAI21_X1 U13498 ( .B1(n10526), .B2(n10525), .A(n10669), .ZN(n10530) );
  INV_X1 U13499 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10527) );
  XNOR2_X1 U13500 ( .A(n10531), .B(n10527), .ZN(n14220) );
  AOI22_X1 U13501 ( .A1(n14220), .A2(n11020), .B1(n12353), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10529) );
  NAND2_X1 U13502 ( .A1(n11057), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n10528) );
  XNOR2_X1 U13503 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n10565), .ZN(
        n19930) );
  INV_X1 U13504 ( .A(n19930), .ZN(n13760) );
  AOI22_X1 U13505 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13506 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U13507 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U13508 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10532) );
  NAND4_X1 U13509 ( .A1(n10535), .A2(n10534), .A3(n10533), .A4(n10532), .ZN(
        n10546) );
  INV_X1 U13510 ( .A(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10879) );
  NAND2_X1 U13511 ( .A1(n11011), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10536) );
  OAI21_X1 U13512 ( .B1(n10879), .B2(n10978), .A(n10536), .ZN(n10540) );
  INV_X1 U13513 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10538) );
  INV_X1 U13514 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10537) );
  OAI22_X1 U13515 ( .A1(n10308), .A2(n10538), .B1(n11039), .B2(n10537), .ZN(
        n10539) );
  NOR2_X1 U13516 ( .A1(n10540), .A2(n10539), .ZN(n10544) );
  AOI22_X1 U13517 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10543) );
  NAND2_X1 U13518 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10542) );
  NAND2_X1 U13519 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10541) );
  NAND4_X1 U13520 ( .A1(n10544), .A2(n10543), .A3(n10542), .A4(n10541), .ZN(
        n10545) );
  OAI21_X1 U13521 ( .B1(n10546), .B2(n10545), .A(n10669), .ZN(n10549) );
  NAND2_X1 U13522 ( .A1(n11057), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n10548) );
  NAND2_X1 U13523 ( .A1(n12353), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10547) );
  NAND3_X1 U13524 ( .A1(n10549), .A2(n10548), .A3(n10547), .ZN(n10550) );
  AOI21_X1 U13525 ( .B1(n13760), .B2(n10780), .A(n10550), .ZN(n13744) );
  AOI22_X1 U13526 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U13527 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U13528 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10552) );
  AOI22_X1 U13529 ( .A1(n10601), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10551) );
  NAND4_X1 U13530 ( .A1(n10554), .A2(n10553), .A3(n10552), .A4(n10551), .ZN(
        n10564) );
  NAND2_X1 U13531 ( .A1(n10154), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10558) );
  NAND2_X1 U13532 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10557) );
  NAND2_X1 U13533 ( .A1(n11011), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10556) );
  NAND2_X1 U13534 ( .A1(n10840), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10555) );
  AND4_X1 U13535 ( .A1(n10558), .A2(n10557), .A3(n10556), .A4(n10555), .ZN(
        n10562) );
  AOI22_X1 U13536 ( .A1(n9586), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10561) );
  NAND2_X1 U13537 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10560) );
  NAND2_X1 U13538 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10559) );
  NAND4_X1 U13539 ( .A1(n10562), .A2(n10561), .A3(n10560), .A4(n10559), .ZN(
        n10563) );
  NOR2_X1 U13540 ( .A1(n10564), .A2(n10563), .ZN(n10568) );
  XNOR2_X1 U13541 ( .A(n10569), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15848) );
  NAND2_X1 U13542 ( .A1(n15848), .A2(n10780), .ZN(n10567) );
  AOI22_X1 U13543 ( .A1(n11057), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12353), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10566) );
  OAI211_X1 U13544 ( .C1(n10568), .C2(n10653), .A(n10567), .B(n10566), .ZN(
        n13735) );
  INV_X1 U13545 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10573) );
  OAI21_X1 U13546 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n10570), .A(
        n10630), .ZN(n15900) );
  NAND2_X1 U13547 ( .A1(n15900), .A2(n10780), .ZN(n10571) );
  OAI21_X1 U13548 ( .B1(n10573), .B2(n10572), .A(n10571), .ZN(n10574) );
  AOI21_X1 U13549 ( .B1(n11057), .B2(P1_EAX_REG_11__SCAN_IN), .A(n10574), .ZN(
        n13763) );
  AOI22_X1 U13550 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10580) );
  AOI22_X1 U13551 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U13552 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10578) );
  AOI22_X1 U13553 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10577) );
  NAND4_X1 U13554 ( .A1(n10580), .A2(n10579), .A3(n10578), .A4(n10577), .ZN(
        n10591) );
  NAND2_X1 U13555 ( .A1(n10154), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10584) );
  NAND2_X1 U13556 ( .A1(n11011), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10583) );
  NAND2_X1 U13557 ( .A1(n9586), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10582) );
  NAND2_X1 U13558 ( .A1(n10840), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10581) );
  AND4_X1 U13559 ( .A1(n10584), .A2(n10583), .A3(n10582), .A4(n10581), .ZN(
        n10589) );
  AOI22_X1 U13560 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10588) );
  NAND2_X1 U13561 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10587) );
  NAND2_X1 U13562 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10586) );
  NAND4_X1 U13563 ( .A1(n10589), .A2(n10588), .A3(n10587), .A4(n10586), .ZN(
        n10590) );
  NOR2_X1 U13564 ( .A1(n10591), .A2(n10590), .ZN(n10592) );
  OR2_X1 U13565 ( .A1(n10653), .A2(n10592), .ZN(n14296) );
  INV_X1 U13566 ( .A(n14296), .ZN(n10593) );
  XNOR2_X1 U13567 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n10650), .ZN(
        n14508) );
  INV_X1 U13568 ( .A(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10596) );
  NAND2_X1 U13569 ( .A1(n9586), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10595) );
  OAI21_X1 U13570 ( .B1(n10596), .B2(n10999), .A(n10595), .ZN(n10600) );
  INV_X1 U13571 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10598) );
  INV_X1 U13572 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10597) );
  OAI22_X1 U13573 ( .A1(n10308), .A2(n10598), .B1(n11039), .B2(n10597), .ZN(
        n10599) );
  NOR2_X1 U13574 ( .A1(n10600), .A2(n10599), .ZN(n10605) );
  AOI22_X1 U13575 ( .A1(n10601), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10604) );
  NAND2_X1 U13576 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10603) );
  NAND2_X1 U13577 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10602) );
  NAND4_X1 U13578 ( .A1(n10605), .A2(n10604), .A3(n10603), .A4(n10602), .ZN(
        n10611) );
  AOI22_X1 U13579 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10609) );
  AOI22_X1 U13580 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10608) );
  AOI22_X1 U13581 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U13582 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10606) );
  NAND4_X1 U13583 ( .A1(n10609), .A2(n10608), .A3(n10607), .A4(n10606), .ZN(
        n10610) );
  OR2_X1 U13584 ( .A1(n10611), .A2(n10610), .ZN(n10612) );
  AOI22_X1 U13585 ( .A1(n10669), .A2(n10612), .B1(n12353), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10614) );
  NAND2_X1 U13586 ( .A1(n11057), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n10613) );
  OAI211_X1 U13587 ( .C1(n14508), .C2(n11055), .A(n10614), .B(n10613), .ZN(
        n14203) );
  INV_X1 U13588 ( .A(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10953) );
  OAI22_X1 U13589 ( .A1(n10978), .A2(n10959), .B1(n10126), .B2(n10953), .ZN(
        n10615) );
  INV_X1 U13590 ( .A(n10615), .ZN(n10619) );
  AOI22_X1 U13591 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10618) );
  AOI22_X1 U13592 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10617) );
  AOI22_X1 U13593 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10616) );
  NAND4_X1 U13594 ( .A1(n10619), .A2(n10618), .A3(n10617), .A4(n10616), .ZN(
        n10629) );
  NAND2_X1 U13595 ( .A1(n10154), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10623) );
  NAND2_X1 U13596 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10622) );
  NAND2_X1 U13597 ( .A1(n11011), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10621) );
  NAND2_X1 U13598 ( .A1(n10840), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10620) );
  AND4_X1 U13599 ( .A1(n10623), .A2(n10622), .A3(n10621), .A4(n10620), .ZN(
        n10627) );
  AOI22_X1 U13600 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10626) );
  NAND2_X1 U13601 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10625) );
  NAND2_X1 U13602 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10624) );
  NAND4_X1 U13603 ( .A1(n10627), .A2(n10626), .A3(n10625), .A4(n10624), .ZN(
        n10628) );
  NOR2_X1 U13604 ( .A1(n10629), .A2(n10628), .ZN(n10634) );
  NAND2_X1 U13605 ( .A1(n11057), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n10633) );
  XNOR2_X1 U13606 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n10630), .ZN(
        n15888) );
  INV_X1 U13607 ( .A(n15888), .ZN(n10631) );
  AOI22_X1 U13608 ( .A1(n12353), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n11020), .B2(n10631), .ZN(n10632) );
  OAI211_X1 U13609 ( .C1(n10653), .C2(n10634), .A(n10633), .B(n10632), .ZN(
        n13765) );
  INV_X1 U13610 ( .A(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10636) );
  NAND2_X1 U13611 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10635) );
  OAI21_X1 U13612 ( .B1(n10636), .B2(n10126), .A(n10635), .ZN(n10639) );
  INV_X1 U13613 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10637) );
  INV_X1 U13614 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11008) );
  OAI22_X1 U13615 ( .A1(n10308), .A2(n10637), .B1(n11039), .B2(n11008), .ZN(
        n10638) );
  NOR2_X1 U13616 ( .A1(n10639), .A2(n10638), .ZN(n10643) );
  AOI22_X1 U13617 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10642) );
  NAND2_X1 U13618 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10641) );
  NAND2_X1 U13619 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10640) );
  NAND4_X1 U13620 ( .A1(n10643), .A2(n10642), .A3(n10641), .A4(n10640), .ZN(
        n10649) );
  AOI22_X1 U13621 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10647) );
  AOI22_X1 U13622 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U13623 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10645) );
  AOI22_X1 U13624 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10644) );
  NAND4_X1 U13625 ( .A1(n10647), .A2(n10646), .A3(n10645), .A4(n10644), .ZN(
        n10648) );
  NOR2_X1 U13626 ( .A1(n10649), .A2(n10648), .ZN(n10654) );
  XNOR2_X1 U13627 ( .A(n10655), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14498) );
  NAND2_X1 U13628 ( .A1(n14498), .A2(n10780), .ZN(n10652) );
  AOI22_X1 U13629 ( .A1(n11057), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n12353), 
        .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10651) );
  OAI211_X1 U13630 ( .C1(n10654), .C2(n10653), .A(n10652), .B(n10651), .ZN(
        n13772) );
  NAND2_X1 U13631 ( .A1(n13769), .A2(n13772), .ZN(n13770) );
  XNOR2_X1 U13632 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n10678), .ZN(
        n15880) );
  INV_X1 U13633 ( .A(n15880), .ZN(n10676) );
  AOI22_X1 U13634 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11034), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10659) );
  AOI22_X1 U13635 ( .A1(n10902), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U13636 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13637 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10656) );
  NAND4_X1 U13638 ( .A1(n10659), .A2(n10658), .A3(n10657), .A4(n10656), .ZN(
        n10671) );
  NAND2_X1 U13639 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10660) );
  OAI21_X1 U13640 ( .B1(n11041), .B2(n10978), .A(n10660), .ZN(n10664) );
  INV_X1 U13641 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10661) );
  OAI22_X1 U13642 ( .A1(n10308), .A2(n10662), .B1(n11039), .B2(n10661), .ZN(
        n10663) );
  NOR2_X1 U13643 ( .A1(n10664), .A2(n10663), .ZN(n10668) );
  AOI22_X1 U13644 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10667) );
  NAND2_X1 U13645 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10666) );
  NAND2_X1 U13646 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10665) );
  NAND4_X1 U13647 ( .A1(n10668), .A2(n10667), .A3(n10666), .A4(n10665), .ZN(
        n10670) );
  OAI21_X1 U13648 ( .B1(n10671), .B2(n10670), .A(n10669), .ZN(n10674) );
  NAND2_X1 U13649 ( .A1(n11057), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n10673) );
  NAND2_X1 U13650 ( .A1(n12353), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10672) );
  NAND3_X1 U13651 ( .A1(n10674), .A2(n10673), .A3(n10672), .ZN(n10675) );
  AOI21_X1 U13652 ( .B1(n10676), .B2(n10780), .A(n10675), .ZN(n14286) );
  INV_X1 U13653 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15808) );
  XNOR2_X1 U13654 ( .A(n10699), .B(n15808), .ZN(n15814) );
  NAND2_X1 U13655 ( .A1(n15814), .A2(n10780), .ZN(n10698) );
  AOI22_X1 U13656 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n11033), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U13657 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U13658 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U13659 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10679) );
  NAND4_X1 U13660 ( .A1(n10682), .A2(n10681), .A3(n10680), .A4(n10679), .ZN(
        n10693) );
  AOI22_X1 U13661 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9623), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10691) );
  NAND2_X1 U13662 ( .A1(n10902), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10683) );
  OAI211_X1 U13663 ( .C1(n10684), .C2(n11039), .A(n10683), .B(n11055), .ZN(
        n10685) );
  INV_X1 U13664 ( .A(n10685), .ZN(n10690) );
  INV_X1 U13665 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10686) );
  OAI22_X1 U13666 ( .A1(n10999), .A2(n10176), .B1(n10308), .B2(n10686), .ZN(
        n10687) );
  INV_X1 U13667 ( .A(n10687), .ZN(n10689) );
  AOI22_X1 U13668 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10688) );
  NAND4_X1 U13669 ( .A1(n10691), .A2(n10690), .A3(n10689), .A4(n10688), .ZN(
        n10692) );
  NAND2_X1 U13670 ( .A1(n11023), .A2(n11055), .ZN(n10820) );
  OAI21_X1 U13671 ( .B1(n10693), .B2(n10692), .A(n10820), .ZN(n10696) );
  NOR2_X1 U13672 ( .A1(n15808), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10694) );
  AOI21_X1 U13673 ( .B1(n11057), .B2(P1_EAX_REG_16__SCAN_IN), .A(n10694), .ZN(
        n10695) );
  NAND2_X1 U13674 ( .A1(n10696), .A2(n10695), .ZN(n10697) );
  NAND2_X1 U13675 ( .A1(n10698), .A2(n10697), .ZN(n14275) );
  XNOR2_X1 U13676 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n10718), .ZN(
        n15872) );
  AOI22_X1 U13677 ( .A1(n11057), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n12353), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13678 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10704) );
  AOI22_X1 U13679 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U13680 ( .A1(n10902), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U13681 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10701) );
  NAND4_X1 U13682 ( .A1(n10704), .A2(n10703), .A3(n10702), .A4(n10701), .ZN(
        n10714) );
  INV_X1 U13683 ( .A(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10883) );
  NAND2_X1 U13684 ( .A1(n9586), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10705) );
  OAI21_X1 U13685 ( .B1(n10978), .B2(n10883), .A(n10705), .ZN(n10708) );
  INV_X1 U13686 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10886) );
  OAI22_X1 U13687 ( .A1(n10308), .A2(n10886), .B1(n11039), .B2(n10706), .ZN(
        n10707) );
  NOR2_X1 U13688 ( .A1(n10708), .A2(n10707), .ZN(n10712) );
  AOI22_X1 U13689 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10711) );
  NAND2_X1 U13690 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10710) );
  NAND2_X1 U13691 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10709) );
  NAND4_X1 U13692 ( .A1(n10712), .A2(n10711), .A3(n10710), .A4(n10709), .ZN(
        n10713) );
  INV_X1 U13693 ( .A(n11023), .ZN(n11052) );
  OAI21_X1 U13694 ( .B1(n10714), .B2(n10713), .A(n11052), .ZN(n10715) );
  OAI211_X1 U13695 ( .C1(n15872), .C2(n11055), .A(n10716), .B(n10715), .ZN(
        n14193) );
  INV_X1 U13696 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15796) );
  XNOR2_X1 U13697 ( .A(n10754), .B(n15796), .ZN(n15803) );
  AOI22_X1 U13698 ( .A1(n11057), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20613), .ZN(n10735) );
  AOI22_X1 U13699 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U13700 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U13701 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U13702 ( .A1(n9586), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10719) );
  NAND4_X1 U13703 ( .A1(n10722), .A2(n10721), .A3(n10720), .A4(n10719), .ZN(
        n10733) );
  AOI22_X1 U13704 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9623), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10731) );
  INV_X1 U13705 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10724) );
  NAND2_X1 U13706 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10723) );
  OAI211_X1 U13707 ( .C1(n10724), .C2(n10308), .A(n10723), .B(n11055), .ZN(
        n10725) );
  INV_X1 U13708 ( .A(n10725), .ZN(n10730) );
  INV_X1 U13709 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10907) );
  OAI22_X1 U13710 ( .A1(n10126), .A2(n10907), .B1(n11039), .B2(n10726), .ZN(
        n10727) );
  INV_X1 U13711 ( .A(n10727), .ZN(n10729) );
  AOI22_X1 U13712 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10728) );
  NAND4_X1 U13713 ( .A1(n10731), .A2(n10730), .A3(n10729), .A4(n10728), .ZN(
        n10732) );
  OAI21_X1 U13714 ( .B1(n10733), .B2(n10732), .A(n10820), .ZN(n10734) );
  AOI22_X1 U13715 ( .A1(n15803), .A2(n10780), .B1(n10735), .B2(n10734), .ZN(
        n14267) );
  NAND2_X1 U13716 ( .A1(n14192), .A2(n14267), .ZN(n14260) );
  NAND2_X1 U13717 ( .A1(n10154), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10739) );
  NAND2_X1 U13718 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10738) );
  NAND2_X1 U13719 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10737) );
  NAND2_X1 U13720 ( .A1(n10840), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10736) );
  AND4_X1 U13721 ( .A1(n10739), .A2(n10738), .A3(n10737), .A4(n10736), .ZN(
        n10743) );
  AOI22_X1 U13722 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10742) );
  NAND2_X1 U13723 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10741) );
  NAND2_X1 U13724 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10740) );
  NAND4_X1 U13725 ( .A1(n10743), .A2(n10742), .A3(n10741), .A4(n10740), .ZN(
        n10749) );
  AOI22_X1 U13726 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U13727 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U13728 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U13729 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10744) );
  NAND4_X1 U13730 ( .A1(n10747), .A2(n10746), .A3(n10745), .A4(n10744), .ZN(
        n10748) );
  NOR2_X1 U13731 ( .A1(n10749), .A2(n10748), .ZN(n10753) );
  NAND2_X1 U13732 ( .A1(n20613), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10750) );
  NAND2_X1 U13733 ( .A1(n11055), .A2(n10750), .ZN(n10751) );
  AOI21_X1 U13734 ( .B1(n11057), .B2(P1_EAX_REG_19__SCAN_IN), .A(n10751), .ZN(
        n10752) );
  OAI21_X1 U13735 ( .B1(n11023), .B2(n10753), .A(n10752), .ZN(n10761) );
  INV_X1 U13736 ( .A(n10802), .ZN(n10759) );
  INV_X1 U13737 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10757) );
  INV_X1 U13738 ( .A(n10755), .ZN(n10756) );
  NAND2_X1 U13739 ( .A1(n10757), .A2(n10756), .ZN(n10758) );
  NAND2_X1 U13740 ( .A1(n10759), .A2(n10758), .ZN(n15862) );
  NAND2_X1 U13741 ( .A1(n10761), .A2(n10760), .ZN(n14261) );
  INV_X1 U13742 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10764) );
  NAND2_X1 U13743 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10763) );
  OAI21_X1 U13744 ( .B1(n10764), .B2(n10999), .A(n10763), .ZN(n10766) );
  INV_X1 U13745 ( .A(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10951) );
  OAI22_X1 U13746 ( .A1(n10308), .A2(n10951), .B1(n11039), .B2(n10125), .ZN(
        n10765) );
  NOR2_X1 U13747 ( .A1(n10766), .A2(n10765), .ZN(n10770) );
  AOI22_X1 U13748 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10769) );
  NAND2_X1 U13749 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10768) );
  NAND2_X1 U13750 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10767) );
  NAND4_X1 U13751 ( .A1(n10770), .A2(n10769), .A3(n10768), .A4(n10767), .ZN(
        n10776) );
  AOI22_X1 U13752 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13753 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U13754 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13755 ( .A1(n11011), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10771) );
  NAND4_X1 U13756 ( .A1(n10774), .A2(n10773), .A3(n10772), .A4(n10771), .ZN(
        n10775) );
  NOR2_X1 U13757 ( .A1(n10776), .A2(n10775), .ZN(n10779) );
  INV_X1 U13758 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14465) );
  AOI21_X1 U13759 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14465), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10777) );
  AOI21_X1 U13760 ( .B1(n11057), .B2(P1_EAX_REG_20__SCAN_IN), .A(n10777), .ZN(
        n10778) );
  OAI21_X1 U13761 ( .B1(n11023), .B2(n10779), .A(n10778), .ZN(n10782) );
  XNOR2_X1 U13762 ( .A(n10802), .B(n14465), .ZN(n15781) );
  NAND2_X1 U13763 ( .A1(n15781), .A2(n10780), .ZN(n10781) );
  INV_X1 U13764 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10977) );
  NAND2_X1 U13765 ( .A1(n9586), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10783) );
  OAI21_X1 U13766 ( .B1(n10977), .B2(n10126), .A(n10783), .ZN(n10787) );
  INV_X1 U13767 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10785) );
  INV_X1 U13768 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10784) );
  OAI22_X1 U13769 ( .A1(n10308), .A2(n10785), .B1(n11039), .B2(n10784), .ZN(
        n10786) );
  NOR2_X1 U13770 ( .A1(n10787), .A2(n10786), .ZN(n10791) );
  AOI22_X1 U13771 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10790) );
  NAND2_X1 U13772 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10789) );
  NAND2_X1 U13773 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10788) );
  NAND4_X1 U13774 ( .A1(n10791), .A2(n10790), .A3(n10789), .A4(n10788), .ZN(
        n10797) );
  AOI22_X1 U13775 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10795) );
  AOI22_X1 U13776 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10858), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U13777 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U13778 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10792) );
  NAND4_X1 U13779 ( .A1(n10795), .A2(n10794), .A3(n10793), .A4(n10792), .ZN(
        n10796) );
  NOR2_X1 U13780 ( .A1(n10797), .A2(n10796), .ZN(n10801) );
  NAND2_X1 U13781 ( .A1(n20613), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10798) );
  NAND2_X1 U13782 ( .A1(n11055), .A2(n10798), .ZN(n10799) );
  AOI21_X1 U13783 ( .B1(n11057), .B2(P1_EAX_REG_21__SCAN_IN), .A(n10799), .ZN(
        n10800) );
  OAI21_X1 U13784 ( .B1(n11023), .B2(n10801), .A(n10800), .ZN(n10808) );
  INV_X1 U13785 ( .A(n10803), .ZN(n10805) );
  INV_X1 U13786 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10804) );
  NAND2_X1 U13787 ( .A1(n10805), .A2(n10804), .ZN(n10806) );
  NAND2_X1 U13788 ( .A1(n10825), .A2(n10806), .ZN(n15776) );
  NAND2_X1 U13789 ( .A1(n10808), .A2(n10807), .ZN(n14250) );
  AOI22_X1 U13790 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11034), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U13791 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11044), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10811) );
  AOI22_X1 U13792 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U13793 ( .A1(n10392), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10809) );
  NAND4_X1 U13794 ( .A1(n10812), .A2(n10811), .A3(n10810), .A4(n10809), .ZN(
        n10822) );
  AOI22_X1 U13795 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9623), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10819) );
  INV_X1 U13796 ( .A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10814) );
  NAND2_X1 U13797 ( .A1(n11003), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10813) );
  OAI211_X1 U13798 ( .C1(n10814), .C2(n10308), .A(n10813), .B(n11055), .ZN(
        n10815) );
  INV_X1 U13799 ( .A(n10815), .ZN(n10818) );
  AOI22_X1 U13800 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10840), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10817) );
  AOI22_X1 U13801 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10816) );
  NAND4_X1 U13802 ( .A1(n10819), .A2(n10818), .A3(n10817), .A4(n10816), .ZN(
        n10821) );
  OAI21_X1 U13803 ( .B1(n10822), .B2(n10821), .A(n10820), .ZN(n10824) );
  AOI22_X1 U13804 ( .A1(n11057), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20613), .ZN(n10823) );
  XNOR2_X1 U13805 ( .A(n10825), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14446) );
  AOI22_X1 U13806 ( .A1(n10824), .A2(n10823), .B1(n11020), .B2(n14446), .ZN(
        n14183) );
  INV_X1 U13807 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10827) );
  NAND2_X1 U13808 ( .A1(n10828), .A2(n10827), .ZN(n10829) );
  NAND2_X1 U13809 ( .A1(n10868), .A2(n10829), .ZN(n14440) );
  INV_X1 U13810 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10839) );
  INV_X1 U13811 ( .A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10831) );
  OAI22_X1 U13812 ( .A1(n10885), .A2(n10831), .B1(n10830), .B2(n10126), .ZN(
        n10836) );
  OAI22_X1 U13813 ( .A1(n10834), .A2(n10882), .B1(n10833), .B2(n10832), .ZN(
        n10835) );
  AOI211_X1 U13814 ( .C1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .C2(n9623), .A(
        n10836), .B(n10835), .ZN(n10838) );
  AOI22_X1 U13815 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n11044), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10837) );
  OAI211_X1 U13816 ( .C1(n10839), .C2(n9619), .A(n10838), .B(n10837), .ZN(
        n10846) );
  AOI22_X1 U13817 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U13818 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n11034), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U13819 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10842) );
  AOI22_X1 U13820 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n10154), .B1(
        n10840), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10841) );
  NAND4_X1 U13821 ( .A1(n10844), .A2(n10843), .A3(n10842), .A4(n10841), .ZN(
        n10845) );
  NOR2_X1 U13822 ( .A1(n10846), .A2(n10845), .ZN(n10869) );
  INV_X1 U13823 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U13824 ( .A1(n10154), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10848) );
  NAND2_X1 U13825 ( .A1(n11003), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10847) );
  OAI211_X1 U13826 ( .C1(n9587), .C2(n11040), .A(n10848), .B(n10847), .ZN(
        n10854) );
  INV_X1 U13827 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10850) );
  OAI22_X1 U13828 ( .A1(n10954), .A2(n11041), .B1(n10882), .B2(n10850), .ZN(
        n10853) );
  INV_X1 U13829 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10851) );
  OAI22_X1 U13830 ( .A1(n10161), .A2(n10851), .B1(n11009), .B2(n11030), .ZN(
        n10852) );
  OR3_X1 U13831 ( .A1(n10854), .A2(n10853), .A3(n10852), .ZN(n10863) );
  INV_X1 U13832 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10855) );
  OAI22_X1 U13833 ( .A1(n10978), .A2(n10855), .B1(n11039), .B2(n10155), .ZN(
        n10857) );
  NOR2_X1 U13834 ( .A1(n9619), .A2(n11038), .ZN(n10856) );
  AOI211_X1 U13835 ( .C1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .C2(n11012), .A(
        n10857), .B(n10856), .ZN(n10861) );
  AOI22_X1 U13836 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10858), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10860) );
  AOI22_X1 U13837 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10859) );
  NAND3_X1 U13838 ( .A1(n10861), .A2(n10860), .A3(n10859), .ZN(n10862) );
  NOR2_X1 U13839 ( .A1(n10863), .A2(n10862), .ZN(n10870) );
  XNOR2_X1 U13840 ( .A(n10869), .B(n10870), .ZN(n10866) );
  AOI21_X1 U13841 ( .B1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20613), .A(
        n11020), .ZN(n10865) );
  NAND2_X1 U13842 ( .A1(n11057), .A2(P1_EAX_REG_23__SCAN_IN), .ZN(n10864) );
  OAI211_X1 U13843 ( .C1(n10866), .C2(n11023), .A(n10865), .B(n10864), .ZN(
        n10867) );
  OAI21_X1 U13844 ( .B1(n11055), .B2(n14440), .A(n10867), .ZN(n14170) );
  XOR2_X1 U13845 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n10895), .Z(
        n14436) );
  INV_X1 U13846 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14432) );
  OAI21_X1 U13847 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14432), .A(n11055), 
        .ZN(n10893) );
  NOR2_X1 U13848 ( .A1(n10870), .A2(n10869), .ZN(n10917) );
  INV_X1 U13849 ( .A(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10872) );
  OAI22_X1 U13850 ( .A1(n10308), .A2(n10872), .B1(n11039), .B2(n10871), .ZN(
        n10876) );
  INV_X1 U13851 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10874) );
  OAI22_X1 U13852 ( .A1(n10978), .A2(n10874), .B1(n10999), .B2(n10873), .ZN(
        n10875) );
  AOI211_X1 U13853 ( .C1(n9623), .C2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n10876), .B(n10875), .ZN(n10878) );
  AOI22_X1 U13854 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10877) );
  OAI211_X1 U13855 ( .C1(n9619), .C2(n10879), .A(n10878), .B(n10877), .ZN(
        n10890) );
  AOI22_X1 U13856 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U13857 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10880) );
  NAND2_X1 U13858 ( .A1(n10881), .A2(n10880), .ZN(n10889) );
  OAI22_X1 U13859 ( .A1(n10954), .A2(n10883), .B1(n10882), .B2(n10538), .ZN(
        n10888) );
  INV_X1 U13860 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10884) );
  OAI22_X1 U13861 ( .A1(n10952), .A2(n10886), .B1(n10885), .B2(n10884), .ZN(
        n10887) );
  XNOR2_X1 U13862 ( .A(n10917), .B(n10916), .ZN(n10891) );
  NOR2_X1 U13863 ( .A1(n10891), .A2(n11023), .ZN(n10892) );
  AOI211_X1 U13864 ( .C1(n11057), .C2(P1_EAX_REG_24__SCAN_IN), .A(n10893), .B(
        n10892), .ZN(n10894) );
  AOI21_X1 U13865 ( .B1(n11020), .B2(n14436), .A(n10894), .ZN(n14160) );
  INV_X1 U13866 ( .A(n10896), .ZN(n10897) );
  OAI21_X1 U13867 ( .B1(n10897), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n10922), .ZN(n14424) );
  NAND2_X1 U13868 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10899) );
  NAND2_X1 U13869 ( .A1(n11033), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10898) );
  OAI211_X1 U13870 ( .C1(n10900), .C2(n11039), .A(n10899), .B(n10898), .ZN(
        n10901) );
  AOI21_X1 U13871 ( .B1(n9623), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A(n10901), .ZN(n10905) );
  AOI22_X1 U13872 ( .A1(n10902), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10904) );
  AOI22_X1 U13873 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10903) );
  NAND3_X1 U13874 ( .A1(n10905), .A2(n10904), .A3(n10903), .ZN(n10915) );
  INV_X1 U13875 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10906) );
  OAI22_X1 U13876 ( .A1(n10978), .A2(n10907), .B1(n10308), .B2(n10906), .ZN(
        n10910) );
  NOR2_X1 U13877 ( .A1(n9619), .A2(n10908), .ZN(n10909) );
  AOI211_X1 U13878 ( .C1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .C2(n11003), .A(
        n10910), .B(n10909), .ZN(n10913) );
  AOI22_X1 U13879 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U13880 ( .A1(n10576), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10911) );
  NAND3_X1 U13881 ( .A1(n10913), .A2(n10912), .A3(n10911), .ZN(n10914) );
  NOR2_X1 U13882 ( .A1(n10915), .A2(n10914), .ZN(n10924) );
  NAND2_X1 U13883 ( .A1(n10917), .A2(n10916), .ZN(n10923) );
  XNOR2_X1 U13884 ( .A(n10924), .B(n10923), .ZN(n10920) );
  AOI21_X1 U13885 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20613), .A(
        n11020), .ZN(n10919) );
  NAND2_X1 U13886 ( .A1(n10457), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n10918) );
  OAI211_X1 U13887 ( .C1(n10920), .C2(n11023), .A(n10919), .B(n10918), .ZN(
        n10921) );
  OAI21_X1 U13888 ( .B1(n11055), .B2(n14424), .A(n10921), .ZN(n14148) );
  XOR2_X1 U13889 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B(n10945), .Z(
        n14417) );
  INV_X1 U13890 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14413) );
  OAI21_X1 U13891 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14413), .A(n11055), 
        .ZN(n10943) );
  NOR2_X1 U13892 ( .A1(n10924), .A2(n10923), .ZN(n10967) );
  INV_X1 U13893 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10926) );
  OAI22_X1 U13894 ( .A1(n10978), .A2(n10926), .B1(n10999), .B2(n10925), .ZN(
        n10930) );
  INV_X1 U13895 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10928) );
  OAI22_X1 U13896 ( .A1(n10308), .A2(n10928), .B1(n11039), .B2(n10927), .ZN(
        n10929) );
  NOR2_X1 U13897 ( .A1(n10930), .A2(n10929), .ZN(n10934) );
  AOI22_X1 U13898 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10933) );
  NAND2_X1 U13899 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10932) );
  NAND2_X1 U13900 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10931) );
  NAND4_X1 U13901 ( .A1(n10934), .A2(n10933), .A3(n10932), .A4(n10931), .ZN(
        n10940) );
  AOI22_X1 U13902 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U13903 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U13904 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10936) );
  AOI22_X1 U13905 ( .A1(n10576), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10935) );
  NAND4_X1 U13906 ( .A1(n10938), .A2(n10937), .A3(n10936), .A4(n10935), .ZN(
        n10939) );
  OR2_X1 U13907 ( .A1(n10940), .A2(n10939), .ZN(n10966) );
  XNOR2_X1 U13908 ( .A(n10967), .B(n10966), .ZN(n10941) );
  NOR2_X1 U13909 ( .A1(n10941), .A2(n11023), .ZN(n10942) );
  AOI211_X1 U13910 ( .C1(n11057), .C2(P1_EAX_REG_26__SCAN_IN), .A(n10943), .B(
        n10942), .ZN(n10944) );
  AOI21_X1 U13911 ( .B1(n11020), .B2(n14417), .A(n10944), .ZN(n14133) );
  NAND2_X1 U13912 ( .A1(n14131), .A2(n14133), .ZN(n14120) );
  INV_X1 U13913 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10946) );
  NAND2_X1 U13914 ( .A1(n10947), .A2(n10946), .ZN(n10948) );
  NAND2_X1 U13915 ( .A1(n10993), .A2(n10948), .ZN(n14406) );
  INV_X1 U13916 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10950) );
  OAI22_X1 U13917 ( .A1(n10308), .A2(n10950), .B1(n11039), .B2(n10949), .ZN(
        n10956) );
  OAI22_X1 U13918 ( .A1(n10954), .A2(n10953), .B1(n10952), .B2(n10951), .ZN(
        n10955) );
  AOI211_X1 U13919 ( .C1(n9623), .C2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n10956), .B(n10955), .ZN(n10958) );
  AOI22_X1 U13920 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10957) );
  OAI211_X1 U13921 ( .C1(n9619), .C2(n10959), .A(n10958), .B(n10957), .ZN(
        n10965) );
  AOI22_X1 U13922 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11032), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10963) );
  AOI22_X1 U13923 ( .A1(n11011), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10962) );
  AOI22_X1 U13924 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U13925 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10960) );
  NAND4_X1 U13926 ( .A1(n10963), .A2(n10962), .A3(n10961), .A4(n10960), .ZN(
        n10964) );
  NOR2_X1 U13927 ( .A1(n10965), .A2(n10964), .ZN(n10974) );
  NAND2_X1 U13928 ( .A1(n10967), .A2(n10966), .ZN(n10973) );
  XNOR2_X1 U13929 ( .A(n10974), .B(n10973), .ZN(n10970) );
  AOI21_X1 U13930 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20613), .A(
        n11020), .ZN(n10969) );
  NAND2_X1 U13931 ( .A1(n10457), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n10968) );
  OAI211_X1 U13932 ( .C1(n10970), .C2(n11023), .A(n10969), .B(n10968), .ZN(
        n10971) );
  OAI21_X1 U13933 ( .B1(n11055), .B2(n14406), .A(n10971), .ZN(n14121) );
  INV_X1 U13934 ( .A(n10993), .ZN(n10972) );
  XOR2_X1 U13935 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B(n10972), .Z(
        n14399) );
  INV_X1 U13936 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14395) );
  AOI21_X1 U13937 ( .B1(n14395), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10991) );
  NOR2_X1 U13938 ( .A1(n10974), .A2(n10973), .ZN(n11019) );
  INV_X1 U13939 ( .A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10976) );
  OAI22_X1 U13940 ( .A1(n10308), .A2(n10976), .B1(n11039), .B2(n10975), .ZN(
        n10980) );
  OAI22_X1 U13941 ( .A1(n10978), .A2(n10977), .B1(n10126), .B2(n10089), .ZN(
        n10979) );
  AOI211_X1 U13942 ( .C1(n9623), .C2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n10980), .B(n10979), .ZN(n10988) );
  AOI22_X1 U13943 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10984) );
  AOI22_X1 U13944 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10902), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10983) );
  AOI22_X1 U13945 ( .A1(n11028), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10982) );
  AOI22_X1 U13946 ( .A1(n10198), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10981) );
  AND4_X1 U13947 ( .A1(n10984), .A2(n10983), .A3(n10982), .A4(n10981), .ZN(
        n10987) );
  AOI22_X1 U13948 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10986) );
  NAND2_X1 U13949 ( .A1(n10585), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10985) );
  NAND4_X1 U13950 ( .A1(n10988), .A2(n10987), .A3(n10986), .A4(n10985), .ZN(
        n11018) );
  XNOR2_X1 U13951 ( .A(n11019), .B(n11018), .ZN(n10989) );
  NOR2_X1 U13952 ( .A1(n10989), .A2(n11023), .ZN(n10990) );
  AOI211_X1 U13953 ( .C1(n11057), .C2(P1_EAX_REG_28__SCAN_IN), .A(n10991), .B(
        n10990), .ZN(n10992) );
  INV_X1 U13954 ( .A(n10994), .ZN(n10996) );
  INV_X1 U13955 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10995) );
  NAND2_X1 U13956 ( .A1(n10996), .A2(n10995), .ZN(n10997) );
  NAND2_X1 U13957 ( .A1(n13621), .A2(n10997), .ZN(n14384) );
  INV_X1 U13958 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10998) );
  OAI22_X1 U13959 ( .A1(n10999), .A2(n10998), .B1(n11039), .B2(n10113), .ZN(
        n11002) );
  INV_X1 U13960 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11000) );
  NOR2_X1 U13961 ( .A1(n9587), .A2(n11000), .ZN(n11001) );
  AOI211_X1 U13962 ( .C1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .C2(n11044), .A(
        n11002), .B(n11001), .ZN(n11006) );
  AOI22_X1 U13963 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U13964 ( .A1(n9586), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11003), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11004) );
  NAND3_X1 U13965 ( .A1(n11006), .A2(n11005), .A3(n11004), .ZN(n11017) );
  AOI22_X1 U13966 ( .A1(n10154), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11007) );
  OAI21_X1 U13967 ( .B1(n11009), .B2(n11008), .A(n11007), .ZN(n11010) );
  AOI21_X1 U13968 ( .B1(n10585), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n11010), .ZN(n11015) );
  AOI22_X1 U13969 ( .A1(n10198), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11014) );
  AOI22_X1 U13970 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11013) );
  NAND3_X1 U13971 ( .A1(n11015), .A2(n11014), .A3(n11013), .ZN(n11016) );
  NOR2_X1 U13972 ( .A1(n11017), .A2(n11016), .ZN(n11027) );
  NAND2_X1 U13973 ( .A1(n11019), .A2(n11018), .ZN(n11026) );
  XNOR2_X1 U13974 ( .A(n11027), .B(n11026), .ZN(n11024) );
  AOI21_X1 U13975 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20613), .A(
        n11020), .ZN(n11022) );
  NAND2_X1 U13976 ( .A1(n10457), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n11021) );
  OAI211_X1 U13977 ( .C1(n11024), .C2(n11023), .A(n11022), .B(n11021), .ZN(
        n11025) );
  OAI21_X1 U13978 ( .B1(n11055), .B2(n14384), .A(n11025), .ZN(n12413) );
  NOR2_X1 U13979 ( .A1(n11027), .A2(n11026), .ZN(n11051) );
  AOI22_X1 U13980 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11028), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11029) );
  OAI21_X1 U13981 ( .B1(n10833), .B2(n11030), .A(n11029), .ZN(n11031) );
  AOI21_X1 U13982 ( .B1(n9623), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A(n11031), .ZN(n11037) );
  AOI22_X1 U13983 ( .A1(n11032), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9586), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11036) );
  AOI22_X1 U13984 ( .A1(n11034), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11033), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11035) );
  NAND3_X1 U13985 ( .A1(n11037), .A2(n11036), .A3(n11035), .ZN(n11049) );
  OAI22_X1 U13986 ( .A1(n10308), .A2(n11040), .B1(n11039), .B2(n11038), .ZN(
        n11043) );
  NOR2_X1 U13987 ( .A1(n9619), .A2(n11041), .ZN(n11042) );
  AOI211_X1 U13988 ( .C1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .C2(n11012), .A(
        n11043), .B(n11042), .ZN(n11047) );
  AOI22_X1 U13989 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11011), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11046) );
  AOI22_X1 U13990 ( .A1(n11044), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10392), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11045) );
  NAND3_X1 U13991 ( .A1(n11047), .A2(n11046), .A3(n11045), .ZN(n11048) );
  NOR2_X1 U13992 ( .A1(n11049), .A2(n11048), .ZN(n11050) );
  XNOR2_X1 U13993 ( .A(n11051), .B(n11050), .ZN(n11053) );
  NAND2_X1 U13994 ( .A1(n11053), .A2(n11052), .ZN(n11060) );
  NAND2_X1 U13995 ( .A1(n20613), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11054) );
  NAND2_X1 U13996 ( .A1(n11055), .A2(n11054), .ZN(n11056) );
  AOI21_X1 U13997 ( .B1(n11057), .B2(P1_EAX_REG_30__SCAN_IN), .A(n11056), .ZN(
        n11059) );
  XNOR2_X1 U13998 ( .A(n13621), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14081) );
  NAND3_X1 U13999 ( .A1(n10259), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16003) );
  INV_X1 U14000 ( .A(n16003), .ZN(n11061) );
  AND3_X1 U14001 ( .A1(n11064), .A2(n11063), .A3(n11128), .ZN(n11065) );
  NOR2_X1 U14002 ( .A1(n9582), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11159) );
  INV_X1 U14003 ( .A(n11066), .ZN(n11091) );
  NAND2_X1 U14004 ( .A1(n11076), .A2(n11075), .ZN(n11090) );
  XNOR2_X1 U14005 ( .A(n11091), .B(n11090), .ZN(n11068) );
  NAND2_X1 U14006 ( .A1(n10223), .A2(n20122), .ZN(n11072) );
  INV_X1 U14007 ( .A(n11072), .ZN(n11067) );
  AOI21_X1 U14008 ( .B1(n11068), .B2(n13252), .A(n11067), .ZN(n11069) );
  OAI21_X1 U14009 ( .B1(n13478), .B2(n9982), .A(n11069), .ZN(n13468) );
  INV_X1 U14010 ( .A(n11075), .ZN(n11071) );
  NAND2_X1 U14011 ( .A1(n13252), .A2(n11071), .ZN(n11073) );
  AND2_X1 U14012 ( .A1(n11073), .A2(n11072), .ZN(n11074) );
  INV_X1 U14013 ( .A(n13252), .ZN(n20771) );
  XNOR2_X1 U14014 ( .A(n11076), .B(n11075), .ZN(n11081) );
  NAND2_X1 U14015 ( .A1(n11077), .A2(n10222), .ZN(n11080) );
  NOR2_X1 U14016 ( .A1(n10221), .A2(n11078), .ZN(n11079) );
  OAI211_X1 U14017 ( .C1(n20771), .C2(n11081), .A(n11080), .B(n11079), .ZN(
        n11083) );
  INV_X1 U14018 ( .A(n11082), .ZN(n11084) );
  NAND2_X1 U14019 ( .A1(n11084), .A2(n11083), .ZN(n11085) );
  INV_X1 U14020 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20071) );
  NAND2_X1 U14021 ( .A1(n11086), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11087) );
  INV_X1 U14022 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20054) );
  NAND2_X1 U14023 ( .A1(n11089), .A2(n11063), .ZN(n11095) );
  NAND2_X1 U14024 ( .A1(n11091), .A2(n11090), .ZN(n11109) );
  INV_X1 U14025 ( .A(n11107), .ZN(n11092) );
  XNOR2_X1 U14026 ( .A(n11109), .B(n11092), .ZN(n11093) );
  NAND2_X1 U14027 ( .A1(n11093), .A2(n13252), .ZN(n11094) );
  NAND2_X1 U14028 ( .A1(n11095), .A2(n11094), .ZN(n13524) );
  NAND2_X1 U14029 ( .A1(n11096), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11097) );
  NAND2_X1 U14030 ( .A1(n13527), .A2(n11097), .ZN(n20028) );
  NAND2_X1 U14031 ( .A1(n11098), .A2(n11063), .ZN(n11102) );
  NAND2_X1 U14032 ( .A1(n11109), .A2(n11107), .ZN(n11099) );
  XNOR2_X1 U14033 ( .A(n11099), .B(n11106), .ZN(n11100) );
  NAND2_X1 U14034 ( .A1(n11100), .A2(n13252), .ZN(n11101) );
  NAND2_X1 U14035 ( .A1(n11102), .A2(n11101), .ZN(n11103) );
  INV_X1 U14036 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20045) );
  XNOR2_X1 U14037 ( .A(n11103), .B(n20045), .ZN(n20027) );
  NAND2_X1 U14038 ( .A1(n11103), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11104) );
  NAND2_X1 U14039 ( .A1(n11105), .A2(n11063), .ZN(n11112) );
  AND2_X1 U14040 ( .A1(n11107), .A2(n11106), .ZN(n11108) );
  NAND2_X1 U14041 ( .A1(n11109), .A2(n11108), .ZN(n11115) );
  XNOR2_X1 U14042 ( .A(n11115), .B(n11116), .ZN(n11110) );
  NAND2_X1 U14043 ( .A1(n11110), .A2(n13252), .ZN(n11111) );
  INV_X1 U14044 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13725) );
  XNOR2_X1 U14045 ( .A(n11113), .B(n13725), .ZN(n15911) );
  NAND3_X1 U14046 ( .A1(n11062), .A2(n11063), .A3(n11114), .ZN(n11120) );
  INV_X1 U14047 ( .A(n11115), .ZN(n11117) );
  NAND2_X1 U14048 ( .A1(n11117), .A2(n11116), .ZN(n11125) );
  XNOR2_X1 U14049 ( .A(n11125), .B(n11126), .ZN(n11118) );
  NAND2_X1 U14050 ( .A1(n11118), .A2(n13252), .ZN(n11119) );
  NAND2_X1 U14051 ( .A1(n11120), .A2(n11119), .ZN(n13719) );
  OR2_X1 U14052 ( .A1(n13719), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11121) );
  NAND2_X1 U14053 ( .A1(n13719), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11122) );
  NAND2_X1 U14054 ( .A1(n9590), .A2(n11122), .ZN(n15901) );
  NAND2_X1 U14055 ( .A1(n11124), .A2(n11063), .ZN(n11131) );
  INV_X1 U14056 ( .A(n11125), .ZN(n11127) );
  NAND2_X1 U14057 ( .A1(n11127), .A2(n11126), .ZN(n11134) );
  XNOR2_X1 U14058 ( .A(n11134), .B(n11128), .ZN(n11129) );
  NAND2_X1 U14059 ( .A1(n11129), .A2(n13252), .ZN(n11130) );
  NAND2_X1 U14060 ( .A1(n11131), .A2(n11130), .ZN(n11132) );
  OR2_X1 U14061 ( .A1(n11132), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15903) );
  NAND2_X1 U14062 ( .A1(n11132), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15902) );
  OR3_X1 U14063 ( .A1(n11134), .A2(n11133), .A3(n20771), .ZN(n11135) );
  NAND2_X1 U14064 ( .A1(n9582), .A2(n11135), .ZN(n13750) );
  OR2_X1 U14065 ( .A1(n13750), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11136) );
  NAND2_X1 U14066 ( .A1(n13750), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11137) );
  INV_X1 U14067 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15980) );
  NAND2_X1 U14068 ( .A1(n9582), .A2(n15980), .ZN(n11139) );
  INV_X1 U14069 ( .A(n14474), .ZN(n11144) );
  INV_X1 U14070 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14540) );
  NAND2_X1 U14071 ( .A1(n9581), .A2(n14540), .ZN(n11140) );
  NAND2_X1 U14072 ( .A1(n14492), .A2(n11140), .ZN(n14507) );
  INV_X1 U14073 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15956) );
  AND2_X1 U14074 ( .A1(n9581), .A2(n15956), .ZN(n14505) );
  NOR2_X1 U14075 ( .A1(n14507), .A2(n14505), .ZN(n14491) );
  INV_X1 U14076 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14673) );
  NAND2_X1 U14077 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14489) );
  OAI21_X1 U14078 ( .B1(n14673), .B2(n14489), .A(n9581), .ZN(n11141) );
  NAND2_X1 U14079 ( .A1(n14491), .A2(n11141), .ZN(n14475) );
  OR2_X1 U14080 ( .A1(n9581), .A2(n14673), .ZN(n11142) );
  NAND2_X1 U14081 ( .A1(n14492), .A2(n11142), .ZN(n11149) );
  INV_X1 U14082 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11145) );
  NOR2_X1 U14083 ( .A1(n9581), .A2(n11145), .ZN(n14479) );
  NOR2_X1 U14084 ( .A1(n11149), .A2(n14479), .ZN(n15864) );
  XNOR2_X1 U14085 ( .A(n9582), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14482) );
  NAND2_X1 U14086 ( .A1(n9582), .A2(n11145), .ZN(n14480) );
  NAND2_X1 U14087 ( .A1(n14482), .A2(n14480), .ZN(n11143) );
  AOI21_X1 U14088 ( .B1(n14475), .B2(n15864), .A(n11143), .ZN(n15865) );
  INV_X1 U14089 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15863) );
  INV_X1 U14090 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11146) );
  AND3_X1 U14091 ( .A1(n15863), .A2(n11146), .A3(n11145), .ZN(n11147) );
  NAND2_X1 U14092 ( .A1(n14474), .A2(n11147), .ZN(n11148) );
  INV_X1 U14093 ( .A(n11149), .ZN(n11151) );
  NOR2_X1 U14094 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14502) );
  AND2_X1 U14095 ( .A1(n14502), .A2(n15956), .ZN(n11150) );
  OR2_X1 U14096 ( .A1(n9581), .A2(n11150), .ZN(n14488) );
  NAND2_X1 U14097 ( .A1(n11151), .A2(n14488), .ZN(n14476) );
  XNOR2_X1 U14098 ( .A(n9581), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14470) );
  NAND2_X1 U14099 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14645) );
  INV_X1 U14100 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14642) );
  NAND2_X1 U14101 ( .A1(n14447), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11155) );
  INV_X1 U14102 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15857) );
  INV_X1 U14103 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14660) );
  INV_X1 U14104 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14463) );
  NAND2_X1 U14105 ( .A1(n14642), .A2(n14463), .ZN(n11154) );
  OAI21_X2 U14106 ( .B1(n14454), .B2(n11154), .A(n15892), .ZN(n14448) );
  NAND2_X1 U14107 ( .A1(n11155), .A2(n14448), .ZN(n14388) );
  NAND3_X1 U14108 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14591) );
  NAND2_X1 U14109 ( .A1(n14388), .A2(n14591), .ZN(n11156) );
  NAND2_X1 U14110 ( .A1(n11155), .A2(n9581), .ZN(n14419) );
  INV_X1 U14111 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14611) );
  INV_X1 U14112 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11157) );
  INV_X1 U14113 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14610) );
  NAND3_X1 U14114 ( .A1(n14611), .A2(n11157), .A3(n14610), .ZN(n14390) );
  OAI21_X1 U14115 ( .B1(n14388), .B2(n14390), .A(n15892), .ZN(n14411) );
  NOR2_X1 U14116 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14572) );
  AND2_X1 U14117 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14571) );
  NAND2_X1 U14118 ( .A1(n9581), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11158) );
  AND2_X1 U14119 ( .A1(n11160), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11161) );
  NOR2_X1 U14120 ( .A1(n14373), .A2(n11161), .ZN(n14559) );
  NAND2_X1 U14121 ( .A1(n20536), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11172) );
  NAND2_X1 U14122 ( .A1(n9875), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11162) );
  NAND2_X1 U14123 ( .A1(n11172), .A2(n11162), .ZN(n11164) );
  OAI21_X1 U14124 ( .B1(n11171), .B2(n11164), .A(n11211), .ZN(n11167) );
  NAND2_X1 U14125 ( .A1(n11078), .A2(n10224), .ZN(n11163) );
  NAND2_X1 U14126 ( .A1(n11163), .A2(n9616), .ZN(n11183) );
  INV_X1 U14127 ( .A(n11164), .ZN(n11165) );
  OAI211_X1 U14128 ( .C1(n10218), .C2(n10223), .A(n11183), .B(n11165), .ZN(
        n11166) );
  XNOR2_X1 U14129 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11173) );
  XNOR2_X1 U14130 ( .A(n11173), .B(n11172), .ZN(n12364) );
  NAND2_X1 U14131 ( .A1(n11078), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11170) );
  NAND2_X1 U14132 ( .A1(n11215), .A2(n10222), .ZN(n11168) );
  OAI211_X1 U14133 ( .C1(n11169), .C2(n12364), .A(n11170), .B(n11168), .ZN(
        n11178) );
  AND3_X1 U14134 ( .A1(n11171), .A2(n10222), .A3(n11170), .ZN(n11193) );
  OAI22_X1 U14135 ( .A1(n11179), .A2(n11178), .B1(n11193), .B2(n12364), .ZN(
        n11192) );
  INV_X1 U14136 ( .A(n11183), .ZN(n11177) );
  INV_X1 U14137 ( .A(n11172), .ZN(n11174) );
  NAND2_X1 U14138 ( .A1(n11174), .A2(n11173), .ZN(n11176) );
  NAND2_X1 U14139 ( .A1(n20505), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11175) );
  NAND2_X1 U14140 ( .A1(n11176), .A2(n11175), .ZN(n11186) );
  XNOR2_X1 U14141 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11185) );
  XNOR2_X1 U14142 ( .A(n11186), .B(n11185), .ZN(n12361) );
  INV_X1 U14143 ( .A(n12361), .ZN(n11182) );
  NAND3_X1 U14144 ( .A1(n11177), .A2(n11215), .A3(n11182), .ZN(n11181) );
  NAND2_X1 U14145 ( .A1(n11179), .A2(n11178), .ZN(n11180) );
  NAND2_X1 U14146 ( .A1(n11215), .A2(n11182), .ZN(n11184) );
  NAND2_X1 U14147 ( .A1(n11184), .A2(n11183), .ZN(n11189) );
  NAND2_X1 U14148 ( .A1(n11186), .A2(n11185), .ZN(n11188) );
  NAND2_X1 U14149 ( .A1(n20425), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11187) );
  NAND2_X1 U14150 ( .A1(n11188), .A2(n11187), .ZN(n11196) );
  XNOR2_X1 U14151 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11195) );
  XNOR2_X1 U14152 ( .A(n11196), .B(n11195), .ZN(n12360) );
  INV_X1 U14153 ( .A(n12360), .ZN(n11198) );
  AOI22_X1 U14154 ( .A1(n11189), .A2(n11198), .B1(n11200), .B2(n12361), .ZN(
        n11190) );
  AOI21_X1 U14155 ( .B1(n11192), .B2(n11191), .A(n11190), .ZN(n11202) );
  INV_X1 U14156 ( .A(n11193), .ZN(n11197) );
  NOR2_X1 U14157 ( .A1(n12996), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11194) );
  AND2_X1 U14158 ( .A1(n11205), .A2(n11208), .ZN(n12362) );
  INV_X1 U14159 ( .A(n12362), .ZN(n11199) );
  OAI22_X1 U14160 ( .A1(n11211), .A2(n11198), .B1(n11197), .B2(n11199), .ZN(
        n11201) );
  OAI22_X1 U14161 ( .A1(n11202), .A2(n11201), .B1(n11200), .B2(n11199), .ZN(
        n11204) );
  NAND2_X1 U14162 ( .A1(n10259), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11203) );
  NAND2_X1 U14163 ( .A1(n11204), .A2(n11203), .ZN(n11213) );
  INV_X1 U14164 ( .A(n11205), .ZN(n11207) );
  NOR2_X1 U14165 ( .A1(n13438), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11206) );
  INV_X1 U14166 ( .A(n11208), .ZN(n11209) );
  NAND2_X1 U14167 ( .A1(n11218), .A2(n13016), .ZN(n11220) );
  INV_X1 U14168 ( .A(n10221), .ZN(n11231) );
  NAND2_X1 U14169 ( .A1(n14692), .A2(n10223), .ZN(n11221) );
  NAND2_X1 U14170 ( .A1(n20622), .A2(n11227), .ZN(n20767) );
  NAND2_X1 U14171 ( .A1(n20767), .A2(n10259), .ZN(n11223) );
  NAND2_X1 U14172 ( .A1(n10259), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11225) );
  NAND2_X1 U14173 ( .A1(n20254), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11224) );
  AND2_X1 U14174 ( .A1(n11225), .A2(n11224), .ZN(n13097) );
  INV_X1 U14175 ( .A(n13097), .ZN(n11226) );
  INV_X1 U14176 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13620) );
  INV_X2 U14177 ( .A(n20065), .ZN(n20024) );
  NAND2_X1 U14178 ( .A1(n20024), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14551) );
  OAI21_X1 U14179 ( .B1(n14484), .B2(n13620), .A(n14551), .ZN(n11228) );
  AOI21_X1 U14180 ( .B1(n14081), .B2(n15889), .A(n11228), .ZN(n11229) );
  OAI211_X1 U14181 ( .C1(n14086), .C2(n20090), .A(n11230), .B(n11229), .ZN(
        P1_U2969) );
  NAND2_X1 U14182 ( .A1(n11231), .A2(n13105), .ZN(n11232) );
  NAND2_X1 U14183 ( .A1(n13008), .A2(n13028), .ZN(n12926) );
  INV_X1 U14184 ( .A(n11233), .ZN(n11234) );
  INV_X1 U14185 ( .A(n10229), .ZN(n14069) );
  AND3_X1 U14186 ( .A1(n13016), .A2(n14069), .A3(n10209), .ZN(n12368) );
  NAND3_X1 U14187 ( .A1(n11234), .A2(n13105), .A3(n12368), .ZN(n11235) );
  NAND2_X1 U14188 ( .A1(n12926), .A2(n11235), .ZN(n11236) );
  NAND2_X1 U14189 ( .A1(n11312), .A2(n20086), .ZN(n11237) );
  OAI211_X1 U14190 ( .C1(n14089), .C2(P1_EBX_REG_1__SCAN_IN), .A(n14087), .B(
        n11237), .ZN(n11238) );
  NAND2_X1 U14191 ( .A1(n11239), .A2(n11238), .ZN(n11241) );
  NAND2_X1 U14192 ( .A1(n11312), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11240) );
  OAI21_X1 U14193 ( .B1(n11320), .B2(P1_EBX_REG_0__SCAN_IN), .A(n11240), .ZN(
        n13022) );
  XNOR2_X1 U14194 ( .A(n11241), .B(n13022), .ZN(n13106) );
  NAND2_X1 U14195 ( .A1(n13106), .A2(n13105), .ZN(n13107) );
  INV_X1 U14196 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n11242) );
  NAND2_X1 U14197 ( .A1(n11312), .A2(n20071), .ZN(n11243) );
  OAI211_X1 U14198 ( .C1(n14089), .C2(P1_EBX_REG_2__SCAN_IN), .A(n14087), .B(
        n11243), .ZN(n11244) );
  AND2_X1 U14199 ( .A1(n11245), .A2(n11244), .ZN(n13473) );
  MUX2_X1 U14200 ( .A(n11310), .B(n14087), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n11249) );
  OAI21_X1 U14201 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14090), .A(
        n11249), .ZN(n13457) );
  MUX2_X1 U14202 ( .A(n11317), .B(n11312), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n11253) );
  INV_X1 U14203 ( .A(n11312), .ZN(n11250) );
  NAND2_X1 U14204 ( .A1(n11250), .A2(n14089), .ZN(n11290) );
  NAND2_X1 U14205 ( .A1(n14089), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11251) );
  AND2_X1 U14206 ( .A1(n11290), .A2(n11251), .ZN(n11252) );
  NAND2_X1 U14207 ( .A1(n11253), .A2(n11252), .ZN(n13542) );
  MUX2_X1 U14208 ( .A(n11310), .B(n14087), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n11254) );
  OAI21_X1 U14209 ( .B1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n14090), .A(
        n11254), .ZN(n13540) );
  MUX2_X1 U14210 ( .A(n11317), .B(n11312), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n11258) );
  NAND2_X1 U14211 ( .A1(n14089), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11256) );
  AND2_X1 U14212 ( .A1(n11290), .A2(n11256), .ZN(n11257) );
  AND2_X1 U14213 ( .A1(n11258), .A2(n11257), .ZN(n13557) );
  INV_X1 U14214 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19937) );
  NAND2_X1 U14215 ( .A1(n11299), .A2(n19937), .ZN(n11261) );
  INV_X1 U14216 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15993) );
  NAND2_X1 U14217 ( .A1(n13105), .A2(n19937), .ZN(n11259) );
  OAI211_X1 U14218 ( .C1(n11320), .C2(n15993), .A(n11259), .B(n11312), .ZN(
        n11260) );
  MUX2_X1 U14219 ( .A(n11317), .B(n11312), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n11264) );
  NAND2_X1 U14220 ( .A1(n14089), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11262) );
  AND2_X1 U14221 ( .A1(n11290), .A2(n11262), .ZN(n11263) );
  NAND2_X1 U14222 ( .A1(n11264), .A2(n11263), .ZN(n13687) );
  NAND2_X1 U14223 ( .A1(n13688), .A2(n13687), .ZN(n15970) );
  INV_X1 U14224 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20002) );
  NAND2_X1 U14225 ( .A1(n11299), .A2(n20002), .ZN(n11267) );
  NAND2_X1 U14226 ( .A1(n13105), .A2(n20002), .ZN(n11265) );
  OAI211_X1 U14227 ( .C1(n11320), .C2(n15980), .A(n11265), .B(n11312), .ZN(
        n11266) );
  NAND2_X1 U14228 ( .A1(n11267), .A2(n11266), .ZN(n15969) );
  INV_X1 U14229 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15845) );
  INV_X1 U14230 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11269) );
  NAND2_X1 U14231 ( .A1(n11312), .A2(n11269), .ZN(n11270) );
  OAI211_X1 U14232 ( .C1(n14089), .C2(P1_EBX_REG_10__SCAN_IN), .A(n14087), .B(
        n11270), .ZN(n11271) );
  AND2_X1 U14233 ( .A1(n11272), .A2(n11271), .ZN(n13740) );
  MUX2_X1 U14234 ( .A(n11299), .B(n11320), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n11274) );
  NOR2_X1 U14235 ( .A1(n14090), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11273) );
  NOR2_X1 U14236 ( .A1(n11274), .A2(n11273), .ZN(n14291) );
  MUX2_X1 U14237 ( .A(n11317), .B(n11312), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n11277) );
  NAND2_X1 U14238 ( .A1(n14089), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11275) );
  AND2_X1 U14239 ( .A1(n11290), .A2(n11275), .ZN(n11276) );
  NAND2_X1 U14240 ( .A1(n11277), .A2(n11276), .ZN(n13767) );
  INV_X1 U14241 ( .A(n13767), .ZN(n14207) );
  MUX2_X1 U14242 ( .A(n11310), .B(n14087), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n11278) );
  OAI21_X1 U14243 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14090), .A(
        n11278), .ZN(n14206) );
  INV_X1 U14244 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n13779) );
  NAND2_X1 U14245 ( .A1(n11312), .A2(n14673), .ZN(n11279) );
  OAI211_X1 U14246 ( .C1(n14089), .C2(P1_EBX_REG_14__SCAN_IN), .A(n14087), .B(
        n11279), .ZN(n11280) );
  MUX2_X1 U14247 ( .A(n11299), .B(n11320), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11283) );
  NOR2_X1 U14248 ( .A1(n14090), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11282) );
  NOR2_X1 U14249 ( .A1(n11283), .A2(n11282), .ZN(n14281) );
  NAND2_X1 U14250 ( .A1(n11312), .A2(n15863), .ZN(n11284) );
  OAI211_X1 U14251 ( .C1(n14089), .C2(P1_EBX_REG_16__SCAN_IN), .A(n14087), .B(
        n11284), .ZN(n11285) );
  OAI21_X1 U14252 ( .B1(n11317), .B2(P1_EBX_REG_16__SCAN_IN), .A(n11285), .ZN(
        n14276) );
  NAND2_X1 U14253 ( .A1(n14284), .A2(n14276), .ZN(n14195) );
  MUX2_X1 U14254 ( .A(n11310), .B(n14087), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n11288) );
  INV_X1 U14255 ( .A(n14090), .ZN(n11286) );
  NAND2_X1 U14256 ( .A1(n11286), .A2(n11146), .ZN(n11287) );
  NAND2_X1 U14257 ( .A1(n11288), .A2(n11287), .ZN(n14196) );
  MUX2_X1 U14258 ( .A(n11317), .B(n11312), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n11292) );
  NAND2_X1 U14259 ( .A1(n14089), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11289) );
  AND2_X1 U14260 ( .A1(n11290), .A2(n11289), .ZN(n11291) );
  NAND2_X1 U14261 ( .A1(n11292), .A2(n11291), .ZN(n14271) );
  INV_X1 U14262 ( .A(n14271), .ZN(n11293) );
  MUX2_X1 U14263 ( .A(n11299), .B(n11320), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n11295) );
  NOR2_X1 U14264 ( .A1(n14090), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11294) );
  NOR2_X1 U14265 ( .A1(n11295), .A2(n11294), .ZN(n14262) );
  MUX2_X1 U14266 ( .A(n11317), .B(n11312), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n11297) );
  NAND2_X1 U14267 ( .A1(n14089), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11296) );
  NAND2_X1 U14268 ( .A1(n11297), .A2(n11296), .ZN(n14256) );
  MUX2_X1 U14269 ( .A(n11310), .B(n14087), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n11298) );
  OAI21_X1 U14270 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n14090), .A(
        n11298), .ZN(n14252) );
  MUX2_X1 U14271 ( .A(n11299), .B(n11320), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n11301) );
  NOR2_X1 U14272 ( .A1(n14090), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11300) );
  NOR2_X1 U14273 ( .A1(n11301), .A2(n11300), .ZN(n14171) );
  MUX2_X1 U14274 ( .A(n11317), .B(n11312), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n11303) );
  NAND2_X1 U14275 ( .A1(n14089), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11302) );
  NAND2_X1 U14276 ( .A1(n11303), .A2(n11302), .ZN(n14184) );
  NAND2_X1 U14277 ( .A1(n11312), .A2(n14610), .ZN(n11304) );
  OAI211_X1 U14278 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n14089), .A(n14087), .B(
        n11304), .ZN(n11305) );
  OAI21_X1 U14279 ( .B1(n11317), .B2(P1_EBX_REG_24__SCAN_IN), .A(n11305), .ZN(
        n14158) );
  NAND2_X1 U14280 ( .A1(n14173), .A2(n14158), .ZN(n14157) );
  MUX2_X1 U14281 ( .A(n11310), .B(n14087), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n11306) );
  OAI21_X1 U14282 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14090), .A(
        n11306), .ZN(n14145) );
  INV_X1 U14283 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14243) );
  INV_X1 U14284 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14542) );
  NAND2_X1 U14285 ( .A1(n11312), .A2(n14542), .ZN(n11307) );
  OAI211_X1 U14286 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n14089), .A(n14087), .B(
        n11307), .ZN(n11308) );
  AND2_X1 U14287 ( .A1(n11309), .A2(n11308), .ZN(n14139) );
  MUX2_X1 U14288 ( .A(n11310), .B(n14087), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n11311) );
  OAI21_X1 U14289 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14090), .A(
        n11311), .ZN(n14128) );
  MUX2_X1 U14290 ( .A(n11317), .B(n11312), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n11314) );
  NAND2_X1 U14291 ( .A1(n14089), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11313) );
  NAND2_X1 U14292 ( .A1(n11314), .A2(n11313), .ZN(n14110) );
  OR2_X1 U14293 ( .A1(n14090), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11316) );
  INV_X1 U14294 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n12416) );
  NAND2_X1 U14295 ( .A1(n13105), .A2(n12416), .ZN(n11315) );
  NAND2_X1 U14296 ( .A1(n11316), .A2(n11315), .ZN(n11318) );
  OAI22_X1 U14297 ( .A1(n11318), .A2(n11320), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n11317), .ZN(n12414) );
  INV_X1 U14298 ( .A(n11318), .ZN(n11319) );
  AOI22_X1 U14299 ( .A1(n9660), .A2(n11320), .B1(n11319), .B2(n14111), .ZN(
        n11321) );
  AOI22_X1 U14300 ( .A1(n14090), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14089), .ZN(n14088) );
  INV_X1 U14301 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n11322) );
  OR2_X1 U14302 ( .A1(n20003), .A2(n11322), .ZN(n11323) );
  INV_X1 U14303 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13947) );
  AND2_X4 U14304 ( .A1(n13348), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11528) );
  AOI22_X1 U14305 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14306 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11408), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11328) );
  INV_X2 U14307 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13349) );
  AND3_X4 U14308 ( .A1(n13349), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U14309 ( .A1(n11349), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11327) );
  NAND3_X1 U14310 ( .A1(n11329), .A2(n11328), .A3(n11327), .ZN(n11336) );
  AOI22_X1 U14311 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14312 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11330) );
  AND3_X1 U14313 ( .A1(n11331), .A2(n11330), .A3(n13115), .ZN(n11334) );
  AOI22_X1 U14314 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11408), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14315 ( .A1(n11349), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11332) );
  NAND3_X1 U14316 ( .A1(n11334), .A2(n11333), .A3(n11332), .ZN(n11335) );
  INV_X2 U14317 ( .A(n11423), .ZN(n12040) );
  AOI22_X1 U14318 ( .A1(n11349), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U14319 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U14320 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11338) );
  AOI22_X1 U14321 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11337) );
  NAND4_X1 U14322 ( .A1(n11340), .A2(n11339), .A3(n11338), .A4(n11337), .ZN(
        n11341) );
  NAND2_X1 U14323 ( .A1(n11341), .A2(n11530), .ZN(n11348) );
  AOI22_X1 U14324 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U14325 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11344) );
  AOI22_X1 U14326 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14327 ( .A1(n11349), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11342) );
  NAND4_X1 U14328 ( .A1(n11345), .A2(n11344), .A3(n11343), .A4(n11342), .ZN(
        n11346) );
  NAND2_X1 U14329 ( .A1(n11346), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11347) );
  AOI22_X1 U14330 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9605), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14331 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11523), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14332 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11351) );
  AOI22_X1 U14333 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n11349), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11350) );
  NAND4_X1 U14334 ( .A1(n11353), .A2(n11352), .A3(n11351), .A4(n11350), .ZN(
        n11354) );
  AOI22_X1 U14335 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14336 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11523), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14337 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U14338 ( .A1(n11349), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11355) );
  NAND4_X1 U14339 ( .A1(n11358), .A2(n11357), .A3(n11356), .A4(n11355), .ZN(
        n11359) );
  NAND3_X1 U14340 ( .A1(n12040), .A2(n12798), .A3(n13675), .ZN(n11381) );
  AOI22_X1 U14341 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11408), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14342 ( .A1(n11349), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14343 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11361) );
  AOI22_X1 U14344 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11360) );
  AOI22_X1 U14345 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11408), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U14346 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11366) );
  AOI22_X1 U14347 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11523), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11365) );
  AOI22_X1 U14348 ( .A1(n11349), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U14349 ( .A1(n11349), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11370) );
  AOI22_X1 U14350 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U14351 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11368) );
  NAND4_X1 U14352 ( .A1(n11371), .A2(n11370), .A3(n11369), .A4(n11368), .ZN(
        n11372) );
  AOI22_X1 U14353 ( .A1(n11349), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14354 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11523), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11373) );
  NAND4_X1 U14355 ( .A1(n11376), .A2(n11375), .A3(n11374), .A4(n11373), .ZN(
        n11377) );
  AOI22_X1 U14356 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11385) );
  AOI22_X1 U14357 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9605), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U14358 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14359 ( .A1(n11349), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11382) );
  NAND4_X1 U14360 ( .A1(n11385), .A2(n11384), .A3(n11383), .A4(n11382), .ZN(
        n11386) );
  AOI22_X1 U14361 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11390) );
  AOI22_X1 U14362 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14363 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11523), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11388) );
  AOI22_X1 U14364 ( .A1(n11349), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11387) );
  NAND4_X1 U14365 ( .A1(n11390), .A2(n11389), .A3(n11388), .A4(n11387), .ZN(
        n11391) );
  AOI22_X1 U14366 ( .A1(n11349), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14367 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14368 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14369 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11394) );
  AOI22_X1 U14370 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14371 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9605), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14372 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11523), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U14373 ( .A1(n11349), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11398) );
  NAND2_X2 U14374 ( .A1(n11895), .A2(n11420), .ZN(n11900) );
  AND3_X2 U14375 ( .A1(n11403), .A2(n12038), .A3(n11402), .ZN(n12030) );
  AOI22_X1 U14376 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U14377 ( .A1(n11349), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11406) );
  AOI22_X1 U14378 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9605), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14379 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11523), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11404) );
  AOI22_X1 U14380 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11528), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14381 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9605), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11411) );
  AOI22_X1 U14382 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11523), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11410) );
  AND2_X2 U14383 ( .A1(n19131), .A2(n11916), .ZN(n12805) );
  NAND2_X1 U14384 ( .A1(n11429), .A2(n11415), .ZN(n11920) );
  INV_X1 U14385 ( .A(n11900), .ZN(n12806) );
  NAND4_X1 U14386 ( .A1(n12806), .A2(n12805), .A3(n11440), .A4(n13679), .ZN(
        n11416) );
  NOR2_X1 U14387 ( .A1(n11737), .A2(n11927), .ZN(n11417) );
  INV_X2 U14388 ( .A(n11521), .ZN(n19119) );
  NAND2_X1 U14389 ( .A1(n13389), .A2(n14757), .ZN(n11419) );
  NAND2_X1 U14390 ( .A1(n9612), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U14391 ( .A1(n11999), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11425) );
  AND2_X1 U14392 ( .A1(n11916), .A2(n12035), .ZN(n11428) );
  INV_X1 U14393 ( .A(n13389), .ZN(n11431) );
  NAND3_X1 U14394 ( .A1(n12069), .A2(n11431), .A3(n11446), .ZN(n11439) );
  NAND3_X1 U14395 ( .A1(n11916), .A2(n13139), .A3(n11737), .ZN(n11434) );
  NAND2_X1 U14396 ( .A1(n11442), .A2(n12035), .ZN(n11436) );
  NAND3_X1 U14397 ( .A1(n11437), .A2(n10019), .A3(n11436), .ZN(n12044) );
  NAND2_X1 U14398 ( .A1(n11442), .A2(n19119), .ZN(n12037) );
  NOR2_X1 U14399 ( .A1(n13368), .A2(n18737), .ZN(n19884) );
  NAND2_X1 U14400 ( .A1(n11442), .A2(n12040), .ZN(n11921) );
  NAND2_X1 U14401 ( .A1(n11440), .A2(n13139), .ZN(n11441) );
  NAND2_X1 U14402 ( .A1(n11442), .A2(n11441), .ZN(n11913) );
  NAND2_X1 U14403 ( .A1(n11913), .A2(n11423), .ZN(n11919) );
  NAND2_X1 U14404 ( .A1(n11443), .A2(n11919), .ZN(n12033) );
  NAND2_X1 U14405 ( .A1(n12033), .A2(n12035), .ZN(n11445) );
  NAND2_X1 U14406 ( .A1(n11445), .A2(n11444), .ZN(n11456) );
  NAND2_X1 U14407 ( .A1(n11456), .A2(n11446), .ZN(n11447) );
  NAND2_X1 U14408 ( .A1(n11467), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11451) );
  NAND2_X1 U14409 ( .A1(n13389), .A2(n13368), .ZN(n12748) );
  NOR2_X1 U14410 ( .A1(n13390), .A2(n19857), .ZN(n11449) );
  AOI21_X1 U14411 ( .B1(n13350), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11449), 
        .ZN(n11450) );
  NAND2_X1 U14412 ( .A1(n9611), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11454) );
  NAND2_X1 U14413 ( .A1(n11999), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n11453) );
  NAND2_X1 U14414 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11452) );
  NAND3_X1 U14415 ( .A1(n11458), .A2(n11455), .A3(n11457), .ZN(n11483) );
  INV_X1 U14416 ( .A(n11459), .ZN(n11461) );
  INV_X1 U14417 ( .A(n13390), .ZN(n11460) );
  AOI22_X1 U14418 ( .A1(n11461), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n11460), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11462) );
  NAND2_X1 U14419 ( .A1(n11463), .A2(n11462), .ZN(n11484) );
  AOI22_X1 U14420 ( .A1(n11999), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11466) );
  NAND2_X1 U14421 ( .A1(n9613), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11465) );
  NAND2_X1 U14422 ( .A1(n11467), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11469) );
  AOI21_X1 U14423 ( .B1(n18737), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11468) );
  NAND2_X1 U14424 ( .A1(n11469), .A2(n11468), .ZN(n11471) );
  NAND2_X1 U14425 ( .A1(n11470), .A2(n11471), .ZN(n11474) );
  NOR2_X1 U14426 ( .A1(n13390), .A2(n19842), .ZN(n11476) );
  NAND2_X1 U14427 ( .A1(n15019), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11482) );
  INV_X1 U14428 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13493) );
  NAND2_X1 U14429 ( .A1(n12014), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11479) );
  NAND2_X1 U14430 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11478) );
  OAI211_X1 U14431 ( .C1(n13493), .C2(n9610), .A(n11479), .B(n11478), .ZN(
        n11480) );
  INV_X1 U14432 ( .A(n11480), .ZN(n11481) );
  BUF_X4 U14433 ( .A(n13077), .Z(n11505) );
  INV_X1 U14434 ( .A(n11484), .ZN(n11485) );
  NAND2_X1 U14435 ( .A1(n18945), .A2(n9600), .ZN(n11512) );
  INV_X1 U14436 ( .A(n11490), .ZN(n11491) );
  NAND2_X1 U14437 ( .A1(n11498), .A2(n11491), .ZN(n11492) );
  INV_X1 U14438 ( .A(n18945), .ZN(n13347) );
  NAND2_X1 U14439 ( .A1(n13355), .A2(n13347), .ZN(n11513) );
  INV_X1 U14440 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11493) );
  OAI22_X1 U14441 ( .A1(n13947), .A2(n19521), .B1(n19419), .B2(n11493), .ZN(
        n11494) );
  INV_X1 U14442 ( .A(n13077), .ZN(n11495) );
  NAND2_X1 U14443 ( .A1(n13057), .A2(n18929), .ZN(n11496) );
  NAND2_X1 U14444 ( .A1(n13057), .A2(n13355), .ZN(n11497) );
  NOR2_X2 U14445 ( .A1(n11518), .A2(n11497), .ZN(n19292) );
  AOI22_X1 U14446 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19360), .B1(
        n19292), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11500) );
  NOR2_X2 U14447 ( .A1(n11514), .A2(n9670), .ZN(n19639) );
  AOI22_X1 U14448 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19458), .B1(
        n19639), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11499) );
  INV_X1 U14449 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13939) );
  NAND2_X1 U14450 ( .A1(n13057), .A2(n11504), .ZN(n11501) );
  INV_X1 U14451 ( .A(n11512), .ZN(n11502) );
  NAND2_X1 U14452 ( .A1(n13057), .A2(n11502), .ZN(n11503) );
  INV_X1 U14453 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13941) );
  OAI22_X1 U14454 ( .A1(n13939), .A2(n19327), .B1(n19389), .B2(n13941), .ZN(
        n11508) );
  INV_X1 U14455 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13938) );
  INV_X1 U14456 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11506) );
  OAI22_X1 U14457 ( .A1(n13938), .A2(n19247), .B1(n11665), .B2(n11506), .ZN(
        n11507) );
  NOR2_X1 U14458 ( .A1(n11508), .A2(n11507), .ZN(n11509) );
  INV_X1 U14459 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13948) );
  INV_X1 U14460 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13949) );
  OAI22_X1 U14461 ( .A1(n13948), .A2(n19591), .B1(n19487), .B2(n13949), .ZN(
        n11517) );
  INV_X1 U14462 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13950) );
  OR2_X2 U14463 ( .A1(n11514), .A2(n11513), .ZN(n19564) );
  INV_X1 U14464 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11515) );
  OAI22_X1 U14465 ( .A1(n13950), .A2(n19684), .B1(n19564), .B2(n11515), .ZN(
        n11516) );
  AND2_X2 U14466 ( .A1(n11522), .A2(n11530), .ZN(n11564) );
  AOI22_X1 U14467 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11564), .B1(
        n11602), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14468 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14469 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11597), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11525) );
  AND2_X2 U14470 ( .A1(n11408), .A2(n13115), .ZN(n13113) );
  AOI22_X1 U14471 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n11611), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11524) );
  NAND4_X1 U14472 ( .A1(n11527), .A2(n11526), .A3(n11525), .A4(n11524), .ZN(
        n11538) );
  AND2_X2 U14473 ( .A1(n11409), .A2(n11530), .ZN(n12120) );
  INV_X1 U14474 ( .A(n9588), .ZN(n13850) );
  AOI22_X1 U14475 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12120), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14476 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n13828), .ZN(n11535) );
  AOI22_X1 U14477 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12170), .B1(
        n12169), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11534) );
  AND2_X2 U14478 ( .A1(n9588), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12139) );
  AOI22_X1 U14479 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11533) );
  NAND4_X1 U14480 ( .A1(n11536), .A2(n11535), .A3(n11534), .A4(n11533), .ZN(
        n11537) );
  INV_X1 U14481 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13895) );
  INV_X1 U14482 ( .A(n19639), .ZN(n19635) );
  INV_X1 U14483 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12142) );
  INV_X1 U14484 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13897) );
  INV_X1 U14485 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11540) );
  OAI22_X1 U14486 ( .A1(n13897), .A2(n19487), .B1(n19419), .B2(n11540), .ZN(
        n11541) );
  NOR2_X1 U14487 ( .A1(n11542), .A2(n11541), .ZN(n11559) );
  INV_X1 U14488 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13889) );
  INV_X1 U14489 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13886) );
  OAI22_X1 U14490 ( .A1(n13889), .A2(n19389), .B1(n19247), .B2(n13886), .ZN(
        n11543) );
  INV_X1 U14491 ( .A(n11543), .ZN(n11547) );
  NAND2_X1 U14492 ( .A1(n19292), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11546) );
  NAND2_X1 U14493 ( .A1(n19360), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11545) );
  NAND2_X1 U14494 ( .A1(n19458), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11544) );
  INV_X1 U14495 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20924) );
  INV_X1 U14496 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11548) );
  OAI21_X1 U14497 ( .B1(n11665), .B2(n11548), .A(n19890), .ZN(n11550) );
  INV_X1 U14498 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13887) );
  NOR2_X1 U14499 ( .A1(n19327), .A2(n13887), .ZN(n11549) );
  NOR2_X1 U14500 ( .A1(n11550), .A2(n11549), .ZN(n11552) );
  NAND2_X1 U14501 ( .A1(n19556), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11551) );
  OAI211_X1 U14502 ( .C1(n11553), .C2(n20924), .A(n11552), .B(n11551), .ZN(
        n11554) );
  INV_X1 U14503 ( .A(n11554), .ZN(n11557) );
  INV_X1 U14504 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13896) );
  OAI22_X1 U14505 ( .A1(n13896), .A2(n19591), .B1(n19684), .B2(n12141), .ZN(
        n11555) );
  AOI21_X1 U14506 ( .B1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n19211), .A(
        n11555), .ZN(n11556) );
  NAND4_X1 U14507 ( .A1(n11559), .A2(n11558), .A3(n11557), .A4(n11556), .ZN(
        n11594) );
  AOI22_X1 U14508 ( .A1(n12120), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13876), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U14509 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12169), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U14510 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14511 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11560) );
  NAND4_X1 U14512 ( .A1(n11563), .A2(n11562), .A3(n11561), .A4(n11560), .ZN(
        n11571) );
  AOI22_X1 U14513 ( .A1(n11564), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11597), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U14514 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U14515 ( .A1(n13113), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13828), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U14516 ( .A1(n13703), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11611), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11566) );
  NAND4_X1 U14517 ( .A1(n11569), .A2(n11568), .A3(n11567), .A4(n11566), .ZN(
        n11570) );
  NOR2_X1 U14518 ( .A1(n11571), .A2(n11570), .ZN(n12761) );
  AOI22_X1 U14519 ( .A1(n13113), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U14520 ( .A1(n12120), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n13828), .ZN(n11574) );
  AOI22_X1 U14521 ( .A1(n13703), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U14522 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11611), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11572) );
  NAND4_X1 U14523 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(
        n11581) );
  AOI22_X1 U14524 ( .A1(n11564), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11597), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14525 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11646), .B1(
        n12169), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14526 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14527 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13876), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11576) );
  NAND4_X1 U14528 ( .A1(n11579), .A2(n11578), .A3(n11577), .A4(n11576), .ZN(
        n11580) );
  NOR2_X1 U14529 ( .A1(n12761), .A2(n12271), .ZN(n11582) );
  NAND2_X1 U14530 ( .A1(n19119), .A2(n11582), .ZN(n12275) );
  AOI22_X1 U14531 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11564), .B1(
        n11602), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U14532 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11597), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U14533 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11646), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14534 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n11611), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11583) );
  NAND4_X1 U14535 ( .A1(n11586), .A2(n11585), .A3(n11584), .A4(n11583), .ZN(
        n11592) );
  AOI22_X1 U14536 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12120), .B1(
        n12139), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U14537 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n13828), .ZN(n11589) );
  AOI22_X1 U14538 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12170), .B1(
        n12169), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U14539 ( .A1(n13703), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11587) );
  NAND4_X1 U14540 ( .A1(n11590), .A2(n11589), .A3(n11588), .A4(n11587), .ZN(
        n11591) );
  NAND2_X1 U14541 ( .A1(n12275), .A2(n12274), .ZN(n11593) );
  AND2_X2 U14542 ( .A1(n11594), .A2(n11593), .ZN(n11596) );
  NAND2_X1 U14543 ( .A1(n11564), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11601) );
  NAND2_X1 U14544 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11600) );
  NAND2_X1 U14545 ( .A1(n12120), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11599) );
  NAND2_X1 U14546 ( .A1(n11597), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11598) );
  NAND2_X1 U14547 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11606) );
  NAND2_X1 U14548 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11605) );
  NAND2_X1 U14549 ( .A1(n13703), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11604) );
  NAND2_X1 U14550 ( .A1(n12170), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11603) );
  NAND2_X1 U14551 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11610) );
  NAND2_X1 U14552 ( .A1(n12169), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11609) );
  NAND2_X1 U14553 ( .A1(n12140), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11608) );
  NAND2_X1 U14554 ( .A1(n13828), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11607) );
  NAND2_X1 U14555 ( .A1(n12121), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11615) );
  NAND2_X1 U14556 ( .A1(n11611), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11614) );
  NAND2_X1 U14557 ( .A1(n13113), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11613) );
  NAND2_X1 U14558 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11612) );
  INV_X1 U14559 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11633) );
  INV_X1 U14560 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n12831) );
  NAND2_X1 U14561 ( .A1(n11633), .A2(n12831), .ZN(n11619) );
  MUX2_X1 U14562 ( .A(n12271), .B(n11619), .S(n12321), .Z(n11639) );
  NAND2_X1 U14563 ( .A1(n19857), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11621) );
  NAND2_X1 U14564 ( .A1(n13349), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11620) );
  NAND2_X1 U14565 ( .A1(n11621), .A2(n11620), .ZN(n11893) );
  NAND2_X1 U14566 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19865), .ZN(
        n11872) );
  NAND2_X1 U14567 ( .A1(n11622), .A2(n11621), .ZN(n11626) );
  NAND2_X1 U14568 ( .A1(n20880), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11627) );
  NAND2_X1 U14569 ( .A1(n9751), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11623) );
  XNOR2_X1 U14570 ( .A(n11626), .B(n11625), .ZN(n11901) );
  INV_X1 U14571 ( .A(n11901), .ZN(n11624) );
  NAND2_X1 U14572 ( .A1(n9602), .A2(n11624), .ZN(n11903) );
  INV_X1 U14573 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12908) );
  NAND2_X1 U14574 ( .A1(n11626), .A2(n11625), .ZN(n11628) );
  NAND2_X1 U14575 ( .A1(n11628), .A2(n11627), .ZN(n11658) );
  XNOR2_X1 U14576 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11657) );
  INV_X1 U14577 ( .A(n11657), .ZN(n11629) );
  XNOR2_X1 U14578 ( .A(n11658), .B(n11629), .ZN(n11867) );
  MUX2_X1 U14579 ( .A(n12100), .B(n11867), .S(n9602), .Z(n11886) );
  INV_X1 U14580 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n11630) );
  MUX2_X1 U14581 ( .A(n11886), .B(n11630), .S(n12321), .Z(n11631) );
  NOR2_X1 U14582 ( .A1(n11637), .A2(n11631), .ZN(n11632) );
  OR2_X1 U14583 ( .A1(n11696), .A2(n11632), .ZN(n14845) );
  OAI21_X1 U14584 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19865), .A(
        n11872), .ZN(n11894) );
  MUX2_X1 U14585 ( .A(n12761), .B(n11894), .S(n9602), .Z(n11634) );
  MUX2_X1 U14586 ( .A(n11634), .B(n11633), .S(n12321), .Z(n18942) );
  OR2_X1 U14587 ( .A1(n18942), .A2(n12758), .ZN(n12767) );
  NAND3_X1 U14588 ( .A1(n12321), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n11635) );
  NAND2_X1 U14589 ( .A1(n11639), .A2(n11635), .ZN(n18924) );
  NOR2_X1 U14590 ( .A1(n12767), .A2(n18924), .ZN(n11636) );
  NAND2_X1 U14591 ( .A1(n12767), .A2(n18924), .ZN(n12766) );
  OAI21_X1 U14592 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n11636), .A(
        n12766), .ZN(n12776) );
  INV_X1 U14593 ( .A(n11637), .ZN(n11641) );
  NAND2_X1 U14594 ( .A1(n11639), .A2(n11638), .ZN(n11640) );
  NAND2_X1 U14595 ( .A1(n11641), .A2(n11640), .ZN(n11642) );
  XNOR2_X1 U14596 ( .A(n11642), .B(n13053), .ZN(n12775) );
  OR2_X1 U14597 ( .A1(n12776), .A2(n12775), .ZN(n12778) );
  INV_X1 U14598 ( .A(n11642), .ZN(n14859) );
  NAND2_X1 U14599 ( .A1(n14859), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11643) );
  NAND2_X1 U14600 ( .A1(n12778), .A2(n11643), .ZN(n13481) );
  NAND2_X1 U14601 ( .A1(n13483), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11644) );
  NAND2_X1 U14602 ( .A1(n11645), .A2(n11644), .ZN(n13563) );
  AOI22_X1 U14603 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11564), .B1(
        n11602), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14604 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14605 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11597), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14606 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n11611), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11647) );
  NAND4_X1 U14607 ( .A1(n11650), .A2(n11649), .A3(n11648), .A4(n11647), .ZN(
        n11656) );
  AOI22_X1 U14608 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12120), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U14609 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n13828), .ZN(n11653) );
  INV_X1 U14610 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n20861) );
  AOI22_X1 U14611 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12170), .B1(
        n12169), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14612 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11651) );
  NAND4_X1 U14613 ( .A1(n11654), .A2(n11653), .A3(n11652), .A4(n11651), .ZN(
        n11655) );
  NAND2_X1 U14614 ( .A1(n11658), .A2(n11657), .ZN(n11660) );
  NAND2_X1 U14615 ( .A1(n19842), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11659) );
  NAND2_X1 U14616 ( .A1(n11660), .A2(n11659), .ZN(n11869) );
  INV_X1 U14617 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15668) );
  NAND2_X1 U14618 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15668), .ZN(
        n11870) );
  OR2_X1 U14619 ( .A1(n11869), .A2(n11870), .ZN(n11885) );
  MUX2_X1 U14620 ( .A(n12282), .B(n11885), .S(n9602), .Z(n11661) );
  INV_X1 U14621 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n18987) );
  MUX2_X1 U14622 ( .A(n11661), .B(n18987), .S(n12321), .Z(n11695) );
  XNOR2_X1 U14623 ( .A(n11696), .B(n11695), .ZN(n11662) );
  XNOR2_X1 U14624 ( .A(n11662), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13562) );
  NAND2_X1 U14625 ( .A1(n13563), .A2(n13562), .ZN(n11664) );
  INV_X1 U14626 ( .A(n11662), .ZN(n18907) );
  NAND2_X1 U14627 ( .A1(n18907), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11663) );
  AOI22_X1 U14628 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19360), .B1(
        n19292), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11673) );
  INV_X1 U14629 ( .A(n19419), .ZN(n19416) );
  AOI22_X1 U14630 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19639), .B1(
        n19416), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11672) );
  INV_X1 U14631 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13994) );
  INV_X1 U14632 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13996) );
  OAI22_X1 U14633 ( .A1(n13994), .A2(n19327), .B1(n19389), .B2(n13996), .ZN(
        n11668) );
  INV_X1 U14634 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13993) );
  INV_X1 U14635 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11666) );
  OAI22_X1 U14636 ( .A1(n13993), .A2(n19247), .B1(n11665), .B2(n11666), .ZN(
        n11667) );
  NOR2_X1 U14637 ( .A1(n11668), .A2(n11667), .ZN(n11671) );
  INV_X1 U14638 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14002) );
  INV_X1 U14639 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14005) );
  OAI22_X1 U14640 ( .A1(n14002), .A2(n19521), .B1(n19684), .B2(n14005), .ZN(
        n11669) );
  INV_X1 U14641 ( .A(n11669), .ZN(n11670) );
  INV_X1 U14642 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14003) );
  INV_X1 U14643 ( .A(n19458), .ZN(n11675) );
  INV_X1 U14644 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11674) );
  OAI22_X1 U14645 ( .A1(n14003), .A2(n19591), .B1(n11675), .B2(n11674), .ZN(
        n11678) );
  INV_X1 U14646 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14004) );
  INV_X1 U14647 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11676) );
  OAI22_X1 U14648 ( .A1(n14004), .A2(n19487), .B1(n19564), .B2(n11676), .ZN(
        n11677) );
  NOR2_X1 U14649 ( .A1(n11678), .A2(n11677), .ZN(n11680) );
  AOI22_X1 U14650 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19211), .B1(
        n19111), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11679) );
  NAND3_X1 U14651 ( .A1(n9664), .A2(n11680), .A3(n11679), .ZN(n11692) );
  AOI22_X1 U14652 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U14653 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14654 ( .A1(n11597), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U14655 ( .A1(n13113), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11611), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11681) );
  NAND4_X1 U14656 ( .A1(n11684), .A2(n11683), .A3(n11682), .A4(n11681), .ZN(
        n11690) );
  AOI22_X1 U14657 ( .A1(n12120), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14658 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13828), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14659 ( .A1(n12169), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U14660 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11685) );
  NAND4_X1 U14661 ( .A1(n11688), .A2(n11687), .A3(n11686), .A4(n11685), .ZN(
        n11689) );
  NAND2_X1 U14662 ( .A1(n11697), .A2(n19119), .ZN(n11691) );
  OR2_X2 U14663 ( .A1(n12281), .A2(n11693), .ZN(n11694) );
  NAND2_X2 U14664 ( .A1(n11694), .A2(n12297), .ZN(n12288) );
  NAND2_X1 U14665 ( .A1(n11696), .A2(n11695), .ZN(n11699) );
  MUX2_X1 U14666 ( .A(n11697), .B(P2_EBX_REG_5__SCAN_IN), .S(n12321), .Z(
        n11698) );
  NAND2_X1 U14667 ( .A1(n11699), .A2(n11698), .ZN(n11700) );
  NAND2_X1 U14668 ( .A1(n11742), .A2(n11700), .ZN(n18893) );
  INV_X1 U14669 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13600) );
  NAND2_X1 U14670 ( .A1(n13587), .A2(n13586), .ZN(n11703) );
  NAND2_X1 U14671 ( .A1(n11701), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11702) );
  AOI22_X1 U14672 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19360), .B1(
        n19292), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14673 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19639), .B1(
        n19458), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11711) );
  INV_X1 U14674 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14015) );
  INV_X1 U14675 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14018) );
  OAI22_X1 U14676 ( .A1(n14015), .A2(n19327), .B1(n19389), .B2(n14018), .ZN(
        n11706) );
  INV_X1 U14677 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14014) );
  INV_X1 U14678 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11704) );
  OAI22_X1 U14679 ( .A1(n14014), .A2(n19247), .B1(n11665), .B2(n11704), .ZN(
        n11705) );
  NOR2_X1 U14680 ( .A1(n11706), .A2(n11705), .ZN(n11710) );
  INV_X1 U14681 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14026) );
  INV_X1 U14682 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11707) );
  OAI22_X1 U14683 ( .A1(n14026), .A2(n19521), .B1(n19419), .B2(n11707), .ZN(
        n11708) );
  INV_X1 U14684 ( .A(n11708), .ZN(n11709) );
  INV_X1 U14685 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14024) );
  INV_X1 U14686 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11713) );
  OAI22_X1 U14687 ( .A1(n14024), .A2(n19487), .B1(n19591), .B2(n11713), .ZN(
        n11716) );
  INV_X1 U14688 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14028) );
  INV_X1 U14689 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11714) );
  OAI22_X1 U14690 ( .A1(n14028), .A2(n19684), .B1(n19564), .B2(n11714), .ZN(
        n11715) );
  NOR2_X1 U14691 ( .A1(n11716), .A2(n11715), .ZN(n11718) );
  AOI22_X1 U14692 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19211), .B1(
        n19111), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11717) );
  NAND3_X1 U14693 ( .A1(n9665), .A2(n11718), .A3(n11717), .ZN(n11730) );
  AOI22_X1 U14694 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11564), .B1(
        n11602), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11722) );
  AOI22_X1 U14695 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11597), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11721) );
  AOI22_X1 U14696 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n13113), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14697 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11646), .B1(
        n11611), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11719) );
  NAND4_X1 U14698 ( .A1(n11722), .A2(n11721), .A3(n11720), .A4(n11719), .ZN(
        n11728) );
  AOI22_X1 U14699 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12120), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U14700 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n13828), .ZN(n11725) );
  AOI22_X1 U14701 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12170), .B1(
        n12169), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11724) );
  AOI22_X1 U14702 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11723) );
  NAND4_X1 U14703 ( .A1(n11726), .A2(n11725), .A3(n11724), .A4(n11723), .ZN(
        n11727) );
  INV_X1 U14704 ( .A(n11731), .ZN(n12111) );
  NAND2_X1 U14705 ( .A1(n12111), .A2(n19119), .ZN(n11729) );
  INV_X1 U14706 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n18891) );
  MUX2_X1 U14707 ( .A(n11731), .B(n18891), .S(n12321), .Z(n11744) );
  INV_X1 U14708 ( .A(n11744), .ZN(n11732) );
  XNOR2_X1 U14709 ( .A(n11742), .B(n11732), .ZN(n18880) );
  INV_X1 U14710 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16198) );
  XNOR2_X1 U14711 ( .A(n11734), .B(n16198), .ZN(n15216) );
  NAND2_X1 U14712 ( .A1(n11734), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11735) );
  INV_X1 U14713 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n11738) );
  MUX2_X1 U14714 ( .A(n11738), .B(n11814), .S(n12077), .Z(n11743) );
  NAND2_X1 U14715 ( .A1(n11744), .A2(n11743), .ZN(n11739) );
  NAND2_X1 U14716 ( .A1(n12321), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11740) );
  OR2_X1 U14717 ( .A1(n11753), .A2(n11740), .ZN(n11741) );
  NAND2_X1 U14718 ( .A1(n11752), .A2(n11741), .ZN(n18858) );
  NOR2_X1 U14719 ( .A1(n18858), .A2(n12300), .ZN(n11747) );
  NAND2_X1 U14720 ( .A1(n11747), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16177) );
  INV_X1 U14721 ( .A(n11742), .ZN(n11745) );
  AOI21_X1 U14722 ( .B1(n11745), .B2(n11744), .A(n11743), .ZN(n11746) );
  OR2_X1 U14723 ( .A1(n11746), .A2(n11753), .ZN(n11749) );
  INV_X1 U14724 ( .A(n11749), .ZN(n18870) );
  NAND2_X1 U14725 ( .A1(n18870), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16178) );
  INV_X1 U14726 ( .A(n11747), .ZN(n11748) );
  INV_X1 U14727 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16199) );
  NAND2_X1 U14728 ( .A1(n11748), .A2(n16199), .ZN(n16176) );
  INV_X1 U14729 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16206) );
  NAND2_X1 U14730 ( .A1(n11749), .A2(n16206), .ZN(n16180) );
  AND2_X1 U14731 ( .A1(n16176), .A2(n16180), .ZN(n11750) );
  NAND2_X1 U14732 ( .A1(n12321), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11751) );
  XNOR2_X1 U14733 ( .A(n11752), .B(n11751), .ZN(n18850) );
  AOI21_X1 U14734 ( .B1(n18850), .B2(n11814), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15502) );
  NAND3_X1 U14735 ( .A1(n11756), .A2(n12321), .A3(P2_EBX_REG_10__SCAN_IN), 
        .ZN(n11754) );
  OAI211_X1 U14736 ( .C1(n11756), .C2(P2_EBX_REG_10__SCAN_IN), .A(n11854), .B(
        n11754), .ZN(n11761) );
  INV_X1 U14737 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11755) );
  OAI21_X1 U14738 ( .B1(n11761), .B2(n12300), .A(n11755), .ZN(n15486) );
  INV_X1 U14739 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13425) );
  NAND2_X1 U14740 ( .A1(n11854), .A2(n11768), .ZN(n11767) );
  INV_X1 U14741 ( .A(n11757), .ZN(n11758) );
  NAND2_X1 U14742 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n11758), .ZN(n11759) );
  NOR2_X1 U14743 ( .A1(n12077), .A2(n11759), .ZN(n11760) );
  NOR2_X1 U14744 ( .A1(n11767), .A2(n11760), .ZN(n18836) );
  AOI21_X1 U14745 ( .B1(n18836), .B2(n11814), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15471) );
  INV_X1 U14746 ( .A(n11761), .ZN(n14835) );
  AND2_X1 U14747 ( .A1(n11814), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11762) );
  NAND2_X1 U14748 ( .A1(n14835), .A2(n11762), .ZN(n15485) );
  AND2_X1 U14749 ( .A1(n11814), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11763) );
  NAND2_X1 U14750 ( .A1(n18850), .A2(n11763), .ZN(n15483) );
  NAND2_X1 U14751 ( .A1(n15485), .A2(n15483), .ZN(n15467) );
  INV_X1 U14752 ( .A(n18836), .ZN(n11765) );
  NAND2_X1 U14753 ( .A1(n11814), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11764) );
  NOR2_X1 U14754 ( .A1(n11765), .A2(n11764), .ZN(n15470) );
  NOR2_X1 U14755 ( .A1(n15467), .A2(n15470), .ZN(n11766) );
  NAND2_X1 U14756 ( .A1(n12321), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11770) );
  INV_X1 U14757 ( .A(n11768), .ZN(n11769) );
  OR2_X1 U14758 ( .A1(n11770), .A2(n11769), .ZN(n11771) );
  NAND2_X1 U14759 ( .A1(n11797), .A2(n11771), .ZN(n14818) );
  INV_X1 U14760 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11772) );
  NOR2_X1 U14761 ( .A1(n11773), .A2(n11772), .ZN(n15454) );
  NAND2_X1 U14762 ( .A1(n11773), .A2(n11772), .ZN(n15452) );
  INV_X1 U14763 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11774) );
  NOR2_X1 U14764 ( .A1(n12077), .A2(n11774), .ZN(n11796) );
  NOR2_X1 U14765 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(P2_EBX_REG_14__SCAN_IN), 
        .ZN(n11775) );
  INV_X1 U14766 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n14788) );
  NAND2_X1 U14767 ( .A1(n12321), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11784) );
  NOR2_X1 U14768 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(P2_EBX_REG_18__SCAN_IN), 
        .ZN(n11776) );
  NOR2_X1 U14769 ( .A1(n12077), .A2(n11776), .ZN(n11777) );
  INV_X1 U14770 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14917) );
  NAND2_X1 U14771 ( .A1(n11834), .A2(n11854), .ZN(n11832) );
  NAND2_X1 U14772 ( .A1(n12321), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11778) );
  NOR2_X1 U14773 ( .A1(n9667), .A2(n11778), .ZN(n11779) );
  NOR2_X1 U14774 ( .A1(n11832), .A2(n11779), .ZN(n14778) );
  INV_X1 U14775 ( .A(n14778), .ZN(n11780) );
  INV_X1 U14776 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15330) );
  OAI21_X1 U14777 ( .B1(n11780), .B2(n12300), .A(n15330), .ZN(n15102) );
  OR2_X1 U14778 ( .A1(n11807), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11809) );
  INV_X1 U14779 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11781) );
  NOR2_X1 U14780 ( .A1(n12077), .A2(n11781), .ZN(n11782) );
  NAND2_X1 U14781 ( .A1(n11809), .A2(n11782), .ZN(n11783) );
  AND2_X1 U14782 ( .A1(n11783), .A2(n11813), .ZN(n11824) );
  INV_X1 U14783 ( .A(n11824), .ZN(n18772) );
  INV_X1 U14784 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15357) );
  OAI21_X1 U14785 ( .B1(n18772), .B2(n12300), .A(n15357), .ZN(n15138) );
  OAI21_X1 U14786 ( .B1(n11785), .B2(n11784), .A(n11807), .ZN(n18797) );
  OR2_X1 U14787 ( .A1(n18797), .A2(n12300), .ZN(n11786) );
  INV_X1 U14788 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15368) );
  NOR2_X1 U14789 ( .A1(n12077), .A2(n14788), .ZN(n11788) );
  INV_X1 U14790 ( .A(n11854), .ZN(n11787) );
  AOI21_X1 U14791 ( .B1(n9661), .B2(n11788), .A(n11787), .ZN(n11789) );
  NAND2_X1 U14792 ( .A1(n11790), .A2(n11789), .ZN(n14791) );
  NAND2_X1 U14793 ( .A1(n11814), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11791) );
  INV_X1 U14794 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15174) );
  OAI21_X1 U14795 ( .B1(n14791), .B2(n12300), .A(n15174), .ZN(n11792) );
  NAND2_X1 U14796 ( .A1(n12321), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11793) );
  MUX2_X1 U14797 ( .A(n12321), .B(n11793), .S(n11799), .Z(n11794) );
  OR2_X1 U14798 ( .A1(n11799), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11803) );
  INV_X1 U14799 ( .A(n11825), .ZN(n11795) );
  INV_X1 U14800 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15422) );
  NAND2_X1 U14801 ( .A1(n11795), .A2(n15422), .ZN(n15416) );
  NAND2_X1 U14802 ( .A1(n11797), .A2(n11796), .ZN(n11798) );
  NAND2_X1 U14803 ( .A1(n11799), .A2(n11798), .ZN(n18819) );
  OR2_X1 U14804 ( .A1(n18819), .A2(n12300), .ZN(n11800) );
  INV_X1 U14805 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15197) );
  NAND2_X1 U14806 ( .A1(n11800), .A2(n15197), .ZN(n15194) );
  INV_X1 U14807 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11801) );
  NOR2_X1 U14808 ( .A1(n12077), .A2(n11801), .ZN(n11802) );
  NAND2_X1 U14809 ( .A1(n11803), .A2(n11802), .ZN(n11804) );
  AND2_X1 U14810 ( .A1(n11804), .A2(n9661), .ZN(n11821) );
  INV_X1 U14811 ( .A(n11821), .ZN(n14802) );
  INV_X1 U14812 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15404) );
  NAND4_X1 U14813 ( .A1(n15167), .A2(n15416), .A3(n15194), .A4(n15182), .ZN(
        n11805) );
  NOR2_X1 U14814 ( .A1(n15107), .A2(n11805), .ZN(n11806) );
  AND2_X1 U14815 ( .A1(n15138), .A2(n11806), .ZN(n11816) );
  NAND2_X1 U14816 ( .A1(n12321), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11808) );
  MUX2_X1 U14817 ( .A(n12321), .B(n11808), .S(n11807), .Z(n11810) );
  NAND2_X1 U14818 ( .A1(n18780), .A2(n11814), .ZN(n11811) );
  INV_X1 U14819 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11993) );
  NAND2_X1 U14820 ( .A1(n11811), .A2(n11993), .ZN(n15148) );
  NAND2_X1 U14821 ( .A1(n12321), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11812) );
  XNOR2_X1 U14822 ( .A(n11813), .B(n11812), .ZN(n18760) );
  NAND2_X1 U14823 ( .A1(n18760), .A2(n11814), .ZN(n11815) );
  INV_X1 U14824 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15342) );
  NAND2_X1 U14825 ( .A1(n11815), .A2(n15342), .ZN(n15120) );
  NAND4_X1 U14826 ( .A1(n15102), .A2(n11816), .A3(n15148), .A4(n15120), .ZN(
        n11830) );
  AND2_X1 U14827 ( .A1(n11814), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11817) );
  NAND2_X1 U14828 ( .A1(n14778), .A2(n11817), .ZN(n15101) );
  AND2_X1 U14829 ( .A1(n11814), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11818) );
  NAND2_X1 U14830 ( .A1(n18780), .A2(n11818), .ZN(n15147) );
  NAND2_X1 U14831 ( .A1(n11814), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11819) );
  OR2_X1 U14832 ( .A1(n18797), .A2(n11819), .ZN(n15108) );
  AND2_X1 U14833 ( .A1(n11814), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11820) );
  NAND2_X1 U14834 ( .A1(n11821), .A2(n11820), .ZN(n15181) );
  NAND2_X1 U14835 ( .A1(n11814), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11822) );
  AND4_X1 U14836 ( .A1(n15108), .A2(n15105), .A3(n15181), .A4(n15193), .ZN(
        n11826) );
  AND2_X1 U14837 ( .A1(n11814), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11823) );
  NAND2_X1 U14838 ( .A1(n11824), .A2(n11823), .ZN(n15137) );
  NAND2_X1 U14839 ( .A1(n11825), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15417) );
  AND4_X1 U14840 ( .A1(n15147), .A2(n11826), .A3(n15137), .A4(n15417), .ZN(
        n11828) );
  AND2_X1 U14841 ( .A1(n11814), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11827) );
  NAND2_X1 U14842 ( .A1(n18760), .A2(n11827), .ZN(n15119) );
  AND3_X1 U14843 ( .A1(n15101), .A2(n11828), .A3(n15119), .ZN(n11829) );
  INV_X1 U14844 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n16105) );
  NOR2_X1 U14845 ( .A1(n12077), .A2(n16105), .ZN(n11833) );
  INV_X1 U14846 ( .A(n11833), .ZN(n11831) );
  NAND2_X1 U14847 ( .A1(n11834), .A2(n11833), .ZN(n11835) );
  NAND2_X1 U14848 ( .A1(n11841), .A2(n11835), .ZN(n15695) );
  INV_X1 U14849 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15321) );
  NAND2_X1 U14850 ( .A1(n11836), .A2(n15321), .ZN(n15309) );
  NAND2_X1 U14851 ( .A1(n15308), .A2(n15309), .ZN(n11837) );
  INV_X1 U14852 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11838) );
  XNOR2_X1 U14853 ( .A(n11841), .B(n9714), .ZN(n16090) );
  NAND2_X1 U14854 ( .A1(n16090), .A2(n11814), .ZN(n11839) );
  XNOR2_X1 U14855 ( .A(n11839), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15096) );
  INV_X1 U14856 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15298) );
  OR2_X1 U14857 ( .A1(n11839), .A2(n15298), .ZN(n11840) );
  NAND3_X1 U14858 ( .A1(n11842), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n12321), 
        .ZN(n11843) );
  NAND2_X1 U14859 ( .A1(n11843), .A2(n11854), .ZN(n11844) );
  OR2_X1 U14860 ( .A1(n9686), .A2(n11844), .ZN(n16082) );
  NOR2_X1 U14861 ( .A1(n16082), .A2(n12300), .ZN(n11845) );
  AND2_X1 U14862 ( .A1(n11845), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15081) );
  INV_X1 U14863 ( .A(n11845), .ZN(n11846) );
  INV_X1 U14864 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n20927) );
  NAND2_X1 U14865 ( .A1(n11846), .A2(n20927), .ZN(n15080) );
  INV_X1 U14866 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n16072) );
  NAND3_X1 U14867 ( .A1(n12321), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n16071), 
        .ZN(n11847) );
  NAND2_X1 U14868 ( .A1(n15006), .A2(n11847), .ZN(n11848) );
  INV_X1 U14869 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15062) );
  OAI21_X1 U14870 ( .B1(n11848), .B2(n12300), .A(n15062), .ZN(n11850) );
  INV_X1 U14871 ( .A(n11848), .ZN(n16054) );
  AND2_X1 U14872 ( .A1(n11814), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11849) );
  NAND2_X1 U14873 ( .A1(n16054), .A2(n11849), .ZN(n11863) );
  NAND2_X1 U14874 ( .A1(n11850), .A2(n11863), .ZN(n15060) );
  NAND2_X1 U14875 ( .A1(n12321), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11852) );
  NAND2_X1 U14876 ( .A1(n11851), .A2(n11852), .ZN(n11859) );
  INV_X1 U14877 ( .A(n11852), .ZN(n11853) );
  NAND2_X1 U14878 ( .A1(n11854), .A2(n11814), .ZN(n11864) );
  INV_X1 U14879 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15276) );
  NAND2_X1 U14880 ( .A1(n11864), .A2(n15276), .ZN(n15069) );
  INV_X1 U14881 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15053) );
  INV_X1 U14882 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15042) );
  INV_X1 U14883 ( .A(n11859), .ZN(n11862) );
  INV_X1 U14884 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11857) );
  NOR2_X1 U14885 ( .A1(n12077), .A2(n11857), .ZN(n11858) );
  INV_X1 U14886 ( .A(n11858), .ZN(n11861) );
  INV_X1 U14887 ( .A(n12320), .ZN(n11860) );
  OAI21_X1 U14888 ( .B1(n11862), .B2(n11861), .A(n11860), .ZN(n16043) );
  NOR2_X1 U14889 ( .A1(n16043), .A2(n12300), .ZN(n15039) );
  INV_X1 U14890 ( .A(n11863), .ZN(n11865) );
  NOR2_X1 U14891 ( .A1(n11864), .A2(n15276), .ZN(n15071) );
  NAND2_X1 U14892 ( .A1(n12321), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12319) );
  XNOR2_X1 U14893 ( .A(n12320), .B(n12319), .ZN(n11866) );
  INV_X1 U14894 ( .A(n11866), .ZN(n16033) );
  NAND3_X1 U14895 ( .A1(n16033), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11814), .ZN(n15000) );
  INV_X1 U14896 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12265) );
  OAI21_X1 U14897 ( .B1(n11866), .B2(n12300), .A(n12265), .ZN(n12325) );
  NAND2_X1 U14898 ( .A1(n11885), .A2(n11867), .ZN(n11909) );
  NOR2_X1 U14899 ( .A1(n11901), .A2(n11909), .ZN(n11874) );
  INV_X1 U14900 ( .A(n11874), .ZN(n11876) );
  INV_X1 U14901 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15759) );
  INV_X1 U14902 ( .A(n11872), .ZN(n11873) );
  XNOR2_X1 U14903 ( .A(n11893), .B(n11873), .ZN(n11896) );
  NAND2_X1 U14904 ( .A1(n11896), .A2(n11874), .ZN(n11875) );
  OAI21_X1 U14905 ( .B1(n11894), .B2(n11876), .A(n13382), .ZN(n11877) );
  INV_X1 U14906 ( .A(n11877), .ZN(n11878) );
  NAND2_X1 U14907 ( .A1(n11878), .A2(n19757), .ZN(n11882) );
  NAND2_X1 U14908 ( .A1(n11531), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11879) );
  NAND2_X1 U14909 ( .A1(n11879), .A2(n15668), .ZN(n15664) );
  INV_X1 U14910 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n11880) );
  OAI21_X1 U14911 ( .B1(n12140), .B2(n15664), .A(n11880), .ZN(n11881) );
  NAND2_X1 U14912 ( .A1(n11881), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19859) );
  NAND2_X1 U14913 ( .A1(n11882), .A2(n19859), .ZN(n19875) );
  NOR2_X1 U14914 ( .A1(n11883), .A2(n19119), .ZN(n11884) );
  NAND2_X1 U14915 ( .A1(n19875), .A2(n11884), .ZN(n11892) );
  NOR2_X1 U14916 ( .A1(n11893), .A2(n11894), .ZN(n11887) );
  OAI211_X1 U14917 ( .C1(n11888), .C2(n11887), .A(n11886), .B(n11885), .ZN(
        n11889) );
  AND2_X1 U14918 ( .A1(n11889), .A2(n11910), .ZN(n19869) );
  INV_X1 U14919 ( .A(n14757), .ZN(n11890) );
  NAND2_X1 U14920 ( .A1(n19869), .A2(n19872), .ZN(n11891) );
  NAND2_X1 U14921 ( .A1(n11892), .A2(n11891), .ZN(n12389) );
  OAI21_X1 U14922 ( .B1(n11894), .B2(n11893), .A(n9808), .ZN(n11899) );
  INV_X1 U14923 ( .A(n11894), .ZN(n11897) );
  OAI211_X1 U14924 ( .C1(n19890), .C2(n11897), .A(n11895), .B(n11896), .ZN(
        n11898) );
  OAI211_X1 U14925 ( .C1(n11900), .C2(n11901), .A(n11899), .B(n11898), .ZN(
        n11907) );
  INV_X1 U14926 ( .A(n11909), .ZN(n11906) );
  NAND2_X1 U14927 ( .A1(n11422), .A2(n19890), .ZN(n11902) );
  NAND2_X1 U14928 ( .A1(n11902), .A2(n11901), .ZN(n11904) );
  NAND2_X1 U14929 ( .A1(n11904), .A2(n11903), .ZN(n11905) );
  NAND3_X1 U14930 ( .A1(n11907), .A2(n11906), .A3(n11905), .ZN(n11912) );
  NAND2_X1 U14931 ( .A1(n11910), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11908) );
  AOI21_X1 U14932 ( .B1(n9808), .B2(n11909), .A(n11908), .ZN(n11911) );
  OR2_X1 U14933 ( .A1(n13377), .A2(n11420), .ZN(n12854) );
  NAND2_X2 U14934 ( .A1(n19813), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19818) );
  INV_X1 U14935 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n18734) );
  NAND2_X1 U14936 ( .A1(n18734), .A2(n19774), .ZN(n19768) );
  NAND2_X1 U14937 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n16228) );
  NAND2_X1 U14938 ( .A1(n19891), .A2(n16228), .ZN(n13388) );
  NOR2_X1 U14939 ( .A1(n12854), .A2(n13388), .ZN(n13127) );
  NAND2_X1 U14940 ( .A1(n13127), .A2(n11927), .ZN(n11931) );
  NAND2_X1 U14941 ( .A1(n13389), .A2(n13382), .ZN(n12852) );
  OAI21_X1 U14942 ( .B1(n11913), .B2(n19157), .A(n14757), .ZN(n12034) );
  OAI21_X1 U14943 ( .B1(n11423), .B2(n19890), .A(n11895), .ZN(n11915) );
  NAND2_X1 U14944 ( .A1(n11915), .A2(n11914), .ZN(n11917) );
  NAND2_X1 U14945 ( .A1(n11917), .A2(n11916), .ZN(n11918) );
  AND3_X1 U14946 ( .A1(n12034), .A2(n11919), .A3(n11918), .ZN(n11924) );
  NAND2_X1 U14947 ( .A1(n11921), .A2(n11916), .ZN(n11922) );
  NAND2_X1 U14948 ( .A1(n11920), .A2(n11922), .ZN(n11923) );
  OAI211_X1 U14949 ( .C1(n12852), .C2(n13388), .A(n11924), .B(n11923), .ZN(
        n11925) );
  INV_X1 U14950 ( .A(n11925), .ZN(n13128) );
  NAND2_X1 U14951 ( .A1(n13377), .A2(n11895), .ZN(n11926) );
  NAND3_X1 U14952 ( .A1(n12854), .A2(n12040), .A3(n11926), .ZN(n11930) );
  MUX2_X1 U14953 ( .A(n13389), .B(n11927), .S(n19119), .Z(n11928) );
  NAND3_X1 U14954 ( .A1(n11928), .A2(n13382), .A3(n16228), .ZN(n11929) );
  NAND4_X1 U14955 ( .A1(n11931), .A2(n13128), .A3(n11930), .A4(n11929), .ZN(
        n11932) );
  NOR2_X1 U14956 ( .A1(n11883), .A2(n9602), .ZN(n19868) );
  NAND2_X2 U14957 ( .A1(n12316), .A2(n19868), .ZN(n16222) );
  NAND2_X1 U14958 ( .A1(n15019), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11939) );
  INV_X1 U14959 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n14817) );
  NAND2_X1 U14960 ( .A1(n12014), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11936) );
  NAND2_X1 U14961 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11935) );
  OAI211_X1 U14962 ( .C1(n14817), .C2(n9610), .A(n11936), .B(n11935), .ZN(
        n11937) );
  INV_X1 U14963 ( .A(n11937), .ZN(n11938) );
  NAND2_X1 U14964 ( .A1(n11939), .A2(n11938), .ZN(n14814) );
  INV_X1 U14965 ( .A(n11942), .ZN(n11944) );
  NAND2_X1 U14966 ( .A1(n11944), .A2(n11943), .ZN(n11945) );
  INV_X1 U14967 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11948) );
  NAND2_X1 U14968 ( .A1(n12014), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11947) );
  NAND2_X1 U14969 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11946) );
  OAI211_X1 U14970 ( .C1(n11948), .C2(n9610), .A(n11947), .B(n11946), .ZN(
        n11949) );
  AOI21_X1 U14971 ( .B1(n15019), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11949), .ZN(n13569) );
  INV_X1 U14972 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13588) );
  NAND2_X1 U14973 ( .A1(n12014), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11952) );
  NAND2_X1 U14974 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11951) );
  OAI211_X1 U14975 ( .C1(n13588), .C2(n9610), .A(n11952), .B(n11951), .ZN(
        n11953) );
  AOI21_X1 U14976 ( .B1(n15019), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11953), .ZN(n13146) );
  INV_X1 U14977 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n15526) );
  NAND2_X1 U14978 ( .A1(n15019), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11955) );
  AOI22_X1 U14979 ( .A1(n12014), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11954) );
  OAI211_X1 U14980 ( .C1(n9610), .C2(n15526), .A(n11955), .B(n11954), .ZN(
        n13166) );
  INV_X1 U14981 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n15210) );
  NAND2_X1 U14982 ( .A1(n12014), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11957) );
  NAND2_X1 U14983 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11956) );
  OAI211_X1 U14984 ( .C1(n15210), .C2(n9610), .A(n11957), .B(n11956), .ZN(
        n11958) );
  AOI21_X1 U14985 ( .B1(n15019), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n11958), .ZN(n13160) );
  NAND2_X1 U14986 ( .A1(n15019), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11964) );
  INV_X1 U14987 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n11961) );
  NAND2_X1 U14988 ( .A1(n12014), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11960) );
  NAND2_X1 U14989 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11959) );
  OAI211_X1 U14990 ( .C1(n11961), .C2(n9610), .A(n11960), .B(n11959), .ZN(
        n11962) );
  INV_X1 U14991 ( .A(n11962), .ZN(n11963) );
  NAND2_X1 U14992 ( .A1(n11964), .A2(n11963), .ZN(n16183) );
  INV_X1 U14993 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n11967) );
  NAND2_X1 U14994 ( .A1(n15019), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11966) );
  AOI22_X1 U14995 ( .A1(n15014), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11965) );
  OAI211_X1 U14996 ( .C1(n9610), .C2(n11967), .A(n11966), .B(n11965), .ZN(
        n13401) );
  INV_X1 U14997 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n11970) );
  NAND2_X1 U14998 ( .A1(n15019), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11969) );
  AOI22_X1 U14999 ( .A1(n15014), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11968) );
  OAI211_X1 U15000 ( .C1(n9610), .C2(n11970), .A(n11969), .B(n11968), .ZN(
        n14829) );
  INV_X1 U15001 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n11973) );
  NAND2_X1 U15002 ( .A1(n12014), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11972) );
  NAND2_X1 U15003 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11971) );
  OAI211_X1 U15004 ( .C1(n11973), .C2(n9610), .A(n11972), .B(n11971), .ZN(
        n11974) );
  AOI21_X1 U15005 ( .B1(n15019), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11974), .ZN(n13423) );
  NAND2_X1 U15006 ( .A1(n14814), .A2(n14813), .ZN(n13514) );
  INV_X1 U15007 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n15199) );
  NAND2_X1 U15008 ( .A1(n12014), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11976) );
  NAND2_X1 U15009 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11975) );
  OAI211_X1 U15010 ( .C1(n15199), .C2(n9610), .A(n11976), .B(n11975), .ZN(
        n11977) );
  AOI21_X1 U15011 ( .B1(n15019), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11977), .ZN(n13515) );
  INV_X1 U15012 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11980) );
  NAND2_X1 U15013 ( .A1(n15014), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11979) );
  NAND2_X1 U15014 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11978) );
  OAI211_X1 U15015 ( .C1(n11980), .C2(n9610), .A(n11979), .B(n11978), .ZN(
        n11981) );
  AOI21_X1 U15016 ( .B1(n15019), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11981), .ZN(n15424) );
  AOI22_X1 U15017 ( .A1(n15014), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11983) );
  NAND2_X1 U15018 ( .A1(n9613), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11982) );
  OAI211_X1 U15019 ( .C1(n12333), .C2(n15404), .A(n11983), .B(n11982), .ZN(
        n13579) );
  INV_X1 U15020 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n11986) );
  NAND2_X1 U15021 ( .A1(n12014), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11985) );
  NAND2_X1 U15022 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11984) );
  OAI211_X1 U15023 ( .C1(n11986), .C2(n9610), .A(n11985), .B(n11984), .ZN(
        n11987) );
  AOI21_X1 U15024 ( .B1(n15019), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11987), .ZN(n14784) );
  INV_X1 U15025 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20892) );
  NAND2_X1 U15026 ( .A1(n11999), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11989) );
  NAND2_X1 U15027 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11988) );
  OAI211_X1 U15028 ( .C1(n20892), .C2(n9610), .A(n11989), .B(n11988), .ZN(
        n11990) );
  AOI21_X1 U15029 ( .B1(n15019), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11990), .ZN(n14927) );
  AOI22_X1 U15030 ( .A1(n15014), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11992) );
  NAND2_X1 U15031 ( .A1(n9613), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11991) );
  OAI211_X1 U15032 ( .C1(n12333), .C2(n11993), .A(n11992), .B(n11991), .ZN(
        n15154) );
  AOI22_X1 U15033 ( .A1(n15014), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11995) );
  NAND2_X1 U15034 ( .A1(n9613), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11994) );
  OAI211_X1 U15035 ( .C1(n12333), .C2(n15357), .A(n11995), .B(n11994), .ZN(
        n14919) );
  INV_X1 U15036 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n15128) );
  NAND2_X1 U15037 ( .A1(n11999), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11997) );
  NAND2_X1 U15038 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11996) );
  OAI211_X1 U15039 ( .C1(n15128), .C2(n9610), .A(n11997), .B(n11996), .ZN(
        n11998) );
  AOI21_X1 U15040 ( .B1(n15019), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11998), .ZN(n15124) );
  NAND2_X1 U15041 ( .A1(n9613), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12001) );
  NAND2_X1 U15042 ( .A1(n11999), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12000) );
  OAI211_X1 U15043 ( .C1(n19757), .C2(n14768), .A(n12001), .B(n12000), .ZN(
        n12002) );
  AOI21_X1 U15044 ( .B1(n15019), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12002), .ZN(n14776) );
  INV_X1 U15045 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n12007) );
  NAND2_X1 U15046 ( .A1(n15014), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12006) );
  NAND2_X1 U15047 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12005) );
  OAI211_X1 U15048 ( .C1(n12007), .C2(n9610), .A(n12006), .B(n12005), .ZN(
        n12008) );
  AOI21_X1 U15049 ( .B1(n15019), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n12008), .ZN(n15312) );
  AOI22_X1 U15050 ( .A1(n15014), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n12010) );
  NAND2_X1 U15051 ( .A1(n9611), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12009) );
  OAI211_X1 U15052 ( .C1(n12333), .C2(n15298), .A(n12010), .B(n12009), .ZN(
        n14910) );
  INV_X1 U15053 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19804) );
  NAND2_X1 U15054 ( .A1(n12014), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12012) );
  NAND2_X1 U15055 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12011) );
  OAI211_X1 U15056 ( .C1(n19804), .C2(n9610), .A(n12012), .B(n12011), .ZN(
        n12013) );
  AOI21_X1 U15057 ( .B1(n15019), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n12013), .ZN(n14902) );
  INV_X1 U15058 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19806) );
  NAND2_X1 U15059 ( .A1(n12014), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12016) );
  NAND2_X1 U15060 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12015) );
  OAI211_X1 U15061 ( .C1(n19806), .C2(n9610), .A(n12016), .B(n12015), .ZN(
        n12017) );
  AOI21_X1 U15062 ( .B1(n15019), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n12017), .ZN(n14894) );
  AOI22_X1 U15063 ( .A1(n15014), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n12019) );
  NAND2_X1 U15064 ( .A1(n9613), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12018) );
  OAI211_X1 U15065 ( .C1(n12333), .C2(n15062), .A(n12019), .B(n12018), .ZN(
        n14887) );
  AOI22_X1 U15066 ( .A1(n15014), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12021) );
  NAND2_X1 U15067 ( .A1(n9612), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12020) );
  OAI211_X1 U15068 ( .C1(n12333), .C2(n15053), .A(n12021), .B(n12020), .ZN(
        n14706) );
  AOI22_X1 U15069 ( .A1(n15014), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12023) );
  NAND2_X1 U15070 ( .A1(n9613), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12022) );
  OAI211_X1 U15071 ( .C1(n12333), .C2(n15042), .A(n12023), .B(n12022), .ZN(
        n14872) );
  AOI22_X1 U15072 ( .A1(n15014), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12025) );
  NAND2_X1 U15073 ( .A1(n9612), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12024) );
  OAI211_X1 U15074 ( .C1(n12333), .C2(n12265), .A(n12025), .B(n12024), .ZN(
        n12027) );
  OAI21_X1 U15075 ( .B1(n12026), .B2(n12027), .A(n15011), .ZN(n15032) );
  INV_X1 U15076 ( .A(n15032), .ZN(n16035) );
  NAND2_X1 U15077 ( .A1(n13350), .A2(n19119), .ZN(n12028) );
  NAND2_X1 U15078 ( .A1(n12028), .A2(n11459), .ZN(n12029) );
  AND3_X1 U15079 ( .A1(n19119), .A2(n11916), .A3(n12077), .ZN(n12032) );
  NAND2_X1 U15080 ( .A1(n12316), .A2(n13378), .ZN(n15381) );
  NAND2_X1 U15081 ( .A1(n12033), .A2(n19890), .ZN(n13341) );
  NAND2_X1 U15082 ( .A1(n13341), .A2(n12034), .ZN(n12036) );
  NAND2_X1 U15083 ( .A1(n12036), .A2(n12035), .ZN(n12043) );
  NAND2_X1 U15084 ( .A1(n12037), .A2(n12049), .ZN(n12039) );
  NAND2_X1 U15085 ( .A1(n12039), .A2(n12038), .ZN(n12041) );
  INV_X1 U15086 ( .A(n12038), .ZN(n12749) );
  AOI22_X1 U15087 ( .A1(n12041), .A2(n12805), .B1(n12749), .B2(n12040), .ZN(
        n12042) );
  NAND2_X1 U15088 ( .A1(n12043), .A2(n12042), .ZN(n12048) );
  INV_X1 U15089 ( .A(n12044), .ZN(n12045) );
  MUX2_X1 U15090 ( .A(n12045), .B(n11916), .S(n13368), .Z(n12046) );
  INV_X1 U15091 ( .A(n12046), .ZN(n12047) );
  NAND2_X1 U15092 ( .A1(n13354), .A2(n12049), .ZN(n12050) );
  NAND2_X1 U15093 ( .A1(n12316), .A2(n12050), .ZN(n15379) );
  NAND3_X1 U15094 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12066) );
  INV_X1 U15095 ( .A(n12066), .ZN(n12061) );
  INV_X1 U15096 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15541) );
  NOR2_X1 U15097 ( .A1(n15541), .A2(n12758), .ZN(n12062) );
  INV_X1 U15098 ( .A(n12316), .ZN(n12051) );
  NAND2_X1 U15099 ( .A1(n19837), .A2(n19757), .ZN(n18736) );
  INV_X1 U15100 ( .A(n13051), .ZN(n18784) );
  INV_X2 U15101 ( .A(n18784), .ZN(n18871) );
  NAND2_X1 U15102 ( .A1(n12051), .A2(n18871), .ZN(n16215) );
  OAI21_X1 U15103 ( .B1(n15379), .B2(n12062), .A(n16215), .ZN(n13055) );
  NOR2_X1 U15104 ( .A1(n15379), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12052) );
  NOR2_X1 U15105 ( .A1(n13055), .A2(n12052), .ZN(n13484) );
  INV_X1 U15106 ( .A(n16216), .ZN(n15523) );
  NOR2_X1 U15107 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12062), .ZN(
        n13048) );
  INV_X1 U15108 ( .A(n13048), .ZN(n13485) );
  INV_X1 U15109 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13567) );
  INV_X1 U15110 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13597) );
  NOR3_X1 U15111 ( .A1(n13567), .A2(n13600), .A3(n13597), .ZN(n15524) );
  INV_X1 U15112 ( .A(n15524), .ZN(n16197) );
  NOR4_X1 U15113 ( .A1(n16199), .A2(n16198), .A3(n16206), .A4(n16197), .ZN(
        n12064) );
  NAND2_X1 U15114 ( .A1(n13485), .A2(n12064), .ZN(n12053) );
  NAND2_X1 U15115 ( .A1(n15523), .A2(n12053), .ZN(n12054) );
  AND2_X1 U15116 ( .A1(n13484), .A2(n12054), .ZN(n15514) );
  NAND2_X1 U15117 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15433) );
  NOR2_X1 U15118 ( .A1(n15433), .A2(n15422), .ZN(n12055) );
  AND3_X1 U15119 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15430) );
  AND2_X1 U15120 ( .A1(n12055), .A2(n15430), .ZN(n12309) );
  OR2_X1 U15121 ( .A1(n16216), .A2(n12309), .ZN(n12056) );
  NAND2_X1 U15122 ( .A1(n15514), .A2(n12056), .ZN(n15409) );
  NAND2_X1 U15123 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15385) );
  NAND2_X1 U15124 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12057) );
  NOR2_X1 U15125 ( .A1(n15385), .A2(n12057), .ZN(n12310) );
  NOR2_X1 U15126 ( .A1(n16216), .A2(n12310), .ZN(n12058) );
  OR2_X1 U15127 ( .A1(n15409), .A2(n12058), .ZN(n15372) );
  AND2_X1 U15128 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12311) );
  NOR2_X1 U15129 ( .A1(n16216), .A2(n12311), .ZN(n12059) );
  NOR2_X1 U15130 ( .A1(n15372), .A2(n12059), .ZN(n15327) );
  NAND3_X1 U15131 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12312) );
  NAND2_X1 U15132 ( .A1(n15523), .A2(n12312), .ZN(n12060) );
  AND2_X1 U15133 ( .A1(n15327), .A2(n12060), .ZN(n15287) );
  OAI21_X1 U15134 ( .B1(n16216), .B2(n12061), .A(n15287), .ZN(n15252) );
  INV_X1 U15135 ( .A(n12062), .ZN(n13091) );
  NOR2_X1 U15136 ( .A1(n13053), .A2(n13091), .ZN(n13047) );
  OAI21_X1 U15137 ( .B1(n13378), .B2(n13047), .A(n13485), .ZN(n12063) );
  NAND2_X1 U15138 ( .A1(n12309), .A2(n15507), .ZN(n15384) );
  INV_X1 U15139 ( .A(n12310), .ZN(n12065) );
  NOR2_X1 U15140 ( .A1(n15384), .A2(n12065), .ZN(n15358) );
  NAND2_X1 U15141 ( .A1(n15331), .A2(n9836), .ZN(n15283) );
  OR2_X1 U15142 ( .A1(n15283), .A2(n12066), .ZN(n15233) );
  NOR2_X1 U15143 ( .A1(n15233), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15250) );
  OR2_X1 U15144 ( .A1(n15252), .A2(n15250), .ZN(n15243) );
  INV_X1 U15145 ( .A(n15243), .ZN(n12068) );
  NAND2_X1 U15146 ( .A1(n15042), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12067) );
  OR2_X1 U15147 ( .A1(n15233), .A2(n12067), .ZN(n15240) );
  AOI21_X1 U15148 ( .B1(n12068), .B2(n15240), .A(n12265), .ZN(n12269) );
  INV_X1 U15149 ( .A(n12069), .ZN(n12070) );
  AND2_X1 U15150 ( .A1(n12070), .A2(n12031), .ZN(n13375) );
  INV_X1 U15151 ( .A(n13375), .ZN(n13117) );
  NAND2_X1 U15152 ( .A1(n12748), .A2(n11920), .ZN(n13374) );
  NAND2_X1 U15153 ( .A1(n13374), .A2(n19890), .ZN(n12071) );
  NAND2_X1 U15154 ( .A1(n13117), .A2(n12071), .ZN(n12072) );
  NOR2_X1 U15155 ( .A1(n13675), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12073) );
  AOI22_X1 U15156 ( .A1(n15224), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12079), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12076) );
  NOR2_X1 U15157 ( .A1(n19890), .A2(n12077), .ZN(n12074) );
  INV_X2 U15158 ( .A(n12208), .ZN(n12119) );
  NAND2_X1 U15159 ( .A1(n12119), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12075) );
  NAND2_X1 U15160 ( .A1(n12076), .A2(n12075), .ZN(n13039) );
  INV_X1 U15161 ( .A(n12817), .ZN(n12809) );
  NAND2_X1 U15162 ( .A1(n12809), .A2(n12079), .ZN(n12096) );
  INV_X1 U15163 ( .A(n12090), .ZN(n12084) );
  NOR2_X1 U15164 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19883), .ZN(
        n19862) );
  INV_X1 U15165 ( .A(n19862), .ZN(n12080) );
  NAND2_X1 U15166 ( .A1(n12084), .A2(n12080), .ZN(n12081) );
  AND2_X1 U15167 ( .A1(n12096), .A2(n12081), .ZN(n12082) );
  INV_X1 U15168 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n20815) );
  OAI21_X1 U15169 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(P2_EAX_REG_0__SCAN_IN), 
        .A(n12084), .ZN(n12086) );
  NAND2_X1 U15170 ( .A1(n19890), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12085) );
  AOI22_X1 U15171 ( .A1(n12073), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12079), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12089) );
  NAND2_X1 U15172 ( .A1(n12119), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12088) );
  NAND2_X1 U15173 ( .A1(n12089), .A2(n12088), .ZN(n12093) );
  OR2_X1 U15174 ( .A1(n12271), .A2(n12112), .ZN(n12092) );
  AOI22_X1 U15175 ( .A1(n12817), .A2(n12090), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12091) );
  NAND2_X1 U15176 ( .A1(n12092), .A2(n12091), .ZN(n12933) );
  NAND2_X1 U15177 ( .A1(n12232), .A2(n12094), .ZN(n12095) );
  OAI211_X1 U15178 ( .C1(n19883), .C2(n20880), .A(n12096), .B(n12095), .ZN(
        n12097) );
  NOR2_X1 U15179 ( .A1(n13039), .A2(n13040), .ZN(n13041) );
  NOR2_X1 U15180 ( .A1(n12098), .A2(n12097), .ZN(n12099) );
  NAND2_X1 U15181 ( .A1(n12119), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U15182 ( .A1(n12079), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12103) );
  NAND2_X1 U15183 ( .A1(n12232), .A2(n12100), .ZN(n12102) );
  NAND2_X1 U15184 ( .A1(n15224), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12101) );
  NAND4_X1 U15185 ( .A1(n12104), .A2(n12103), .A3(n12102), .A4(n12101), .ZN(
        n13240) );
  AOI22_X1 U15186 ( .A1(n15224), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12079), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12107) );
  NAND2_X1 U15187 ( .A1(n12119), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12106) );
  NAND2_X1 U15188 ( .A1(n12232), .A2(n12282), .ZN(n12105) );
  AOI22_X1 U15189 ( .A1(n12119), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n15224), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12110) );
  AOI22_X1 U15190 ( .A1(n12232), .A2(n12108), .B1(n12079), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12109) );
  NAND2_X1 U15191 ( .A1(n12110), .A2(n12109), .ZN(n13599) );
  AOI22_X1 U15192 ( .A1(n15224), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12079), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12115) );
  NAND2_X1 U15193 ( .A1(n12119), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12114) );
  NAND2_X1 U15194 ( .A1(n12115), .A2(n12114), .ZN(n12999) );
  INV_X1 U15195 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19035) );
  OAI222_X1 U15196 ( .A1(n16206), .A2(n12118), .B1(n12117), .B2(n19035), .C1(
        n12208), .C2(n15210), .ZN(n13037) );
  AOI22_X1 U15197 ( .A1(n15224), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12079), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12134) );
  NAND2_X1 U15198 ( .A1(n12119), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15199 ( .A1(n12120), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12125) );
  AOI22_X1 U15200 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11597), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12124) );
  AOI22_X1 U15201 ( .A1(n12121), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15202 ( .A1(n11646), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11611), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12122) );
  NAND4_X1 U15203 ( .A1(n12125), .A2(n12124), .A3(n12123), .A4(n12122), .ZN(
        n12131) );
  AOI22_X1 U15204 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15205 ( .A1(n12170), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13828), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12128) );
  AOI22_X1 U15206 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15207 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12169), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12126) );
  NAND4_X1 U15208 ( .A1(n12129), .A2(n12128), .A3(n12127), .A4(n12126), .ZN(
        n12130) );
  NAND2_X1 U15209 ( .A1(n12232), .A2(n13399), .ZN(n12132) );
  AOI22_X1 U15210 ( .A1(n12119), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U15211 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n11564), .B1(
        n11602), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15212 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U15213 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11597), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U15214 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11611), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12135) );
  NAND4_X1 U15215 ( .A1(n12138), .A2(n12137), .A3(n12136), .A4(n12135), .ZN(
        n12149) );
  AOI22_X1 U15216 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12120), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12147) );
  AOI22_X1 U15217 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n13828), .ZN(n12146) );
  AOI22_X1 U15218 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12170), .B1(
        n12169), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12145) );
  INV_X1 U15219 ( .A(n12139), .ZN(n13831) );
  INV_X1 U15220 ( .A(n12140), .ZN(n13830) );
  INV_X1 U15221 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12141) );
  OAI22_X1 U15222 ( .A1(n13831), .A2(n12142), .B1(n13830), .B2(n12141), .ZN(
        n12143) );
  INV_X1 U15223 ( .A(n12143), .ZN(n12144) );
  NAND4_X1 U15224 ( .A1(n12147), .A2(n12146), .A3(n12145), .A4(n12144), .ZN(
        n12148) );
  AOI22_X1 U15225 ( .A1(n12232), .A2(n18970), .B1(n15224), .B2(
        P2_EAX_REG_9__SCAN_IN), .ZN(n12150) );
  NAND2_X1 U15226 ( .A1(n12151), .A2(n12150), .ZN(n15505) );
  AOI22_X1 U15227 ( .A1(n15224), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12164) );
  NAND2_X1 U15228 ( .A1(n12119), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15229 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n11564), .B1(
        n11602), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12155) );
  AOI22_X1 U15230 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11597), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U15231 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n12121), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U15232 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11611), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12152) );
  NAND4_X1 U15233 ( .A1(n12155), .A2(n12154), .A3(n12153), .A4(n12152), .ZN(
        n12161) );
  AOI22_X1 U15234 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12120), .B1(
        n12139), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15235 ( .A1(n12169), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n13828), .ZN(n12158) );
  AOI22_X1 U15236 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n13876), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U15237 ( .A1(n13703), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12156) );
  NAND4_X1 U15238 ( .A1(n12159), .A2(n12158), .A3(n12157), .A4(n12156), .ZN(
        n12160) );
  NAND2_X1 U15239 ( .A1(n12232), .A2(n18969), .ZN(n12162) );
  AOI22_X1 U15240 ( .A1(n12119), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U15241 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n11564), .B1(
        n11602), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15242 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15243 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11597), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U15244 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11611), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12165) );
  NAND4_X1 U15245 ( .A1(n12168), .A2(n12167), .A3(n12166), .A4(n12165), .ZN(
        n12180) );
  AOI22_X1 U15246 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12120), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15247 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n13828), .ZN(n12177) );
  INV_X1 U15248 ( .A(n12169), .ZN(n12173) );
  INV_X1 U15249 ( .A(n12170), .ZN(n12172) );
  INV_X1 U15250 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12171) );
  OAI22_X1 U15251 ( .A1(n11515), .A2(n12173), .B1(n12172), .B2(n12171), .ZN(
        n12174) );
  INV_X1 U15252 ( .A(n12174), .ZN(n12176) );
  AOI22_X1 U15253 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12175) );
  NAND4_X1 U15254 ( .A1(n12178), .A2(n12177), .A3(n12176), .A4(n12175), .ZN(
        n12179) );
  AOI22_X1 U15255 ( .A1(n12232), .A2(n18964), .B1(n15224), .B2(
        P2_EAX_REG_11__SCAN_IN), .ZN(n12181) );
  NAND2_X1 U15256 ( .A1(n12182), .A2(n12181), .ZN(n13432) );
  AOI22_X1 U15257 ( .A1(n15224), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12195) );
  NAND2_X1 U15258 ( .A1(n12119), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15259 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11564), .B1(
        n11602), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15260 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12185) );
  AOI22_X1 U15261 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11597), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U15262 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11611), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12183) );
  NAND4_X1 U15263 ( .A1(n12186), .A2(n12185), .A3(n12184), .A4(n12183), .ZN(
        n12192) );
  AOI22_X1 U15264 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12120), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15265 ( .A1(n12140), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n13828), .ZN(n12189) );
  AOI22_X1 U15266 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12169), .B1(
        n13876), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U15267 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12187) );
  NAND4_X1 U15268 ( .A1(n12190), .A2(n12189), .A3(n12188), .A4(n12187), .ZN(
        n12191) );
  NAND2_X1 U15269 ( .A1(n12232), .A2(n18963), .ZN(n12193) );
  AOI22_X1 U15270 ( .A1(n15224), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15271 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15272 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15273 ( .A1(n11597), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U15274 ( .A1(n13113), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11611), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12196) );
  NAND4_X1 U15275 ( .A1(n12199), .A2(n12198), .A3(n12197), .A4(n12196), .ZN(
        n12205) );
  AOI22_X1 U15276 ( .A1(n12120), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15277 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13828), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U15278 ( .A1(n12169), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12201) );
  AOI22_X1 U15279 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12200) );
  NAND4_X1 U15280 ( .A1(n12203), .A2(n12202), .A3(n12201), .A4(n12200), .ZN(
        n12204) );
  NAND2_X1 U15281 ( .A1(n12232), .A2(n13513), .ZN(n12206) );
  OAI211_X1 U15282 ( .C1(n12208), .C2(n15199), .A(n12207), .B(n12206), .ZN(
        n13523) );
  AOI22_X1 U15283 ( .A1(n15224), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12221) );
  NAND2_X1 U15284 ( .A1(n12119), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15285 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12120), .B1(
        n11602), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15286 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11597), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U15287 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n12121), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15288 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11611), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12209) );
  NAND4_X1 U15289 ( .A1(n12212), .A2(n12211), .A3(n12210), .A4(n12209), .ZN(
        n12218) );
  AOI22_X1 U15290 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n11564), .B1(
        n12139), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15291 ( .A1(n12169), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n13828), .ZN(n12215) );
  AOI22_X1 U15292 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12170), .B1(
        n13876), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U15293 ( .A1(n13703), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12213) );
  NAND4_X1 U15294 ( .A1(n12216), .A2(n12215), .A3(n12214), .A4(n12213), .ZN(
        n12217) );
  NAND2_X1 U15295 ( .A1(n12232), .A2(n13577), .ZN(n12219) );
  AOI22_X1 U15296 ( .A1(n12119), .A2(P2_REIP_REG_15__SCAN_IN), .B1(n15224), 
        .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U15297 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n11564), .B1(
        n11602), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15298 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15299 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n11597), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15300 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11611), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12222) );
  NAND4_X1 U15301 ( .A1(n12225), .A2(n12224), .A3(n12223), .A4(n12222), .ZN(
        n12231) );
  AOI22_X1 U15302 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12120), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15303 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n13828), .ZN(n12228) );
  AOI22_X1 U15304 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12170), .B1(
        n12169), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15305 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12226) );
  NAND4_X1 U15306 ( .A1(n12229), .A2(n12228), .A3(n12227), .A4(n12226), .ZN(
        n12230) );
  AOI22_X1 U15307 ( .A1(n12232), .A2(n13578), .B1(n12079), .B2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12233) );
  NAND2_X1 U15308 ( .A1(n12234), .A2(n12233), .ZN(n13613) );
  NAND2_X1 U15309 ( .A1(n13611), .A2(n13613), .ZN(n13612) );
  AOI22_X1 U15310 ( .A1(n15224), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12236) );
  NAND2_X1 U15311 ( .A1(n12119), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12235) );
  NAND2_X1 U15312 ( .A1(n12236), .A2(n12235), .ZN(n13691) );
  AOI22_X1 U15313 ( .A1(n15224), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12238) );
  NAND2_X1 U15314 ( .A1(n12119), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12237) );
  NAND2_X1 U15315 ( .A1(n12238), .A2(n12237), .ZN(n13692) );
  NAND2_X1 U15316 ( .A1(n13691), .A2(n13692), .ZN(n12239) );
  AOI22_X1 U15317 ( .A1(n15224), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12241) );
  NAND2_X1 U15318 ( .A1(n12119), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12240) );
  NAND2_X1 U15319 ( .A1(n12241), .A2(n12240), .ZN(n15366) );
  AOI22_X1 U15320 ( .A1(n15224), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12243) );
  NAND2_X1 U15321 ( .A1(n12119), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12242) );
  AOI222_X1 U15322 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n12119), .B1(n15224), 
        .B2(P2_EAX_REG_20__SCAN_IN), .C1(n12079), .C2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15341) );
  AOI22_X1 U15323 ( .A1(n15224), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12245) );
  NAND2_X1 U15324 ( .A1(n12119), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12244) );
  NAND2_X1 U15325 ( .A1(n12245), .A2(n12244), .ZN(n14767) );
  AOI22_X1 U15326 ( .A1(n15224), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12247) );
  NAND2_X1 U15327 ( .A1(n12119), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12246) );
  NAND2_X1 U15328 ( .A1(n12247), .A2(n12246), .ZN(n15317) );
  AOI22_X1 U15329 ( .A1(n15224), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12249) );
  NAND2_X1 U15330 ( .A1(n12119), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12248) );
  NOR2_X2 U15331 ( .A1(n14986), .A2(n14985), .ZN(n14976) );
  AOI22_X1 U15332 ( .A1(n15224), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12251) );
  NAND2_X1 U15333 ( .A1(n12119), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12250) );
  NAND2_X1 U15334 ( .A1(n12251), .A2(n12250), .ZN(n14975) );
  AOI22_X1 U15335 ( .A1(n15224), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12253) );
  NAND2_X1 U15336 ( .A1(n12119), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15337 ( .A1(n12073), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12255) );
  NAND2_X1 U15338 ( .A1(n12119), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12254) );
  AND2_X1 U15339 ( .A1(n12255), .A2(n12254), .ZN(n14955) );
  AOI22_X1 U15340 ( .A1(n12073), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12257) );
  NAND2_X1 U15341 ( .A1(n12119), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12256) );
  AND2_X1 U15342 ( .A1(n12257), .A2(n12256), .ZN(n14754) );
  NOR2_X4 U15343 ( .A1(n14958), .A2(n14754), .ZN(n14941) );
  AOI22_X1 U15344 ( .A1(n12073), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12259) );
  NAND2_X1 U15345 ( .A1(n12119), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12258) );
  NAND2_X1 U15346 ( .A1(n12259), .A2(n12258), .ZN(n14940) );
  AOI22_X1 U15347 ( .A1(n12073), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12261) );
  NAND2_X1 U15348 ( .A1(n12119), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12260) );
  NAND2_X1 U15349 ( .A1(n12261), .A2(n12260), .ZN(n12263) );
  NOR2_X1 U15350 ( .A1(n12262), .A2(n12263), .ZN(n12264) );
  NAND2_X1 U15351 ( .A1(n19090), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15028) );
  INV_X1 U15352 ( .A(n15233), .ZN(n12266) );
  AND2_X1 U15353 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12314) );
  NAND3_X1 U15354 ( .A1(n12266), .A2(n12314), .A3(n12265), .ZN(n12267) );
  OAI211_X1 U15355 ( .C1(n16204), .C2(n14935), .A(n15028), .B(n12267), .ZN(
        n12268) );
  AOI211_X1 U15356 ( .C1(n16035), .C2(n16218), .A(n12269), .B(n12268), .ZN(
        n12318) );
  NAND2_X1 U15357 ( .A1(n12761), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12760) );
  NOR2_X1 U15358 ( .A1(n12271), .A2(n12760), .ZN(n12273) );
  INV_X1 U15359 ( .A(n12761), .ZN(n12270) );
  NOR2_X1 U15360 ( .A1(n12270), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12272) );
  XNOR2_X1 U15361 ( .A(n12272), .B(n12271), .ZN(n12770) );
  NOR2_X1 U15362 ( .A1(n15541), .A2(n12770), .ZN(n12769) );
  NOR2_X1 U15363 ( .A1(n12273), .A2(n12769), .ZN(n12277) );
  XNOR2_X1 U15364 ( .A(n13053), .B(n12277), .ZN(n12781) );
  INV_X1 U15365 ( .A(n12781), .ZN(n12276) );
  XNOR2_X1 U15366 ( .A(n12275), .B(n12274), .ZN(n12779) );
  NAND2_X1 U15367 ( .A1(n12276), .A2(n12779), .ZN(n12783) );
  OR2_X1 U15368 ( .A1(n12277), .A2(n13053), .ZN(n12278) );
  NAND2_X1 U15369 ( .A1(n12783), .A2(n12278), .ZN(n12279) );
  XNOR2_X1 U15370 ( .A(n12279), .B(n13567), .ZN(n13490) );
  NAND2_X1 U15371 ( .A1(n12279), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12280) );
  INV_X1 U15372 ( .A(n12281), .ZN(n12285) );
  NAND2_X1 U15373 ( .A1(n12283), .A2(n9991), .ZN(n12284) );
  NAND2_X1 U15374 ( .A1(n12285), .A2(n12284), .ZN(n13564) );
  AND2_X1 U15375 ( .A1(n12288), .A2(n13600), .ZN(n13590) );
  INV_X1 U15376 ( .A(n13590), .ZN(n12286) );
  OR2_X2 U15377 ( .A1(n12288), .A2(n13600), .ZN(n12290) );
  INV_X1 U15378 ( .A(n12294), .ZN(n12293) );
  INV_X1 U15379 ( .A(n12290), .ZN(n13591) );
  INV_X1 U15380 ( .A(n12298), .ZN(n12291) );
  NAND2_X1 U15381 ( .A1(n12295), .A2(n12294), .ZN(n12296) );
  XNOR2_X1 U15382 ( .A(n12306), .B(n12300), .ZN(n15204) );
  NAND2_X1 U15383 ( .A1(n15204), .A2(n16206), .ZN(n12301) );
  NAND2_X1 U15384 ( .A1(n15206), .A2(n12301), .ZN(n12304) );
  INV_X1 U15385 ( .A(n15204), .ZN(n12302) );
  NAND2_X1 U15386 ( .A1(n12302), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12303) );
  XNOR2_X1 U15387 ( .A(n12305), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16185) );
  NAND2_X1 U15388 ( .A1(n16186), .A2(n16185), .ZN(n12308) );
  AND2_X2 U15389 ( .A1(n15196), .A2(n12309), .ZN(n15421) );
  INV_X1 U15390 ( .A(n12313), .ZN(n15063) );
  NOR2_X1 U15391 ( .A1(n15063), .A2(n15053), .ZN(n15052) );
  AOI21_X1 U15392 ( .B1(n15052), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12315) );
  NAND2_X1 U15393 ( .A1(n12314), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15231) );
  NAND2_X1 U15394 ( .A1(n15034), .A2(n16192), .ZN(n12317) );
  OAI211_X1 U15395 ( .C1(n15036), .C2(n16222), .A(n12318), .B(n12317), .ZN(
        P2_U3017) );
  NAND2_X1 U15396 ( .A1(n12320), .A2(n12319), .ZN(n15004) );
  NAND2_X1 U15397 ( .A1(n12321), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12322) );
  AOI21_X1 U15398 ( .B1(n16026), .B2(n11814), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15002) );
  INV_X1 U15399 ( .A(n16026), .ZN(n12323) );
  INV_X1 U15400 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15232) );
  INV_X1 U15401 ( .A(n15001), .ZN(n12324) );
  NOR2_X1 U15402 ( .A1(n15002), .A2(n12324), .ZN(n12328) );
  NAND2_X1 U15403 ( .A1(n15003), .A2(n15000), .ZN(n12327) );
  XNOR2_X1 U15404 ( .A(n12328), .B(n12327), .ZN(n12412) );
  NOR2_X1 U15405 ( .A1(n12391), .A2(n16227), .ZN(n12335) );
  AOI22_X1 U15406 ( .A1(n15014), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12332) );
  NAND2_X1 U15407 ( .A1(n9613), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12331) );
  OAI211_X1 U15408 ( .C1(n12333), .C2(n15232), .A(n12332), .B(n12331), .ZN(
        n15012) );
  XOR2_X1 U15409 ( .A(n15012), .B(n15011), .Z(n16032) );
  INV_X1 U15410 ( .A(n16032), .ZN(n12398) );
  AND2_X1 U15411 ( .A1(n12398), .A2(n16218), .ZN(n12334) );
  OR2_X1 U15412 ( .A1(n15523), .A2(n13055), .ZN(n15263) );
  AOI21_X1 U15413 ( .B1(n15231), .B2(n15263), .A(n15252), .ZN(n15229) );
  AOI22_X1 U15414 ( .A1(n12073), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12337) );
  NAND2_X1 U15415 ( .A1(n12119), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12336) );
  NAND2_X1 U15416 ( .A1(n12337), .A2(n12336), .ZN(n12339) );
  INV_X1 U15417 ( .A(n12338), .ZN(n12341) );
  INV_X1 U15418 ( .A(n12339), .ZN(n12340) );
  NAND2_X1 U15419 ( .A1(n12341), .A2(n12340), .ZN(n12342) );
  NOR2_X1 U15420 ( .A1(n15233), .A2(n10034), .ZN(n12344) );
  INV_X1 U15421 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n12343) );
  NOR2_X1 U15422 ( .A1(n13051), .A2(n12343), .ZN(n12404) );
  INV_X1 U15423 ( .A(n12346), .ZN(n12347) );
  OAI21_X1 U15424 ( .B1(n15229), .B2(n15232), .A(n12347), .ZN(n12348) );
  INV_X1 U15425 ( .A(n12348), .ZN(n12349) );
  OAI211_X1 U15426 ( .C1(n12412), .C2(n16222), .A(n12350), .B(n12349), .ZN(
        P2_U3016) );
  AOI22_X1 U15427 ( .A1(n10457), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12353), .ZN(n12354) );
  INV_X1 U15428 ( .A(n12354), .ZN(n12355) );
  NAND2_X1 U15429 ( .A1(n12918), .A2(n13624), .ZN(n13015) );
  NAND2_X1 U15430 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20768) );
  INV_X1 U15431 ( .A(n12359), .ZN(n12912) );
  NOR3_X1 U15432 ( .A1(n12362), .A2(n12361), .A3(n12360), .ZN(n12363) );
  NAND2_X1 U15433 ( .A1(n12364), .A2(n12363), .ZN(n12365) );
  NAND2_X1 U15434 ( .A1(n12366), .A2(n12365), .ZN(n12843) );
  NOR2_X1 U15435 ( .A1(n12843), .A2(n20687), .ZN(n13002) );
  NAND2_X1 U15436 ( .A1(n12912), .A2(n13002), .ZN(n12923) );
  NAND2_X1 U15437 ( .A1(n12367), .A2(n12368), .ZN(n12369) );
  NOR4_X1 U15438 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n12375) );
  NOR4_X1 U15439 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12374) );
  NOR4_X1 U15440 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n12373) );
  NOR4_X1 U15441 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12372) );
  AND4_X1 U15442 ( .A1(n12375), .A2(n12374), .A3(n12373), .A4(n12372), .ZN(
        n12380) );
  NOR4_X1 U15443 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_27__SCAN_IN), .A4(
        P1_ADDRESS_REG_0__SCAN_IN), .ZN(n12378) );
  NOR4_X1 U15444 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n12377) );
  NOR4_X1 U15445 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n12376) );
  AND4_X1 U15446 ( .A1(n12378), .A2(n12377), .A3(n12376), .A4(n20698), .ZN(
        n12379) );
  NAND2_X1 U15447 ( .A1(n12380), .A2(n12379), .ZN(n12381) );
  AOI22_X1 U15448 ( .A1(n14355), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14366), .ZN(n12382) );
  INV_X1 U15449 ( .A(n12382), .ZN(n12385) );
  INV_X1 U15450 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16300) );
  NOR2_X1 U15451 ( .A1(n12385), .A2(n12384), .ZN(n12386) );
  AND2_X1 U15452 ( .A1(n13368), .A2(n12850), .ZN(n12388) );
  INV_X1 U15453 ( .A(n12757), .ZN(n12390) );
  NOR2_X1 U15454 ( .A1(n12391), .A2(n16169), .ZN(n12410) );
  NAND2_X1 U15455 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n18737), .ZN(n13134) );
  INV_X1 U15456 ( .A(n13134), .ZN(n12392) );
  OAI21_X1 U15457 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n18737), .ZN(n19885) );
  INV_X1 U15458 ( .A(n19885), .ZN(n12395) );
  INV_X1 U15459 ( .A(n13133), .ZN(n12394) );
  NOR2_X1 U15460 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19833) );
  OR2_X1 U15461 ( .A1(n19837), .A2(n19833), .ZN(n19849) );
  NAND2_X1 U15462 ( .A1(n19849), .A2(n18737), .ZN(n12399) );
  INV_X1 U15463 ( .A(n13076), .ZN(n12401) );
  NAND2_X1 U15464 ( .A1(n19630), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12400) );
  NAND2_X1 U15465 ( .A1(n12401), .A2(n12400), .ZN(n12762) );
  NAND2_X1 U15466 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n13494), .ZN(
        n14719) );
  INV_X1 U15467 ( .A(n14716), .ZN(n14723) );
  NAND2_X1 U15468 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n14726), .ZN(
        n14715) );
  AND2_X1 U15469 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12402) );
  INV_X1 U15470 ( .A(n14736), .ZN(n12403) );
  INV_X1 U15471 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14759) );
  INV_X1 U15472 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15043) );
  INV_X1 U15473 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15029) );
  XNOR2_X1 U15474 ( .A(n15027), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16028) );
  AOI21_X1 U15475 ( .B1(n16156), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n12404), .ZN(n12405) );
  OAI21_X1 U15476 ( .B1(n16166), .B2(n16028), .A(n12405), .ZN(n12406) );
  INV_X1 U15477 ( .A(n12406), .ZN(n12407) );
  OAI21_X1 U15478 ( .B1(n12412), .B2(n16168), .A(n12411), .ZN(P2_U2984) );
  INV_X1 U15479 ( .A(n14386), .ZN(n14305) );
  OR2_X1 U15480 ( .A1(n14111), .A2(n12414), .ZN(n12415) );
  NAND2_X1 U15481 ( .A1(n9660), .A2(n12415), .ZN(n14564) );
  INV_X1 U15482 ( .A(n9579), .ZN(n15592) );
  BUF_X4 U15483 ( .A(n12469), .Z(n17055) );
  AOI22_X1 U15484 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12424) );
  INV_X4 U15485 ( .A(n12438), .ZN(n17012) );
  AOI22_X1 U15486 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12423) );
  INV_X2 U15487 ( .A(n12588), .ZN(n17060) );
  AOI22_X1 U15488 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12422) );
  AOI22_X1 U15489 ( .A1(n16965), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15627), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12421) );
  NAND4_X1 U15490 ( .A1(n12424), .A2(n12423), .A3(n12422), .A4(n12421), .ZN(
        n12437) );
  NOR2_X2 U15491 ( .A1(n12428), .A2(n12430), .ZN(n17065) );
  INV_X4 U15492 ( .A(n15641), .ZN(n17041) );
  AOI22_X1 U15493 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12435) );
  AOI22_X1 U15494 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12434) );
  NOR2_X2 U15495 ( .A1(n12429), .A2(n12428), .ZN(n12495) );
  AOI22_X1 U15496 ( .A1(n17034), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12433) );
  INV_X2 U15497 ( .A(n10014), .ZN(n17066) );
  AOI22_X1 U15498 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12432) );
  NAND4_X1 U15499 ( .A1(n12435), .A2(n12434), .A3(n12433), .A4(n12432), .ZN(
        n12436) );
  INV_X2 U15500 ( .A(n15614), .ZN(n16806) );
  INV_X2 U15501 ( .A(n12588), .ZN(n15612) );
  AOI22_X1 U15502 ( .A1(n16806), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15612), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12442) );
  AOI22_X1 U15503 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12441) );
  INV_X2 U15505 ( .A(n10022), .ZN(n15626) );
  AOI22_X1 U15506 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15626), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12440) );
  AOI22_X1 U15507 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12439) );
  NAND4_X1 U15508 ( .A1(n12442), .A2(n12441), .A3(n12440), .A4(n12439), .ZN(
        n12448) );
  AOI22_X1 U15509 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15615), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12446) );
  AOI22_X1 U15510 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15627), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12445) );
  AOI22_X1 U15511 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12444) );
  INV_X2 U15512 ( .A(n10014), .ZN(n16983) );
  AOI22_X1 U15513 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12443) );
  NAND4_X1 U15514 ( .A1(n12446), .A2(n12445), .A3(n12444), .A4(n12443), .ZN(
        n12447) );
  AOI22_X1 U15515 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15626), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12452) );
  AOI22_X1 U15516 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15615), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12451) );
  AOI22_X1 U15517 ( .A1(n17065), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U15518 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12449) );
  NAND4_X1 U15519 ( .A1(n12452), .A2(n12451), .A3(n12450), .A4(n12449), .ZN(
        n12458) );
  INV_X2 U15520 ( .A(n16883), .ZN(n17051) );
  AOI22_X1 U15521 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12456) );
  AOI22_X1 U15522 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15612), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U15523 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U15524 ( .A1(n17034), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15627), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12453) );
  NAND4_X1 U15525 ( .A1(n12456), .A2(n12455), .A3(n12454), .A4(n12453), .ZN(
        n12457) );
  AOI22_X1 U15526 ( .A1(n12515), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12495), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U15527 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9579), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12461) );
  AOI22_X1 U15528 ( .A1(n12469), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15612), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12460) );
  AOI22_X1 U15529 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12475), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12459) );
  NAND4_X1 U15530 ( .A1(n12462), .A2(n12461), .A3(n12460), .A4(n12459), .ZN(
        n12468) );
  AOI22_X1 U15531 ( .A1(n17065), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15615), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12466) );
  AOI22_X1 U15532 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n16806), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12465) );
  AOI22_X1 U15533 ( .A1(n12470), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15627), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15534 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n15626), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12463) );
  NAND4_X1 U15535 ( .A1(n12466), .A2(n12465), .A3(n12464), .A4(n12463), .ZN(
        n12467) );
  AOI22_X1 U15536 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12469), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12484) );
  AOI22_X1 U15537 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15626), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12483) );
  INV_X1 U15538 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17095) );
  AOI22_X1 U15539 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15615), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12471) );
  OAI21_X1 U15540 ( .B1(n12472), .B2(n17095), .A(n12471), .ZN(n12481) );
  AOI22_X1 U15541 ( .A1(n12497), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12473), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12479) );
  AOI22_X1 U15542 ( .A1(n12427), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9579), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U15543 ( .A1(n12515), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12495), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U15544 ( .A1(n17065), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12475), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12476) );
  NAND4_X1 U15545 ( .A1(n12479), .A2(n12478), .A3(n12477), .A4(n12476), .ZN(
        n12480) );
  NAND3_X1 U15546 ( .A1(n12484), .A2(n12483), .A3(n12482), .ZN(n17237) );
  NAND2_X1 U15547 ( .A1(n17246), .A2(n17237), .ZN(n12526) );
  AOI22_X1 U15548 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15615), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12494) );
  INV_X2 U15549 ( .A(n10022), .ZN(n17064) );
  AOI22_X1 U15550 ( .A1(n17034), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17064), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12493) );
  INV_X1 U15551 ( .A(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n20839) );
  AOI22_X1 U15552 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12485) );
  OAI21_X1 U15553 ( .B1(n10015), .B2(n20839), .A(n12485), .ZN(n12491) );
  AOI22_X1 U15554 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12489) );
  AOI22_X1 U15555 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U15556 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U15557 ( .A1(n17065), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15627), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12486) );
  NAND4_X1 U15558 ( .A1(n12489), .A2(n12488), .A3(n12487), .A4(n12486), .ZN(
        n12490) );
  AOI211_X1 U15559 ( .C1(n16813), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n12491), .B(n12490), .ZN(n12492) );
  NAND3_X1 U15560 ( .A1(n12494), .A2(n12493), .A3(n12492), .ZN(n12701) );
  NAND2_X1 U15561 ( .A1(n12530), .A2(n12701), .ZN(n12508) );
  AOI22_X1 U15562 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U15563 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12505) );
  INV_X1 U15564 ( .A(n12495), .ZN(n16883) );
  INV_X2 U15565 ( .A(n15614), .ZN(n17034) );
  AOI22_X1 U15566 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12496) );
  OAI21_X1 U15567 ( .B1(n16883), .B2(n20820), .A(n12496), .ZN(n12503) );
  AOI22_X1 U15568 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12501) );
  AOI22_X1 U15569 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U15570 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12499) );
  AOI22_X1 U15571 ( .A1(n16965), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12498) );
  NAND4_X1 U15572 ( .A1(n12501), .A2(n12500), .A3(n12499), .A4(n12498), .ZN(
        n12502) );
  AOI211_X1 U15573 ( .C1(n17041), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n12503), .B(n12502), .ZN(n12504) );
  NAND3_X1 U15574 ( .A1(n12506), .A2(n12505), .A3(n12504), .ZN(n12702) );
  INV_X1 U15575 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18676) );
  NOR2_X1 U15576 ( .A1(n17608), .A2(n18676), .ZN(n12565) );
  INV_X1 U15577 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17752) );
  INV_X1 U15578 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17764) );
  INV_X1 U15579 ( .A(n12702), .ZN(n17222) );
  XNOR2_X1 U15580 ( .A(n12507), .B(n17222), .ZN(n12533) );
  NAND2_X1 U15581 ( .A1(n12533), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12534) );
  INV_X1 U15582 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17988) );
  XOR2_X1 U15583 ( .A(n12508), .B(n17226), .Z(n17674) );
  XNOR2_X1 U15584 ( .A(n12523), .B(n12510), .ZN(n17717) );
  AOI22_X1 U15585 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12514) );
  AOI22_X1 U15586 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16806), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12513) );
  AOI22_X1 U15587 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12512) );
  AOI22_X1 U15588 ( .A1(n17065), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12475), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12511) );
  NAND4_X1 U15589 ( .A1(n12514), .A2(n12513), .A3(n12512), .A4(n12511), .ZN(
        n12521) );
  AOI22_X1 U15590 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17064), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12519) );
  AOI22_X1 U15591 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12518) );
  AOI22_X1 U15592 ( .A1(n12515), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12517) );
  AOI22_X1 U15593 ( .A1(n12495), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12469), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12516) );
  NAND4_X1 U15594 ( .A1(n12519), .A2(n12518), .A3(n12517), .A4(n12516), .ZN(
        n12520) );
  NOR2_X1 U15595 ( .A1(n12521), .A2(n12520), .ZN(n17734) );
  INV_X1 U15596 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18694) );
  NOR2_X1 U15597 ( .A1(n17734), .A2(n18694), .ZN(n17733) );
  NAND2_X1 U15598 ( .A1(n17733), .A2(n17725), .ZN(n17724) );
  NAND2_X1 U15599 ( .A1(n12522), .A2(n17724), .ZN(n17716) );
  NAND2_X1 U15600 ( .A1(n17717), .A2(n17716), .ZN(n17715) );
  NAND2_X1 U15601 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12523), .ZN(
        n12524) );
  XOR2_X1 U15602 ( .A(n12526), .B(n17233), .Z(n17706) );
  NAND2_X1 U15603 ( .A1(n17705), .A2(n17706), .ZN(n17704) );
  NAND2_X1 U15604 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12527), .ZN(
        n12528) );
  NAND2_X2 U15605 ( .A1(n17704), .A2(n12528), .ZN(n12531) );
  XNOR2_X2 U15606 ( .A(n12531), .B(n12529), .ZN(n17694) );
  INV_X1 U15607 ( .A(n12701), .ZN(n17229) );
  XNOR2_X1 U15608 ( .A(n12530), .B(n17229), .ZN(n17695) );
  NAND2_X1 U15609 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12531), .ZN(
        n12532) );
  INV_X1 U15610 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17985) );
  XNOR2_X1 U15611 ( .A(n17985), .B(n12533), .ZN(n17667) );
  AOI21_X1 U15612 ( .B1(n15689), .B2(n12535), .A(n17608), .ZN(n12538) );
  NAND2_X1 U15613 ( .A1(n12538), .A2(n12537), .ZN(n12539) );
  NAND2_X1 U15614 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17926) );
  NOR2_X1 U15615 ( .A1(n17926), .A2(n17591), .ZN(n17929) );
  NAND2_X1 U15616 ( .A1(n17929), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17563) );
  NOR2_X1 U15617 ( .A1(n17563), .A2(n17573), .ZN(n17887) );
  NAND2_X1 U15618 ( .A1(n17887), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17555) );
  NOR2_X1 U15619 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17559) );
  NOR2_X1 U15620 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17873) );
  NOR2_X1 U15621 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17612) );
  NAND4_X1 U15622 ( .A1(n17559), .A2(n17873), .A3(n17612), .A4(n17591), .ZN(
        n12543) );
  OAI21_X1 U15623 ( .B1(n12542), .B2(n12543), .A(n17639), .ZN(n12546) );
  INV_X1 U15624 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17865) );
  INV_X1 U15625 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17853) );
  NAND2_X1 U15626 ( .A1(n12546), .A2(n12545), .ZN(n17450) );
  NAND2_X1 U15627 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17842) );
  INV_X1 U15628 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17850) );
  NOR2_X1 U15629 ( .A1(n17842), .A2(n17850), .ZN(n17474) );
  INV_X1 U15630 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17478) );
  NOR2_X1 U15631 ( .A1(n17839), .A2(n17478), .ZN(n17815) );
  NAND2_X1 U15632 ( .A1(n17474), .A2(n17815), .ZN(n17469) );
  INV_X1 U15633 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17472) );
  INV_X1 U15634 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17811) );
  INV_X1 U15635 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17792) );
  NOR2_X1 U15636 ( .A1(n16279), .A2(n17792), .ZN(n17423) );
  NAND2_X1 U15637 ( .A1(n17450), .A2(n17423), .ZN(n12548) );
  NOR2_X1 U15638 ( .A1(n17608), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17506) );
  NAND2_X1 U15639 ( .A1(n17506), .A2(n17839), .ZN(n12547) );
  NOR2_X1 U15640 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12547), .ZN(
        n17467) );
  NAND2_X1 U15641 ( .A1(n17467), .A2(n17472), .ZN(n17452) );
  NOR2_X2 U15642 ( .A1(n17425), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17424) );
  NAND3_X1 U15643 ( .A1(n17815), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15685) );
  INV_X1 U15644 ( .A(n15685), .ZN(n15681) );
  INV_X1 U15645 ( .A(n17842), .ZN(n12550) );
  NAND2_X1 U15646 ( .A1(n12550), .A2(n17450), .ZN(n17466) );
  NAND2_X2 U15647 ( .A1(n17476), .A2(n17466), .ZN(n17507) );
  NAND3_X1 U15648 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15681), .A3(
        n17507), .ZN(n17431) );
  NOR3_X2 U15649 ( .A1(n17424), .A2(n17792), .A3(n17431), .ZN(n12552) );
  INV_X1 U15650 ( .A(n12552), .ZN(n17415) );
  NOR2_X1 U15651 ( .A1(n17608), .A2(n17424), .ZN(n17414) );
  AOI221_X2 U15652 ( .B1(n17608), .B2(n17764), .C1(n17415), .C2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n17414), .ZN(n17401) );
  INV_X1 U15653 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17404) );
  NAND2_X1 U15654 ( .A1(n17401), .A2(n17404), .ZN(n17400) );
  NAND2_X1 U15655 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17744) );
  INV_X1 U15656 ( .A(n17744), .ZN(n12551) );
  NAND2_X1 U15657 ( .A1(n12552), .A2(n12551), .ZN(n12553) );
  NAND2_X1 U15658 ( .A1(n17752), .A2(n12555), .ZN(n16286) );
  INV_X1 U15659 ( .A(n16286), .ZN(n17383) );
  INV_X1 U15660 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16281) );
  NAND2_X1 U15661 ( .A1(n17383), .A2(n16281), .ZN(n15690) );
  NOR2_X2 U15662 ( .A1(n15690), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15745) );
  NOR2_X1 U15663 ( .A1(n17608), .A2(n15745), .ZN(n12562) );
  NAND2_X1 U15664 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16252) );
  INV_X1 U15665 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16265) );
  NOR2_X1 U15666 ( .A1(n16252), .A2(n16265), .ZN(n16267) );
  INV_X1 U15667 ( .A(n16267), .ZN(n15750) );
  AND2_X1 U15668 ( .A1(n18676), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12556) );
  NOR2_X1 U15669 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18676), .ZN(
        n16273) );
  INV_X1 U15670 ( .A(n16273), .ZN(n12557) );
  OAI21_X1 U15671 ( .B1(n12562), .B2(n12558), .A(n12557), .ZN(n12559) );
  NAND2_X1 U15672 ( .A1(n12559), .A2(n10026), .ZN(n12564) );
  AOI22_X1 U15673 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17608), .B1(
        n12560), .B2(n18676), .ZN(n12561) );
  OAI21_X1 U15674 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n12562), .A(
        n12561), .ZN(n12563) );
  OAI21_X1 U15675 ( .B1(n12565), .B2(n12564), .A(n12563), .ZN(n16274) );
  OAI21_X1 U15676 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18682), .A(
        n12567), .ZN(n12568) );
  NOR2_X1 U15677 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18545), .ZN(
        n12569) );
  NAND2_X1 U15678 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12568), .ZN(
        n12573) );
  AOI22_X1 U15679 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12574), .B1(
        n12569), .B2(n12573), .ZN(n12577) );
  OAI21_X1 U15680 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18533), .A(
        n12679), .ZN(n12678) );
  NOR2_X1 U15681 ( .A1(n12680), .A2(n12678), .ZN(n12576) );
  OAI21_X1 U15682 ( .B1(n12572), .B2(n12571), .A(n12577), .ZN(n12570) );
  AOI22_X1 U15683 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n15626), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12581) );
  AOI22_X1 U15684 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12580) );
  AOI22_X1 U15685 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U15686 ( .A1(n16965), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12578) );
  NAND4_X1 U15687 ( .A1(n12581), .A2(n12580), .A3(n12579), .A4(n12578), .ZN(
        n12587) );
  AOI22_X1 U15688 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U15689 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12584) );
  AOI22_X1 U15690 ( .A1(n16813), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U15691 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12582) );
  NAND4_X1 U15692 ( .A1(n12585), .A2(n12584), .A3(n12583), .A4(n12582), .ZN(
        n12586) );
  AOI22_X1 U15693 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12592) );
  AOI22_X1 U15694 ( .A1(n16813), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U15695 ( .A1(n16806), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12590) );
  AOI22_X1 U15696 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12589) );
  NAND4_X1 U15697 ( .A1(n12592), .A2(n12591), .A3(n12590), .A4(n12589), .ZN(
        n12598) );
  AOI22_X1 U15698 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U15699 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17064), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U15700 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12594) );
  AOI22_X1 U15701 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12593) );
  NAND4_X1 U15702 ( .A1(n12596), .A2(n12595), .A3(n12594), .A4(n12593), .ZN(
        n12597) );
  NAND2_X1 U15703 ( .A1(n18062), .A2(n16410), .ZN(n12689) );
  NOR2_X1 U15704 ( .A1(n16410), .A2(n18062), .ZN(n12663) );
  INV_X1 U15705 ( .A(n12663), .ZN(n12599) );
  NAND2_X1 U15706 ( .A1(n12689), .A2(n12599), .ZN(n18728) );
  AOI22_X1 U15707 ( .A1(n16813), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12603) );
  AOI22_X1 U15708 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12602) );
  AOI22_X1 U15709 ( .A1(n16806), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12601) );
  AOI22_X1 U15710 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17064), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12600) );
  NAND4_X1 U15711 ( .A1(n12603), .A2(n12602), .A3(n12601), .A4(n12600), .ZN(
        n12609) );
  AOI22_X1 U15712 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12607) );
  AOI22_X1 U15713 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12606) );
  AOI22_X1 U15714 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12605) );
  AOI22_X1 U15715 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16965), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12604) );
  NAND4_X1 U15716 ( .A1(n12607), .A2(n12606), .A3(n12605), .A4(n12604), .ZN(
        n12608) );
  AOI22_X1 U15717 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15612), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12619) );
  AOI22_X1 U15718 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16965), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U15719 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12610) );
  OAI21_X1 U15720 ( .B1(n15592), .B2(n20820), .A(n12610), .ZN(n12616) );
  AOI22_X1 U15721 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n15626), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U15722 ( .A1(n16813), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12613) );
  AOI22_X1 U15723 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12612) );
  AOI22_X1 U15724 ( .A1(n17052), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12611) );
  NAND4_X1 U15725 ( .A1(n12614), .A2(n12613), .A3(n12612), .A4(n12611), .ZN(
        n12615) );
  AOI211_X1 U15726 ( .C1(n17066), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n12616), .B(n12615), .ZN(n12617) );
  NAND3_X1 U15727 ( .A1(n12619), .A2(n12618), .A3(n12617), .ZN(n12686) );
  NOR2_X1 U15728 ( .A1(n18081), .A2(n12686), .ZN(n18510) );
  AOI22_X1 U15729 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U15730 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12628) );
  INV_X1 U15731 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n20893) );
  AOI22_X1 U15732 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15612), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12620) );
  OAI21_X1 U15733 ( .B1(n12438), .B2(n20893), .A(n12620), .ZN(n12626) );
  AOI22_X1 U15734 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12624) );
  AOI22_X1 U15735 ( .A1(n16813), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12623) );
  AOI22_X1 U15736 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16965), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12622) );
  AOI22_X1 U15737 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12621) );
  NAND4_X1 U15738 ( .A1(n12624), .A2(n12623), .A3(n12622), .A4(n12621), .ZN(
        n12625) );
  NAND2_X1 U15739 ( .A1(n18089), .A2(n17111), .ZN(n18528) );
  AOI22_X1 U15740 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12633) );
  AOI22_X1 U15741 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15615), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12632) );
  AOI22_X1 U15742 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U15743 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12630) );
  NAND4_X1 U15744 ( .A1(n12633), .A2(n12632), .A3(n12631), .A4(n12630), .ZN(
        n12639) );
  AOI22_X1 U15745 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15612), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12637) );
  AOI22_X1 U15746 ( .A1(n16806), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12636) );
  AOI22_X1 U15747 ( .A1(n16813), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15627), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12635) );
  AOI22_X1 U15748 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15626), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12634) );
  NAND4_X1 U15749 ( .A1(n12637), .A2(n12636), .A3(n12635), .A4(n12634), .ZN(
        n12638) );
  AOI22_X1 U15750 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n16806), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12643) );
  AOI22_X1 U15751 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17012), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12642) );
  AOI22_X1 U15752 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17060), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n9579), .ZN(n12641) );
  AOI22_X1 U15753 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17036), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12640) );
  NAND4_X1 U15754 ( .A1(n12643), .A2(n12642), .A3(n12641), .A4(n12640), .ZN(
        n12649) );
  AOI22_X1 U15755 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17052), .ZN(n12647) );
  AOI22_X1 U15756 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17064), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12646) );
  AOI22_X1 U15757 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n16965), .ZN(n12645) );
  INV_X2 U15758 ( .A(n10015), .ZN(n17035) );
  AOI22_X1 U15759 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17055), .ZN(n12644) );
  NAND4_X1 U15760 ( .A1(n12647), .A2(n12646), .A3(n12645), .A4(n12644), .ZN(
        n12648) );
  AOI22_X1 U15761 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17053), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12653) );
  AOI22_X1 U15762 ( .A1(n16813), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12652) );
  AOI22_X1 U15763 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15612), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12651) );
  AOI22_X1 U15764 ( .A1(n16965), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12650) );
  NAND4_X1 U15765 ( .A1(n12653), .A2(n12652), .A3(n12651), .A4(n12650), .ZN(
        n12659) );
  AOI22_X1 U15766 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12657) );
  AOI22_X1 U15767 ( .A1(n16806), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12656) );
  AOI22_X1 U15768 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15627), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U15769 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15626), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12654) );
  NAND4_X1 U15770 ( .A1(n12657), .A2(n12656), .A3(n12655), .A4(n12654), .ZN(
        n12658) );
  NOR2_X1 U15771 ( .A1(n9615), .A2(n18076), .ZN(n12674) );
  NAND2_X1 U15772 ( .A1(n18072), .A2(n12674), .ZN(n12660) );
  AOI21_X1 U15773 ( .B1(n15557), .B2(n18528), .A(n12660), .ZN(n12690) );
  NAND2_X1 U15774 ( .A1(n18510), .A2(n12690), .ZN(n15554) );
  NOR2_X2 U15775 ( .A1(n18728), .A2(n15554), .ZN(n18519) );
  NAND2_X1 U15776 ( .A1(n18062), .A2(n17185), .ZN(n12666) );
  NAND2_X1 U15777 ( .A1(n12687), .A2(n18509), .ZN(n15556) );
  NOR2_X1 U15778 ( .A1(n12666), .A2(n15556), .ZN(n12662) );
  NOR3_X1 U15779 ( .A1(n18062), .A2(n15557), .A3(n12660), .ZN(n12661) );
  NAND3_X1 U15780 ( .A1(n18089), .A2(n18085), .A3(n12661), .ZN(n15649) );
  NAND3_X1 U15781 ( .A1(n18081), .A2(n12686), .A3(n17111), .ZN(n12664) );
  NAND2_X1 U15782 ( .A1(n12673), .A2(n12685), .ZN(n15651) );
  NAND2_X1 U15783 ( .A1(n15649), .A2(n15651), .ZN(n16392) );
  NOR3_X1 U15784 ( .A1(n18510), .A2(n12687), .A3(n12685), .ZN(n12667) );
  NOR2_X1 U15785 ( .A1(n18085), .A2(n12685), .ZN(n15675) );
  OAI21_X1 U15786 ( .B1(n18094), .B2(n15763), .A(n12663), .ZN(n15654) );
  OAI21_X1 U15787 ( .B1(n12667), .B2(n15675), .A(n15654), .ZN(n12671) );
  INV_X1 U15788 ( .A(n12664), .ZN(n12670) );
  OAI211_X1 U15789 ( .C1(n18510), .C2(n18085), .A(n12689), .B(n17185), .ZN(
        n12665) );
  INV_X1 U15790 ( .A(n12665), .ZN(n12669) );
  AOI22_X1 U15791 ( .A1(n18062), .A2(n12667), .B1(n18076), .B2(n12666), .ZN(
        n12668) );
  OAI221_X1 U15792 ( .B1(n12670), .B2(n18072), .C1(n12670), .C2(n12669), .A(
        n12668), .ZN(n15652) );
  AOI21_X1 U15793 ( .B1(n12672), .B2(n12671), .A(n15652), .ZN(n12677) );
  NAND2_X1 U15794 ( .A1(n12673), .A2(n12677), .ZN(n15657) );
  INV_X1 U15795 ( .A(n12674), .ZN(n12675) );
  NAND3_X1 U15796 ( .A1(n12675), .A2(n16410), .A3(n15650), .ZN(n12676) );
  NAND2_X1 U15797 ( .A1(n12677), .A2(n12676), .ZN(n18508) );
  AOI21_X2 U15798 ( .B1(n18509), .B2(n18515), .A(n18508), .ZN(n18529) );
  INV_X1 U15799 ( .A(n12678), .ZN(n12683) );
  XOR2_X1 U15800 ( .A(n12680), .B(n12679), .Z(n12682) );
  INV_X1 U15801 ( .A(n18498), .ZN(n15672) );
  NOR2_X1 U15802 ( .A1(n18716), .A2(n12685), .ZN(n15671) );
  NAND2_X1 U15803 ( .A1(n15671), .A2(n12686), .ZN(n15676) );
  INV_X1 U15804 ( .A(n12687), .ZN(n12688) );
  NAND3_X1 U15805 ( .A1(n12690), .A2(n12689), .A3(n12688), .ZN(n15653) );
  NAND2_X1 U15806 ( .A1(n18675), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18566) );
  NAND2_X1 U15807 ( .A1(n16274), .A2(n17615), .ZN(n12731) );
  NOR2_X1 U15808 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18693) );
  INV_X1 U15809 ( .A(n18693), .ZN(n12695) );
  NAND2_X1 U15810 ( .A1(n18563), .A2(n18667), .ZN(n16389) );
  NAND2_X1 U15811 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17632) );
  NAND2_X1 U15812 ( .A1(n17683), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17662) );
  NAND2_X1 U15813 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17634) );
  NOR2_X1 U15814 ( .A1(n17634), .A2(n17621), .ZN(n17593) );
  NAND2_X1 U15815 ( .A1(n16424), .A2(n12691), .ZN(n17512) );
  NAND3_X1 U15816 ( .A1(n17487), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16420) );
  INV_X1 U15817 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12692) );
  XNOR2_X2 U15818 ( .A(n12694), .B(n12693), .ZN(n16723) );
  INV_X1 U15819 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18649) );
  INV_X1 U15820 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n12696) );
  NAND2_X2 U15821 ( .A1(n18730), .A2(n12696), .ZN(n18048) );
  NOR2_X1 U15822 ( .A1(n18649), .A2(n18048), .ZN(n16272) );
  NOR2_X1 U15823 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18720) );
  AOI21_X1 U15824 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n18720), .ZN(n18570) );
  INV_X1 U15825 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18715) );
  INV_X1 U15826 ( .A(n17579), .ZN(n17527) );
  OR2_X1 U15827 ( .A1(n9716), .A2(n17527), .ZN(n16240) );
  XOR2_X1 U15828 ( .A(n12693), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n12698) );
  NOR2_X1 U15829 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17482), .ZN(
        n16255) );
  NAND2_X1 U15830 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16257), .ZN(
        n16413) );
  AOI22_X1 U15831 ( .A1(n17489), .A2(n16413), .B1(n18374), .B2(n9716), .ZN(
        n12697) );
  NAND2_X1 U15832 ( .A1(n12697), .A2(n17735), .ZN(n16256) );
  NOR2_X1 U15833 ( .A1(n16255), .A2(n16256), .ZN(n16239) );
  OAI22_X1 U15834 ( .A1(n16240), .A2(n12698), .B1(n16239), .B2(n12693), .ZN(
        n12699) );
  AOI211_X1 U15835 ( .C1(n17582), .C2(n16723), .A(n16272), .B(n12699), .ZN(
        n12730) );
  NAND2_X1 U15836 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17742) );
  NOR2_X1 U15837 ( .A1(n17742), .A2(n17744), .ZN(n15686) );
  INV_X1 U15838 ( .A(n15686), .ZN(n16280) );
  NOR2_X1 U15839 ( .A1(n16279), .A2(n16280), .ZN(n17749) );
  NAND2_X1 U15840 ( .A1(n17871), .A2(n17749), .ZN(n17745) );
  NOR2_X1 U15841 ( .A1(n17745), .A2(n15750), .ZN(n16243) );
  NAND2_X1 U15842 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16243), .ZN(
        n12700) );
  XNOR2_X1 U15843 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12700), .ZN(
        n16275) );
  NOR2_X1 U15844 ( .A1(n12710), .A2(n17237), .ZN(n12708) );
  NOR2_X1 U15845 ( .A1(n17233), .A2(n12708), .ZN(n12707) );
  NAND2_X1 U15846 ( .A1(n12707), .A2(n12701), .ZN(n12705) );
  NOR2_X1 U15847 ( .A1(n17226), .A2(n12705), .ZN(n12704) );
  NAND2_X1 U15848 ( .A1(n12704), .A2(n12702), .ZN(n12703) );
  NOR2_X1 U15849 ( .A1(n15689), .A2(n12703), .ZN(n12725) );
  XNOR2_X1 U15850 ( .A(n17217), .B(n12703), .ZN(n17655) );
  XNOR2_X1 U15851 ( .A(n17222), .B(n12704), .ZN(n12718) );
  XOR2_X1 U15852 ( .A(n17226), .B(n12705), .Z(n12706) );
  NAND2_X1 U15853 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12706), .ZN(
        n12717) );
  XNOR2_X1 U15854 ( .A(n17988), .B(n12706), .ZN(n17679) );
  XNOR2_X1 U15855 ( .A(n17229), .B(n12707), .ZN(n17689) );
  XOR2_X1 U15856 ( .A(n17233), .B(n12708), .Z(n12709) );
  NAND2_X1 U15857 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12709), .ZN(
        n12715) );
  XNOR2_X1 U15858 ( .A(n12525), .B(n12709), .ZN(n17703) );
  XNOR2_X1 U15859 ( .A(n17237), .B(n12710), .ZN(n12711) );
  NAND2_X1 U15860 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12711), .ZN(
        n12714) );
  XOR2_X1 U15861 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12711), .Z(
        n17714) );
  INV_X1 U15862 ( .A(n17734), .ZN(n15764) );
  AOI21_X1 U15863 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17246), .A(
        n15764), .ZN(n12713) );
  NOR2_X1 U15864 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17246), .ZN(
        n12712) );
  AOI221_X1 U15865 ( .B1(n15764), .B2(n17246), .C1(n12713), .C2(n18694), .A(
        n12712), .ZN(n17713) );
  NAND2_X1 U15866 ( .A1(n17714), .A2(n17713), .ZN(n17712) );
  NAND2_X1 U15867 ( .A1(n12714), .A2(n17712), .ZN(n17702) );
  NAND2_X1 U15868 ( .A1(n17703), .A2(n17702), .ZN(n17701) );
  NAND2_X1 U15869 ( .A1(n12715), .A2(n17701), .ZN(n17690) );
  NAND2_X1 U15870 ( .A1(n17689), .A2(n17690), .ZN(n17688) );
  NOR2_X1 U15871 ( .A1(n17689), .A2(n17690), .ZN(n12716) );
  AOI21_X1 U15872 ( .B1(n12529), .B2(n17688), .A(n12716), .ZN(n17678) );
  NAND2_X1 U15873 ( .A1(n17679), .A2(n17678), .ZN(n17677) );
  NAND2_X1 U15874 ( .A1(n12717), .A2(n17677), .ZN(n12719) );
  NAND2_X1 U15875 ( .A1(n12718), .A2(n12719), .ZN(n12720) );
  XOR2_X1 U15876 ( .A(n12719), .B(n12718), .Z(n17661) );
  NAND2_X1 U15877 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17661), .ZN(
        n17660) );
  NAND2_X1 U15878 ( .A1(n12720), .A2(n17660), .ZN(n17654) );
  NOR2_X1 U15879 ( .A1(n17655), .A2(n17654), .ZN(n17653) );
  INV_X1 U15880 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17970) );
  NOR2_X1 U15881 ( .A1(n17653), .A2(n17970), .ZN(n12721) );
  NAND2_X1 U15882 ( .A1(n12725), .A2(n12721), .ZN(n12726) );
  INV_X1 U15883 ( .A(n12721), .ZN(n12724) );
  NAND2_X1 U15884 ( .A1(n17655), .A2(n17654), .ZN(n12723) );
  NAND2_X1 U15885 ( .A1(n12725), .A2(n12724), .ZN(n12722) );
  OAI211_X1 U15886 ( .C1(n12725), .C2(n12724), .A(n12723), .B(n12722), .ZN(
        n17641) );
  NAND2_X1 U15887 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17641), .ZN(
        n17640) );
  NAND2_X1 U15888 ( .A1(n17749), .A2(n17870), .ZN(n17746) );
  NAND3_X1 U15889 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16250), .A3(
        n16267), .ZN(n12727) );
  XOR2_X1 U15890 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12727), .Z(
        n16278) );
  NAND2_X1 U15891 ( .A1(n12731), .A2(n10021), .ZN(P3_U2799) );
  NOR2_X1 U15892 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12733) );
  NOR4_X1 U15893 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12732) );
  NAND4_X1 U15894 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12733), .A4(n12732), .ZN(n12746) );
  INV_X1 U15895 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n20778) );
  INV_X1 U15896 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20764) );
  NOR4_X1 U15897 ( .A1(n20778), .A2(n20764), .A3(P1_BE_N_REG_1__SCAN_IN), .A4(
        P1_BE_N_REG_3__SCAN_IN), .ZN(n12735) );
  NOR4_X1 U15898 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_2__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12734) );
  NAND3_X1 U15899 ( .A1(n20091), .A2(n12735), .A3(n12734), .ZN(U214) );
  NOR4_X1 U15900 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_16__SCAN_IN), .A3(P2_ADDRESS_REG_19__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n12739) );
  NOR4_X1 U15901 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_15__SCAN_IN), .A4(
        P2_ADDRESS_REG_0__SCAN_IN), .ZN(n12738) );
  NOR4_X1 U15902 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n12737) );
  NOR4_X1 U15903 ( .A1(P2_ADDRESS_REG_21__SCAN_IN), .A2(
        P2_ADDRESS_REG_24__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12736) );
  NAND4_X1 U15904 ( .A1(n12739), .A2(n12738), .A3(n12737), .A4(n12736), .ZN(
        n12744) );
  NOR4_X1 U15905 ( .A1(P2_ADDRESS_REG_3__SCAN_IN), .A2(
        P2_ADDRESS_REG_4__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n12742) );
  NOR4_X1 U15906 ( .A1(P2_ADDRESS_REG_8__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_6__SCAN_IN), .A4(
        P2_ADDRESS_REG_5__SCAN_IN), .ZN(n12741) );
  NOR4_X1 U15907 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12740) );
  NAND4_X1 U15908 ( .A1(n12742), .A2(n12741), .A3(n12740), .A4(n19786), .ZN(
        n12743) );
  NOR2_X1 U15909 ( .A1(n19101), .A2(n12746), .ZN(n16299) );
  NAND2_X1 U15910 ( .A1(n16299), .A2(U214), .ZN(U212) );
  NAND2_X1 U15911 ( .A1(n13382), .A2(n12850), .ZN(n12747) );
  NOR2_X1 U15912 ( .A1(n11920), .A2(n12747), .ZN(n18948) );
  INV_X1 U15913 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19899) );
  OAI211_X1 U15914 ( .C1(n18948), .C2(n19899), .A(n18736), .B(n14746), .ZN(
        P2_U2814) );
  NAND2_X1 U15915 ( .A1(n13374), .A2(n13382), .ZN(n12802) );
  NOR2_X1 U15916 ( .A1(n19878), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n12750)
         );
  AOI22_X1 U15917 ( .A1(n12750), .A2(n18736), .B1(n12749), .B2(n19878), .ZN(
        P2_U3612) );
  INV_X1 U15918 ( .A(n12843), .ZN(n12752) );
  AND2_X1 U15919 ( .A1(n12751), .A2(n12752), .ZN(n12833) );
  NAND2_X1 U15920 ( .A1(n12833), .A2(n13012), .ZN(n12791) );
  INV_X1 U15921 ( .A(n12791), .ZN(n12755) );
  INV_X1 U15922 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n20832) );
  AND2_X1 U15923 ( .A1(n20624), .A2(n15734), .ZN(n13777) );
  INV_X1 U15924 ( .A(n13777), .ZN(n12754) );
  OAI211_X1 U15925 ( .C1(n12755), .C2(n20832), .A(n13254), .B(n12754), .ZN(
        P1_U2801) );
  NAND2_X1 U15926 ( .A1(n12038), .A2(n16228), .ZN(n12801) );
  NAND2_X1 U15927 ( .A1(n12801), .A2(n13388), .ZN(n12756) );
  OR2_X1 U15928 ( .A1(n12802), .A2(n12756), .ZN(n13373) );
  AND2_X1 U15929 ( .A1(n13373), .A2(n12850), .ZN(n19876) );
  OAI21_X1 U15930 ( .B1(n11880), .B2(n19876), .A(n12757), .ZN(P2_U2819) );
  NAND2_X1 U15931 ( .A1(n18942), .A2(n12758), .ZN(n12759) );
  NAND2_X1 U15932 ( .A1(n12767), .A2(n12759), .ZN(n16221) );
  OAI22_X1 U15933 ( .A1(n19102), .A2(n13347), .B1(n16168), .B2(n16221), .ZN(
        n12765) );
  OAI21_X1 U15934 ( .B1(n12761), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12760), .ZN(n16226) );
  OAI21_X1 U15935 ( .B1(n16156), .B2(n12762), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12763) );
  OR2_X1 U15936 ( .A1(n18871), .A2(n20815), .ZN(n16224) );
  OAI211_X1 U15937 ( .C1(n16169), .C2(n16226), .A(n12763), .B(n16224), .ZN(
        n12764) );
  OR2_X1 U15938 ( .A1(n12765), .A2(n12764), .ZN(P2_U3014) );
  OAI21_X1 U15939 ( .B1(n12767), .B2(n18924), .A(n12766), .ZN(n12768) );
  XNOR2_X1 U15940 ( .A(n12768), .B(n15541), .ZN(n13096) );
  AOI21_X1 U15941 ( .B1(n15541), .B2(n12770), .A(n12769), .ZN(n13090) );
  INV_X1 U15942 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19776) );
  NOR2_X1 U15943 ( .A1(n18871), .A2(n19776), .ZN(n13089) );
  AOI21_X1 U15944 ( .B1(n19091), .B2(n13090), .A(n13089), .ZN(n12772) );
  NAND2_X1 U15945 ( .A1(n19089), .A2(n18930), .ZN(n12771) );
  OAI211_X1 U15946 ( .C1(n18930), .C2(n19100), .A(n12772), .B(n12771), .ZN(
        n12773) );
  AOI21_X1 U15947 ( .B1(n19094), .B2(n18929), .A(n12773), .ZN(n12774) );
  OAI21_X1 U15948 ( .B1(n13096), .B2(n16168), .A(n12774), .ZN(P2_U3013) );
  NAND2_X1 U15949 ( .A1(n12776), .A2(n12775), .ZN(n12777) );
  NAND2_X1 U15950 ( .A1(n12778), .A2(n12777), .ZN(n13044) );
  INV_X1 U15951 ( .A(n12779), .ZN(n12780) );
  NAND2_X1 U15952 ( .A1(n12781), .A2(n12780), .ZN(n12782) );
  NAND2_X1 U15953 ( .A1(n12783), .A2(n12782), .ZN(n13043) );
  AOI22_X1 U15954 ( .A1(n16156), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n19090), .ZN(n12786) );
  AOI21_X1 U15955 ( .B1(n12784), .B2(n18930), .A(n13494), .ZN(n14855) );
  NAND2_X1 U15956 ( .A1(n19089), .A2(n14855), .ZN(n12785) );
  OAI211_X1 U15957 ( .C1(n13043), .C2(n16169), .A(n12786), .B(n12785), .ZN(
        n12787) );
  AOI21_X1 U15958 ( .B1(n19094), .B2(n13057), .A(n12787), .ZN(n12788) );
  OAI21_X1 U15959 ( .B1(n16168), .B2(n13044), .A(n12788), .ZN(P2_U3012) );
  NAND2_X1 U15960 ( .A1(n12751), .A2(n10222), .ZN(n15706) );
  AND2_X1 U15961 ( .A1(n15706), .A2(n12753), .ZN(n12789) );
  INV_X1 U15962 ( .A(n20766), .ZN(n12793) );
  OAI21_X1 U15963 ( .B1(n13777), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n12793), 
        .ZN(n12792) );
  OAI21_X1 U15964 ( .B1(n12794), .B2(n12793), .A(n12792), .ZN(P1_U3487) );
  NAND2_X1 U15965 ( .A1(n13139), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12795) );
  AOI22_X1 U15966 ( .A1(n13081), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19837), .B2(n19865), .ZN(n12796) );
  NAND2_X1 U15967 ( .A1(n19890), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12799) );
  AND4_X1 U15968 ( .A1(n12798), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n12799), 
        .A4(n19883), .ZN(n12800) );
  INV_X1 U15969 ( .A(n13377), .ZN(n13376) );
  NAND2_X1 U15970 ( .A1(n13376), .A2(n13378), .ZN(n12804) );
  OR2_X1 U15971 ( .A1(n12802), .A2(n12801), .ZN(n12803) );
  NAND3_X1 U15972 ( .A1(n12829), .A2(n12806), .A3(n12805), .ZN(n12807) );
  NAND2_X1 U15973 ( .A1(n13131), .A2(n12807), .ZN(n12808) );
  AOI21_X1 U15974 ( .B1(n19861), .B2(n20791), .A(n18989), .ZN(n12822) );
  INV_X1 U15975 ( .A(n12810), .ZN(n12816) );
  INV_X1 U15976 ( .A(n12811), .ZN(n12814) );
  INV_X1 U15977 ( .A(n12812), .ZN(n12813) );
  NAND2_X1 U15978 ( .A1(n12814), .A2(n12813), .ZN(n12815) );
  NAND2_X1 U15979 ( .A1(n12816), .A2(n12815), .ZN(n12932) );
  AND2_X1 U15980 ( .A1(n12817), .A2(n13675), .ZN(n12818) );
  AOI22_X1 U15981 ( .A1(n19103), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19101), .ZN(n19109) );
  NOR2_X1 U15982 ( .A1(n13614), .A2(n19109), .ZN(n12820) );
  INV_X1 U15983 ( .A(n12932), .ZN(n18938) );
  NOR3_X1 U15984 ( .A1(n19861), .A2(n18938), .A3(n14996), .ZN(n12819) );
  AOI211_X1 U15985 ( .C1(P2_EAX_REG_0__SCAN_IN), .C2(n20780), .A(n12820), .B(
        n12819), .ZN(n12821) );
  OAI21_X1 U15986 ( .B1(n12822), .B2(n12932), .A(n12821), .ZN(P2_U2919) );
  NAND2_X1 U15987 ( .A1(n13081), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12824) );
  INV_X1 U15988 ( .A(n19519), .ZN(n13356) );
  NAND2_X1 U15989 ( .A1(n19857), .A2(n19865), .ZN(n19555) );
  AND2_X1 U15990 ( .A1(n13356), .A2(n19555), .ZN(n19286) );
  NAND2_X1 U15991 ( .A1(n19286), .A2(n19837), .ZN(n19489) );
  NAND2_X1 U15992 ( .A1(n12824), .A2(n19489), .ZN(n12825) );
  NAND2_X1 U15993 ( .A1(n13354), .A2(n12829), .ZN(n13112) );
  NAND2_X1 U15994 ( .A1(n13375), .A2(n13377), .ZN(n13129) );
  NAND2_X1 U15995 ( .A1(n13112), .A2(n13129), .ZN(n12830) );
  MUX2_X1 U15996 ( .A(n13355), .B(n12831), .S(n18983), .Z(n12832) );
  OAI21_X1 U15997 ( .B1(n19280), .B2(n18984), .A(n12832), .ZN(P2_U2886) );
  INV_X1 U15998 ( .A(n13008), .ZN(n12835) );
  INV_X1 U15999 ( .A(n12753), .ZN(n12834) );
  OAI22_X1 U16000 ( .A1(n12835), .A2(n13624), .B1(n12834), .B2(n12833), .ZN(
        n19902) );
  INV_X1 U16001 ( .A(n12836), .ZN(n12838) );
  INV_X1 U16002 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n12837) );
  NAND2_X1 U16003 ( .A1(n12838), .A2(n12837), .ZN(n15754) );
  INV_X1 U16004 ( .A(n15754), .ZN(n15732) );
  NOR3_X1 U16005 ( .A1(n13624), .A2(n13105), .A3(n15732), .ZN(n12839) );
  NOR2_X1 U16006 ( .A1(n12839), .A2(n20687), .ZN(n20770) );
  NOR2_X1 U16007 ( .A1(n19902), .A2(n20770), .ZN(n15722) );
  NOR2_X1 U16008 ( .A1(n15722), .A2(n19901), .ZN(n19910) );
  INV_X1 U16009 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n12849) );
  NAND3_X1 U16010 ( .A1(n12840), .A2(n13016), .A3(n10224), .ZN(n12841) );
  NAND3_X1 U16011 ( .A1(n13015), .A2(n15724), .A3(n12841), .ZN(n12842) );
  NAND2_X1 U16012 ( .A1(n13008), .A2(n12842), .ZN(n12845) );
  NAND2_X1 U16013 ( .A1(n12751), .A2(n12843), .ZN(n12844) );
  OAI211_X1 U16014 ( .C1(n13008), .C2(n12966), .A(n12845), .B(n12844), .ZN(
        n12846) );
  NAND2_X1 U16015 ( .A1(n12846), .A2(n10229), .ZN(n15723) );
  INV_X1 U16016 ( .A(n15723), .ZN(n12847) );
  NAND2_X1 U16017 ( .A1(n19910), .A2(n12847), .ZN(n12848) );
  OAI21_X1 U16018 ( .B1(n19910), .B2(n12849), .A(n12848), .ZN(P1_U3484) );
  INV_X1 U16019 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n12857) );
  INV_X1 U16020 ( .A(n11920), .ZN(n15665) );
  NAND2_X1 U16021 ( .A1(n15665), .A2(n12850), .ZN(n12853) );
  NAND2_X1 U16022 ( .A1(n14757), .A2(n12850), .ZN(n12851) );
  OAI21_X1 U16023 ( .B1(n12854), .B2(n12853), .A(n12897), .ZN(n12855) );
  NAND2_X1 U16024 ( .A1(n18737), .A2(n13133), .ZN(n19880) );
  INV_X2 U16025 ( .A(n19880), .ZN(n19045) );
  AOI22_X1 U16026 ( .A1(n19045), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12856) );
  OAI21_X1 U16027 ( .B1(n12857), .B2(n19014), .A(n12856), .ZN(P2_U2933) );
  INV_X1 U16028 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n12859) );
  AOI22_X1 U16029 ( .A1(n19045), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12858) );
  OAI21_X1 U16030 ( .B1(n12859), .B2(n19014), .A(n12858), .ZN(P2_U2934) );
  INV_X1 U16031 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14950) );
  AOI22_X1 U16032 ( .A1(n19045), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12860) );
  OAI21_X1 U16033 ( .B1(n14950), .B2(n19014), .A(n12860), .ZN(P2_U2924) );
  INV_X1 U16034 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n12862) );
  AOI22_X1 U16035 ( .A1(n19045), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12861) );
  OAI21_X1 U16036 ( .B1(n12862), .B2(n19014), .A(n12861), .ZN(P2_U2929) );
  INV_X1 U16037 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n12864) );
  AOI22_X1 U16038 ( .A1(n19045), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12863) );
  OAI21_X1 U16039 ( .B1(n12864), .B2(n19014), .A(n12863), .ZN(P2_U2932) );
  INV_X1 U16040 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n12866) );
  AOI22_X1 U16041 ( .A1(n19045), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12865) );
  OAI21_X1 U16042 ( .B1(n12866), .B2(n19014), .A(n12865), .ZN(P2_U2931) );
  INV_X1 U16043 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13677) );
  AOI22_X1 U16044 ( .A1(n19045), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n12867) );
  OAI21_X1 U16045 ( .B1(n13677), .B2(n19014), .A(n12867), .ZN(P2_U2935) );
  INV_X1 U16046 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U16047 ( .A1(n19045), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12868) );
  OAI21_X1 U16048 ( .B1(n12890), .B2(n19014), .A(n12868), .ZN(P2_U2925) );
  INV_X1 U16049 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n12870) );
  AOI22_X1 U16050 ( .A1(n19045), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12869) );
  OAI21_X1 U16051 ( .B1(n12870), .B2(n19014), .A(n12869), .ZN(P2_U2928) );
  INV_X1 U16052 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14978) );
  AOI22_X1 U16053 ( .A1(n19045), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12871) );
  OAI21_X1 U16054 ( .B1(n14978), .B2(n19014), .A(n12871), .ZN(P2_U2927) );
  INV_X1 U16055 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14966) );
  AOI22_X1 U16056 ( .A1(n19045), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12872) );
  OAI21_X1 U16057 ( .B1(n14966), .B2(n19014), .A(n12872), .ZN(P2_U2926) );
  INV_X1 U16058 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n12874) );
  AOI22_X1 U16059 ( .A1(n19045), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12873) );
  OAI21_X1 U16060 ( .B1(n12874), .B2(n19014), .A(n12873), .ZN(P2_U2930) );
  INV_X1 U16061 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n12876) );
  AOI22_X1 U16062 ( .A1(n19045), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12875) );
  OAI21_X1 U16063 ( .B1(n12876), .B2(n19014), .A(n12875), .ZN(P2_U2922) );
  INV_X1 U16064 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12887) );
  AOI22_X1 U16065 ( .A1(n19045), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12877) );
  OAI21_X1 U16066 ( .B1(n12887), .B2(n19014), .A(n12877), .ZN(P2_U2921) );
  NAND2_X1 U16067 ( .A1(n19413), .A2(n18954), .ZN(n12879) );
  NAND2_X1 U16068 ( .A1(n18945), .A2(n18988), .ZN(n12878) );
  OAI211_X1 U16069 ( .C1(n18988), .C2(n11633), .A(n12879), .B(n12878), .ZN(
        P2_U2887) );
  INV_X1 U16070 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19031) );
  NAND2_X1 U16071 ( .A1(n19890), .A2(n16228), .ZN(n12880) );
  NAND2_X1 U16072 ( .A1(n19081), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n12882) );
  INV_X1 U16073 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16330) );
  NOR2_X1 U16074 ( .A1(n19101), .A2(n16330), .ZN(n12881) );
  AOI21_X1 U16075 ( .B1(n19101), .B2(BUF2_REG_9__SCAN_IN), .A(n12881), .ZN(
        n14968) );
  INV_X1 U16076 ( .A(n14968), .ZN(n19001) );
  NAND2_X1 U16077 ( .A1(n19063), .A2(n19001), .ZN(n12891) );
  OAI211_X1 U16078 ( .C1(n19031), .C2(n12897), .A(n12882), .B(n12891), .ZN(
        P2_U2976) );
  NAND2_X1 U16079 ( .A1(n19081), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12886) );
  INV_X1 U16080 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n12883) );
  OR2_X1 U16081 ( .A1(n19101), .A2(n12883), .ZN(n12885) );
  NAND2_X1 U16082 ( .A1(n19101), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12884) );
  NAND2_X1 U16083 ( .A1(n12885), .A2(n12884), .ZN(n18993) );
  NAND2_X1 U16084 ( .A1(n19063), .A2(n18993), .ZN(n12893) );
  OAI211_X1 U16085 ( .C1(n12887), .C2(n12897), .A(n12886), .B(n12893), .ZN(
        P2_U2966) );
  NAND2_X1 U16086 ( .A1(n19081), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12889) );
  INV_X1 U16087 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16328) );
  NOR2_X1 U16088 ( .A1(n19101), .A2(n16328), .ZN(n12888) );
  AOI21_X1 U16089 ( .B1(n19101), .B2(BUF2_REG_10__SCAN_IN), .A(n12888), .ZN(
        n14959) );
  INV_X1 U16090 ( .A(n14959), .ZN(n18998) );
  NAND2_X1 U16091 ( .A1(n19063), .A2(n18998), .ZN(n12895) );
  OAI211_X1 U16092 ( .C1(n12890), .C2(n12897), .A(n12889), .B(n12895), .ZN(
        P2_U2962) );
  NAND2_X1 U16093 ( .A1(n19081), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n12892) );
  OAI211_X1 U16094 ( .C1(n12897), .C2(n14966), .A(n12892), .B(n12891), .ZN(
        P2_U2961) );
  INV_X1 U16095 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19021) );
  NAND2_X1 U16096 ( .A1(n19081), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n12894) );
  OAI211_X1 U16097 ( .C1(n19021), .C2(n12897), .A(n12894), .B(n12893), .ZN(
        P2_U2981) );
  INV_X1 U16098 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19029) );
  NAND2_X1 U16099 ( .A1(n19081), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12896) );
  OAI211_X1 U16100 ( .C1(n19029), .C2(n12897), .A(n12896), .B(n12895), .ZN(
        P2_U2977) );
  XNOR2_X1 U16101 ( .A(n13356), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19287) );
  AOI22_X1 U16102 ( .A1(n13081), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19837), .B2(n19287), .ZN(n12899) );
  INV_X1 U16103 ( .A(n12901), .ZN(n15534) );
  NAND2_X1 U16104 ( .A1(n15534), .A2(n12902), .ZN(n12903) );
  NAND2_X1 U16105 ( .A1(n12906), .A2(n12905), .ZN(n13074) );
  INV_X1 U16106 ( .A(n19281), .ZN(n19845) );
  MUX2_X1 U16107 ( .A(n14861), .B(n12908), .S(n18983), .Z(n12909) );
  OAI21_X1 U16108 ( .B1(n19845), .B2(n18984), .A(n12909), .ZN(P2_U2885) );
  NOR2_X1 U16109 ( .A1(n12910), .A2(n9846), .ZN(n12911) );
  XOR2_X1 U16110 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n12911), .Z(
        n19969) );
  NAND2_X1 U16111 ( .A1(n19969), .A2(n12912), .ZN(n13435) );
  OAI21_X1 U16112 ( .B1(n20687), .B2(n15754), .A(n12913), .ZN(n12916) );
  NAND3_X1 U16113 ( .A1(n15706), .A2(n12914), .A3(n13015), .ZN(n12915) );
  NAND2_X1 U16114 ( .A1(n12916), .A2(n12915), .ZN(n12917) );
  OR2_X1 U16115 ( .A1(n13008), .A2(n12917), .ZN(n12925) );
  INV_X1 U16116 ( .A(n12751), .ZN(n12921) );
  INV_X1 U16117 ( .A(n12918), .ZN(n12920) );
  INV_X1 U16118 ( .A(n12945), .ZN(n12919) );
  AOI21_X1 U16119 ( .B1(n12921), .B2(n12920), .A(n12919), .ZN(n13010) );
  NAND2_X1 U16120 ( .A1(n13630), .A2(n10211), .ZN(n12922) );
  AND3_X1 U16121 ( .A1(n13010), .A2(n12923), .A3(n12922), .ZN(n12924) );
  INV_X1 U16122 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19909) );
  NAND2_X1 U16123 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16008), .ZN(n16009) );
  OAI22_X1 U16124 ( .A1(n13434), .A2(n19901), .B1(n19909), .B2(n16009), .ZN(
        n12927) );
  NAND2_X1 U16125 ( .A1(n12994), .A2(n12927), .ZN(n12928) );
  NOR2_X1 U16126 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20510), .ZN(n20097) );
  NOR2_X1 U16127 ( .A1(n20097), .A2(n12927), .ZN(n12995) );
  INV_X1 U16128 ( .A(n12995), .ZN(n14702) );
  OAI22_X1 U16129 ( .A1(n13435), .A2(n12928), .B1(n13438), .B2(n14702), .ZN(
        P1_U3468) );
  NOR2_X1 U16130 ( .A1(n12751), .A2(n9616), .ZN(n12929) );
  INV_X1 U16131 ( .A(n16008), .ZN(n13450) );
  NOR2_X1 U16132 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13450), .ZN(n20769) );
  INV_X2 U16133 ( .A(n20769), .ZN(n20011) );
  INV_X1 U16134 ( .A(n13238), .ZN(n20008) );
  AOI222_X1 U16135 ( .A1(n20009), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n20008), 
        .B2(P1_EAX_REG_4__SCAN_IN), .C1(n20769), .C2(P1_LWORD_REG_4__SCAN_IN), 
        .ZN(n12931) );
  INV_X1 U16136 ( .A(n12931), .ZN(P1_U2932) );
  NOR2_X1 U16137 ( .A1(n19861), .A2(n12932), .ZN(n12936) );
  XNOR2_X1 U16138 ( .A(n12934), .B(n12933), .ZN(n19855) );
  INV_X1 U16139 ( .A(n19855), .ZN(n18926) );
  NAND2_X1 U16140 ( .A1(n19280), .A2(n18926), .ZN(n13060) );
  OAI21_X1 U16141 ( .B1(n19280), .B2(n18926), .A(n13060), .ZN(n12935) );
  NOR2_X1 U16142 ( .A1(n12935), .A2(n12936), .ZN(n13062) );
  AOI21_X1 U16143 ( .B1(n12936), .B2(n12935), .A(n13062), .ZN(n12940) );
  AOI22_X1 U16144 ( .A1(n19103), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19101), .ZN(n19121) );
  INV_X1 U16145 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n12937) );
  OAI22_X1 U16146 ( .A1(n13614), .A2(n19121), .B1(n14979), .B2(n12937), .ZN(
        n12938) );
  AOI21_X1 U16147 ( .B1(n18989), .B2(n19855), .A(n12938), .ZN(n12939) );
  OAI21_X1 U16148 ( .B1(n12940), .B2(n14996), .A(n12939), .ZN(P2_U2918) );
  NAND2_X1 U16149 ( .A1(n12941), .A2(n10242), .ZN(n12942) );
  NAND2_X1 U16150 ( .A1(n12942), .A2(n10222), .ZN(n12943) );
  AND3_X1 U16151 ( .A1(n12945), .A2(n12944), .A3(n12943), .ZN(n13032) );
  INV_X1 U16152 ( .A(n12367), .ZN(n12946) );
  NAND2_X1 U16153 ( .A1(n12946), .A2(n12914), .ZN(n12950) );
  NAND2_X1 U16154 ( .A1(n10246), .A2(n12947), .ZN(n12949) );
  AND2_X1 U16155 ( .A1(n10218), .A2(n13630), .ZN(n12948) );
  OR2_X1 U16156 ( .A1(n12949), .A2(n12948), .ZN(n13029) );
  NOR2_X1 U16157 ( .A1(n12950), .A2(n13029), .ZN(n12951) );
  NAND3_X1 U16158 ( .A1(n12359), .A2(n13032), .A3(n12951), .ZN(n14694) );
  INV_X1 U16159 ( .A(n14692), .ZN(n13007) );
  AOI22_X1 U16160 ( .A1(n13631), .A2(n14694), .B1(n13007), .B2(n9875), .ZN(
        n15705) );
  INV_X1 U16161 ( .A(n12994), .ZN(n14701) );
  INV_X1 U16162 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20058) );
  AOI22_X1 U16163 ( .A1(n15739), .A2(n9875), .B1(n20058), .B2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n12952) );
  OAI21_X1 U16164 ( .B1(n15705), .B2(n14701), .A(n12952), .ZN(n12954) );
  OAI21_X1 U16165 ( .B1(n15706), .B2(n14701), .A(n14702), .ZN(n12953) );
  AOI22_X1 U16166 ( .A1(n12954), .A2(n14702), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n12953), .ZN(n12955) );
  INV_X1 U16167 ( .A(n12955), .ZN(P1_U3474) );
  INV_X1 U16168 ( .A(n12956), .ZN(n12960) );
  INV_X1 U16169 ( .A(n12957), .ZN(n12959) );
  OAI21_X1 U16170 ( .B1(n12960), .B2(n12959), .A(n12958), .ZN(n13615) );
  NAND2_X1 U16171 ( .A1(n12961), .A2(n10229), .ZN(n12962) );
  INV_X1 U16172 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n13181) );
  INV_X1 U16173 ( .A(n12962), .ZN(n12963) );
  INV_X1 U16174 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16348) );
  NAND2_X1 U16175 ( .A1(n20091), .A2(n16348), .ZN(n12964) );
  OAI21_X1 U16176 ( .B1(n20091), .B2(DATAI_0_), .A(n12964), .ZN(n20105) );
  OAI222_X1 U16177 ( .A1(n13615), .A2(n14370), .B1(n14365), .B2(n13181), .C1(
        n14364), .C2(n20105), .ZN(P1_U2904) );
  INV_X1 U16178 ( .A(n12965), .ZN(n20103) );
  XNOR2_X1 U16179 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12974) );
  NAND2_X1 U16180 ( .A1(n13015), .A2(n12966), .ZN(n12984) );
  INV_X1 U16181 ( .A(n12967), .ZN(n12969) );
  INV_X1 U16182 ( .A(n12968), .ZN(n14690) );
  NAND2_X1 U16183 ( .A1(n14690), .A2(n10059), .ZN(n12982) );
  NAND2_X1 U16184 ( .A1(n12969), .A2(n12982), .ZN(n12971) );
  NAND2_X1 U16185 ( .A1(n12984), .A2(n12971), .ZN(n12973) );
  NOR2_X1 U16186 ( .A1(n12970), .A2(n10242), .ZN(n12986) );
  INV_X1 U16187 ( .A(n12971), .ZN(n12976) );
  NAND3_X1 U16188 ( .A1(n13007), .A2(n12986), .A3(n12976), .ZN(n12972) );
  OAI211_X1 U16189 ( .C1(n12974), .C2(n15706), .A(n12973), .B(n12972), .ZN(
        n12975) );
  AOI21_X1 U16190 ( .B1(n20103), .B2(n14694), .A(n12975), .ZN(n13442) );
  INV_X1 U16191 ( .A(n13442), .ZN(n12977) );
  NOR2_X1 U16192 ( .A1(n15734), .A2(n20058), .ZN(n14698) );
  AOI22_X1 U16193 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20086), .B2(n14374), .ZN(
        n14696) );
  AOI222_X1 U16194 ( .A1(n12977), .A2(n12994), .B1(n14698), .B2(n14696), .C1(
        n12976), .C2(n15739), .ZN(n12979) );
  NAND2_X1 U16195 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n12995), .ZN(
        n12978) );
  OAI21_X1 U16196 ( .B1(n12979), .B2(n12995), .A(n12978), .ZN(P1_U3472) );
  NAND2_X1 U16197 ( .A1(n9603), .A2(n14694), .ZN(n12992) );
  XNOR2_X1 U16198 ( .A(n12981), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12989) );
  XNOR2_X1 U16199 ( .A(n12982), .B(n12996), .ZN(n12983) );
  NAND2_X1 U16200 ( .A1(n12984), .A2(n12983), .ZN(n12988) );
  NOR2_X1 U16201 ( .A1(n12967), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12985) );
  NOR2_X1 U16202 ( .A1(n9623), .A2(n12985), .ZN(n12993) );
  NAND3_X1 U16203 ( .A1(n13007), .A2(n12986), .A3(n12993), .ZN(n12987) );
  OAI211_X1 U16204 ( .C1(n12989), .C2(n15706), .A(n12988), .B(n12987), .ZN(
        n12990) );
  INV_X1 U16205 ( .A(n12990), .ZN(n12991) );
  NAND2_X1 U16206 ( .A1(n12992), .A2(n12991), .ZN(n13440) );
  AOI22_X1 U16207 ( .A1(n13440), .A2(n12994), .B1(n12993), .B2(n15739), .ZN(
        n12997) );
  MUX2_X1 U16208 ( .A(n12997), .B(n12996), .S(n12995), .Z(n12998) );
  INV_X1 U16209 ( .A(n12998), .ZN(P1_U3469) );
  XOR2_X1 U16210 ( .A(n13000), .B(n12999), .Z(n15530) );
  INV_X1 U16211 ( .A(n15530), .ZN(n18886) );
  AND2_X1 U16212 ( .A1(n14996), .A2(n20787), .ZN(n19012) );
  OAI22_X1 U16213 ( .A1(n19101), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19103), .ZN(n19152) );
  INV_X1 U16214 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19037) );
  OAI222_X1 U16215 ( .A1(n18886), .A2(n19012), .B1(n13614), .B2(n19152), .C1(
        n19037), .C2(n14979), .ZN(P2_U2913) );
  OAI21_X1 U16216 ( .B1(n13001), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n11082), .ZN(n13098) );
  OAI21_X1 U16217 ( .B1(n9616), .B2(n15732), .A(n13002), .ZN(n13006) );
  OAI21_X1 U16218 ( .B1(n10222), .B2(n15732), .A(n20768), .ZN(n13627) );
  OAI211_X1 U16219 ( .C1(n12914), .C2(n13627), .A(n10224), .B(n10207), .ZN(
        n13003) );
  INV_X1 U16220 ( .A(n13003), .ZN(n13004) );
  OR2_X1 U16221 ( .A1(n13008), .A2(n13004), .ZN(n13005) );
  MUX2_X1 U16222 ( .A(n13006), .B(n13005), .S(n10211), .Z(n13011) );
  NAND3_X1 U16223 ( .A1(n13008), .A2(n13007), .A3(n10222), .ZN(n13009) );
  NAND3_X1 U16224 ( .A1(n13011), .A2(n13010), .A3(n13009), .ZN(n13013) );
  OAI211_X1 U16225 ( .C1(n13016), .C2(n13014), .A(n15724), .B(n13015), .ZN(
        n13017) );
  OR2_X1 U16226 ( .A1(n13018), .A2(n13017), .ZN(n13019) );
  OAI22_X1 U16227 ( .A1(n20127), .A2(n13014), .B1(n12753), .B2(n10222), .ZN(
        n13020) );
  OR2_X1 U16228 ( .A1(n14090), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13021) );
  NAND2_X1 U16229 ( .A1(n13022), .A2(n13021), .ZN(n13634) );
  INV_X1 U16230 ( .A(n13634), .ZN(n13027) );
  INV_X1 U16231 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13023) );
  NOR2_X1 U16232 ( .A1(n20065), .A2(n13023), .ZN(n13100) );
  INV_X1 U16233 ( .A(n13034), .ZN(n13024) );
  INV_X1 U16234 ( .A(n13722), .ZN(n13025) );
  NAND2_X1 U16235 ( .A1(n20065), .A2(n13024), .ZN(n20085) );
  AOI21_X1 U16236 ( .B1(n13025), .B2(n20085), .A(n20058), .ZN(n13026) );
  AOI211_X1 U16237 ( .C1(n20048), .C2(n13027), .A(n13100), .B(n13026), .ZN(
        n13035) );
  INV_X1 U16238 ( .A(n20057), .ZN(n13729) );
  OAI21_X1 U16239 ( .B1(n10223), .B2(n10221), .A(n13029), .ZN(n13030) );
  NAND3_X1 U16240 ( .A1(n13032), .A2(n13031), .A3(n13030), .ZN(n13033) );
  NAND2_X1 U16241 ( .A1(n13034), .A2(n13033), .ZN(n13728) );
  OAI21_X1 U16242 ( .B1(n13729), .B2(n13721), .A(n20058), .ZN(n20084) );
  OAI211_X1 U16243 ( .C1(n13098), .C2(n20073), .A(n13035), .B(n20084), .ZN(
        P1_U3031) );
  AOI22_X1 U16244 ( .A1(n19103), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19101), .ZN(n19161) );
  OAI21_X1 U16245 ( .B1(n13038), .B2(n13037), .A(n13036), .ZN(n18875) );
  OAI222_X1 U16246 ( .A1(n13614), .A2(n19161), .B1(n18875), .B2(n19012), .C1(
        n19035), .C2(n14979), .ZN(P2_U2912) );
  NAND2_X1 U16247 ( .A1(n13040), .A2(n13039), .ZN(n13042) );
  NAND2_X1 U16248 ( .A1(n13042), .A2(n9736), .ZN(n19847) );
  INV_X1 U16249 ( .A(n19847), .ZN(n13063) );
  INV_X1 U16250 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19777) );
  OAI22_X1 U16251 ( .A1(n13044), .A2(n16222), .B1(n16227), .B2(n13043), .ZN(
        n13045) );
  INV_X1 U16252 ( .A(n13045), .ZN(n13050) );
  INV_X1 U16253 ( .A(n15381), .ZN(n13046) );
  OAI21_X1 U16254 ( .B1(n13048), .B2(n13047), .A(n13046), .ZN(n13049) );
  OAI211_X1 U16255 ( .C1(n13051), .C2(n19777), .A(n13050), .B(n13049), .ZN(
        n13052) );
  INV_X1 U16256 ( .A(n13052), .ZN(n13059) );
  NOR2_X1 U16257 ( .A1(n15379), .A2(n13091), .ZN(n13054) );
  MUX2_X1 U16258 ( .A(n13055), .B(n13054), .S(n13053), .Z(n13056) );
  AOI21_X1 U16259 ( .B1(n16218), .B2(n13057), .A(n13056), .ZN(n13058) );
  OAI211_X1 U16260 ( .C1(n13063), .C2(n16204), .A(n13059), .B(n13058), .ZN(
        P2_U3044) );
  INV_X1 U16261 ( .A(n13060), .ZN(n13061) );
  NOR2_X1 U16262 ( .A1(n13062), .A2(n13061), .ZN(n13065) );
  NAND2_X1 U16263 ( .A1(n19845), .A2(n13063), .ZN(n13244) );
  OAI21_X1 U16264 ( .B1(n19845), .B2(n13063), .A(n13244), .ZN(n13064) );
  NOR2_X1 U16265 ( .A1(n13064), .A2(n13065), .ZN(n13246) );
  AOI21_X1 U16266 ( .B1(n13065), .B2(n13064), .A(n13246), .ZN(n13068) );
  INV_X1 U16267 ( .A(n13614), .ZN(n19005) );
  INV_X1 U16268 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16342) );
  INV_X1 U16269 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18071) );
  AOI22_X1 U16270 ( .A1(n19103), .A2(n16342), .B1(n18071), .B2(n19101), .ZN(
        n19126) );
  AOI22_X1 U16271 ( .A1(n19005), .A2(n19126), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n20780), .ZN(n13067) );
  NAND2_X1 U16272 ( .A1(n19847), .A2(n18989), .ZN(n13066) );
  OAI211_X1 U16273 ( .C1(n13068), .C2(n14996), .A(n13067), .B(n13066), .ZN(
        P2_U2917) );
  INV_X1 U16274 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13069) );
  OAI222_X1 U16275 ( .A1(n13634), .A2(n14298), .B1(n13069), .B2(n20003), .C1(
        n13615), .C2(n14297), .ZN(P1_U2872) );
  INV_X1 U16276 ( .A(n13070), .ZN(n13071) );
  NAND2_X1 U16277 ( .A1(n13072), .A2(n13071), .ZN(n13073) );
  INV_X1 U16278 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13075) );
  NOR2_X1 U16279 ( .A1(n13958), .A2(n13075), .ZN(n13084) );
  NAND2_X1 U16280 ( .A1(n13077), .A2(n13076), .ZN(n13083) );
  NAND2_X1 U16281 ( .A1(n19842), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19356) );
  INV_X1 U16282 ( .A(n19356), .ZN(n13078) );
  NAND2_X1 U16283 ( .A1(n19519), .A2(n13078), .ZN(n19423) );
  NOR2_X1 U16284 ( .A1(n19842), .A2(n20880), .ZN(n19589) );
  NAND2_X1 U16285 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19589), .ZN(
        n19693) );
  NOR2_X2 U16286 ( .A1(n19865), .A2(n19693), .ZN(n19739) );
  INV_X1 U16287 ( .A(n19739), .ZN(n13079) );
  NAND2_X1 U16288 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13079), .ZN(
        n13080) );
  NAND2_X1 U16289 ( .A1(n19423), .A2(n13080), .ZN(n19559) );
  AOI21_X1 U16290 ( .B1(n13081), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19554), .ZN(n13082) );
  NAND2_X1 U16291 ( .A1(n13142), .A2(n13084), .ZN(n13406) );
  OAI21_X1 U16292 ( .B1(n13084), .B2(n13142), .A(n13406), .ZN(n13085) );
  INV_X1 U16293 ( .A(n13085), .ZN(n13138) );
  INV_X1 U16294 ( .A(n19450), .ZN(n19839) );
  MUX2_X1 U16295 ( .A(n14847), .B(P2_EBX_REG_3__SCAN_IN), .S(n18983), .Z(
        n13086) );
  AOI21_X1 U16296 ( .B1(n19839), .B2(n18954), .A(n13086), .ZN(n13087) );
  INV_X1 U16297 ( .A(n13087), .ZN(P2_U2884) );
  NOR2_X1 U16298 ( .A1(n16215), .A2(n15541), .ZN(n13088) );
  AOI211_X1 U16299 ( .C1(n13090), .C2(n16192), .A(n13089), .B(n13088), .ZN(
        n13093) );
  OAI211_X1 U16300 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15523), .B(n13091), .ZN(n13092) );
  OAI211_X1 U16301 ( .C1(n13355), .C2(n15521), .A(n13093), .B(n13092), .ZN(
        n13094) );
  AOI21_X1 U16302 ( .B1(n16217), .B2(n19855), .A(n13094), .ZN(n13095) );
  OAI21_X1 U16303 ( .B1(n13096), .B2(n16222), .A(n13095), .ZN(P2_U3045) );
  NAND2_X1 U16304 ( .A1(n13097), .A2(n14484), .ZN(n13101) );
  NOR2_X1 U16305 ( .A1(n13098), .A2(n19908), .ZN(n13099) );
  AOI211_X1 U16306 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n13101), .A(
        n13100), .B(n13099), .ZN(n13102) );
  OAI21_X1 U16307 ( .B1(n20090), .B2(n13615), .A(n13102), .ZN(P1_U2999) );
  OAI21_X1 U16308 ( .B1(n13104), .B2(n13103), .A(n13463), .ZN(n13655) );
  OR2_X1 U16309 ( .A1(n13106), .A2(n13105), .ZN(n13108) );
  AND2_X1 U16310 ( .A1(n13108), .A2(n13107), .ZN(n20080) );
  INV_X1 U16311 ( .A(n20080), .ZN(n13109) );
  AOI22_X1 U16312 ( .A1(n12418), .A2(n13109), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14288), .ZN(n13110) );
  OAI21_X1 U16313 ( .B1(n13655), .B2(n14290), .A(n13110), .ZN(P1_U2871) );
  INV_X1 U16314 ( .A(n13354), .ZN(n13111) );
  NAND2_X1 U16315 ( .A1(n14847), .A2(n13111), .ZN(n13126) );
  NAND2_X1 U16316 ( .A1(n13112), .A2(n11459), .ZN(n13337) );
  INV_X1 U16317 ( .A(n13113), .ZN(n13114) );
  OAI21_X1 U16318 ( .B1(n11408), .B2(n13115), .A(n13114), .ZN(n13124) );
  INV_X1 U16319 ( .A(n13378), .ZN(n13116) );
  NAND2_X1 U16320 ( .A1(n13117), .A2(n13116), .ZN(n13335) );
  NOR2_X1 U16321 ( .A1(n13118), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13331) );
  XNOR2_X1 U16322 ( .A(n13331), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13119) );
  NAND2_X1 U16323 ( .A1(n13335), .A2(n13119), .ZN(n13122) );
  XNOR2_X1 U16324 ( .A(n11531), .B(n11530), .ZN(n13120) );
  NAND2_X1 U16325 ( .A1(n13350), .A2(n13120), .ZN(n13121) );
  NAND2_X1 U16326 ( .A1(n13122), .A2(n13121), .ZN(n13123) );
  AOI21_X1 U16327 ( .B1(n13337), .B2(n13124), .A(n13123), .ZN(n13125) );
  NAND2_X1 U16328 ( .A1(n13126), .A2(n13125), .ZN(n13360) );
  AOI22_X1 U16329 ( .A1(n19839), .A2(n10024), .B1(n19833), .B2(n13360), .ZN(
        n13136) );
  NAND2_X1 U16330 ( .A1(n13127), .A2(n15665), .ZN(n13132) );
  AND2_X1 U16331 ( .A1(n13129), .A2(n13128), .ZN(n13130) );
  NAND2_X1 U16332 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13133), .ZN(n15758) );
  INV_X1 U16333 ( .A(n15758), .ZN(n16231) );
  NAND2_X1 U16334 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(n16231), .ZN(n15757) );
  OAI211_X1 U16335 ( .C1(n13367), .C2(n16236), .A(n13134), .B(n15757), .ZN(
        n15669) );
  NAND2_X1 U16336 ( .A1(n15552), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13135) );
  OAI21_X1 U16337 ( .B1(n13136), .B2(n15552), .A(n13135), .ZN(P2_U3596) );
  NAND2_X1 U16338 ( .A1(n13138), .A2(n13137), .ZN(n13141) );
  NAND2_X1 U16339 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13139), .ZN(
        n13140) );
  AND2_X1 U16340 ( .A1(n13142), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13144) );
  INV_X1 U16341 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13143) );
  NOR2_X1 U16342 ( .A1(n13958), .A2(n13143), .ZN(n13407) );
  XOR2_X1 U16343 ( .A(n13159), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13149)
         );
  INV_X1 U16344 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n18905) );
  AND2_X1 U16345 ( .A1(n13572), .A2(n13146), .ZN(n13147) );
  NOR2_X1 U16346 ( .A1(n13145), .A2(n13147), .ZN(n13604) );
  INV_X1 U16347 ( .A(n13604), .ZN(n18899) );
  MUX2_X1 U16348 ( .A(n18905), .B(n18899), .S(n18988), .Z(n13148) );
  OAI21_X1 U16349 ( .B1(n13149), .B2(n18984), .A(n13148), .ZN(P2_U2882) );
  INV_X1 U16350 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13649) );
  INV_X1 U16351 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n14227) );
  OR2_X1 U16352 ( .A1(n20065), .A2(n14227), .ZN(n20077) );
  OAI21_X1 U16353 ( .B1(n14484), .B2(n13649), .A(n20077), .ZN(n13150) );
  AOI21_X1 U16354 ( .B1(n15889), .B2(n13649), .A(n13150), .ZN(n13155) );
  NOR2_X1 U16355 ( .A1(n9596), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20074) );
  INV_X1 U16356 ( .A(n20074), .ZN(n13153) );
  NAND3_X1 U16357 ( .A1(n13153), .A2(n20032), .A3(n13152), .ZN(n13154) );
  OAI211_X1 U16358 ( .C1(n13655), .C2(n20090), .A(n13155), .B(n13154), .ZN(
        P1_U2998) );
  AOI22_X1 U16359 ( .A1(n19103), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n19101), .ZN(n19076) );
  AOI21_X1 U16360 ( .B1(n13157), .B2(n13036), .A(n15506), .ZN(n18863) );
  INV_X1 U16361 ( .A(n18863), .ZN(n13158) );
  INV_X1 U16362 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19033) );
  OAI222_X1 U16363 ( .A1(n13614), .A2(n19076), .B1(n13158), .B2(n19012), .C1(
        n19033), .C2(n14979), .ZN(P2_U2911) );
  XNOR2_X1 U16364 ( .A(n13398), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13165) );
  NAND2_X1 U16365 ( .A1(n13160), .A2(n13167), .ZN(n13163) );
  INV_X1 U16366 ( .A(n13161), .ZN(n13162) );
  NAND2_X1 U16367 ( .A1(n13163), .A2(n13162), .ZN(n18874) );
  MUX2_X1 U16368 ( .A(n11738), .B(n18874), .S(n18988), .Z(n13164) );
  OAI21_X1 U16369 ( .B1(n13165), .B2(n18984), .A(n13164), .ZN(P2_U2880) );
  OR2_X1 U16370 ( .A1(n13145), .A2(n13166), .ZN(n13168) );
  NAND2_X1 U16371 ( .A1(n13168), .A2(n13167), .ZN(n18885) );
  NOR2_X1 U16372 ( .A1(n13159), .A2(n13829), .ZN(n13170) );
  INV_X1 U16373 ( .A(n13398), .ZN(n13169) );
  OAI211_X1 U16374 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13170), .A(
        n13169), .B(n18954), .ZN(n13172) );
  NAND2_X1 U16375 ( .A1(n18983), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13171) );
  OAI211_X1 U16376 ( .C1(n18885), .C2(n18983), .A(n13172), .B(n13171), .ZN(
        P2_U2881) );
  INV_X1 U16377 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n13174) );
  INV_X1 U16378 ( .A(P1_LWORD_REG_5__SCAN_IN), .ZN(n13173) );
  OAI222_X1 U16379 ( .A1(n13174), .A2(n20007), .B1(n13238), .B2(n13289), .C1(
        n13173), .C2(n20011), .ZN(P1_U2931) );
  INV_X1 U16380 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n13176) );
  INV_X1 U16381 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n13187) );
  INV_X1 U16382 ( .A(P1_LWORD_REG_1__SCAN_IN), .ZN(n13175) );
  OAI222_X1 U16383 ( .A1(n13176), .A2(n20007), .B1(n13238), .B2(n13187), .C1(
        n13175), .C2(n20011), .ZN(P1_U2935) );
  INV_X1 U16384 ( .A(P1_LWORD_REG_7__SCAN_IN), .ZN(n13177) );
  OAI222_X1 U16385 ( .A1(n20902), .A2(n20007), .B1(n13238), .B2(n13297), .C1(
        n13177), .C2(n20011), .ZN(P1_U2929) );
  INV_X1 U16386 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n13179) );
  INV_X1 U16387 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20865) );
  INV_X1 U16388 ( .A(P1_LWORD_REG_3__SCAN_IN), .ZN(n13178) );
  OAI222_X1 U16389 ( .A1(n13179), .A2(n20007), .B1(n13238), .B2(n20865), .C1(
        n13178), .C2(n20011), .ZN(P1_U2933) );
  INV_X1 U16390 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n13182) );
  INV_X1 U16391 ( .A(P1_LWORD_REG_0__SCAN_IN), .ZN(n13180) );
  OAI222_X1 U16392 ( .A1(n13182), .A2(n20007), .B1(n13238), .B2(n13181), .C1(
        n13180), .C2(n20011), .ZN(P1_U2936) );
  INV_X1 U16393 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n13184) );
  INV_X1 U16394 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n13502) );
  INV_X1 U16395 ( .A(P1_LWORD_REG_2__SCAN_IN), .ZN(n13183) );
  OAI222_X1 U16396 ( .A1(n13184), .A2(n20007), .B1(n13238), .B2(n13502), .C1(
        n13183), .C2(n20011), .ZN(P1_U2934) );
  NAND2_X1 U16397 ( .A1(n20089), .A2(DATAI_1_), .ZN(n13186) );
  NAND2_X1 U16398 ( .A1(n20091), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13185) );
  OAI222_X1 U16399 ( .A1(n14370), .A2(n13655), .B1(n14365), .B2(n13187), .C1(
        n14364), .C2(n20114), .ZN(P1_U2903) );
  INV_X1 U16400 ( .A(P1_UWORD_REG_5__SCAN_IN), .ZN(n13190) );
  NOR2_X1 U16401 ( .A1(n13238), .A2(n10223), .ZN(n20004) );
  INV_X1 U16402 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13189) );
  INV_X1 U16403 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n13188) );
  OAI222_X1 U16404 ( .A1(n13190), .A2(n20011), .B1(n13235), .B2(n13189), .C1(
        n20007), .C2(n13188), .ZN(P1_U2915) );
  INV_X1 U16405 ( .A(P1_UWORD_REG_8__SCAN_IN), .ZN(n13192) );
  INV_X1 U16406 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13313) );
  INV_X1 U16407 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13191) );
  OAI222_X1 U16408 ( .A1(n13192), .A2(n20011), .B1(n13235), .B2(n13313), .C1(
        n20007), .C2(n13191), .ZN(P1_U2912) );
  INV_X1 U16409 ( .A(P1_UWORD_REG_11__SCAN_IN), .ZN(n13194) );
  INV_X1 U16410 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13324) );
  INV_X1 U16411 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13193) );
  OAI222_X1 U16412 ( .A1(n13194), .A2(n20011), .B1(n13235), .B2(n13324), .C1(
        n20007), .C2(n13193), .ZN(P1_U2909) );
  INV_X1 U16413 ( .A(P1_UWORD_REG_6__SCAN_IN), .ZN(n13197) );
  INV_X1 U16414 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13196) );
  INV_X1 U16415 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n13195) );
  OAI222_X1 U16416 ( .A1(n13197), .A2(n20011), .B1(n13235), .B2(n13196), .C1(
        n20007), .C2(n13195), .ZN(P1_U2914) );
  INV_X1 U16417 ( .A(P1_UWORD_REG_14__SCAN_IN), .ZN(n13199) );
  INV_X1 U16418 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13317) );
  INV_X1 U16419 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13198) );
  OAI222_X1 U16420 ( .A1(n13199), .A2(n20011), .B1(n13235), .B2(n13317), .C1(
        n20007), .C2(n13198), .ZN(P1_U2906) );
  INV_X1 U16421 ( .A(P1_UWORD_REG_4__SCAN_IN), .ZN(n13202) );
  INV_X1 U16422 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13201) );
  INV_X1 U16423 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n13200) );
  OAI222_X1 U16424 ( .A1(n13202), .A2(n20011), .B1(n13235), .B2(n13201), .C1(
        n20007), .C2(n13200), .ZN(P1_U2916) );
  INV_X1 U16425 ( .A(P1_UWORD_REG_3__SCAN_IN), .ZN(n13205) );
  INV_X1 U16426 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13204) );
  INV_X1 U16427 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n13203) );
  OAI222_X1 U16428 ( .A1(n13205), .A2(n20011), .B1(n13235), .B2(n13204), .C1(
        n20007), .C2(n13203), .ZN(P1_U2917) );
  INV_X1 U16429 ( .A(P1_UWORD_REG_2__SCAN_IN), .ZN(n13208) );
  INV_X1 U16430 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13207) );
  INV_X1 U16431 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n13206) );
  OAI222_X1 U16432 ( .A1(n13208), .A2(n20011), .B1(n13235), .B2(n13207), .C1(
        n20007), .C2(n13206), .ZN(P1_U2918) );
  INV_X1 U16433 ( .A(P1_UWORD_REG_1__SCAN_IN), .ZN(n13211) );
  INV_X1 U16434 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13210) );
  INV_X1 U16435 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n13209) );
  OAI222_X1 U16436 ( .A1(n13211), .A2(n20011), .B1(n13235), .B2(n13210), .C1(
        n20007), .C2(n13209), .ZN(P1_U2919) );
  INV_X1 U16437 ( .A(P1_UWORD_REG_12__SCAN_IN), .ZN(n13213) );
  INV_X1 U16438 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13260) );
  INV_X1 U16439 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13212) );
  OAI222_X1 U16440 ( .A1(n13213), .A2(n20011), .B1(n13235), .B2(n13260), .C1(
        n20007), .C2(n13212), .ZN(P1_U2908) );
  INV_X1 U16441 ( .A(P1_LWORD_REG_14__SCAN_IN), .ZN(n13215) );
  INV_X1 U16442 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n13320) );
  INV_X1 U16443 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n13214) );
  OAI222_X1 U16444 ( .A1(n13215), .A2(n20011), .B1(n13238), .B2(n13320), .C1(
        n20007), .C2(n13214), .ZN(P1_U2922) );
  INV_X1 U16445 ( .A(P1_UWORD_REG_10__SCAN_IN), .ZN(n13217) );
  INV_X1 U16446 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13263) );
  INV_X1 U16447 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13216) );
  OAI222_X1 U16448 ( .A1(n13217), .A2(n20011), .B1(n13235), .B2(n13263), .C1(
        n20007), .C2(n13216), .ZN(P1_U2910) );
  INV_X1 U16449 ( .A(P1_LWORD_REG_12__SCAN_IN), .ZN(n13219) );
  INV_X1 U16450 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n13282) );
  INV_X1 U16451 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n13218) );
  OAI222_X1 U16452 ( .A1(n13219), .A2(n20011), .B1(n13238), .B2(n13282), .C1(
        n20007), .C2(n13218), .ZN(P1_U2924) );
  INV_X1 U16453 ( .A(P1_LWORD_REG_11__SCAN_IN), .ZN(n13221) );
  INV_X1 U16454 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n13327) );
  INV_X1 U16455 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n13220) );
  OAI222_X1 U16456 ( .A1(n13221), .A2(n20011), .B1(n13238), .B2(n13327), .C1(
        n20007), .C2(n13220), .ZN(P1_U2925) );
  INV_X1 U16457 ( .A(P1_LWORD_REG_10__SCAN_IN), .ZN(n13223) );
  INV_X1 U16458 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13303) );
  INV_X1 U16459 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n13222) );
  OAI222_X1 U16460 ( .A1(n13223), .A2(n20011), .B1(n13238), .B2(n13303), .C1(
        n20007), .C2(n13222), .ZN(P1_U2926) );
  INV_X1 U16461 ( .A(P1_UWORD_REG_9__SCAN_IN), .ZN(n13225) );
  INV_X1 U16462 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13294) );
  INV_X1 U16463 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13224) );
  OAI222_X1 U16464 ( .A1(n13225), .A2(n20011), .B1(n13235), .B2(n13294), .C1(
        n20007), .C2(n13224), .ZN(P1_U2911) );
  INV_X1 U16465 ( .A(P1_LWORD_REG_8__SCAN_IN), .ZN(n13227) );
  INV_X1 U16466 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13330) );
  INV_X1 U16467 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n13226) );
  OAI222_X1 U16468 ( .A1(n13227), .A2(n20011), .B1(n13238), .B2(n13330), .C1(
        n20007), .C2(n13226), .ZN(P1_U2928) );
  INV_X1 U16469 ( .A(P1_UWORD_REG_7__SCAN_IN), .ZN(n13230) );
  INV_X1 U16470 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13229) );
  INV_X1 U16471 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n13228) );
  OAI222_X1 U16472 ( .A1(n13230), .A2(n20011), .B1(n13235), .B2(n13229), .C1(
        n20007), .C2(n13228), .ZN(P1_U2913) );
  INV_X1 U16473 ( .A(P1_LWORD_REG_6__SCAN_IN), .ZN(n13232) );
  INV_X1 U16474 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n13231) );
  OAI222_X1 U16475 ( .A1(n13232), .A2(n20011), .B1(n13238), .B2(n13584), .C1(
        n20007), .C2(n13231), .ZN(P1_U2930) );
  INV_X1 U16476 ( .A(P1_UWORD_REG_0__SCAN_IN), .ZN(n13236) );
  INV_X1 U16477 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13234) );
  INV_X1 U16478 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n13233) );
  OAI222_X1 U16479 ( .A1(n13236), .A2(n20011), .B1(n13235), .B2(n13234), .C1(
        n20007), .C2(n13233), .ZN(P1_U2920) );
  INV_X1 U16480 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13239) );
  INV_X1 U16481 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14359) );
  INV_X1 U16482 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n13237) );
  OAI222_X1 U16483 ( .A1(n13239), .A2(n20011), .B1(n13238), .B2(n14359), .C1(
        n13237), .C2(n20007), .ZN(P1_U2921) );
  OR2_X1 U16484 ( .A1(n13241), .A2(n13240), .ZN(n13243) );
  NAND2_X1 U16485 ( .A1(n13243), .A2(n13242), .ZN(n14849) );
  XNOR2_X1 U16486 ( .A(n19450), .B(n14849), .ZN(n13248) );
  INV_X1 U16487 ( .A(n13244), .ZN(n13245) );
  NOR2_X1 U16488 ( .A1(n13246), .A2(n13245), .ZN(n13247) );
  NOR2_X1 U16489 ( .A1(n13247), .A2(n13248), .ZN(n13416) );
  AOI21_X1 U16490 ( .B1(n13248), .B2(n13247), .A(n13416), .ZN(n13251) );
  AOI22_X1 U16491 ( .A1(n19103), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19101), .ZN(n19133) );
  INV_X1 U16492 ( .A(n19133), .ZN(n20781) );
  AOI22_X1 U16493 ( .A1(n19005), .A2(n20781), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n20780), .ZN(n13250) );
  INV_X1 U16494 ( .A(n14849), .ZN(n19838) );
  NAND2_X1 U16495 ( .A1(n19838), .A2(n18989), .ZN(n13249) );
  OAI211_X1 U16496 ( .C1(n13251), .C2(n14996), .A(n13250), .B(n13249), .ZN(
        P2_U2916) );
  NOR2_X1 U16497 ( .A1(n13252), .A2(n20768), .ZN(n13253) );
  OR2_X2 U16498 ( .A1(n13254), .A2(n13253), .ZN(n20020) );
  NOR2_X1 U16499 ( .A1(n20020), .A2(n10222), .ZN(n20021) );
  NAND2_X1 U16500 ( .A1(n20089), .A2(DATAI_3_), .ZN(n13256) );
  NAND2_X1 U16501 ( .A1(n20091), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13255) );
  AND2_X1 U16502 ( .A1(n13256), .A2(n13255), .ZN(n20124) );
  NOR2_X1 U16503 ( .A1(n13396), .A2(n20124), .ZN(n13283) );
  AOI21_X1 U16504 ( .B1(P1_UWORD_REG_3__SCAN_IN), .B2(n20020), .A(n13283), 
        .ZN(n13257) );
  OAI21_X1 U16505 ( .B1(n13204), .B2(n13397), .A(n13257), .ZN(P1_U2940) );
  INV_X1 U16506 ( .A(DATAI_12_), .ZN(n13258) );
  INV_X1 U16507 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16325) );
  MUX2_X1 U16508 ( .A(n13258), .B(n16325), .S(n20091), .Z(n14363) );
  NOR2_X1 U16509 ( .A1(n13396), .A2(n14363), .ZN(n13280) );
  AOI21_X1 U16510 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(n20020), .A(n13280), 
        .ZN(n13259) );
  OAI21_X1 U16511 ( .B1(n13260), .B2(n13397), .A(n13259), .ZN(P1_U2949) );
  INV_X1 U16512 ( .A(DATAI_10_), .ZN(n13261) );
  MUX2_X1 U16513 ( .A(n13261), .B(n16328), .S(n20091), .Z(n14313) );
  NOR2_X1 U16514 ( .A1(n13396), .A2(n14313), .ZN(n13301) );
  AOI21_X1 U16515 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n20020), .A(n13301), 
        .ZN(n13262) );
  OAI21_X1 U16516 ( .B1(n13263), .B2(n13397), .A(n13262), .ZN(P1_U2947) );
  NOR2_X1 U16517 ( .A1(n13396), .A2(n20105), .ZN(n13285) );
  AOI21_X1 U16518 ( .B1(P1_LWORD_REG_0__SCAN_IN), .B2(n20020), .A(n13285), 
        .ZN(n13264) );
  OAI21_X1 U16519 ( .B1(n13181), .B2(n13397), .A(n13264), .ZN(P1_U2952) );
  NAND2_X1 U16520 ( .A1(n20089), .A2(DATAI_7_), .ZN(n13266) );
  NAND2_X1 U16521 ( .A1(n20091), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13265) );
  NOR2_X1 U16522 ( .A1(n13396), .A2(n20145), .ZN(n13295) );
  AOI21_X1 U16523 ( .B1(P1_UWORD_REG_7__SCAN_IN), .B2(n20020), .A(n13295), 
        .ZN(n13267) );
  OAI21_X1 U16524 ( .B1(n13229), .B2(n13397), .A(n13267), .ZN(P1_U2944) );
  NAND2_X1 U16525 ( .A1(n20089), .A2(DATAI_2_), .ZN(n13269) );
  NAND2_X1 U16526 ( .A1(n20091), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13268) );
  AND2_X1 U16527 ( .A1(n13269), .A2(n13268), .ZN(n20119) );
  NOR2_X1 U16528 ( .A1(n13396), .A2(n20119), .ZN(n13304) );
  AOI21_X1 U16529 ( .B1(P1_UWORD_REG_2__SCAN_IN), .B2(n20020), .A(n13304), 
        .ZN(n13270) );
  OAI21_X1 U16530 ( .B1(n13207), .B2(n13397), .A(n13270), .ZN(P1_U2939) );
  NAND2_X1 U16531 ( .A1(n20089), .A2(DATAI_6_), .ZN(n13272) );
  NAND2_X1 U16532 ( .A1(n20091), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13271) );
  AND2_X1 U16533 ( .A1(n13272), .A2(n13271), .ZN(n20138) );
  NOR2_X1 U16534 ( .A1(n13396), .A2(n20138), .ZN(n13306) );
  AOI21_X1 U16535 ( .B1(P1_UWORD_REG_6__SCAN_IN), .B2(n20020), .A(n13306), 
        .ZN(n13273) );
  OAI21_X1 U16536 ( .B1(n13196), .B2(n13397), .A(n13273), .ZN(P1_U2943) );
  NAND2_X1 U16537 ( .A1(n20089), .A2(DATAI_5_), .ZN(n13275) );
  NAND2_X1 U16538 ( .A1(n20091), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13274) );
  AND2_X1 U16539 ( .A1(n13275), .A2(n13274), .ZN(n20134) );
  NOR2_X1 U16540 ( .A1(n13396), .A2(n20134), .ZN(n13287) );
  AOI21_X1 U16541 ( .B1(P1_UWORD_REG_5__SCAN_IN), .B2(n20020), .A(n13287), 
        .ZN(n13276) );
  OAI21_X1 U16542 ( .B1(n13189), .B2(n13397), .A(n13276), .ZN(P1_U2942) );
  NOR2_X1 U16543 ( .A1(n13396), .A2(n20114), .ZN(n13278) );
  AOI21_X1 U16544 ( .B1(P1_LWORD_REG_1__SCAN_IN), .B2(n20020), .A(n13278), 
        .ZN(n13277) );
  OAI21_X1 U16545 ( .B1(n13187), .B2(n13397), .A(n13277), .ZN(P1_U2953) );
  AOI21_X1 U16546 ( .B1(P1_UWORD_REG_1__SCAN_IN), .B2(n20020), .A(n13278), 
        .ZN(n13279) );
  OAI21_X1 U16547 ( .B1(n13210), .B2(n13397), .A(n13279), .ZN(P1_U2938) );
  AOI21_X1 U16548 ( .B1(P1_LWORD_REG_12__SCAN_IN), .B2(n20020), .A(n13280), 
        .ZN(n13281) );
  OAI21_X1 U16549 ( .B1(n13282), .B2(n13397), .A(n13281), .ZN(P1_U2964) );
  AOI21_X1 U16550 ( .B1(P1_LWORD_REG_3__SCAN_IN), .B2(n20020), .A(n13283), 
        .ZN(n13284) );
  OAI21_X1 U16551 ( .B1(n20865), .B2(n13397), .A(n13284), .ZN(P1_U2955) );
  AOI21_X1 U16552 ( .B1(P1_UWORD_REG_0__SCAN_IN), .B2(n20020), .A(n13285), 
        .ZN(n13286) );
  OAI21_X1 U16553 ( .B1(n13234), .B2(n13397), .A(n13286), .ZN(P1_U2937) );
  AOI21_X1 U16554 ( .B1(P1_LWORD_REG_5__SCAN_IN), .B2(n20020), .A(n13287), 
        .ZN(n13288) );
  OAI21_X1 U16555 ( .B1(n13289), .B2(n13397), .A(n13288), .ZN(P1_U2957) );
  INV_X1 U16556 ( .A(DATAI_9_), .ZN(n13291) );
  NAND2_X1 U16557 ( .A1(n20091), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13290) );
  OAI21_X1 U16558 ( .B1(n20091), .B2(n13291), .A(n13290), .ZN(n14317) );
  INV_X1 U16559 ( .A(n14317), .ZN(n13292) );
  NOR2_X1 U16560 ( .A1(n13396), .A2(n13292), .ZN(n20017) );
  AOI21_X1 U16561 ( .B1(P1_UWORD_REG_9__SCAN_IN), .B2(n20020), .A(n20017), 
        .ZN(n13293) );
  OAI21_X1 U16562 ( .B1(n13294), .B2(n13397), .A(n13293), .ZN(P1_U2946) );
  AOI21_X1 U16563 ( .B1(P1_LWORD_REG_7__SCAN_IN), .B2(n20020), .A(n13295), 
        .ZN(n13296) );
  OAI21_X1 U16564 ( .B1(n13297), .B2(n13397), .A(n13296), .ZN(P1_U2959) );
  INV_X1 U16565 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n13519) );
  NAND2_X1 U16566 ( .A1(n20089), .A2(DATAI_4_), .ZN(n13299) );
  NAND2_X1 U16567 ( .A1(n20091), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13298) );
  AND2_X1 U16568 ( .A1(n13299), .A2(n13298), .ZN(n20129) );
  NOR2_X1 U16569 ( .A1(n13396), .A2(n20129), .ZN(n13308) );
  AOI21_X1 U16570 ( .B1(P1_LWORD_REG_4__SCAN_IN), .B2(n20020), .A(n13308), 
        .ZN(n13300) );
  OAI21_X1 U16571 ( .B1(n13519), .B2(n13397), .A(n13300), .ZN(P1_U2956) );
  AOI21_X1 U16572 ( .B1(P1_LWORD_REG_10__SCAN_IN), .B2(n20020), .A(n13301), 
        .ZN(n13302) );
  OAI21_X1 U16573 ( .B1(n13303), .B2(n13397), .A(n13302), .ZN(P1_U2962) );
  AOI21_X1 U16574 ( .B1(P1_LWORD_REG_2__SCAN_IN), .B2(n20020), .A(n13304), 
        .ZN(n13305) );
  OAI21_X1 U16575 ( .B1(n13502), .B2(n13397), .A(n13305), .ZN(P1_U2954) );
  AOI21_X1 U16576 ( .B1(P1_LWORD_REG_6__SCAN_IN), .B2(n20020), .A(n13306), 
        .ZN(n13307) );
  OAI21_X1 U16577 ( .B1(n13584), .B2(n13397), .A(n13307), .ZN(P1_U2958) );
  AOI21_X1 U16578 ( .B1(P1_UWORD_REG_4__SCAN_IN), .B2(n20020), .A(n13308), 
        .ZN(n13309) );
  OAI21_X1 U16579 ( .B1(n13201), .B2(n13397), .A(n13309), .ZN(P1_U2941) );
  NAND2_X1 U16580 ( .A1(n20020), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13312) );
  INV_X1 U16581 ( .A(DATAI_8_), .ZN(n13311) );
  NAND2_X1 U16582 ( .A1(n20091), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13310) );
  OAI21_X1 U16583 ( .B1(n20091), .B2(n13311), .A(n13310), .ZN(n14322) );
  NAND2_X1 U16584 ( .A1(n20014), .A2(n14322), .ZN(n13329) );
  OAI211_X1 U16585 ( .C1(n13397), .C2(n13313), .A(n13312), .B(n13329), .ZN(
        P1_U2945) );
  NAND2_X1 U16586 ( .A1(n20020), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13316) );
  INV_X1 U16587 ( .A(DATAI_14_), .ZN(n13315) );
  NAND2_X1 U16588 ( .A1(n20091), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13314) );
  OAI21_X1 U16589 ( .B1(n20091), .B2(n13315), .A(n13314), .ZN(n14070) );
  NAND2_X1 U16590 ( .A1(n20014), .A2(n14070), .ZN(n13319) );
  OAI211_X1 U16591 ( .C1(n13397), .C2(n13317), .A(n13316), .B(n13319), .ZN(
        P1_U2951) );
  NAND2_X1 U16592 ( .A1(n20020), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n13318) );
  OAI211_X1 U16593 ( .C1(n13397), .C2(n13320), .A(n13319), .B(n13318), .ZN(
        P1_U2966) );
  NAND2_X1 U16594 ( .A1(n20020), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13323) );
  INV_X1 U16595 ( .A(DATAI_11_), .ZN(n13322) );
  NAND2_X1 U16596 ( .A1(n20091), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13321) );
  OAI21_X1 U16597 ( .B1(n20091), .B2(n13322), .A(n13321), .ZN(n14367) );
  NAND2_X1 U16598 ( .A1(n20014), .A2(n14367), .ZN(n13326) );
  OAI211_X1 U16599 ( .C1(n13397), .C2(n13324), .A(n13323), .B(n13326), .ZN(
        P1_U2948) );
  NAND2_X1 U16600 ( .A1(n20020), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n13325) );
  OAI211_X1 U16601 ( .C1(n13397), .C2(n13327), .A(n13326), .B(n13325), .ZN(
        P1_U2963) );
  NAND2_X1 U16602 ( .A1(n20020), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13328) );
  OAI211_X1 U16603 ( .C1(n13397), .C2(n13330), .A(n13329), .B(n13328), .ZN(
        P1_U2960) );
  INV_X1 U16604 ( .A(n13367), .ZN(n13340) );
  AOI22_X1 U16605 ( .A1(n13367), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n13360), .B2(n13340), .ZN(n13366) );
  NOR2_X1 U16606 ( .A1(n13331), .A2(n11408), .ZN(n13336) );
  INV_X1 U16607 ( .A(n13336), .ZN(n13334) );
  NOR2_X1 U16608 ( .A1(n13332), .A2(n11531), .ZN(n13333) );
  AOI22_X1 U16609 ( .A1(n13335), .A2(n13334), .B1(n13333), .B2(n13350), .ZN(
        n13339) );
  NAND2_X1 U16610 ( .A1(n13337), .A2(n13336), .ZN(n13338) );
  OAI211_X1 U16611 ( .C1(n14861), .C2(n13354), .A(n13339), .B(n13338), .ZN(
        n15549) );
  AOI22_X1 U16612 ( .A1(n13367), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15549), .B2(n13340), .ZN(n13365) );
  INV_X1 U16613 ( .A(n13366), .ZN(n13363) );
  INV_X1 U16614 ( .A(n13350), .ZN(n13345) );
  INV_X1 U16615 ( .A(n12031), .ZN(n13342) );
  NAND2_X1 U16616 ( .A1(n13342), .A2(n13341), .ZN(n13352) );
  INV_X1 U16617 ( .A(n13352), .ZN(n13344) );
  MUX2_X1 U16618 ( .A(n13345), .B(n13344), .S(n13343), .Z(n13346) );
  OAI21_X1 U16619 ( .B1(n13347), .B2(n13354), .A(n13346), .ZN(n15535) );
  INV_X1 U16620 ( .A(n13348), .ZN(n13351) );
  AOI22_X1 U16621 ( .A1(n13352), .A2(n13351), .B1(n13350), .B2(n13349), .ZN(
        n13353) );
  OAI22_X1 U16622 ( .A1(n13355), .A2(n13354), .B1(n13118), .B2(n13353), .ZN(
        n15544) );
  OAI21_X1 U16623 ( .B1(n13356), .B2(n15535), .A(n15544), .ZN(n13358) );
  OAI21_X1 U16624 ( .B1(n15535), .B2(n19865), .A(n19857), .ZN(n13357) );
  AOI21_X1 U16625 ( .B1(n13358), .B2(n13357), .A(n13367), .ZN(n13359) );
  OAI21_X1 U16626 ( .B1(n19842), .B2(n13360), .A(n13359), .ZN(n13361) );
  NAND2_X1 U16627 ( .A1(n19842), .A2(n20880), .ZN(n19212) );
  AOI222_X1 U16628 ( .A1(n13365), .A2(n13361), .B1(n13365), .B2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C1(n13361), .C2(n19212), .ZN(
        n13362) );
  AOI21_X1 U16629 ( .B1(n19842), .B2(n13363), .A(n13362), .ZN(n13364) );
  OAI22_X1 U16630 ( .A1(n13366), .A2(n13365), .B1(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n13364), .ZN(n13387) );
  NAND2_X1 U16631 ( .A1(n13367), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13385) );
  NOR2_X1 U16632 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n13372) );
  NAND3_X1 U16633 ( .A1(n15665), .A2(n19119), .A3(n15664), .ZN(n13371) );
  INV_X1 U16634 ( .A(n11883), .ZN(n13369) );
  NAND2_X1 U16635 ( .A1(n13369), .A2(n13368), .ZN(n13370) );
  OAI211_X1 U16636 ( .C1(n13373), .C2(n13372), .A(n13371), .B(n13370), .ZN(
        n13383) );
  INV_X1 U16637 ( .A(n13374), .ZN(n13381) );
  NAND2_X1 U16638 ( .A1(n13376), .A2(n13375), .ZN(n13380) );
  NAND2_X1 U16639 ( .A1(n13378), .A2(n13377), .ZN(n13379) );
  OAI211_X1 U16640 ( .C1(n13382), .C2(n13381), .A(n13380), .B(n13379), .ZN(
        n19870) );
  NOR2_X1 U16641 ( .A1(n13383), .A2(n19870), .ZN(n13384) );
  NAND2_X1 U16642 ( .A1(n13385), .A2(n13384), .ZN(n13386) );
  NOR2_X1 U16643 ( .A1(n13387), .A2(n13386), .ZN(n16237) );
  AOI21_X1 U16644 ( .B1(n16237), .B2(n19757), .A(n18737), .ZN(n13392) );
  NOR2_X1 U16645 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13388), .ZN(n14756) );
  AND3_X1 U16646 ( .A1(n13389), .A2(n14757), .A3(n14756), .ZN(n13391) );
  NAND2_X1 U16647 ( .A1(n13390), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19882) );
  NOR3_X1 U16648 ( .A1(n13392), .A2(n13391), .A3(n19882), .ZN(n16232) );
  OAI21_X1 U16649 ( .B1(n16232), .B2(n18737), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13393) );
  NAND2_X1 U16650 ( .A1(n13393), .A2(n15758), .ZN(P2_U3593) );
  INV_X1 U16651 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13394) );
  NOR2_X1 U16652 ( .A1(n20089), .A2(n13394), .ZN(n13395) );
  AOI21_X1 U16653 ( .B1(DATAI_15_), .B2(n20089), .A(n13395), .ZN(n14358) );
  OAI222_X1 U16654 ( .A1(n13397), .A2(n14359), .B1(n13396), .B2(n14358), .C1(
        n20019), .C2(n13239), .ZN(P1_U2967) );
  INV_X1 U16655 ( .A(n18976), .ZN(n13400) );
  NAND2_X1 U16656 ( .A1(n13400), .A2(n13399), .ZN(n13422) );
  INV_X1 U16657 ( .A(n13422), .ZN(n18977) );
  XNOR2_X1 U16658 ( .A(n18977), .B(n18970), .ZN(n13405) );
  NOR2_X1 U16659 ( .A1(n9709), .A2(n13401), .ZN(n13402) );
  OR2_X1 U16660 ( .A1(n9711), .A2(n13402), .ZN(n18852) );
  INV_X1 U16661 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13403) );
  MUX2_X1 U16662 ( .A(n18852), .B(n13403), .S(n18983), .Z(n13404) );
  OAI21_X1 U16663 ( .B1(n13405), .B2(n18984), .A(n13404), .ZN(P2_U2878) );
  INV_X1 U16664 ( .A(n13407), .ZN(n13408) );
  NAND2_X1 U16665 ( .A1(n13406), .A2(n13408), .ZN(n13409) );
  OR2_X1 U16666 ( .A1(n13410), .A2(n13409), .ZN(n13411) );
  NAND2_X1 U16667 ( .A1(n13159), .A2(n13411), .ZN(n19006) );
  NOR2_X1 U16668 ( .A1(n19839), .A2(n19838), .ZN(n13415) );
  NAND2_X1 U16669 ( .A1(n13412), .A2(n13242), .ZN(n13414) );
  NAND2_X1 U16670 ( .A1(n13414), .A2(n9739), .ZN(n18908) );
  OAI21_X1 U16671 ( .B1(n13416), .B2(n13415), .A(n18908), .ZN(n19008) );
  XOR2_X1 U16672 ( .A(n19006), .B(n19008), .Z(n13420) );
  OAI22_X1 U16673 ( .A1(n19101), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19103), .ZN(n19139) );
  INV_X1 U16674 ( .A(n19139), .ZN(n16119) );
  INV_X1 U16675 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n13417) );
  OAI22_X1 U16676 ( .A1(n20787), .A2(n18908), .B1(n14979), .B2(n13417), .ZN(
        n13418) );
  AOI21_X1 U16677 ( .B1(n19005), .B2(n16119), .A(n13418), .ZN(n13419) );
  OAI21_X1 U16678 ( .B1(n13420), .B2(n14996), .A(n13419), .ZN(P2_U2915) );
  NAND2_X1 U16679 ( .A1(n18970), .A2(n18969), .ZN(n13421) );
  XNOR2_X1 U16680 ( .A(n13511), .B(n18964), .ZN(n13428) );
  NAND2_X1 U16681 ( .A1(n13423), .A2(n14830), .ZN(n13424) );
  AND2_X1 U16682 ( .A1(n13424), .A2(n9785), .ZN(n18838) );
  NOR2_X1 U16683 ( .A1(n18988), .A2(n13425), .ZN(n13426) );
  AOI21_X1 U16684 ( .B1(n18838), .B2(n18988), .A(n13426), .ZN(n13427) );
  OAI21_X1 U16685 ( .B1(n13428), .B2(n18984), .A(n13427), .ZN(P2_U2876) );
  INV_X1 U16686 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13429) );
  OR2_X1 U16687 ( .A1(n19101), .A2(n13429), .ZN(n13431) );
  NAND2_X1 U16688 ( .A1(n19101), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13430) );
  AND2_X1 U16689 ( .A1(n13431), .A2(n13430), .ZN(n19078) );
  INV_X1 U16690 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19027) );
  OAI21_X1 U16691 ( .B1(n13433), .B2(n13432), .A(n14809), .ZN(n18834) );
  OAI222_X1 U16692 ( .A1(n13614), .A2(n19078), .B1(n14979), .B2(n19027), .C1(
        n19012), .C2(n18834), .ZN(P2_U2908) );
  NOR2_X1 U16693 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n15734), .ZN(n13443) );
  INV_X1 U16694 ( .A(n13443), .ZN(n13439) );
  AOI21_X1 U16695 ( .B1(n13435), .B2(n15708), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n13436) );
  OAI21_X1 U16696 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n15708), .A(
        n13436), .ZN(n13437) );
  OAI21_X1 U16697 ( .B1(n13439), .B2(n13438), .A(n13437), .ZN(n15704) );
  MUX2_X1 U16698 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13440), .S(
        n15708), .Z(n15717) );
  AOI22_X1 U16699 ( .A1(n15717), .A2(n15734), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13443), .ZN(n13445) );
  NOR2_X1 U16700 ( .A1(n15708), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13441) );
  AOI21_X1 U16701 ( .B1(n13442), .B2(n15708), .A(n13441), .ZN(n15713) );
  AOI22_X1 U16702 ( .A1(n13443), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15713), .B2(n15734), .ZN(n13444) );
  NOR2_X1 U16703 ( .A1(n13445), .A2(n13444), .ZN(n15727) );
  INV_X1 U16704 ( .A(n15727), .ZN(n13447) );
  NOR2_X1 U16705 ( .A1(n13447), .A2(n13446), .ZN(n13451) );
  NOR3_X1 U16706 ( .A1(n15704), .A2(n13451), .A3(P1_FLUSH_REG_SCAN_IN), .ZN(
        n13449) );
  NOR3_X1 U16707 ( .A1(n15704), .A2(n13451), .A3(n13450), .ZN(n15735) );
  INV_X1 U16708 ( .A(n13631), .ZN(n20214) );
  NAND2_X1 U16709 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20510), .ZN(n13477) );
  INV_X1 U16710 ( .A(n13477), .ZN(n13452) );
  OAI22_X1 U16711 ( .A1(n11070), .A2(n20622), .B1(n20214), .B2(n13452), .ZN(
        n13453) );
  OAI21_X1 U16712 ( .B1(n15735), .B2(n13453), .A(n20087), .ZN(n13454) );
  OAI21_X1 U16713 ( .B1(n20087), .B2(n20536), .A(n13454), .ZN(P1_U3478) );
  OAI21_X1 U16714 ( .B1(n13456), .B2(n13455), .A(n13534), .ZN(n19991) );
  NOR2_X1 U16715 ( .A1(n13543), .A2(n9717), .ZN(n20047) );
  AOI22_X1 U16716 ( .A1(n12418), .A2(n20047), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14288), .ZN(n13458) );
  OAI21_X1 U16717 ( .B1(n19991), .B2(n14297), .A(n13458), .ZN(P1_U2869) );
  NAND2_X1 U16718 ( .A1(n13459), .A2(n13460), .ZN(n13464) );
  INV_X1 U16719 ( .A(n13461), .ZN(n13462) );
  AOI21_X1 U16720 ( .B1(n13464), .B2(n13463), .A(n13462), .ZN(n13472) );
  AOI22_X1 U16721 ( .A1(n20025), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20024), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13465) );
  OAI21_X1 U16722 ( .B1(n20036), .B2(n14230), .A(n13465), .ZN(n13466) );
  AOI21_X1 U16723 ( .B1(n13472), .B2(n20031), .A(n13466), .ZN(n13471) );
  OR2_X1 U16724 ( .A1(n13467), .A2(n13468), .ZN(n20063) );
  NAND3_X1 U16725 ( .A1(n20063), .A2(n20032), .A3(n13469), .ZN(n13470) );
  NAND2_X1 U16726 ( .A1(n13471), .A2(n13470), .ZN(P1_U2997) );
  OAI222_X1 U16727 ( .A1(n14370), .A2(n19991), .B1(n14365), .B2(n20865), .C1(
        n14364), .C2(n20124), .ZN(P1_U2901) );
  INV_X1 U16728 ( .A(n13472), .ZN(n14236) );
  NAND2_X1 U16729 ( .A1(n13474), .A2(n13473), .ZN(n13475) );
  AOI22_X1 U16730 ( .A1(n12418), .A2(n20064), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n14288), .ZN(n13476) );
  OAI21_X1 U16731 ( .B1(n14236), .B2(n14297), .A(n13476), .ZN(P1_U2870) );
  NAND2_X1 U16732 ( .A1(n20087), .A2(n13477), .ZN(n13790) );
  NAND2_X1 U16733 ( .A1(n20087), .A2(n20624), .ZN(n13785) );
  NAND2_X1 U16734 ( .A1(n13479), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20618) );
  XNOR2_X1 U16735 ( .A(n20093), .B(n20618), .ZN(n13480) );
  OAI222_X1 U16736 ( .A1(n13790), .A2(n12965), .B1(n20087), .B2(n20425), .C1(
        n13785), .C2(n13480), .ZN(P1_U3476) );
  XNOR2_X1 U16737 ( .A(n13481), .B(n13567), .ZN(n13482) );
  XNOR2_X1 U16738 ( .A(n13483), .B(n13482), .ZN(n13501) );
  OAI21_X1 U16739 ( .B1(n15381), .B2(n13485), .A(n13484), .ZN(n15522) );
  INV_X1 U16740 ( .A(n15522), .ZN(n13486) );
  MUX2_X1 U16741 ( .A(n16196), .B(n13486), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n13487) );
  OAI21_X1 U16742 ( .B1(n13493), .B2(n18871), .A(n13487), .ZN(n13489) );
  NOR2_X1 U16743 ( .A1(n14849), .A2(n16204), .ZN(n13488) );
  AOI211_X1 U16744 ( .C1(n16218), .C2(n14847), .A(n13489), .B(n13488), .ZN(
        n13492) );
  OR2_X1 U16745 ( .A1(n9663), .A2(n13490), .ZN(n13498) );
  NAND3_X1 U16746 ( .A1(n13498), .A2(n16192), .A3(n13497), .ZN(n13491) );
  OAI211_X1 U16747 ( .C1(n13501), .C2(n16222), .A(n13492), .B(n13491), .ZN(
        P2_U3043) );
  NOR2_X1 U16748 ( .A1(n18871), .A2(n13493), .ZN(n13496) );
  INV_X1 U16749 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14841) );
  OAI21_X1 U16750 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13494), .A(
        n14719), .ZN(n14839) );
  OAI22_X1 U16751 ( .A1(n14841), .A2(n19100), .B1(n16166), .B2(n14839), .ZN(
        n13495) );
  AOI211_X1 U16752 ( .C1(n19094), .C2(n14847), .A(n13496), .B(n13495), .ZN(
        n13500) );
  NAND3_X1 U16753 ( .A1(n13498), .A2(n19091), .A3(n13497), .ZN(n13499) );
  OAI211_X1 U16754 ( .C1(n13501), .C2(n16168), .A(n13500), .B(n13499), .ZN(
        P2_U3011) );
  OAI222_X1 U16755 ( .A1(n14370), .A2(n14236), .B1(n14365), .B2(n13502), .C1(
        n14364), .C2(n20119), .ZN(P1_U2902) );
  INV_X1 U16756 ( .A(n9603), .ZN(n13509) );
  INV_X1 U16757 ( .A(n13785), .ZN(n13507) );
  OR2_X1 U16758 ( .A1(n13479), .A2(n20254), .ZN(n20541) );
  OAI22_X1 U16759 ( .A1(n20343), .A2(n20618), .B1(n20539), .B2(n20541), .ZN(
        n13505) );
  INV_X1 U16760 ( .A(n11089), .ZN(n13504) );
  AOI22_X1 U16761 ( .A1(n13505), .A2(n20481), .B1(n13504), .B2(n20254), .ZN(
        n13506) );
  INV_X1 U16762 ( .A(n20087), .ZN(n13788) );
  AOI22_X1 U16763 ( .A1(n13507), .A2(n13506), .B1(n13788), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13508) );
  OAI21_X1 U16764 ( .B1(n13509), .B2(n13790), .A(n13508), .ZN(P1_U3475) );
  AND2_X1 U16765 ( .A1(n18964), .A2(n18963), .ZN(n13510) );
  OAI211_X1 U16766 ( .C1(n13512), .C2(n13513), .A(n13671), .B(n18954), .ZN(
        n13518) );
  NAND2_X1 U16767 ( .A1(n13514), .A2(n13515), .ZN(n13516) );
  AND2_X1 U16768 ( .A1(n15425), .A2(n13516), .ZN(n18824) );
  NAND2_X1 U16769 ( .A1(n18824), .A2(n18988), .ZN(n13517) );
  OAI211_X1 U16770 ( .C1(n18988), .C2(n11774), .A(n13518), .B(n13517), .ZN(
        P2_U2874) );
  XOR2_X1 U16771 ( .A(n13534), .B(n13533), .Z(n20030) );
  INV_X1 U16772 ( .A(n20030), .ZN(n13546) );
  OAI222_X1 U16773 ( .A1(n14364), .A2(n20129), .B1(n14370), .B2(n13546), .C1(
        n13519), .C2(n14365), .ZN(P1_U2900) );
  INV_X1 U16774 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14299) );
  OR2_X1 U16775 ( .A1(n19101), .A2(n14299), .ZN(n13521) );
  NAND2_X1 U16776 ( .A1(n19101), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13520) );
  AND2_X1 U16777 ( .A1(n13521), .A2(n13520), .ZN(n19083) );
  OAI21_X1 U16778 ( .B1(n13523), .B2(n13522), .A(n15428), .ZN(n18825) );
  INV_X1 U16779 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19023) );
  OAI222_X1 U16780 ( .A1(n13614), .A2(n19083), .B1(n18825), .B2(n19012), .C1(
        n19023), .C2(n14979), .ZN(P2_U2906) );
  OR2_X1 U16781 ( .A1(n13525), .A2(n13524), .ZN(n13526) );
  AND2_X1 U16782 ( .A1(n13527), .A2(n13526), .ZN(n20051) );
  NAND2_X1 U16783 ( .A1(n20051), .A2(n20032), .ZN(n13532) );
  INV_X1 U16784 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13528) );
  NOR2_X1 U16785 ( .A1(n20065), .A2(n13528), .ZN(n20046) );
  NOR2_X1 U16786 ( .A1(n14484), .A2(n13529), .ZN(n13530) );
  AOI211_X1 U16787 ( .C1(n15889), .C2(n19994), .A(n20046), .B(n13530), .ZN(
        n13531) );
  OAI211_X1 U16788 ( .C1(n20090), .C2(n19991), .A(n13532), .B(n13531), .ZN(
        P1_U2996) );
  OR2_X1 U16789 ( .A1(n13534), .A2(n13533), .ZN(n13535) );
  AND2_X1 U16790 ( .A1(n13536), .A2(n13535), .ZN(n13538) );
  OR2_X1 U16791 ( .A1(n13538), .A2(n13537), .ZN(n15914) );
  INV_X1 U16792 ( .A(n13558), .ZN(n13539) );
  AOI21_X1 U16793 ( .B1(n13540), .B2(n13545), .A(n13539), .ZN(n19960) );
  AOI22_X1 U16794 ( .A1(n12418), .A2(n19960), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14288), .ZN(n13541) );
  OAI21_X1 U16795 ( .B1(n15914), .B2(n14290), .A(n13541), .ZN(P1_U2867) );
  OR2_X1 U16796 ( .A1(n13543), .A2(n13542), .ZN(n13544) );
  NAND2_X1 U16797 ( .A1(n13545), .A2(n13544), .ZN(n20039) );
  INV_X1 U16798 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13547) );
  OAI222_X1 U16799 ( .A1(n20039), .A2(n14298), .B1(n13547), .B2(n20003), .C1(
        n14297), .C2(n13546), .ZN(P1_U2868) );
  OAI222_X1 U16800 ( .A1(n14370), .A2(n15914), .B1(n14365), .B2(n13289), .C1(
        n14364), .C2(n20134), .ZN(P1_U2899) );
  NAND2_X1 U16801 ( .A1(n13549), .A2(n13550), .ZN(n13551) );
  AND2_X1 U16802 ( .A1(n13548), .A2(n13551), .ZN(n19944) );
  INV_X1 U16803 ( .A(n19944), .ZN(n13583) );
  INV_X1 U16804 ( .A(n13552), .ZN(n13554) );
  INV_X1 U16805 ( .A(n13560), .ZN(n13553) );
  AOI21_X1 U16806 ( .B1(n13554), .B2(n13553), .A(n13688), .ZN(n19935) );
  AOI22_X1 U16807 ( .A1(n19935), .A2(n12418), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n14288), .ZN(n13555) );
  OAI21_X1 U16808 ( .B1(n13583), .B2(n14290), .A(n13555), .ZN(P1_U2865) );
  XOR2_X1 U16809 ( .A(n13537), .B(n13556), .Z(n19956) );
  INV_X1 U16810 ( .A(n19956), .ZN(n13585) );
  AND2_X1 U16811 ( .A1(n13558), .A2(n13557), .ZN(n13559) );
  NOR2_X1 U16812 ( .A1(n13560), .A2(n13559), .ZN(n19948) );
  AOI22_X1 U16813 ( .A1(n12418), .A2(n19948), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14288), .ZN(n13561) );
  OAI21_X1 U16814 ( .B1(n13585), .B2(n14297), .A(n13561), .ZN(P1_U2866) );
  XOR2_X1 U16815 ( .A(n13563), .B(n13562), .Z(n19096) );
  INV_X1 U16816 ( .A(n19096), .ZN(n13576) );
  XNOR2_X1 U16817 ( .A(n13564), .B(n13597), .ZN(n13566) );
  XNOR2_X1 U16818 ( .A(n13566), .B(n13565), .ZN(n19092) );
  NAND2_X1 U16819 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15525), .ZN(
        n13596) );
  OAI21_X1 U16820 ( .B1(n15522), .B2(n13567), .A(n15263), .ZN(n13601) );
  NAND2_X1 U16821 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19090), .ZN(n13568) );
  OAI221_X1 U16822 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13596), .C1(
        n13597), .C2(n13601), .A(n13568), .ZN(n13574) );
  NAND2_X1 U16823 ( .A1(n13570), .A2(n13569), .ZN(n13571) );
  AND2_X1 U16824 ( .A1(n13572), .A2(n13571), .ZN(n19093) );
  INV_X1 U16825 ( .A(n19093), .ZN(n18982) );
  OAI22_X1 U16826 ( .A1(n18982), .A2(n15521), .B1(n16204), .B2(n18908), .ZN(
        n13573) );
  AOI211_X1 U16827 ( .C1(n19092), .C2(n16192), .A(n13574), .B(n13573), .ZN(
        n13575) );
  OAI21_X1 U16828 ( .B1(n13576), .B2(n16222), .A(n13575), .ZN(P2_U3042) );
  INV_X1 U16829 ( .A(n13577), .ZN(n18958) );
  OR2_X1 U16830 ( .A1(n13671), .A2(n18958), .ZN(n18959) );
  INV_X1 U16831 ( .A(n13578), .ZN(n13672) );
  XNOR2_X1 U16832 ( .A(n18959), .B(n13672), .ZN(n13582) );
  OR2_X1 U16833 ( .A1(n15426), .A2(n13579), .ZN(n13580) );
  NAND2_X1 U16834 ( .A1(n14785), .A2(n13580), .ZN(n15407) );
  MUX2_X1 U16835 ( .A(n15407), .B(n11801), .S(n18983), .Z(n13581) );
  OAI21_X1 U16836 ( .B1(n13582), .B2(n18984), .A(n13581), .ZN(P2_U2872) );
  OAI222_X1 U16837 ( .A1(n14370), .A2(n13583), .B1(n14365), .B2(n13297), .C1(
        n14364), .C2(n20145), .ZN(P1_U2897) );
  OAI222_X1 U16838 ( .A1(n14364), .A2(n20138), .B1(n14370), .B2(n13585), .C1(
        n13584), .C2(n14365), .ZN(P1_U2898) );
  XNOR2_X1 U16839 ( .A(n13587), .B(n9598), .ZN(n13610) );
  NOR2_X1 U16840 ( .A1(n18871), .A2(n13588), .ZN(n13603) );
  OAI21_X1 U16841 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n14718), .A(
        n14717), .ZN(n18898) );
  OAI22_X1 U16842 ( .A1(n19100), .A2(n9898), .B1(n16166), .B2(n18898), .ZN(
        n13589) );
  AOI211_X1 U16843 ( .C1(n13604), .C2(n19094), .A(n13603), .B(n13589), .ZN(
        n13595) );
  NOR2_X1 U16844 ( .A1(n13591), .A2(n13590), .ZN(n13593) );
  XNOR2_X1 U16845 ( .A(n13593), .B(n13592), .ZN(n13608) );
  NAND2_X1 U16846 ( .A1(n13608), .A2(n19091), .ZN(n13594) );
  OAI211_X1 U16847 ( .C1(n13610), .C2(n16168), .A(n13595), .B(n13594), .ZN(
        P2_U3009) );
  AOI221_X1 U16848 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n13600), .C2(n13597), .A(
        n13596), .ZN(n13607) );
  OAI21_X1 U16849 ( .B1(n13413), .B2(n13599), .A(n13598), .ZN(n19011) );
  NOR2_X1 U16850 ( .A1(n13601), .A2(n13600), .ZN(n13602) );
  AOI211_X1 U16851 ( .C1(n13604), .C2(n16218), .A(n13603), .B(n13602), .ZN(
        n13605) );
  OAI21_X1 U16852 ( .B1(n19011), .B2(n16204), .A(n13605), .ZN(n13606) );
  AOI211_X1 U16853 ( .C1(n13608), .C2(n16192), .A(n13607), .B(n13606), .ZN(
        n13609) );
  OAI21_X1 U16854 ( .B1(n16222), .B2(n13610), .A(n13609), .ZN(P2_U3041) );
  AOI22_X1 U16855 ( .A1(n19103), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19101), .ZN(n19087) );
  OAI21_X1 U16856 ( .B1(n13611), .B2(n13613), .A(n13695), .ZN(n15411) );
  INV_X1 U16857 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19019) );
  OAI222_X1 U16858 ( .A1(n13614), .A2(n19087), .B1(n15411), .B2(n19012), .C1(
        n19019), .C2(n14979), .ZN(P2_U2904) );
  INV_X1 U16859 ( .A(n13615), .ZN(n13642) );
  NOR2_X1 U16860 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15734), .ZN(n13616) );
  AND2_X1 U16861 ( .A1(n11020), .A2(n13616), .ZN(n13619) );
  NAND2_X1 U16862 ( .A1(n19904), .A2(n20772), .ZN(n13617) );
  NOR2_X1 U16863 ( .A1(n13617), .A2(n20097), .ZN(n13618) );
  INV_X1 U16864 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14093) );
  NOR2_X1 U16865 ( .A1(n14377), .A2(n15734), .ZN(n13623) );
  NAND2_X1 U16866 ( .A1(n20766), .A2(n13624), .ZN(n13625) );
  NAND2_X1 U16867 ( .A1(n15810), .A2(n13625), .ZN(n19978) );
  NAND2_X1 U16868 ( .A1(n20766), .A2(n10224), .ZN(n13637) );
  AND2_X1 U16869 ( .A1(n20768), .A2(n20254), .ZN(n15731) );
  NAND2_X1 U16870 ( .A1(n10222), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13626) );
  INV_X1 U16871 ( .A(n13626), .ZN(n13629) );
  OR2_X1 U16872 ( .A1(n13627), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13636) );
  INV_X1 U16873 ( .A(n13636), .ZN(n13628) );
  NAND2_X1 U16874 ( .A1(n19982), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13633) );
  AND2_X1 U16875 ( .A1(n20766), .A2(n13630), .ZN(n19987) );
  NAND2_X1 U16876 ( .A1(n19987), .A2(n13631), .ZN(n13632) );
  OAI211_X1 U16877 ( .C1(n13634), .C2(n19971), .A(n13633), .B(n13632), .ZN(
        n13641) );
  OAI21_X1 U16878 ( .B1(n19986), .B2(n19993), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13639) );
  NAND2_X1 U16879 ( .A1(n15838), .A2(n14217), .ZN(n15834) );
  NAND2_X1 U16880 ( .A1(n15834), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13638) );
  NAND2_X1 U16881 ( .A1(n13639), .A2(n13638), .ZN(n13640) );
  AOI211_X1 U16882 ( .C1(n13642), .C2(n19978), .A(n13641), .B(n13640), .ZN(
        n13643) );
  INV_X1 U16883 ( .A(n13643), .ZN(P1_U2840) );
  INV_X1 U16884 ( .A(n19978), .ZN(n19990) );
  OAI22_X1 U16885 ( .A1(n15838), .A2(P1_REIP_REG_1__SCAN_IN), .B1(n19971), 
        .B2(n20080), .ZN(n13646) );
  INV_X1 U16886 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13644) );
  OAI22_X1 U16887 ( .A1(n19936), .A2(n13644), .B1(n14217), .B2(n14227), .ZN(
        n13645) );
  NOR2_X1 U16888 ( .A1(n13646), .A2(n13645), .ZN(n13653) );
  INV_X1 U16889 ( .A(n13648), .ZN(n20564) );
  NAND2_X1 U16890 ( .A1(n20564), .A2(n19987), .ZN(n13652) );
  NAND2_X1 U16891 ( .A1(n19993), .A2(n13649), .ZN(n13651) );
  NAND2_X1 U16892 ( .A1(n19986), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13650) );
  AND4_X1 U16893 ( .A1(n13653), .A2(n13652), .A3(n13651), .A4(n13650), .ZN(
        n13654) );
  OAI21_X1 U16894 ( .B1(n13655), .B2(n19990), .A(n13654), .ZN(P1_U2839) );
  INV_X1 U16895 ( .A(n13657), .ZN(n13658) );
  AOI21_X1 U16896 ( .B1(n13659), .B2(n13548), .A(n13658), .ZN(n13754) );
  INV_X1 U16897 ( .A(n13754), .ZN(n14226) );
  INV_X1 U16898 ( .A(n14364), .ZN(n14368) );
  AOI22_X1 U16899 ( .A1(n14368), .A2(n14322), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14366), .ZN(n13660) );
  OAI21_X1 U16900 ( .B1(n14226), .B2(n14370), .A(n13660), .ZN(P1_U2896) );
  XNOR2_X1 U16901 ( .A(n13695), .B(n13691), .ZN(n15398) );
  INV_X1 U16902 ( .A(n15398), .ZN(n14796) );
  AOI22_X1 U16903 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13664) );
  AOI22_X1 U16904 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13663) );
  AOI22_X1 U16905 ( .A1(n11597), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13662) );
  AOI22_X1 U16906 ( .A1(n13113), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11611), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13661) );
  NAND4_X1 U16907 ( .A1(n13664), .A2(n13663), .A3(n13662), .A4(n13661), .ZN(
        n13670) );
  AOI22_X1 U16908 ( .A1(n12120), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13668) );
  AOI22_X1 U16909 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13828), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13667) );
  AOI22_X1 U16910 ( .A1(n12169), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13666) );
  AOI22_X1 U16911 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13665) );
  NAND4_X1 U16912 ( .A1(n13668), .A2(n13667), .A3(n13666), .A4(n13665), .ZN(
        n13669) );
  NOR2_X1 U16913 ( .A1(n13670), .A2(n13669), .ZN(n13674) );
  AOI21_X1 U16914 ( .B1(n13674), .B2(n13673), .A(n13710), .ZN(n18955) );
  AND2_X1 U16915 ( .A1(n12321), .A2(n13675), .ZN(n13676) );
  INV_X1 U16916 ( .A(n20782), .ZN(n14980) );
  OAI22_X1 U16917 ( .A1(n14980), .A2(n19109), .B1(n14979), .B2(n13677), .ZN(
        n13685) );
  AND2_X1 U16918 ( .A1(n13679), .A2(n19101), .ZN(n13678) );
  INV_X1 U16919 ( .A(n20784), .ZN(n14969) );
  INV_X1 U16920 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n13683) );
  AND2_X1 U16921 ( .A1(n13679), .A2(n19103), .ZN(n13680) );
  INV_X1 U16922 ( .A(n20783), .ZN(n13682) );
  INV_X1 U16923 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n13681) );
  OAI22_X1 U16924 ( .A1(n14969), .A2(n13683), .B1(n13682), .B2(n13681), .ZN(
        n13684) );
  AOI211_X1 U16925 ( .C1(n18955), .C2(n20791), .A(n13685), .B(n13684), .ZN(
        n13686) );
  OAI21_X1 U16926 ( .B1(n14796), .B2(n20787), .A(n13686), .ZN(P2_U2903) );
  INV_X1 U16927 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13690) );
  OR2_X1 U16928 ( .A1(n13688), .A2(n13687), .ZN(n13689) );
  NAND2_X1 U16929 ( .A1(n15970), .A2(n13689), .ZN(n15984) );
  OAI222_X1 U16930 ( .A1(n14226), .A2(n14297), .B1(n20003), .B2(n13690), .C1(
        n15984), .C2(n14298), .ZN(P1_U2864) );
  INV_X1 U16931 ( .A(n13691), .ZN(n13694) );
  INV_X1 U16932 ( .A(n13692), .ZN(n13693) );
  OAI21_X1 U16933 ( .B1(n13695), .B2(n13694), .A(n13693), .ZN(n13696) );
  INV_X1 U16934 ( .A(n13696), .ZN(n13698) );
  OR2_X1 U16935 ( .A1(n13698), .A2(n13697), .ZN(n18801) );
  AOI22_X1 U16936 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11564), .B1(
        n11602), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13702) );
  AOI22_X1 U16937 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13701) );
  AOI22_X1 U16938 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11597), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13700) );
  AOI22_X1 U16939 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11611), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13699) );
  NAND4_X1 U16940 ( .A1(n13702), .A2(n13701), .A3(n13700), .A4(n13699), .ZN(
        n13709) );
  AOI22_X1 U16941 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12120), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13707) );
  AOI22_X1 U16942 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n13828), .ZN(n13706) );
  AOI22_X1 U16943 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12170), .B1(
        n12169), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13705) );
  AOI22_X1 U16944 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13704) );
  NAND4_X1 U16945 ( .A1(n13707), .A2(n13706), .A3(n13705), .A4(n13704), .ZN(
        n13708) );
  NAND2_X1 U16946 ( .A1(n13710), .A2(n13711), .ZN(n13791) );
  OR2_X1 U16947 ( .A1(n13710), .A2(n13711), .ZN(n13712) );
  NAND2_X1 U16948 ( .A1(n13791), .A2(n13712), .ZN(n14932) );
  INV_X1 U16949 ( .A(n19121), .ZN(n13713) );
  AOI22_X1 U16950 ( .A1(n20782), .A2(n13713), .B1(n20780), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n13715) );
  AOI22_X1 U16951 ( .A1(n20784), .A2(BUF2_REG_17__SCAN_IN), .B1(n20783), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n13714) );
  OAI211_X1 U16952 ( .C1(n14932), .C2(n14996), .A(n13715), .B(n13714), .ZN(
        n13716) );
  INV_X1 U16953 ( .A(n13716), .ZN(n13717) );
  OAI21_X1 U16954 ( .B1(n18801), .B2(n20787), .A(n13717), .ZN(P2_U2902) );
  XNOR2_X1 U16955 ( .A(n13719), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13720) );
  XNOR2_X1 U16956 ( .A(n9576), .B(n13720), .ZN(n15907) );
  INV_X1 U16957 ( .A(n15907), .ZN(n13734) );
  NOR2_X1 U16958 ( .A1(n20071), .A2(n20086), .ZN(n13726) );
  NAND2_X1 U16959 ( .A1(n20056), .A2(n13726), .ZN(n13731) );
  OAI21_X1 U16960 ( .B1(n20058), .B2(n20086), .A(n20071), .ZN(n20037) );
  INV_X1 U16961 ( .A(n20037), .ZN(n13723) );
  OR2_X1 U16962 ( .A1(n20057), .A2(n13723), .ZN(n13724) );
  NOR2_X1 U16963 ( .A1(n20045), .A2(n20054), .ZN(n20040) );
  INV_X1 U16964 ( .A(n20040), .ZN(n13727) );
  NAND2_X1 U16965 ( .A1(n20040), .A2(n13725), .ZN(n15999) );
  INV_X1 U16966 ( .A(n13726), .ZN(n20038) );
  NOR2_X1 U16967 ( .A1(n13727), .A2(n20038), .ZN(n14522) );
  NAND3_X1 U16968 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20040), .A3(
        n20037), .ZN(n14537) );
  OAI21_X1 U16969 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13728), .A(
        n20085), .ZN(n20059) );
  AOI21_X1 U16970 ( .B1(n13729), .B2(n14537), .A(n20059), .ZN(n15946) );
  OAI21_X1 U16971 ( .B1(n14681), .B2(n14522), .A(n15946), .ZN(n15995) );
  INV_X1 U16972 ( .A(n15995), .ZN(n13730) );
  OAI211_X1 U16973 ( .C1(n13731), .C2(n15999), .A(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n13730), .ZN(n15981) );
  OAI21_X1 U16974 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15983), .A(
        n15981), .ZN(n13733) );
  AOI22_X1 U16975 ( .A1(n20048), .A2(n19948), .B1(n20024), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n13732) );
  OAI211_X1 U16976 ( .C1(n13734), .C2(n20073), .A(n13733), .B(n13732), .ZN(
        P1_U3025) );
  INV_X1 U16977 ( .A(n13735), .ZN(n13739) );
  INV_X1 U16978 ( .A(n13736), .ZN(n13738) );
  AOI21_X1 U16979 ( .B1(n13739), .B2(n13738), .A(n13737), .ZN(n15850) );
  AND2_X1 U16980 ( .A1(n15972), .A2(n13740), .ZN(n13741) );
  OR2_X1 U16981 ( .A1(n14292), .A2(n13741), .ZN(n15846) );
  OAI22_X1 U16982 ( .A1(n15846), .A2(n14298), .B1(n15845), .B2(n20003), .ZN(
        n13742) );
  AOI21_X1 U16983 ( .B1(n15850), .B2(n19999), .A(n13742), .ZN(n13743) );
  INV_X1 U16984 ( .A(n13743), .ZN(P1_U2862) );
  AND2_X1 U16985 ( .A1(n13657), .A2(n13744), .ZN(n13745) );
  NOR2_X1 U16986 ( .A1(n13736), .A2(n13745), .ZN(n20000) );
  INV_X1 U16987 ( .A(n20000), .ZN(n13747) );
  AOI22_X1 U16988 ( .A1(n14368), .A2(n14317), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14366), .ZN(n13746) );
  OAI21_X1 U16989 ( .B1(n13747), .B2(n14370), .A(n13746), .ZN(P1_U2895) );
  INV_X1 U16990 ( .A(n15850), .ZN(n13748) );
  OAI222_X1 U16991 ( .A1(n14370), .A2(n13748), .B1(n14364), .B2(n14313), .C1(
        n13303), .C2(n14365), .ZN(P1_U2894) );
  XNOR2_X1 U16992 ( .A(n13750), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13751) );
  XNOR2_X1 U16993 ( .A(n9597), .B(n13751), .ZN(n15987) );
  INV_X1 U16994 ( .A(n15987), .ZN(n13756) );
  AOI22_X1 U16995 ( .A1(n20025), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20024), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13752) );
  OAI21_X1 U16996 ( .B1(n20036), .B2(n14220), .A(n13752), .ZN(n13753) );
  AOI21_X1 U16997 ( .B1(n13754), .B2(n20031), .A(n13753), .ZN(n13755) );
  OAI21_X1 U16998 ( .B1(n13756), .B2(n19908), .A(n13755), .ZN(P1_U2991) );
  XNOR2_X1 U16999 ( .A(n9582), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13758) );
  XNOR2_X1 U17000 ( .A(n13757), .B(n13758), .ZN(n15974) );
  AOI22_X1 U17001 ( .A1(n20025), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n20024), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n13759) );
  OAI21_X1 U17002 ( .B1(n20036), .B2(n13760), .A(n13759), .ZN(n13761) );
  AOI21_X1 U17003 ( .B1(n20000), .B2(n20031), .A(n13761), .ZN(n13762) );
  OAI21_X1 U17004 ( .B1(n15974), .B2(n19908), .A(n13762), .ZN(P1_U2990) );
  OAI21_X1 U17005 ( .B1(n13737), .B2(n10575), .A(n13764), .ZN(n14295) );
  OAI21_X1 U17006 ( .B1(n14295), .B2(n14296), .A(n13764), .ZN(n13766) );
  NAND2_X1 U17007 ( .A1(n13766), .A2(n13765), .ZN(n14205) );
  OAI21_X1 U17008 ( .B1(n13766), .B2(n13765), .A(n14205), .ZN(n15825) );
  XNOR2_X1 U17009 ( .A(n14294), .B(n13767), .ZN(n15951) );
  AOI22_X1 U17010 ( .A1(n15951), .A2(n12418), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n14288), .ZN(n13768) );
  OAI21_X1 U17011 ( .B1(n15825), .B2(n14290), .A(n13768), .ZN(P1_U2860) );
  OAI21_X1 U17012 ( .B1(n13769), .B2(n13772), .A(n13771), .ZN(n14496) );
  AOI22_X1 U17013 ( .A1(n14368), .A2(n14070), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14366), .ZN(n13773) );
  OAI21_X1 U17014 ( .B1(n14496), .B2(n14370), .A(n13773), .ZN(P1_U2890) );
  AOI21_X1 U17015 ( .B1(n13774), .B2(n14208), .A(n14282), .ZN(n14670) );
  AOI22_X1 U17016 ( .A1(n14670), .A2(n12418), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n14288), .ZN(n13775) );
  OAI21_X1 U17017 ( .B1(n14496), .B2(n14290), .A(n13775), .ZN(P1_U2858) );
  INV_X1 U17018 ( .A(n14498), .ZN(n13776) );
  AOI22_X1 U17019 ( .A1(n13776), .A2(n19993), .B1(n19986), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n13778) );
  NAND2_X1 U17020 ( .A1(n14217), .A2(n13777), .ZN(n19962) );
  OAI211_X1 U17021 ( .C1(n13779), .C2(n19936), .A(n13778), .B(n19962), .ZN(
        n13780) );
  AOI21_X1 U17022 ( .B1(n14670), .B2(n19983), .A(n13780), .ZN(n13784) );
  NAND4_X1 U17023 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(P1_REIP_REG_14__SCAN_IN), .A4(P1_REIP_REG_13__SCAN_IN), .ZN(n14075) );
  INV_X1 U17024 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20697) );
  NAND2_X1 U17025 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n19984) );
  NOR3_X1 U17026 ( .A1(n14227), .A2(n20697), .A3(n19984), .ZN(n19924) );
  INV_X1 U17027 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20706) );
  INV_X1 U17028 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20704) );
  NAND2_X1 U17029 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19941) );
  NOR3_X1 U17030 ( .A1(n20706), .A2(n20704), .A3(n19941), .ZN(n19926) );
  NAND4_X1 U17031 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(n19924), .A4(n19926), .ZN(n15837) );
  INV_X1 U17032 ( .A(n14217), .ZN(n14228) );
  OR2_X1 U17033 ( .A1(n15837), .A2(n14228), .ZN(n15833) );
  OAI21_X1 U17034 ( .B1(n14075), .B2(n15833), .A(n15834), .ZN(n13781) );
  INV_X1 U17035 ( .A(n13781), .ZN(n15820) );
  INV_X1 U17036 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20714) );
  INV_X1 U17037 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20710) );
  NOR3_X1 U17038 ( .A1(n15838), .A2(n15837), .A3(n20710), .ZN(n15828) );
  NAND2_X1 U17039 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n15828), .ZN(n14213) );
  INV_X1 U17040 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20716) );
  OAI21_X1 U17041 ( .B1(n20714), .B2(n14213), .A(n20716), .ZN(n13782) );
  NAND2_X1 U17042 ( .A1(n15820), .A2(n13782), .ZN(n13783) );
  OAI211_X1 U17043 ( .C1(n14496), .C2(n15810), .A(n13784), .B(n13783), .ZN(
        P1_U2826) );
  INV_X1 U17044 ( .A(n13479), .ZN(n13786) );
  INV_X1 U17045 ( .A(n20618), .ZN(n20217) );
  AOI211_X1 U17046 ( .C1(n13786), .C2(n20254), .A(n20217), .B(n13785), .ZN(
        n13787) );
  AOI21_X1 U17047 ( .B1(n13788), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n13787), .ZN(n13789) );
  OAI21_X1 U17048 ( .B1(n13648), .B2(n13790), .A(n13789), .ZN(P1_U3477) );
  INV_X1 U17049 ( .A(n13791), .ZN(n13803) );
  AOI22_X1 U17050 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n11564), .B1(
        n11602), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13795) );
  AOI22_X1 U17051 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13794) );
  AOI22_X1 U17052 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11597), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13793) );
  AOI22_X1 U17053 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11611), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13792) );
  NAND4_X1 U17054 ( .A1(n13795), .A2(n13794), .A3(n13793), .A4(n13792), .ZN(
        n13801) );
  AOI22_X1 U17055 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12120), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13799) );
  AOI22_X1 U17056 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n13828), .ZN(n13798) );
  AOI22_X1 U17057 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12170), .B1(
        n12169), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13797) );
  AOI22_X1 U17058 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13796) );
  NAND4_X1 U17059 ( .A1(n13799), .A2(n13798), .A3(n13797), .A4(n13796), .ZN(
        n13800) );
  NOR2_X1 U17060 ( .A1(n13801), .A2(n13800), .ZN(n16111) );
  NAND2_X1 U17061 ( .A1(n13803), .A2(n13802), .ZN(n14921) );
  AOI22_X1 U17062 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n11564), .B1(
        n11602), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13807) );
  AOI22_X1 U17063 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13806) );
  AOI22_X1 U17064 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11597), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13805) );
  AOI22_X1 U17065 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11611), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13804) );
  NAND4_X1 U17066 ( .A1(n13807), .A2(n13806), .A3(n13805), .A4(n13804), .ZN(
        n13813) );
  AOI22_X1 U17067 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12120), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13811) );
  AOI22_X1 U17068 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n13828), .ZN(n13810) );
  AOI22_X1 U17069 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12170), .B1(
        n12169), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13809) );
  AOI22_X1 U17070 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13808) );
  NAND4_X1 U17071 ( .A1(n13811), .A2(n13810), .A3(n13809), .A4(n13808), .ZN(
        n13812) );
  NOR2_X1 U17072 ( .A1(n13813), .A2(n13812), .ZN(n14923) );
  AOI22_X1 U17073 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11564), .B1(
        n11602), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13817) );
  AOI22_X1 U17074 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13816) );
  AOI22_X1 U17075 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11597), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13815) );
  AOI22_X1 U17076 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11611), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13814) );
  NAND4_X1 U17077 ( .A1(n13817), .A2(n13816), .A3(n13815), .A4(n13814), .ZN(
        n13823) );
  AOI22_X1 U17078 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12120), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13821) );
  AOI22_X1 U17079 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n13828), .ZN(n13820) );
  AOI22_X1 U17080 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12170), .B1(
        n12169), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13819) );
  AOI22_X1 U17081 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13818) );
  NAND4_X1 U17082 ( .A1(n13821), .A2(n13820), .A3(n13819), .A4(n13818), .ZN(
        n13822) );
  OR2_X1 U17083 ( .A1(n13823), .A2(n13822), .ZN(n16106) );
  AOI22_X1 U17084 ( .A1(n11602), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13827) );
  AOI22_X1 U17085 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13826) );
  AOI22_X1 U17086 ( .A1(n11597), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13825) );
  AOI22_X1 U17087 ( .A1(n13113), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11611), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13824) );
  NAND4_X1 U17088 ( .A1(n13827), .A2(n13826), .A3(n13825), .A4(n13824), .ZN(
        n13838) );
  AOI22_X1 U17089 ( .A1(n12120), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13836) );
  AOI22_X1 U17090 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13828), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13835) );
  AOI22_X1 U17091 ( .A1(n12169), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13834) );
  INV_X1 U17092 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13829) );
  OAI22_X1 U17093 ( .A1(n13831), .A2(n14005), .B1(n13830), .B2(n13829), .ZN(
        n13832) );
  INV_X1 U17094 ( .A(n13832), .ZN(n13833) );
  NAND4_X1 U17095 ( .A1(n13836), .A2(n13835), .A3(n13834), .A4(n13833), .ZN(
        n13837) );
  OR2_X1 U17096 ( .A1(n13838), .A2(n13837), .ZN(n14915) );
  AOI22_X1 U17097 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11564), .B1(
        n11602), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13842) );
  AOI22_X1 U17098 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13841) );
  AOI22_X1 U17099 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11597), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13840) );
  AOI22_X1 U17100 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11611), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13839) );
  NAND4_X1 U17101 ( .A1(n13842), .A2(n13841), .A3(n13840), .A4(n13839), .ZN(
        n13848) );
  AOI22_X1 U17102 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12120), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13846) );
  AOI22_X1 U17103 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n13828), .ZN(n13845) );
  AOI22_X1 U17104 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12170), .B1(
        n12169), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13844) );
  AOI22_X1 U17105 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13843) );
  NAND4_X1 U17106 ( .A1(n13846), .A2(n13845), .A3(n13844), .A4(n13843), .ZN(
        n13847) );
  NOR2_X1 U17107 ( .A1(n13848), .A2(n13847), .ZN(n16103) );
  INV_X1 U17108 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13852) );
  INV_X1 U17109 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13851) );
  OAI22_X1 U17110 ( .A1(n13849), .A2(n13852), .B1(n13850), .B2(n13851), .ZN(
        n13857) );
  INV_X1 U17111 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13855) );
  INV_X1 U17112 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n19466) );
  OAI22_X1 U17113 ( .A1(n13853), .A2(n13855), .B1(n13854), .B2(n19466), .ZN(
        n13856) );
  NOR2_X1 U17114 ( .A1(n13857), .A2(n13856), .ZN(n13860) );
  XNOR2_X1 U17115 ( .A(n13115), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14050) );
  AOI22_X1 U17116 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13859) );
  AOI22_X1 U17117 ( .A1(n14052), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11408), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13858) );
  NAND4_X1 U17118 ( .A1(n13860), .A2(n14050), .A3(n13859), .A4(n13858), .ZN(
        n13871) );
  INV_X1 U17119 ( .A(n11409), .ZN(n14016) );
  INV_X1 U17120 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13862) );
  INV_X1 U17121 ( .A(n11523), .ZN(n14025) );
  INV_X1 U17122 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13861) );
  OAI22_X1 U17123 ( .A1(n14016), .A2(n13862), .B1(n14025), .B2(n13861), .ZN(
        n13866) );
  INV_X1 U17124 ( .A(n14052), .ZN(n14029) );
  INV_X1 U17125 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13864) );
  INV_X1 U17126 ( .A(n11408), .ZN(n14027) );
  INV_X1 U17127 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13863) );
  OAI22_X1 U17128 ( .A1(n14029), .A2(n13864), .B1(n14027), .B2(n13863), .ZN(
        n13865) );
  NOR2_X1 U17129 ( .A1(n13866), .A2(n13865), .ZN(n13869) );
  AOI22_X1 U17130 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13868) );
  AOI22_X1 U17131 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13867) );
  INV_X1 U17132 ( .A(n14050), .ZN(n14046) );
  NAND4_X1 U17133 ( .A1(n13869), .A2(n13868), .A3(n13867), .A4(n14046), .ZN(
        n13870) );
  NAND2_X1 U17134 ( .A1(n13871), .A2(n13870), .ZN(n13905) );
  NOR2_X1 U17135 ( .A1(n11420), .A2(n13905), .ZN(n13883) );
  AOI22_X1 U17136 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11564), .B1(
        n11602), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13875) );
  AOI22_X1 U17137 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11646), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13874) );
  AOI22_X1 U17138 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11597), .B1(
        n12121), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13873) );
  AOI22_X1 U17139 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11611), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13872) );
  NAND4_X1 U17140 ( .A1(n13875), .A2(n13874), .A3(n13873), .A4(n13872), .ZN(
        n13882) );
  AOI22_X1 U17141 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12120), .B1(
        n13703), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13880) );
  AOI22_X1 U17142 ( .A1(n13876), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n13828), .ZN(n13879) );
  AOI22_X1 U17143 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12170), .B1(
        n12169), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13878) );
  AOI22_X1 U17144 ( .A1(n12139), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12140), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13877) );
  NAND4_X1 U17145 ( .A1(n13880), .A2(n13879), .A3(n13878), .A4(n13877), .ZN(
        n13881) );
  OR2_X1 U17146 ( .A1(n13882), .A2(n13881), .ZN(n13907) );
  XNOR2_X1 U17147 ( .A(n13883), .B(n13907), .ZN(n13884) );
  XNOR2_X1 U17148 ( .A(n16102), .B(n13884), .ZN(n14907) );
  NOR2_X1 U17149 ( .A1(n19890), .A2(n13905), .ZN(n14909) );
  NAND2_X1 U17150 ( .A1(n14907), .A2(n14909), .ZN(n14908) );
  INV_X1 U17151 ( .A(n16102), .ZN(n13885) );
  OAI22_X1 U17152 ( .A1(n14016), .A2(n13887), .B1(n14027), .B2(n13886), .ZN(
        n13891) );
  INV_X1 U17153 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13888) );
  OAI22_X1 U17154 ( .A1(n14029), .A2(n13889), .B1(n14025), .B2(n13888), .ZN(
        n13890) );
  NOR2_X1 U17155 ( .A1(n13891), .A2(n13890), .ZN(n13894) );
  AOI22_X1 U17156 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13893) );
  AOI22_X1 U17157 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13892) );
  NAND4_X1 U17158 ( .A1(n13894), .A2(n13893), .A3(n13892), .A4(n14046), .ZN(
        n13904) );
  OAI22_X1 U17159 ( .A1(n14016), .A2(n13896), .B1(n14027), .B2(n13895), .ZN(
        n13899) );
  OAI22_X1 U17160 ( .A1(n14029), .A2(n12141), .B1(n14025), .B2(n13897), .ZN(
        n13898) );
  NOR2_X1 U17161 ( .A1(n13899), .A2(n13898), .ZN(n13902) );
  AOI22_X1 U17162 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13901) );
  AOI22_X1 U17163 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13900) );
  NAND4_X1 U17164 ( .A1(n13902), .A2(n14050), .A3(n13901), .A4(n13900), .ZN(
        n13903) );
  NAND2_X1 U17165 ( .A1(n13904), .A2(n13903), .ZN(n13911) );
  INV_X1 U17166 ( .A(n13905), .ZN(n13906) );
  NAND2_X1 U17167 ( .A1(n13907), .A2(n13906), .ZN(n13912) );
  INV_X1 U17168 ( .A(n13912), .ZN(n13908) );
  NAND2_X1 U17169 ( .A1(n13987), .A2(n13908), .ZN(n13910) );
  NOR3_X1 U17170 ( .A1(n19119), .A2(n13912), .A3(n13911), .ZN(n13909) );
  AOI21_X1 U17171 ( .B1(n13911), .B2(n13910), .A(n13909), .ZN(n14899) );
  NOR2_X1 U17172 ( .A1(n13912), .A2(n13911), .ZN(n13933) );
  INV_X1 U17173 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13914) );
  INV_X1 U17174 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13913) );
  OAI22_X1 U17175 ( .A1(n14016), .A2(n13914), .B1(n14027), .B2(n13913), .ZN(
        n13918) );
  INV_X1 U17176 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13916) );
  INV_X1 U17177 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13915) );
  OAI22_X1 U17178 ( .A1(n14029), .A2(n13916), .B1(n14025), .B2(n13915), .ZN(
        n13917) );
  NOR2_X1 U17179 ( .A1(n13918), .A2(n13917), .ZN(n13921) );
  AOI22_X1 U17180 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13920) );
  AOI22_X1 U17181 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13919) );
  NAND4_X1 U17182 ( .A1(n13921), .A2(n13920), .A3(n13919), .A4(n14046), .ZN(
        n13932) );
  INV_X1 U17183 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13923) );
  INV_X1 U17184 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13922) );
  OAI22_X1 U17185 ( .A1(n14016), .A2(n13923), .B1(n14027), .B2(n13922), .ZN(
        n13927) );
  INV_X1 U17186 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13925) );
  INV_X1 U17187 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13924) );
  OAI22_X1 U17188 ( .A1(n14029), .A2(n13925), .B1(n14025), .B2(n13924), .ZN(
        n13926) );
  NOR2_X1 U17189 ( .A1(n13927), .A2(n13926), .ZN(n13930) );
  AOI22_X1 U17190 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13929) );
  AOI22_X1 U17191 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13928) );
  NAND4_X1 U17192 ( .A1(n13930), .A2(n14050), .A3(n13929), .A4(n13928), .ZN(
        n13931) );
  AND2_X1 U17193 ( .A1(n13932), .A2(n13931), .ZN(n13935) );
  NAND2_X1 U17194 ( .A1(n13933), .A2(n13935), .ZN(n13959) );
  OAI211_X1 U17195 ( .C1(n13933), .C2(n13935), .A(n13987), .B(n13959), .ZN(
        n13937) );
  INV_X1 U17196 ( .A(n13937), .ZN(n13934) );
  INV_X1 U17197 ( .A(n13935), .ZN(n13936) );
  NOR2_X1 U17198 ( .A1(n19890), .A2(n13936), .ZN(n14893) );
  NAND2_X1 U17199 ( .A1(n14891), .A2(n14893), .ZN(n14892) );
  OAI22_X1 U17200 ( .A1(n14016), .A2(n13939), .B1(n14027), .B2(n13938), .ZN(
        n13943) );
  INV_X1 U17201 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13940) );
  OAI22_X1 U17202 ( .A1(n14029), .A2(n13941), .B1(n14025), .B2(n13940), .ZN(
        n13942) );
  NOR2_X1 U17203 ( .A1(n13943), .A2(n13942), .ZN(n13946) );
  AOI22_X1 U17204 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13945) );
  AOI22_X1 U17205 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13944) );
  NAND4_X1 U17206 ( .A1(n13946), .A2(n13945), .A3(n13944), .A4(n14046), .ZN(
        n13957) );
  OAI22_X1 U17207 ( .A1(n14016), .A2(n13948), .B1(n14027), .B2(n13947), .ZN(
        n13952) );
  OAI22_X1 U17208 ( .A1(n14029), .A2(n13950), .B1(n14025), .B2(n13949), .ZN(
        n13951) );
  NOR2_X1 U17209 ( .A1(n13952), .A2(n13951), .ZN(n13955) );
  AOI22_X1 U17210 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13954) );
  AOI22_X1 U17211 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13953) );
  NAND4_X1 U17212 ( .A1(n13955), .A2(n14050), .A3(n13954), .A4(n13953), .ZN(
        n13956) );
  NAND2_X1 U17213 ( .A1(n13957), .A2(n13956), .ZN(n13962) );
  AOI21_X1 U17214 ( .B1(n13959), .B2(n13962), .A(n13958), .ZN(n13960) );
  NAND2_X1 U17215 ( .A1(n13960), .A2(n13986), .ZN(n13965) );
  INV_X1 U17216 ( .A(n13965), .ZN(n13961) );
  INV_X1 U17217 ( .A(n13962), .ZN(n13963) );
  NAND2_X1 U17218 ( .A1(n19119), .A2(n13963), .ZN(n14884) );
  INV_X1 U17219 ( .A(n13964), .ZN(n13966) );
  INV_X1 U17220 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13968) );
  INV_X1 U17221 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13967) );
  OAI22_X1 U17222 ( .A1(n14016), .A2(n13968), .B1(n14027), .B2(n13967), .ZN(
        n13972) );
  INV_X1 U17223 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13970) );
  INV_X1 U17224 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13969) );
  OAI22_X1 U17225 ( .A1(n14029), .A2(n13970), .B1(n14025), .B2(n13969), .ZN(
        n13971) );
  NOR2_X1 U17226 ( .A1(n13972), .A2(n13971), .ZN(n13975) );
  AOI22_X1 U17227 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13974) );
  AOI22_X1 U17228 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13973) );
  NAND4_X1 U17229 ( .A1(n13975), .A2(n13974), .A3(n13973), .A4(n14046), .ZN(
        n13985) );
  INV_X1 U17230 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13976) );
  OAI22_X1 U17231 ( .A1(n14016), .A2(n13976), .B1(n14027), .B2(n20861), .ZN(
        n13980) );
  INV_X1 U17232 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13978) );
  INV_X1 U17233 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13977) );
  OAI22_X1 U17234 ( .A1(n14029), .A2(n13978), .B1(n14025), .B2(n13977), .ZN(
        n13979) );
  NOR2_X1 U17235 ( .A1(n13980), .A2(n13979), .ZN(n13983) );
  AOI22_X1 U17236 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13982) );
  AOI22_X1 U17237 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13981) );
  NAND4_X1 U17238 ( .A1(n13983), .A2(n14050), .A3(n13982), .A4(n13981), .ZN(
        n13984) );
  NAND2_X1 U17239 ( .A1(n13985), .A2(n13984), .ZN(n13991) );
  INV_X1 U17240 ( .A(n13991), .ZN(n13989) );
  INV_X1 U17241 ( .A(n13986), .ZN(n13988) );
  OR2_X1 U17242 ( .A1(n13986), .A2(n13991), .ZN(n14037) );
  OAI211_X1 U17243 ( .C1(n13989), .C2(n13988), .A(n14037), .B(n13987), .ZN(
        n13990) );
  NOR2_X1 U17244 ( .A1(n19890), .A2(n13991), .ZN(n14879) );
  NAND2_X1 U17245 ( .A1(n14876), .A2(n14879), .ZN(n14878) );
  INV_X1 U17246 ( .A(n13992), .ZN(n14013) );
  OAI22_X1 U17247 ( .A1(n14016), .A2(n13994), .B1(n14027), .B2(n13993), .ZN(
        n13998) );
  INV_X1 U17248 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13995) );
  OAI22_X1 U17249 ( .A1(n14029), .A2(n13996), .B1(n14025), .B2(n13995), .ZN(
        n13997) );
  NOR2_X1 U17250 ( .A1(n13998), .A2(n13997), .ZN(n14001) );
  AOI22_X1 U17251 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14000) );
  AOI22_X1 U17252 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13999) );
  NAND4_X1 U17253 ( .A1(n14001), .A2(n14000), .A3(n13999), .A4(n14046), .ZN(
        n14012) );
  OAI22_X1 U17254 ( .A1(n14016), .A2(n14003), .B1(n14027), .B2(n14002), .ZN(
        n14007) );
  OAI22_X1 U17255 ( .A1(n14029), .A2(n14005), .B1(n14025), .B2(n14004), .ZN(
        n14006) );
  NOR2_X1 U17256 ( .A1(n14007), .A2(n14006), .ZN(n14010) );
  AOI22_X1 U17257 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14009) );
  AOI22_X1 U17258 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14008) );
  NAND4_X1 U17259 ( .A1(n14010), .A2(n14050), .A3(n14009), .A4(n14008), .ZN(
        n14011) );
  NAND2_X1 U17260 ( .A1(n14012), .A2(n14011), .ZN(n14870) );
  OAI22_X1 U17261 ( .A1(n14016), .A2(n14015), .B1(n14027), .B2(n14014), .ZN(
        n14020) );
  INV_X1 U17262 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14017) );
  OAI22_X1 U17263 ( .A1(n14029), .A2(n14018), .B1(n14025), .B2(n14017), .ZN(
        n14019) );
  NOR2_X1 U17264 ( .A1(n14020), .A2(n14019), .ZN(n14023) );
  AOI22_X1 U17265 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14022) );
  AOI22_X1 U17266 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14021) );
  NAND4_X1 U17267 ( .A1(n14023), .A2(n14022), .A3(n14021), .A4(n14046), .ZN(
        n14036) );
  OAI22_X1 U17268 ( .A1(n13849), .A2(n11714), .B1(n14025), .B2(n14024), .ZN(
        n14031) );
  OAI22_X1 U17269 ( .A1(n14029), .A2(n14028), .B1(n14027), .B2(n14026), .ZN(
        n14030) );
  NOR2_X1 U17270 ( .A1(n14031), .A2(n14030), .ZN(n14034) );
  INV_X1 U17271 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n20921) );
  AOI22_X1 U17272 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14033) );
  AOI22_X1 U17273 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14032) );
  NAND4_X1 U17274 ( .A1(n14034), .A2(n14050), .A3(n14033), .A4(n14032), .ZN(
        n14035) );
  NAND2_X1 U17275 ( .A1(n14036), .A2(n14035), .ZN(n14041) );
  INV_X1 U17276 ( .A(n14037), .ZN(n14869) );
  INV_X1 U17277 ( .A(n14870), .ZN(n14038) );
  AND2_X1 U17278 ( .A1(n19890), .A2(n14038), .ZN(n14039) );
  NAND2_X1 U17279 ( .A1(n14869), .A2(n14039), .ZN(n14040) );
  NOR2_X1 U17280 ( .A1(n14040), .A2(n14041), .ZN(n14042) );
  AOI21_X1 U17281 ( .B1(n14041), .B2(n14040), .A(n14042), .ZN(n14865) );
  INV_X1 U17282 ( .A(n14042), .ZN(n14043) );
  AOI22_X1 U17283 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14052), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14045) );
  AOI22_X1 U17284 ( .A1(n11408), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14044) );
  NAND2_X1 U17285 ( .A1(n14045), .A2(n14044), .ZN(n14058) );
  AOI22_X1 U17286 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14048) );
  AOI22_X1 U17287 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14047) );
  NAND3_X1 U17288 ( .A1(n14048), .A2(n14047), .A3(n14046), .ZN(n14057) );
  AOI22_X1 U17289 ( .A1(n11409), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9588), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14051) );
  AOI22_X1 U17290 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11529), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14049) );
  NAND3_X1 U17291 ( .A1(n14051), .A2(n14050), .A3(n14049), .ZN(n14056) );
  AOI22_X1 U17292 ( .A1(n11522), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14052), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14054) );
  AOI22_X1 U17293 ( .A1(n11408), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9607), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14053) );
  NAND2_X1 U17294 ( .A1(n14054), .A2(n14053), .ZN(n14055) );
  OAI22_X1 U17295 ( .A1(n14058), .A2(n14057), .B1(n14056), .B2(n14055), .ZN(
        n14059) );
  INV_X1 U17296 ( .A(n14059), .ZN(n14060) );
  NOR2_X1 U17297 ( .A1(n16032), .A2(n18983), .ZN(n14062) );
  AOI21_X1 U17298 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n18983), .A(n14062), .ZN(
        n14063) );
  OAI21_X1 U17299 ( .B1(n14068), .B2(n18984), .A(n14063), .ZN(P2_U2857) );
  AOI22_X1 U17300 ( .A1(n20782), .A2(n18993), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n20780), .ZN(n14065) );
  AOI22_X1 U17301 ( .A1(n20784), .A2(BUF2_REG_30__SCAN_IN), .B1(n20783), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n14064) );
  OAI211_X1 U17302 ( .C1(n16023), .C2(n20787), .A(n14065), .B(n14064), .ZN(
        n14066) );
  INV_X1 U17303 ( .A(n14066), .ZN(n14067) );
  OAI21_X1 U17304 ( .B1(n14068), .B2(n14996), .A(n14067), .ZN(P2_U2889) );
  INV_X1 U17305 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14072) );
  NOR3_X1 U17306 ( .A1(n14366), .A2(n14069), .A3(n20132), .ZN(n14323) );
  AOI22_X1 U17307 ( .A1(n14323), .A2(n14070), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n14366), .ZN(n14071) );
  OAI21_X1 U17308 ( .B1(n14072), .B2(n14326), .A(n14071), .ZN(n14073) );
  AOI21_X1 U17309 ( .B1(n14355), .B2(DATAI_30_), .A(n14073), .ZN(n14074) );
  OAI21_X1 U17310 ( .B1(n14086), .B2(n14370), .A(n14074), .ZN(P1_U2874) );
  NAND2_X1 U17311 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14094) );
  INV_X1 U17312 ( .A(n14094), .ZN(n14077) );
  AND2_X1 U17313 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14079) );
  INV_X1 U17314 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20731) );
  INV_X1 U17315 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20727) );
  INV_X1 U17316 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20724) );
  INV_X1 U17317 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20721) );
  NAND2_X1 U17318 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15806) );
  NOR4_X1 U17319 ( .A1(n20721), .A2(n15837), .A3(n14075), .A4(n15806), .ZN(
        n15787) );
  NAND2_X1 U17320 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15787), .ZN(n15786) );
  NOR2_X1 U17321 ( .A1(n20724), .A2(n15786), .ZN(n15777) );
  NAND2_X1 U17322 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n15777), .ZN(n15767) );
  NOR2_X1 U17323 ( .A1(n20727), .A2(n15767), .ZN(n14185) );
  NAND2_X1 U17324 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n14185), .ZN(n14175) );
  NOR2_X1 U17325 ( .A1(n20731), .A2(n14175), .ZN(n14162) );
  AND2_X1 U17326 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n14162), .ZN(n14150) );
  AND2_X1 U17327 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n14150), .ZN(n14134) );
  NAND2_X1 U17328 ( .A1(n14134), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14078) );
  INV_X1 U17329 ( .A(n14078), .ZN(n14122) );
  NAND3_X1 U17330 ( .A1(n14217), .A2(n14079), .A3(n14122), .ZN(n14076) );
  NAND2_X1 U17331 ( .A1(n15834), .A2(n14076), .ZN(n14116) );
  OAI21_X1 U17332 ( .B1(n14077), .B2(n15838), .A(n14116), .ZN(n14097) );
  NOR2_X1 U17333 ( .A1(n15838), .A2(n14078), .ZN(n14123) );
  NAND2_X1 U17334 ( .A1(n14123), .A2(n14079), .ZN(n14101) );
  INV_X1 U17335 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20743) );
  INV_X1 U17336 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14080) );
  OAI21_X1 U17337 ( .B1(n14101), .B2(n20743), .A(n14080), .ZN(n14085) );
  INV_X1 U17338 ( .A(n14081), .ZN(n14083) );
  AOI22_X1 U17339 ( .A1(P1_EBX_REG_30__SCAN_IN), .A2(n19982), .B1(n19986), 
        .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14082) );
  OAI21_X1 U17340 ( .B1(n14083), .B2(n19981), .A(n14082), .ZN(n14084) );
  MUX2_X1 U17341 ( .A(n14088), .B(n14087), .S(n9660), .Z(n14092) );
  AOI22_X1 U17342 ( .A1(n14090), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n14089), .ZN(n14091) );
  NAND2_X1 U17343 ( .A1(n14379), .A2(n19955), .ZN(n14099) );
  INV_X1 U17344 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14240) );
  OAI22_X1 U17345 ( .A1(n19928), .A2(n14093), .B1(n14240), .B2(n19936), .ZN(
        n14096) );
  NOR3_X1 U17346 ( .A1(n14101), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14094), 
        .ZN(n14095) );
  AOI211_X1 U17347 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14097), .A(n14096), 
        .B(n14095), .ZN(n14098) );
  OAI211_X1 U17348 ( .C1(n14534), .C2(n19971), .A(n14099), .B(n14098), .ZN(
        P1_U2809) );
  NAND2_X1 U17349 ( .A1(n14386), .A2(n19955), .ZN(n14106) );
  INV_X1 U17350 ( .A(n14116), .ZN(n14104) );
  AOI22_X1 U17351 ( .A1(n19982), .A2(P1_EBX_REG_29__SCAN_IN), .B1(n19986), 
        .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14100) );
  OAI21_X1 U17352 ( .B1(n14384), .B2(n19981), .A(n14100), .ZN(n14103) );
  NOR2_X1 U17353 ( .A1(n14101), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14102) );
  AOI211_X1 U17354 ( .C1(n14104), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14103), 
        .B(n14102), .ZN(n14105) );
  OAI211_X1 U17355 ( .C1(n19971), .C2(n14564), .A(n14106), .B(n14105), .ZN(
        P1_U2811) );
  OAI21_X2 U17356 ( .B1(n14107), .B2(n14109), .A(n14108), .ZN(n14396) );
  INV_X1 U17357 ( .A(n14110), .ZN(n14113) );
  INV_X1 U17358 ( .A(n14127), .ZN(n14112) );
  AOI21_X1 U17359 ( .B1(n14113), .B2(n14112), .A(n14111), .ZN(n14575) );
  AOI21_X1 U17360 ( .B1(n14123), .B2(P1_REIP_REG_27__SCAN_IN), .A(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14117) );
  AOI22_X1 U17361 ( .A1(n19982), .A2(P1_EBX_REG_28__SCAN_IN), .B1(n19986), 
        .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14115) );
  NAND2_X1 U17362 ( .A1(n19993), .A2(n14399), .ZN(n14114) );
  OAI211_X1 U17363 ( .C1(n14117), .C2(n14116), .A(n14115), .B(n14114), .ZN(
        n14118) );
  AOI21_X1 U17364 ( .B1(n14575), .B2(n19983), .A(n14118), .ZN(n14119) );
  OAI21_X1 U17365 ( .B1(n14396), .B2(n15810), .A(n14119), .ZN(P1_U2812) );
  AOI21_X1 U17366 ( .B1(n14121), .B2(n14132), .A(n14107), .ZN(n14408) );
  INV_X1 U17367 ( .A(n14408), .ZN(n14312) );
  OR2_X1 U17368 ( .A1(n15838), .A2(n14122), .ZN(n14137) );
  NAND2_X1 U17369 ( .A1(n14137), .A2(n14217), .ZN(n14143) );
  AOI22_X1 U17370 ( .A1(n19982), .A2(P1_EBX_REG_27__SCAN_IN), .B1(n19986), 
        .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14125) );
  INV_X1 U17371 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20738) );
  NAND2_X1 U17372 ( .A1(n14123), .A2(n20738), .ZN(n14124) );
  OAI211_X1 U17373 ( .C1(n19981), .C2(n14406), .A(n14125), .B(n14124), .ZN(
        n14126) );
  AOI21_X1 U17374 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n14143), .A(n14126), 
        .ZN(n14130) );
  AOI21_X1 U17375 ( .B1(n14128), .B2(n9681), .A(n14127), .ZN(n14583) );
  NAND2_X1 U17376 ( .A1(n14583), .A2(n19983), .ZN(n14129) );
  OAI211_X1 U17377 ( .C1(n14312), .C2(n15810), .A(n14130), .B(n14129), .ZN(
        P1_U2813) );
  OAI21_X1 U17378 ( .B1(n14131), .B2(n14133), .A(n14132), .ZN(n14414) );
  INV_X1 U17379 ( .A(n14134), .ZN(n14138) );
  OAI22_X1 U17380 ( .A1(n19928), .A2(n14413), .B1(n19936), .B2(n14243), .ZN(
        n14135) );
  AOI21_X1 U17381 ( .B1(n14417), .B2(n19993), .A(n14135), .ZN(n14136) );
  OAI21_X1 U17382 ( .B1(n14138), .B2(n14137), .A(n14136), .ZN(n14142) );
  NAND2_X1 U17383 ( .A1(n9626), .A2(n14139), .ZN(n14140) );
  NAND2_X1 U17384 ( .A1(n9681), .A2(n14140), .ZN(n14588) );
  NOR2_X1 U17385 ( .A1(n14588), .A2(n19971), .ZN(n14141) );
  AOI211_X1 U17386 ( .C1(P1_REIP_REG_26__SCAN_IN), .C2(n14143), .A(n14142), 
        .B(n14141), .ZN(n14144) );
  OAI21_X1 U17387 ( .B1(n14414), .B2(n15810), .A(n14144), .ZN(P1_U2814) );
  NAND2_X1 U17388 ( .A1(n14157), .A2(n14145), .ZN(n14146) );
  NAND2_X1 U17389 ( .A1(n9626), .A2(n14146), .ZN(n14598) );
  AOI21_X1 U17390 ( .B1(n14148), .B2(n14147), .A(n14131), .ZN(n14426) );
  NAND2_X1 U17391 ( .A1(n14426), .A2(n19955), .ZN(n14156) );
  INV_X1 U17392 ( .A(n15834), .ZN(n14218) );
  AOI21_X1 U17393 ( .B1(n14162), .B2(n14217), .A(n14218), .ZN(n14176) );
  NAND2_X1 U17394 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14149) );
  OAI21_X1 U17395 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n14150), .A(n14149), 
        .ZN(n14151) );
  INV_X1 U17396 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14244) );
  OAI22_X1 U17397 ( .A1(n15838), .A2(n14151), .B1(n19936), .B2(n14244), .ZN(
        n14154) );
  OAI22_X1 U17398 ( .A1(n14152), .A2(n19928), .B1(n19981), .B2(n14424), .ZN(
        n14153) );
  AOI211_X1 U17399 ( .C1(n14176), .C2(P1_REIP_REG_25__SCAN_IN), .A(n14154), 
        .B(n14153), .ZN(n14155) );
  OAI211_X1 U17400 ( .C1(n19971), .C2(n14598), .A(n14156), .B(n14155), .ZN(
        P1_U2815) );
  OAI21_X1 U17401 ( .B1(n14173), .B2(n14158), .A(n14157), .ZN(n14606) );
  OAI21_X1 U17402 ( .B1(n14159), .B2(n14160), .A(n14147), .ZN(n14433) );
  INV_X1 U17403 ( .A(n14433), .ZN(n14161) );
  NAND2_X1 U17404 ( .A1(n14161), .A2(n19955), .ZN(n14168) );
  INV_X1 U17405 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20734) );
  NAND2_X1 U17406 ( .A1(n20734), .A2(n14162), .ZN(n14163) );
  INV_X1 U17407 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14245) );
  OAI22_X1 U17408 ( .A1(n15838), .A2(n14163), .B1(n19936), .B2(n14245), .ZN(
        n14166) );
  INV_X1 U17409 ( .A(n14436), .ZN(n14164) );
  OAI22_X1 U17410 ( .A1(n14432), .A2(n19928), .B1(n19981), .B2(n14164), .ZN(
        n14165) );
  AOI211_X1 U17411 ( .C1(n14176), .C2(P1_REIP_REG_24__SCAN_IN), .A(n14166), 
        .B(n14165), .ZN(n14167) );
  OAI211_X1 U17412 ( .C1(n19971), .C2(n14606), .A(n14168), .B(n14167), .ZN(
        P1_U2816) );
  AOI21_X1 U17413 ( .B1(n14170), .B2(n14169), .A(n14159), .ZN(n14442) );
  INV_X1 U17414 ( .A(n14442), .ZN(n14332) );
  INV_X1 U17415 ( .A(n14254), .ZN(n14172) );
  AOI21_X1 U17416 ( .B1(n14172), .B2(n14184), .A(n14171), .ZN(n14174) );
  NOR2_X1 U17417 ( .A1(n14174), .A2(n14173), .ZN(n14621) );
  NOR2_X1 U17418 ( .A1(n15838), .A2(n14175), .ZN(n14177) );
  OAI21_X1 U17419 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(n14177), .A(n14176), 
        .ZN(n14179) );
  AOI22_X1 U17420 ( .A1(n19982), .A2(P1_EBX_REG_23__SCAN_IN), .B1(n19986), 
        .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14178) );
  OAI211_X1 U17421 ( .C1(n19981), .C2(n14440), .A(n14179), .B(n14178), .ZN(
        n14180) );
  AOI21_X1 U17422 ( .B1(n14621), .B2(n19983), .A(n14180), .ZN(n14181) );
  OAI21_X1 U17423 ( .B1(n14332), .B2(n15810), .A(n14181), .ZN(P1_U2817) );
  OAI21_X1 U17424 ( .B1(n14182), .B2(n14183), .A(n14169), .ZN(n14452) );
  XNOR2_X1 U17425 ( .A(n14254), .B(n14184), .ZN(n14631) );
  AOI21_X1 U17426 ( .B1(n19925), .B2(n15767), .A(n14228), .ZN(n15785) );
  NAND2_X1 U17427 ( .A1(n19925), .A2(n20727), .ZN(n15768) );
  INV_X1 U17428 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20729) );
  AOI21_X1 U17429 ( .B1(n15785), .B2(n15768), .A(n20729), .ZN(n14190) );
  NAND2_X1 U17430 ( .A1(n19925), .A2(n14185), .ZN(n14188) );
  AOI22_X1 U17431 ( .A1(n19982), .A2(P1_EBX_REG_22__SCAN_IN), .B1(n19986), 
        .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14187) );
  NAND2_X1 U17432 ( .A1(n19993), .A2(n14446), .ZN(n14186) );
  OAI211_X1 U17433 ( .C1(n14188), .C2(P1_REIP_REG_22__SCAN_IN), .A(n14187), 
        .B(n14186), .ZN(n14189) );
  AOI211_X1 U17434 ( .C1(n14631), .C2(n19983), .A(n14190), .B(n14189), .ZN(
        n14191) );
  OAI21_X1 U17435 ( .B1(n14452), .B2(n15810), .A(n14191), .ZN(P1_U2818) );
  NOR2_X1 U17436 ( .A1(n9656), .A2(n14193), .ZN(n14194) );
  OR3_X1 U17437 ( .A1(n20716), .A2(n20714), .A3(n14213), .ZN(n15824) );
  OAI21_X1 U17438 ( .B1(n15806), .B2(n15824), .A(n20721), .ZN(n14201) );
  OAI21_X1 U17439 ( .B1(n15838), .B2(n15787), .A(n14217), .ZN(n15799) );
  NAND2_X1 U17440 ( .A1(n14195), .A2(n14196), .ZN(n14197) );
  NAND2_X1 U17441 ( .A1(n14268), .A2(n14197), .ZN(n15925) );
  NOR2_X1 U17442 ( .A1(n15925), .A2(n19971), .ZN(n14200) );
  INV_X1 U17443 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n20838) );
  AOI22_X1 U17444 ( .A1(n19986), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n19993), .B2(n15872), .ZN(n14198) );
  OAI211_X1 U17445 ( .C1(n20838), .C2(n19936), .A(n14198), .B(n19962), .ZN(
        n14199) );
  AOI211_X1 U17446 ( .C1(n14201), .C2(n15799), .A(n14200), .B(n14199), .ZN(
        n14202) );
  OAI21_X1 U17447 ( .B1(n15871), .B2(n15810), .A(n14202), .ZN(P1_U2823) );
  INV_X1 U17448 ( .A(n14203), .ZN(n14204) );
  AOI21_X1 U17449 ( .B1(n14205), .B2(n14204), .A(n13769), .ZN(n14512) );
  INV_X1 U17450 ( .A(n14512), .ZN(n14362) );
  OAI21_X1 U17451 ( .B1(n14294), .B2(n14207), .A(n14206), .ZN(n14209) );
  AND2_X1 U17452 ( .A1(n14209), .A2(n14208), .ZN(n15941) );
  AOI22_X1 U17453 ( .A1(n15941), .A2(n19983), .B1(n19982), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14210) );
  OAI211_X1 U17454 ( .C1(n19928), .C2(n14211), .A(n14210), .B(n19962), .ZN(
        n14215) );
  NAND2_X1 U17455 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14212) );
  OAI21_X1 U17456 ( .B1(n14212), .B2(n15833), .A(n15834), .ZN(n15826) );
  AOI22_X1 U17457 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n15826), .B1(n14213), 
        .B2(n20714), .ZN(n14214) );
  AOI211_X1 U17458 ( .C1(n14508), .C2(n19993), .A(n14215), .B(n14214), .ZN(
        n14216) );
  OAI21_X1 U17459 ( .B1(n14362), .B2(n15810), .A(n14216), .ZN(P1_U2827) );
  NAND2_X1 U17460 ( .A1(n19924), .A2(n14217), .ZN(n14219) );
  NAND2_X1 U17461 ( .A1(n15834), .A2(n14219), .ZN(n19975) );
  OAI21_X1 U17462 ( .B1(n19926), .B2(n14218), .A(n19975), .ZN(n15844) );
  OAI21_X1 U17463 ( .B1(n19941), .B2(n14219), .A(n15834), .ZN(n19950) );
  NAND2_X1 U17464 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19950), .ZN(n19942) );
  NAND2_X1 U17465 ( .A1(n20706), .A2(n19942), .ZN(n14224) );
  OAI22_X1 U17466 ( .A1(n10527), .A2(n19928), .B1(n19981), .B2(n14220), .ZN(
        n14221) );
  AOI211_X1 U17467 ( .C1(n19982), .C2(P1_EBX_REG_8__SCAN_IN), .A(n19973), .B(
        n14221), .ZN(n14222) );
  OAI21_X1 U17468 ( .B1(n19971), .B2(n15984), .A(n14222), .ZN(n14223) );
  AOI21_X1 U17469 ( .B1(n15844), .B2(n14224), .A(n14223), .ZN(n14225) );
  OAI21_X1 U17470 ( .B1(n14226), .B2(n15810), .A(n14225), .ZN(P1_U2832) );
  NOR2_X1 U17471 ( .A1(n15838), .A2(n14227), .ZN(n19985) );
  INV_X1 U17472 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20695) );
  NAND2_X1 U17473 ( .A1(n19985), .A2(n20695), .ZN(n14235) );
  AOI22_X1 U17474 ( .A1(n19983), .A2(n20064), .B1(n19986), .B2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14234) );
  AOI21_X1 U17475 ( .B1(n19925), .B2(n14227), .A(n14228), .ZN(n19997) );
  OAI22_X1 U17476 ( .A1(n19936), .A2(n11242), .B1(n20695), .B2(n19997), .ZN(
        n14229) );
  INV_X1 U17477 ( .A(n14229), .ZN(n14233) );
  INV_X1 U17478 ( .A(n14230), .ZN(n14231) );
  NAND2_X1 U17479 ( .A1(n19993), .A2(n14231), .ZN(n14232) );
  NAND4_X1 U17480 ( .A1(n14235), .A2(n14234), .A3(n14233), .A4(n14232), .ZN(
        n14238) );
  NOR2_X1 U17481 ( .A1(n14236), .A2(n19990), .ZN(n14237) );
  AOI211_X1 U17482 ( .C1(n19987), .C2(n20103), .A(n14238), .B(n14237), .ZN(
        n14239) );
  INV_X1 U17483 ( .A(n14239), .ZN(P1_U2838) );
  OAI22_X1 U17484 ( .A1(n14534), .A2(n14298), .B1(n20003), .B2(n14240), .ZN(
        P1_U2841) );
  AOI22_X1 U17485 ( .A1(n14575), .A2(n12418), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n14288), .ZN(n14241) );
  OAI21_X1 U17486 ( .B1(n14396), .B2(n14297), .A(n14241), .ZN(P1_U2844) );
  AOI22_X1 U17487 ( .A1(n14583), .A2(n12418), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n14288), .ZN(n14242) );
  OAI21_X1 U17488 ( .B1(n14312), .B2(n14290), .A(n14242), .ZN(P1_U2845) );
  OAI222_X1 U17489 ( .A1(n14297), .A2(n14414), .B1(n14243), .B2(n20003), .C1(
        n14588), .C2(n14298), .ZN(P1_U2846) );
  INV_X1 U17490 ( .A(n14426), .ZN(n14321) );
  OAI222_X1 U17491 ( .A1(n14297), .A2(n14321), .B1(n14244), .B2(n20003), .C1(
        n14598), .C2(n14298), .ZN(P1_U2847) );
  OAI222_X1 U17492 ( .A1(n14297), .A2(n14433), .B1(n14245), .B2(n20003), .C1(
        n14606), .C2(n14298), .ZN(P1_U2848) );
  AOI22_X1 U17493 ( .A1(n14621), .A2(n12418), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n14288), .ZN(n14246) );
  OAI21_X1 U17494 ( .B1(n14332), .B2(n14297), .A(n14246), .ZN(P1_U2849) );
  AOI22_X1 U17495 ( .A1(n14631), .A2(n12418), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n14288), .ZN(n14247) );
  OAI21_X1 U17496 ( .B1(n14452), .B2(n14290), .A(n14247), .ZN(P1_U2850) );
  AND2_X1 U17497 ( .A1(n14249), .A2(n14250), .ZN(n14251) );
  OR2_X1 U17498 ( .A1(n14251), .A2(n14182), .ZN(n15772) );
  INV_X1 U17499 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14255) );
  NAND2_X1 U17500 ( .A1(n14258), .A2(n14252), .ZN(n14253) );
  NAND2_X1 U17501 ( .A1(n14254), .A2(n14253), .ZN(n15771) );
  OAI222_X1 U17502 ( .A1(n14297), .A2(n15772), .B1(n14255), .B2(n20003), .C1(
        n15771), .C2(n14298), .ZN(P1_U2851) );
  OAI21_X1 U17503 ( .B1(n9657), .B2(n10016), .A(n14249), .ZN(n15779) );
  INV_X1 U17504 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14259) );
  OR2_X1 U17505 ( .A1(n14264), .A2(n14256), .ZN(n14257) );
  NAND2_X1 U17506 ( .A1(n14258), .A2(n14257), .ZN(n15778) );
  OAI222_X1 U17507 ( .A1(n15779), .A2(n14290), .B1(n20003), .B2(n14259), .C1(
        n15778), .C2(n14298), .ZN(P1_U2852) );
  AOI21_X1 U17508 ( .B1(n14261), .B2(n14266), .A(n9657), .ZN(n15859) );
  INV_X1 U17509 ( .A(n15859), .ZN(n14345) );
  INV_X1 U17510 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14265) );
  NOR2_X1 U17511 ( .A1(n14269), .A2(n14262), .ZN(n14263) );
  OR2_X1 U17512 ( .A1(n14264), .A2(n14263), .ZN(n15792) );
  OAI222_X1 U17513 ( .A1(n14297), .A2(n14345), .B1(n14265), .B2(n20003), .C1(
        n15792), .C2(n14298), .ZN(P1_U2853) );
  OAI21_X1 U17514 ( .B1(n14192), .B2(n14267), .A(n14266), .ZN(n15801) );
  INV_X1 U17515 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14273) );
  INV_X1 U17516 ( .A(n14268), .ZN(n14272) );
  INV_X1 U17517 ( .A(n14269), .ZN(n14270) );
  OAI21_X1 U17518 ( .B1(n14272), .B2(n14271), .A(n14270), .ZN(n15805) );
  OAI222_X1 U17519 ( .A1(n15801), .A2(n14290), .B1(n20003), .B2(n14273), .C1(
        n15805), .C2(n14298), .ZN(P1_U2854) );
  OAI222_X1 U17520 ( .A1(n15925), .A2(n14298), .B1(n20003), .B2(n20838), .C1(
        n15871), .C2(n14297), .ZN(P1_U2855) );
  AOI21_X1 U17521 ( .B1(n14275), .B2(n14274), .A(n9656), .ZN(n14486) );
  INV_X1 U17522 ( .A(n14486), .ZN(n15811) );
  OR2_X1 U17523 ( .A1(n14284), .A2(n14276), .ZN(n14277) );
  NAND2_X1 U17524 ( .A1(n14195), .A2(n14277), .ZN(n15809) );
  INV_X1 U17525 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14278) );
  OAI22_X1 U17526 ( .A1(n15809), .A2(n14298), .B1(n14278), .B2(n20003), .ZN(
        n14279) );
  INV_X1 U17527 ( .A(n14279), .ZN(n14280) );
  OAI21_X1 U17528 ( .B1(n15811), .B2(n14290), .A(n14280), .ZN(P1_U2856) );
  NOR2_X1 U17529 ( .A1(n14282), .A2(n14281), .ZN(n14283) );
  OR2_X1 U17530 ( .A1(n14284), .A2(n14283), .ZN(n15821) );
  INV_X1 U17531 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14287) );
  INV_X1 U17532 ( .A(n14274), .ZN(n14285) );
  AOI21_X1 U17533 ( .B1(n14286), .B2(n13771), .A(n14285), .ZN(n15881) );
  INV_X1 U17534 ( .A(n15881), .ZN(n14360) );
  OAI222_X1 U17535 ( .A1(n15821), .A2(n14298), .B1(n14287), .B2(n20003), .C1(
        n14360), .C2(n14297), .ZN(P1_U2857) );
  AOI22_X1 U17536 ( .A1(n15941), .A2(n12418), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14288), .ZN(n14289) );
  OAI21_X1 U17537 ( .B1(n14362), .B2(n14290), .A(n14289), .ZN(P1_U2859) );
  OR2_X1 U17538 ( .A1(n14292), .A2(n14291), .ZN(n14293) );
  NAND2_X1 U17539 ( .A1(n14294), .A2(n14293), .ZN(n15960) );
  INV_X1 U17540 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15835) );
  XOR2_X1 U17541 ( .A(n14296), .B(n14295), .Z(n15897) );
  INV_X1 U17542 ( .A(n15897), .ZN(n14371) );
  OAI222_X1 U17543 ( .A1(n15960), .A2(n14298), .B1(n15835), .B2(n20003), .C1(
        n14371), .C2(n14297), .ZN(P1_U2861) );
  INV_X1 U17544 ( .A(DATAI_13_), .ZN(n14300) );
  MUX2_X1 U17545 ( .A(n14300), .B(n14299), .S(n20091), .Z(n20012) );
  INV_X1 U17546 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14301) );
  OAI22_X1 U17547 ( .A1(n14352), .A2(n20012), .B1(n14365), .B2(n14301), .ZN(
        n14302) );
  AOI21_X1 U17548 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n14354), .A(n14302), .ZN(
        n14304) );
  NAND2_X1 U17549 ( .A1(n14355), .A2(DATAI_29_), .ZN(n14303) );
  OAI211_X1 U17550 ( .C1(n14305), .C2(n14370), .A(n14304), .B(n14303), .ZN(
        P1_U2875) );
  OAI22_X1 U17551 ( .A1(n14352), .A2(n14363), .B1(n14365), .B2(n13260), .ZN(
        n14306) );
  AOI21_X1 U17552 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14354), .A(n14306), .ZN(
        n14308) );
  NAND2_X1 U17553 ( .A1(n14355), .A2(DATAI_28_), .ZN(n14307) );
  OAI211_X1 U17554 ( .C1(n14396), .C2(n14370), .A(n14308), .B(n14307), .ZN(
        P1_U2876) );
  INV_X1 U17555 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16306) );
  AOI22_X1 U17556 ( .A1(n14323), .A2(n14367), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n14366), .ZN(n14309) );
  OAI21_X1 U17557 ( .B1(n16306), .B2(n14326), .A(n14309), .ZN(n14310) );
  AOI21_X1 U17558 ( .B1(n14355), .B2(DATAI_27_), .A(n14310), .ZN(n14311) );
  OAI21_X1 U17559 ( .B1(n14312), .B2(n14370), .A(n14311), .ZN(P1_U2877) );
  OAI22_X1 U17560 ( .A1(n14352), .A2(n14313), .B1(n14365), .B2(n13263), .ZN(
        n14314) );
  AOI21_X1 U17561 ( .B1(n14354), .B2(BUF1_REG_26__SCAN_IN), .A(n14314), .ZN(
        n14316) );
  NAND2_X1 U17562 ( .A1(n14355), .A2(DATAI_26_), .ZN(n14315) );
  OAI211_X1 U17563 ( .C1(n14414), .C2(n14370), .A(n14316), .B(n14315), .ZN(
        P1_U2878) );
  INV_X1 U17564 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n19118) );
  AOI22_X1 U17565 ( .A1(n14323), .A2(n14317), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n14366), .ZN(n14318) );
  OAI21_X1 U17566 ( .B1(n14326), .B2(n19118), .A(n14318), .ZN(n14319) );
  AOI21_X1 U17567 ( .B1(n14355), .B2(DATAI_25_), .A(n14319), .ZN(n14320) );
  OAI21_X1 U17568 ( .B1(n14321), .B2(n14370), .A(n14320), .ZN(P1_U2879) );
  INV_X1 U17569 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n14325) );
  AOI22_X1 U17570 ( .A1(n14323), .A2(n14322), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n14366), .ZN(n14324) );
  OAI21_X1 U17571 ( .B1(n14326), .B2(n14325), .A(n14324), .ZN(n14327) );
  AOI21_X1 U17572 ( .B1(n14355), .B2(DATAI_24_), .A(n14327), .ZN(n14328) );
  OAI21_X1 U17573 ( .B1(n14433), .B2(n14370), .A(n14328), .ZN(P1_U2880) );
  OAI22_X1 U17574 ( .A1(n14352), .A2(n20145), .B1(n14365), .B2(n13229), .ZN(
        n14329) );
  AOI21_X1 U17575 ( .B1(n14354), .B2(BUF1_REG_23__SCAN_IN), .A(n14329), .ZN(
        n14331) );
  NAND2_X1 U17576 ( .A1(n14355), .A2(DATAI_23_), .ZN(n14330) );
  OAI211_X1 U17577 ( .C1(n14332), .C2(n14370), .A(n14331), .B(n14330), .ZN(
        P1_U2881) );
  OAI22_X1 U17578 ( .A1(n14352), .A2(n20138), .B1(n14365), .B2(n13196), .ZN(
        n14333) );
  AOI21_X1 U17579 ( .B1(n14354), .B2(BUF1_REG_22__SCAN_IN), .A(n14333), .ZN(
        n14335) );
  NAND2_X1 U17580 ( .A1(n14355), .A2(DATAI_22_), .ZN(n14334) );
  OAI211_X1 U17581 ( .C1(n14452), .C2(n14370), .A(n14335), .B(n14334), .ZN(
        P1_U2882) );
  OAI22_X1 U17582 ( .A1(n14352), .A2(n20134), .B1(n14365), .B2(n13189), .ZN(
        n14336) );
  AOI21_X1 U17583 ( .B1(n14354), .B2(BUF1_REG_21__SCAN_IN), .A(n14336), .ZN(
        n14338) );
  NAND2_X1 U17584 ( .A1(n14355), .A2(DATAI_21_), .ZN(n14337) );
  OAI211_X1 U17585 ( .C1(n15772), .C2(n14370), .A(n14338), .B(n14337), .ZN(
        P1_U2883) );
  OAI22_X1 U17586 ( .A1(n14352), .A2(n20129), .B1(n14365), .B2(n13201), .ZN(
        n14339) );
  AOI21_X1 U17587 ( .B1(n14354), .B2(BUF1_REG_20__SCAN_IN), .A(n14339), .ZN(
        n14341) );
  NAND2_X1 U17588 ( .A1(n14355), .A2(DATAI_20_), .ZN(n14340) );
  OAI211_X1 U17589 ( .C1(n15779), .C2(n14370), .A(n14341), .B(n14340), .ZN(
        P1_U2884) );
  OAI22_X1 U17590 ( .A1(n14352), .A2(n20124), .B1(n14365), .B2(n13204), .ZN(
        n14342) );
  AOI21_X1 U17591 ( .B1(n14354), .B2(BUF1_REG_19__SCAN_IN), .A(n14342), .ZN(
        n14344) );
  NAND2_X1 U17592 ( .A1(n14355), .A2(DATAI_19_), .ZN(n14343) );
  OAI211_X1 U17593 ( .C1(n14345), .C2(n14370), .A(n14344), .B(n14343), .ZN(
        P1_U2885) );
  OAI22_X1 U17594 ( .A1(n14352), .A2(n20119), .B1(n14365), .B2(n13207), .ZN(
        n14346) );
  AOI21_X1 U17595 ( .B1(n14354), .B2(BUF1_REG_18__SCAN_IN), .A(n14346), .ZN(
        n14348) );
  NAND2_X1 U17596 ( .A1(n14355), .A2(DATAI_18_), .ZN(n14347) );
  OAI211_X1 U17597 ( .C1(n15801), .C2(n14370), .A(n14348), .B(n14347), .ZN(
        P1_U2886) );
  OAI22_X1 U17598 ( .A1(n14352), .A2(n20114), .B1(n14365), .B2(n13210), .ZN(
        n14349) );
  AOI21_X1 U17599 ( .B1(n14354), .B2(BUF1_REG_17__SCAN_IN), .A(n14349), .ZN(
        n14351) );
  NAND2_X1 U17600 ( .A1(n14355), .A2(DATAI_17_), .ZN(n14350) );
  OAI211_X1 U17601 ( .C1(n15871), .C2(n14370), .A(n14351), .B(n14350), .ZN(
        P1_U2887) );
  OAI22_X1 U17602 ( .A1(n14352), .A2(n20105), .B1(n14365), .B2(n13234), .ZN(
        n14353) );
  AOI21_X1 U17603 ( .B1(n14354), .B2(BUF1_REG_16__SCAN_IN), .A(n14353), .ZN(
        n14357) );
  NAND2_X1 U17604 ( .A1(n14355), .A2(DATAI_16_), .ZN(n14356) );
  OAI211_X1 U17605 ( .C1(n15811), .C2(n14370), .A(n14357), .B(n14356), .ZN(
        P1_U2888) );
  OAI222_X1 U17606 ( .A1(n14370), .A2(n14360), .B1(n14365), .B2(n14359), .C1(
        n14364), .C2(n14358), .ZN(P1_U2889) );
  INV_X1 U17607 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14361) );
  OAI222_X1 U17608 ( .A1(n14370), .A2(n14362), .B1(n14364), .B2(n20012), .C1(
        n14361), .C2(n14365), .ZN(P1_U2891) );
  OAI222_X1 U17609 ( .A1(n15825), .A2(n14370), .B1(n13282), .B2(n14365), .C1(
        n14364), .C2(n14363), .ZN(P1_U2892) );
  AOI22_X1 U17610 ( .A1(n14368), .A2(n14367), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14366), .ZN(n14369) );
  OAI21_X1 U17611 ( .B1(n14371), .B2(n14370), .A(n14369), .ZN(P1_U2893) );
  XNOR2_X1 U17612 ( .A(n14375), .B(n14374), .ZN(n14549) );
  INV_X1 U17613 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20747) );
  NOR2_X1 U17614 ( .A1(n20065), .A2(n20747), .ZN(n14545) );
  AOI21_X1 U17615 ( .B1(n20025), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14545), .ZN(n14376) );
  OAI21_X1 U17616 ( .B1(n20036), .B2(n14377), .A(n14376), .ZN(n14378) );
  OAI21_X1 U17617 ( .B1(n14549), .B2(n19908), .A(n14380), .ZN(P1_U2968) );
  NOR2_X1 U17618 ( .A1(n20065), .A2(n20743), .ZN(n14560) );
  AOI21_X1 U17619 ( .B1(n20025), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14560), .ZN(n14383) );
  OAI21_X1 U17620 ( .B1(n20036), .B2(n14384), .A(n14383), .ZN(n14385) );
  AOI21_X1 U17621 ( .B1(n14386), .B2(n20031), .A(n14385), .ZN(n14387) );
  OAI21_X1 U17622 ( .B1(n19908), .B2(n14568), .A(n14387), .ZN(P1_U2970) );
  NAND2_X1 U17624 ( .A1(n9582), .A2(n14591), .ZN(n14410) );
  NAND2_X1 U17625 ( .A1(n14389), .A2(n14410), .ZN(n14393) );
  OAI21_X1 U17626 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14390), .A(
        n14393), .ZN(n14392) );
  INV_X1 U17627 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14403) );
  MUX2_X1 U17628 ( .A(n14403), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n9581), .Z(n14391) );
  OAI211_X1 U17629 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14393), .A(
        n14392), .B(n14391), .ZN(n14394) );
  XOR2_X1 U17630 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14394), .Z(
        n14579) );
  NAND2_X1 U17631 ( .A1(n20024), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14569) );
  OAI21_X1 U17632 ( .B1(n14484), .B2(n14395), .A(n14569), .ZN(n14398) );
  NOR2_X1 U17633 ( .A1(n14396), .A2(n20090), .ZN(n14397) );
  OAI21_X1 U17634 ( .B1(n19908), .B2(n14579), .A(n14400), .ZN(P1_U2971) );
  MUX2_X1 U17635 ( .A(n14402), .B(n14401), .S(n15892), .Z(n14404) );
  XNOR2_X1 U17636 ( .A(n14404), .B(n14403), .ZN(n14587) );
  NOR2_X1 U17637 ( .A1(n20065), .A2(n20738), .ZN(n14582) );
  AOI21_X1 U17638 ( .B1(n20025), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14582), .ZN(n14405) );
  OAI21_X1 U17639 ( .B1(n20036), .B2(n14406), .A(n14405), .ZN(n14407) );
  AOI21_X1 U17640 ( .B1(n14408), .B2(n20031), .A(n14407), .ZN(n14409) );
  OAI21_X1 U17641 ( .B1(n19908), .B2(n14587), .A(n14409), .ZN(P1_U2972) );
  OAI211_X1 U17642 ( .C1(n15892), .C2(n14389), .A(n14411), .B(n14410), .ZN(
        n14412) );
  XNOR2_X1 U17643 ( .A(n14412), .B(n14542), .ZN(n14597) );
  NAND2_X1 U17644 ( .A1(n20024), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14589) );
  OAI21_X1 U17645 ( .B1(n14484), .B2(n14413), .A(n14589), .ZN(n14416) );
  NOR2_X1 U17646 ( .A1(n14414), .A2(n20090), .ZN(n14415) );
  OAI21_X1 U17647 ( .B1(n19908), .B2(n14597), .A(n14418), .ZN(P1_U2973) );
  NAND2_X1 U17648 ( .A1(n14419), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14429) );
  NOR2_X1 U17649 ( .A1(n14429), .A2(n14610), .ZN(n14421) );
  NOR3_X1 U17650 ( .A1(n14389), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14420) );
  MUX2_X1 U17651 ( .A(n14421), .B(n14420), .S(n15892), .Z(n14422) );
  XNOR2_X1 U17652 ( .A(n14422), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14605) );
  INV_X1 U17653 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20732) );
  NOR2_X1 U17654 ( .A1(n20065), .A2(n20732), .ZN(n14600) );
  AOI21_X1 U17655 ( .B1(n20025), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14600), .ZN(n14423) );
  OAI21_X1 U17656 ( .B1(n20036), .B2(n14424), .A(n14423), .ZN(n14425) );
  AOI21_X1 U17657 ( .B1(n14426), .B2(n20031), .A(n14425), .ZN(n14427) );
  OAI21_X1 U17658 ( .B1(n19908), .B2(n14605), .A(n14427), .ZN(P1_U2974) );
  INV_X1 U17659 ( .A(n14389), .ZN(n14428) );
  NAND2_X1 U17660 ( .A1(n14429), .A2(n14428), .ZN(n14430) );
  MUX2_X1 U17661 ( .A(n14430), .B(n14429), .S(n9582), .Z(n14431) );
  XNOR2_X1 U17662 ( .A(n14431), .B(n14610), .ZN(n14617) );
  NAND2_X1 U17663 ( .A1(n20024), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14607) );
  OAI21_X1 U17664 ( .B1(n14484), .B2(n14432), .A(n14607), .ZN(n14435) );
  NOR2_X1 U17665 ( .A1(n14433), .A2(n20090), .ZN(n14434) );
  AOI211_X1 U17666 ( .C1(n15889), .C2(n14436), .A(n14435), .B(n14434), .ZN(
        n14437) );
  OAI21_X1 U17667 ( .B1(n19908), .B2(n14617), .A(n14437), .ZN(P1_U2975) );
  XNOR2_X1 U17668 ( .A(n9582), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14438) );
  XNOR2_X1 U17669 ( .A(n14389), .B(n14438), .ZN(n14625) );
  NOR2_X1 U17670 ( .A1(n20065), .A2(n20731), .ZN(n14620) );
  AOI21_X1 U17671 ( .B1(n20025), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n14620), .ZN(n14439) );
  OAI21_X1 U17672 ( .B1(n20036), .B2(n14440), .A(n14439), .ZN(n14441) );
  AOI21_X1 U17673 ( .B1(n14442), .B2(n20031), .A(n14441), .ZN(n14443) );
  OAI21_X1 U17674 ( .B1(n14625), .B2(n19908), .A(n14443), .ZN(P1_U2976) );
  NOR2_X1 U17675 ( .A1(n20065), .A2(n20729), .ZN(n14627) );
  INV_X1 U17676 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14444) );
  NOR2_X1 U17677 ( .A1(n14484), .A2(n14444), .ZN(n14445) );
  AOI211_X1 U17678 ( .C1(n15889), .C2(n14446), .A(n14627), .B(n14445), .ZN(
        n14451) );
  NAND2_X1 U17679 ( .A1(n14448), .A2(n14447), .ZN(n14449) );
  XNOR2_X1 U17680 ( .A(n14449), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14626) );
  NAND2_X1 U17681 ( .A1(n14626), .A2(n20032), .ZN(n14450) );
  OAI211_X1 U17682 ( .C1(n14452), .C2(n20090), .A(n14451), .B(n14450), .ZN(
        P1_U2977) );
  NOR3_X1 U17683 ( .A1(n14453), .A2(n15892), .A3(n15857), .ZN(n14464) );
  OR2_X1 U17684 ( .A1(n14454), .A2(n9582), .ZN(n14459) );
  NOR2_X1 U17685 ( .A1(n14459), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14462) );
  AOI21_X1 U17686 ( .B1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n14464), .A(
        n14462), .ZN(n14455) );
  XNOR2_X1 U17687 ( .A(n14455), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14635) );
  NAND2_X1 U17688 ( .A1(n14635), .A2(n20032), .ZN(n14458) );
  AND2_X1 U17689 ( .A1(n20024), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14638) );
  NOR2_X1 U17690 ( .A1(n20036), .A2(n15776), .ZN(n14456) );
  AOI211_X1 U17691 ( .C1(n20025), .C2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n14638), .B(n14456), .ZN(n14457) );
  OAI211_X1 U17692 ( .C1(n15772), .C2(n20090), .A(n14458), .B(n14457), .ZN(
        P1_U2978) );
  INV_X1 U17693 ( .A(n14459), .ZN(n14460) );
  NOR3_X1 U17694 ( .A1(n14464), .A2(n14463), .A3(n14460), .ZN(n14461) );
  AOI211_X1 U17695 ( .C1(n14464), .C2(n14463), .A(n14462), .B(n14461), .ZN(
        n14651) );
  NAND2_X1 U17696 ( .A1(n20024), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14648) );
  OAI21_X1 U17697 ( .B1(n14484), .B2(n14465), .A(n14648), .ZN(n14467) );
  NOR2_X1 U17698 ( .A1(n15779), .A2(n20090), .ZN(n14466) );
  AOI211_X1 U17699 ( .C1(n15889), .C2(n15781), .A(n14467), .B(n14466), .ZN(
        n14468) );
  OAI21_X1 U17700 ( .B1(n14651), .B2(n19908), .A(n14468), .ZN(P1_U2979) );
  NAND2_X1 U17701 ( .A1(n20024), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14654) );
  OAI21_X1 U17702 ( .B1(n14484), .B2(n15796), .A(n14654), .ZN(n14469) );
  AOI21_X1 U17703 ( .B1(n15803), .B2(n15889), .A(n14469), .ZN(n14473) );
  OR2_X1 U17704 ( .A1(n14471), .A2(n14470), .ZN(n14652) );
  NAND3_X1 U17705 ( .A1(n14652), .A2(n14453), .A3(n20032), .ZN(n14472) );
  OAI211_X1 U17706 ( .C1(n15801), .C2(n20090), .A(n14473), .B(n14472), .ZN(
        P1_U2981) );
  INV_X1 U17707 ( .A(n14475), .ZN(n14477) );
  AOI21_X1 U17708 ( .B1(n11144), .B2(n14477), .A(n14476), .ZN(n15878) );
  INV_X1 U17709 ( .A(n14480), .ZN(n14478) );
  NOR2_X1 U17710 ( .A1(n14479), .A2(n14478), .ZN(n15877) );
  NAND2_X1 U17711 ( .A1(n15878), .A2(n15877), .ZN(n15876) );
  NAND2_X1 U17712 ( .A1(n15876), .A2(n14480), .ZN(n14481) );
  XOR2_X1 U17713 ( .A(n14482), .B(n14481), .Z(n14668) );
  NAND2_X1 U17714 ( .A1(n15889), .A2(n15814), .ZN(n14483) );
  NAND2_X1 U17715 ( .A1(n20024), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n14664) );
  OAI211_X1 U17716 ( .C1(n14484), .C2(n15808), .A(n14483), .B(n14664), .ZN(
        n14485) );
  AOI21_X1 U17717 ( .B1(n14486), .B2(n20031), .A(n14485), .ZN(n14487) );
  OAI21_X1 U17718 ( .B1(n14668), .B2(n19908), .A(n14487), .ZN(P1_U2983) );
  NAND2_X1 U17719 ( .A1(n15893), .A2(n14488), .ZN(n15867) );
  AND2_X1 U17720 ( .A1(n9582), .A2(n14489), .ZN(n14503) );
  INV_X1 U17721 ( .A(n14503), .ZN(n14490) );
  NAND3_X1 U17722 ( .A1(n15867), .A2(n14491), .A3(n14490), .ZN(n14493) );
  NAND2_X1 U17723 ( .A1(n14493), .A2(n14492), .ZN(n14495) );
  XNOR2_X1 U17724 ( .A(n9581), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14494) );
  XNOR2_X1 U17725 ( .A(n14495), .B(n14494), .ZN(n14678) );
  INV_X1 U17726 ( .A(n14496), .ZN(n14500) );
  NAND2_X1 U17727 ( .A1(n20024), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n14672) );
  NAND2_X1 U17728 ( .A1(n20025), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14497) );
  OAI211_X1 U17729 ( .C1(n20036), .C2(n14498), .A(n14672), .B(n14497), .ZN(
        n14499) );
  AOI21_X1 U17730 ( .B1(n14500), .B2(n20031), .A(n14499), .ZN(n14501) );
  OAI21_X1 U17731 ( .B1(n14678), .B2(n19908), .A(n14501), .ZN(P1_U2985) );
  OAI22_X1 U17732 ( .A1(n15893), .A2(n14503), .B1(n14502), .B2(n9582), .ZN(
        n15886) );
  INV_X1 U17733 ( .A(n14505), .ZN(n14504) );
  OAI21_X1 U17734 ( .B1(n9581), .B2(n15956), .A(n14504), .ZN(n15885) );
  NOR2_X1 U17735 ( .A1(n15886), .A2(n15885), .ZN(n15884) );
  NOR2_X1 U17736 ( .A1(n15884), .A2(n14505), .ZN(n14506) );
  XOR2_X1 U17737 ( .A(n14507), .B(n14506), .Z(n15940) );
  INV_X1 U17738 ( .A(n14508), .ZN(n14510) );
  AOI22_X1 U17739 ( .A1(n20025), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n20024), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14509) );
  OAI21_X1 U17740 ( .B1(n20036), .B2(n14510), .A(n14509), .ZN(n14511) );
  AOI21_X1 U17741 ( .B1(n14512), .B2(n20031), .A(n14511), .ZN(n14513) );
  OAI21_X1 U17742 ( .B1(n15940), .B2(n19908), .A(n14513), .ZN(P1_U2986) );
  AND2_X1 U17743 ( .A1(n14514), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14516) );
  XNOR2_X1 U17744 ( .A(n15893), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14515) );
  MUX2_X1 U17745 ( .A(n14516), .B(n14515), .S(n9581), .Z(n14517) );
  NOR3_X1 U17746 ( .A1(n14514), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n9581), .ZN(n15894) );
  NOR2_X1 U17747 ( .A1(n14517), .A2(n15894), .ZN(n14689) );
  INV_X1 U17748 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14518) );
  NOR2_X1 U17749 ( .A1(n20065), .A2(n14518), .ZN(n14686) );
  AOI21_X1 U17750 ( .B1(n20025), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n14686), .ZN(n14519) );
  OAI21_X1 U17751 ( .B1(n20036), .B2(n15848), .A(n14519), .ZN(n14520) );
  AOI21_X1 U17752 ( .B1(n15850), .B2(n20031), .A(n14520), .ZN(n14521) );
  OAI21_X1 U17753 ( .B1(n14689), .B2(n19908), .A(n14521), .ZN(P1_U2989) );
  INV_X1 U17754 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14561) );
  NAND2_X1 U17755 ( .A1(n20057), .A2(n14681), .ZN(n20075) );
  INV_X1 U17756 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14554) );
  INV_X1 U17757 ( .A(n20075), .ZN(n14662) );
  NAND2_X1 U17758 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14532) );
  AND3_X1 U17759 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14679) );
  NAND3_X1 U17760 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n14679), .ZN(n14523) );
  NAND2_X1 U17761 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14522), .ZN(
        n14535) );
  OR2_X1 U17762 ( .A1(n14523), .A2(n14535), .ZN(n15949) );
  NAND3_X1 U17763 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14669) );
  AOI221_X1 U17764 ( .B1(n15949), .B2(n20061), .C1(n14669), .C2(n20061), .A(
        n20059), .ZN(n14527) );
  INV_X1 U17765 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15966) );
  NOR2_X1 U17766 ( .A1(n15966), .A2(n14523), .ZN(n15947) );
  NAND2_X1 U17767 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15947), .ZN(
        n14536) );
  NOR2_X1 U17768 ( .A1(n14537), .A2(n14536), .ZN(n14524) );
  AND2_X1 U17769 ( .A1(n14524), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14525) );
  OR2_X1 U17770 ( .A1(n20057), .A2(n14525), .ZN(n14526) );
  NAND4_X1 U17771 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14653) );
  NOR2_X1 U17772 ( .A1(n14660), .A2(n14653), .ZN(n14644) );
  AND2_X1 U17773 ( .A1(n14644), .A2(n11153), .ZN(n14528) );
  NAND2_X1 U17774 ( .A1(n14674), .A2(n14528), .ZN(n14529) );
  NAND2_X1 U17775 ( .A1(n14529), .A2(n15982), .ZN(n14643) );
  NAND2_X1 U17776 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14541) );
  NAND2_X1 U17777 ( .A1(n20075), .A2(n14541), .ZN(n14530) );
  NAND2_X1 U17778 ( .A1(n14643), .A2(n14530), .ZN(n14622) );
  AOI21_X1 U17779 ( .B1(n15982), .B2(n14532), .A(n14602), .ZN(n14576) );
  OAI21_X1 U17780 ( .B1(n14571), .B2(n14662), .A(n14576), .ZN(n14566) );
  INV_X1 U17781 ( .A(n15982), .ZN(n14533) );
  NOR3_X1 U17782 ( .A1(n14552), .A2(n14533), .A3(n14374), .ZN(n14547) );
  NOR2_X1 U17783 ( .A1(n14534), .A2(n20079), .ZN(n14546) );
  INV_X1 U17784 ( .A(n14535), .ZN(n14680) );
  NAND2_X1 U17785 ( .A1(n20056), .A2(n14680), .ZN(n14538) );
  AOI211_X1 U17786 ( .C1(n20057), .C2(n14538), .A(n14537), .B(n14536), .ZN(
        n14539) );
  INV_X1 U17787 ( .A(n14539), .ZN(n15945) );
  NAND2_X1 U17788 ( .A1(n14644), .A2(n14661), .ZN(n15922) );
  NOR2_X1 U17789 ( .A1(n14636), .A2(n14541), .ZN(n14590) );
  NOR2_X1 U17790 ( .A1(n14591), .A2(n14542), .ZN(n14543) );
  AND2_X1 U17791 ( .A1(n14590), .A2(n14543), .ZN(n14570) );
  NAND3_X1 U17792 ( .A1(n14570), .A2(n14571), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14553) );
  NOR3_X1 U17793 ( .A1(n14553), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14554), .ZN(n14544) );
  OAI21_X1 U17794 ( .B1(n14549), .B2(n20073), .A(n14548), .ZN(P1_U3000) );
  INV_X1 U17795 ( .A(n14550), .ZN(n14557) );
  INV_X1 U17796 ( .A(n14551), .ZN(n14556) );
  AOI21_X1 U17797 ( .B1(n14554), .B2(n14553), .A(n14552), .ZN(n14555) );
  AOI211_X1 U17798 ( .C1(n20048), .C2(n14557), .A(n14556), .B(n14555), .ZN(
        n14558) );
  OAI21_X1 U17799 ( .B1(n14559), .B2(n20073), .A(n14558), .ZN(P1_U3001) );
  INV_X1 U17800 ( .A(n14560), .ZN(n14563) );
  NAND3_X1 U17801 ( .A1(n14570), .A2(n14571), .A3(n14561), .ZN(n14562) );
  OAI211_X1 U17802 ( .C1(n14564), .C2(n20079), .A(n14563), .B(n14562), .ZN(
        n14565) );
  AOI21_X1 U17803 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n14566), .A(
        n14565), .ZN(n14567) );
  OAI21_X1 U17804 ( .B1(n14568), .B2(n20073), .A(n14567), .ZN(P1_U3002) );
  INV_X1 U17805 ( .A(n14569), .ZN(n14574) );
  INV_X1 U17806 ( .A(n14570), .ZN(n14580) );
  NOR3_X1 U17807 ( .A1(n14580), .A2(n14572), .A3(n14571), .ZN(n14573) );
  AOI211_X1 U17808 ( .C1(n14575), .C2(n20048), .A(n14574), .B(n14573), .ZN(
        n14578) );
  INV_X1 U17809 ( .A(n14576), .ZN(n14584) );
  NAND2_X1 U17810 ( .A1(n14584), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14577) );
  OAI211_X1 U17811 ( .C1(n14579), .C2(n20073), .A(n14578), .B(n14577), .ZN(
        P1_U3003) );
  NOR2_X1 U17812 ( .A1(n14580), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14581) );
  AOI211_X1 U17813 ( .C1(n14583), .C2(n20048), .A(n14582), .B(n14581), .ZN(
        n14586) );
  NAND2_X1 U17814 ( .A1(n14584), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14585) );
  OAI211_X1 U17815 ( .C1(n14587), .C2(n20073), .A(n14586), .B(n14585), .ZN(
        P1_U3004) );
  INV_X1 U17816 ( .A(n14588), .ZN(n14594) );
  INV_X1 U17817 ( .A(n14589), .ZN(n14593) );
  INV_X1 U17818 ( .A(n14590), .ZN(n14618) );
  NOR3_X1 U17819 ( .A1(n14618), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14591), .ZN(n14592) );
  AOI211_X1 U17820 ( .C1(n14594), .C2(n20048), .A(n14593), .B(n14592), .ZN(
        n14596) );
  NOR4_X1 U17821 ( .A1(n14618), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n14611), .A4(n14610), .ZN(n14599) );
  OAI21_X1 U17822 ( .B1(n14602), .B2(n14599), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14595) );
  OAI211_X1 U17823 ( .C1(n14597), .C2(n20073), .A(n14596), .B(n14595), .ZN(
        P1_U3005) );
  INV_X1 U17824 ( .A(n14598), .ZN(n14601) );
  AOI211_X1 U17825 ( .C1(n14601), .C2(n20048), .A(n14600), .B(n14599), .ZN(
        n14604) );
  NAND2_X1 U17826 ( .A1(n14602), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14603) );
  OAI211_X1 U17827 ( .C1(n14605), .C2(n20073), .A(n14604), .B(n14603), .ZN(
        P1_U3006) );
  INV_X1 U17828 ( .A(n14606), .ZN(n14609) );
  INV_X1 U17829 ( .A(n14607), .ZN(n14608) );
  AOI21_X1 U17830 ( .B1(n14609), .B2(n20048), .A(n14608), .ZN(n14616) );
  AOI21_X1 U17831 ( .B1(n15950), .B2(n20057), .A(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14613) );
  OAI21_X1 U17832 ( .B1(n14618), .B2(n14611), .A(n14610), .ZN(n14612) );
  OAI21_X1 U17833 ( .B1(n14614), .B2(n14613), .A(n14612), .ZN(n14615) );
  OAI211_X1 U17834 ( .C1(n14617), .C2(n20073), .A(n14616), .B(n14615), .ZN(
        P1_U3007) );
  NOR2_X1 U17835 ( .A1(n14618), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14619) );
  AOI211_X1 U17836 ( .C1(n14621), .C2(n20048), .A(n14620), .B(n14619), .ZN(
        n14624) );
  NAND2_X1 U17837 ( .A1(n14622), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14623) );
  OAI211_X1 U17838 ( .C1(n14625), .C2(n20073), .A(n14624), .B(n14623), .ZN(
        P1_U3008) );
  INV_X1 U17839 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14634) );
  NAND2_X1 U17840 ( .A1(n14626), .A2(n20062), .ZN(n14633) );
  XNOR2_X1 U17841 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14629) );
  INV_X1 U17842 ( .A(n14627), .ZN(n14628) );
  OAI21_X1 U17843 ( .B1(n14636), .B2(n14629), .A(n14628), .ZN(n14630) );
  AOI21_X1 U17844 ( .B1(n14631), .B2(n20048), .A(n14630), .ZN(n14632) );
  OAI211_X1 U17845 ( .C1(n14643), .C2(n14634), .A(n14633), .B(n14632), .ZN(
        P1_U3009) );
  NAND2_X1 U17846 ( .A1(n14635), .A2(n20062), .ZN(n14641) );
  INV_X1 U17847 ( .A(n15771), .ZN(n14639) );
  NOR2_X1 U17848 ( .A1(n14636), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14637) );
  AOI211_X1 U17849 ( .C1(n14639), .C2(n20048), .A(n14638), .B(n14637), .ZN(
        n14640) );
  OAI211_X1 U17850 ( .C1(n14643), .C2(n14642), .A(n14641), .B(n14640), .ZN(
        P1_U3010) );
  OAI21_X1 U17851 ( .B1(n14662), .B2(n14644), .A(n14674), .ZN(n15917) );
  INV_X1 U17852 ( .A(n15922), .ZN(n14646) );
  OAI211_X1 U17853 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n14646), .B(n14645), .ZN(
        n14647) );
  OAI211_X1 U17854 ( .C1(n15778), .C2(n20079), .A(n14648), .B(n14647), .ZN(
        n14649) );
  AOI21_X1 U17855 ( .B1(n15917), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14649), .ZN(n14650) );
  OAI21_X1 U17856 ( .B1(n14651), .B2(n20073), .A(n14650), .ZN(P1_U3011) );
  INV_X1 U17857 ( .A(n14674), .ZN(n15939) );
  AOI21_X1 U17858 ( .B1(n14653), .B2(n20075), .A(n15939), .ZN(n15924) );
  NAND3_X1 U17859 ( .A1(n14652), .A2(n14453), .A3(n20062), .ZN(n14659) );
  NOR2_X1 U17860 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14653), .ZN(
        n14657) );
  INV_X1 U17861 ( .A(n14654), .ZN(n14656) );
  NOR2_X1 U17862 ( .A1(n15805), .A2(n20079), .ZN(n14655) );
  AOI211_X1 U17863 ( .C1(n14661), .C2(n14657), .A(n14656), .B(n14655), .ZN(
        n14658) );
  OAI211_X1 U17864 ( .C1(n15924), .C2(n14660), .A(n14659), .B(n14658), .ZN(
        P1_U3013) );
  NAND2_X1 U17865 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14661), .ZN(
        n15933) );
  AOI21_X1 U17866 ( .B1(n11145), .B2(n15863), .A(n15933), .ZN(n14666) );
  NAND2_X1 U17867 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15923) );
  OAI21_X1 U17868 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14662), .A(
        n14674), .ZN(n15932) );
  NAND2_X1 U17869 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15932), .ZN(
        n14663) );
  OAI211_X1 U17870 ( .C1(n15809), .C2(n20079), .A(n14664), .B(n14663), .ZN(
        n14665) );
  AOI21_X1 U17871 ( .B1(n14666), .B2(n15923), .A(n14665), .ZN(n14667) );
  OAI21_X1 U17872 ( .B1(n14668), .B2(n20073), .A(n14667), .ZN(P1_U3015) );
  NAND2_X1 U17873 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14683) );
  NAND2_X1 U17874 ( .A1(n14679), .A2(n15983), .ZN(n15968) );
  NOR2_X1 U17875 ( .A1(n14683), .A2(n15968), .ZN(n15962) );
  NOR2_X1 U17876 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14669), .ZN(
        n14676) );
  NAND2_X1 U17877 ( .A1(n14670), .A2(n20048), .ZN(n14671) );
  OAI211_X1 U17878 ( .C1(n14674), .C2(n14673), .A(n14672), .B(n14671), .ZN(
        n14675) );
  AOI21_X1 U17879 ( .B1(n15962), .B2(n14676), .A(n14675), .ZN(n14677) );
  OAI21_X1 U17880 ( .B1(n14678), .B2(n20073), .A(n14677), .ZN(P1_U3017) );
  INV_X1 U17881 ( .A(n15846), .ZN(n14687) );
  OAI211_X1 U17882 ( .C1(n14681), .C2(n14680), .A(n14679), .B(n15946), .ZN(
        n14682) );
  NAND2_X1 U17883 ( .A1(n15982), .A2(n14682), .ZN(n15979) );
  OAI21_X1 U17884 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n14683), .ZN(n14684) );
  OAI22_X1 U17885 ( .A1(n11269), .A2(n15979), .B1(n15968), .B2(n14684), .ZN(
        n14685) );
  AOI211_X1 U17886 ( .C1(n20048), .C2(n14687), .A(n14686), .B(n14685), .ZN(
        n14688) );
  OAI21_X1 U17887 ( .B1(n14689), .B2(n20073), .A(n14688), .ZN(P1_U3021) );
  INV_X1 U17888 ( .A(n13446), .ZN(n14691) );
  NAND2_X1 U17889 ( .A1(n14691), .A2(n14690), .ZN(n14695) );
  OAI22_X1 U17890 ( .A1(n15706), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n14695), .B2(n14692), .ZN(n14693) );
  AOI21_X1 U17891 ( .B1(n20564), .B2(n14694), .A(n14693), .ZN(n15707) );
  INV_X1 U17892 ( .A(n14695), .ZN(n14699) );
  INV_X1 U17893 ( .A(n14696), .ZN(n14697) );
  AOI22_X1 U17894 ( .A1(n15739), .A2(n14699), .B1(n14698), .B2(n14697), .ZN(
        n14700) );
  OAI21_X1 U17895 ( .B1(n15707), .B2(n14701), .A(n14700), .ZN(n14703) );
  MUX2_X1 U17896 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14703), .S(
        n14702), .Z(P1_U3473) );
  NOR2_X1 U17897 ( .A1(n14705), .A2(n14706), .ZN(n14707) );
  INV_X1 U17898 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14710) );
  INV_X1 U17899 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14708) );
  NAND2_X1 U17900 ( .A1(n14768), .A2(n14713), .ZN(n14712) );
  AND2_X1 U17901 ( .A1(n14712), .A2(n9888), .ZN(n14771) );
  OAI21_X1 U17902 ( .B1(n14734), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14713), .ZN(n15130) );
  INV_X1 U17903 ( .A(n15130), .ZN(n18761) );
  AOI21_X1 U17904 ( .B1(n14731), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14714) );
  OR2_X1 U17905 ( .A1(n14732), .A2(n14714), .ZN(n15157) );
  INV_X1 U17906 ( .A(n15157), .ZN(n18786) );
  AOI21_X1 U17907 ( .B1(n15169), .B2(n14729), .A(n14731), .ZN(n14783) );
  OAI21_X1 U17908 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n14726), .A(
        n14715), .ZN(n18808) );
  INV_X1 U17909 ( .A(n18808), .ZN(n14728) );
  OAI21_X1 U17910 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n9682), .A(
        n14727), .ZN(n16150) );
  INV_X1 U17911 ( .A(n16150), .ZN(n14811) );
  OAI21_X1 U17912 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n14722), .A(
        n14725), .ZN(n16165) );
  INV_X1 U17913 ( .A(n16165), .ZN(n14827) );
  AOI21_X1 U17914 ( .B1(n16189), .B2(n14720), .A(n14716), .ZN(n18862) );
  AOI21_X1 U17915 ( .B1(n15217), .B2(n14717), .A(n14721), .ZN(n18884) );
  AOI21_X1 U17916 ( .B1(n19099), .B2(n14719), .A(n14718), .ZN(n19088) );
  AOI22_X1 U17917 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18737), .ZN(n15540) );
  AOI22_X1 U17918 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18930), .B2(n18737), .ZN(
        n15539) );
  NAND2_X1 U17919 ( .A1(n15540), .A2(n15539), .ZN(n15538) );
  NOR2_X1 U17920 ( .A1(n14855), .A2(n15538), .ZN(n14838) );
  NAND2_X1 U17921 ( .A1(n14838), .A2(n14839), .ZN(n18914) );
  NOR2_X1 U17922 ( .A1(n19088), .A2(n18914), .ZN(n18895) );
  NAND2_X1 U17923 ( .A1(n18895), .A2(n18898), .ZN(n18882) );
  NOR2_X1 U17924 ( .A1(n18884), .A2(n18882), .ZN(n18867) );
  OAI21_X1 U17925 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n14721), .A(
        n14720), .ZN(n18869) );
  NAND2_X1 U17926 ( .A1(n18867), .A2(n18869), .ZN(n18860) );
  NOR2_X1 U17927 ( .A1(n18862), .A2(n18860), .ZN(n18847) );
  AOI21_X1 U17928 ( .B1(n16175), .B2(n14723), .A(n14722), .ZN(n18848) );
  INV_X1 U17929 ( .A(n18848), .ZN(n14724) );
  NAND2_X1 U17930 ( .A1(n18847), .A2(n14724), .ZN(n14825) );
  NOR2_X1 U17931 ( .A1(n14827), .A2(n14825), .ZN(n18842) );
  AOI21_X1 U17932 ( .B1(n18831), .B2(n14725), .A(n9682), .ZN(n18837) );
  INV_X1 U17933 ( .A(n18837), .ZN(n18841) );
  NAND2_X1 U17934 ( .A1(n18842), .A2(n18841), .ZN(n18840) );
  NOR2_X1 U17935 ( .A1(n14811), .A2(n18840), .ZN(n18821) );
  AOI21_X1 U17936 ( .B1(n18818), .B2(n14727), .A(n14726), .ZN(n18823) );
  INV_X1 U17937 ( .A(n18823), .ZN(n15200) );
  NAND2_X1 U17938 ( .A1(n18821), .A2(n15200), .ZN(n18806) );
  NOR2_X1 U17939 ( .A1(n14728), .A2(n18806), .ZN(n14798) );
  OAI21_X1 U17940 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n14730), .A(
        n14729), .ZN(n15186) );
  NAND2_X1 U17941 ( .A1(n14798), .A2(n15186), .ZN(n14792) );
  NOR2_X1 U17942 ( .A1(n14783), .A2(n14792), .ZN(n18793) );
  XNOR2_X1 U17943 ( .A(n14731), .B(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18794) );
  NAND2_X1 U17944 ( .A1(n18793), .A2(n18794), .ZN(n18785) );
  NOR2_X1 U17945 ( .A1(n18786), .A2(n18785), .ZN(n18768) );
  NOR2_X1 U17946 ( .A1(n14732), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14733) );
  NOR2_X1 U17947 ( .A1(n14734), .A2(n14733), .ZN(n18770) );
  INV_X1 U17948 ( .A(n18770), .ZN(n15141) );
  NAND2_X1 U17949 ( .A1(n18768), .A2(n15141), .ZN(n18758) );
  NOR2_X1 U17950 ( .A1(n18761), .A2(n18758), .ZN(n14770) );
  NOR2_X1 U17951 ( .A1(n18896), .A2(n14770), .ZN(n14769) );
  OAI21_X1 U17952 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n14735), .A(
        n14736), .ZN(n16136) );
  NAND2_X1 U17953 ( .A1(n15699), .A2(n16136), .ZN(n15698) );
  NAND2_X1 U17954 ( .A1(n18915), .A2(n15698), .ZN(n16094) );
  INV_X1 U17955 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15092) );
  AOI21_X1 U17956 ( .B1(n15092), .B2(n14736), .A(n14737), .ZN(n15095) );
  INV_X1 U17957 ( .A(n15095), .ZN(n16095) );
  NAND2_X1 U17958 ( .A1(n16094), .A2(n16095), .ZN(n16093) );
  NAND2_X1 U17959 ( .A1(n18915), .A2(n16093), .ZN(n16085) );
  OAI21_X1 U17960 ( .B1(n14737), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14738), .ZN(n16086) );
  NAND2_X1 U17961 ( .A1(n16085), .A2(n16086), .ZN(n16084) );
  NAND2_X1 U17962 ( .A1(n18915), .A2(n16084), .ZN(n16069) );
  AOI21_X1 U17963 ( .B1(n15075), .B2(n14738), .A(n9706), .ZN(n15073) );
  INV_X1 U17964 ( .A(n15073), .ZN(n16070) );
  NAND2_X1 U17965 ( .A1(n16069), .A2(n16070), .ZN(n16068) );
  NAND2_X1 U17966 ( .A1(n18915), .A2(n16068), .ZN(n16059) );
  OR2_X1 U17967 ( .A1(n9706), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14739) );
  NAND2_X1 U17968 ( .A1(n14740), .A2(n14739), .ZN(n16060) );
  NAND2_X1 U17969 ( .A1(n16059), .A2(n16060), .ZN(n16058) );
  NAND2_X1 U17970 ( .A1(n18915), .A2(n16058), .ZN(n14743) );
  NAND2_X1 U17971 ( .A1(n14740), .A2(n14759), .ZN(n14741) );
  NAND2_X1 U17972 ( .A1(n15044), .A2(n14741), .ZN(n15054) );
  NOR4_X1 U17973 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n19757), .ZN(n14742) );
  NAND2_X1 U17974 ( .A1(n14743), .A2(n15054), .ZN(n16011) );
  OAI211_X1 U17975 ( .C1(n14743), .C2(n15054), .A(n18901), .B(n16011), .ZN(
        n14765) );
  INV_X1 U17976 ( .A(n14744), .ZN(n14763) );
  AND2_X1 U17977 ( .A1(n16228), .A2(n19630), .ZN(n14745) );
  NOR2_X1 U17978 ( .A1(n14746), .A2(n14745), .ZN(n14748) );
  AND2_X1 U17979 ( .A1(n19890), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14747) );
  INV_X1 U17980 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16100) );
  NAND2_X1 U17981 ( .A1(n14748), .A2(n16100), .ZN(n14750) );
  INV_X1 U17982 ( .A(n14756), .ZN(n14749) );
  NAND2_X1 U17983 ( .A1(n19084), .A2(n14749), .ZN(n16015) );
  INV_X1 U17984 ( .A(n18935), .ZN(n18909) );
  INV_X1 U17985 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n14753) );
  INV_X1 U17986 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19811) );
  NAND2_X1 U17987 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19491), .ZN(n19751) );
  INV_X1 U17988 ( .A(n19751), .ZN(n19593) );
  AND2_X1 U17989 ( .A1(n19752), .A2(n19593), .ZN(n16229) );
  INV_X1 U17990 ( .A(n16229), .ZN(n14751) );
  NAND2_X1 U17991 ( .A1(n18934), .A2(n14751), .ZN(n14752) );
  OAI22_X1 U17992 ( .A1(n18909), .A2(n14753), .B1(n19811), .B2(n18873), .ZN(
        n14762) );
  AND2_X1 U17993 ( .A1(n14958), .A2(n14754), .ZN(n14755) );
  NOR2_X1 U17994 ( .A1(n14941), .A2(n14755), .ZN(n15251) );
  INV_X1 U17995 ( .A(n15251), .ZN(n14760) );
  AND2_X1 U17996 ( .A1(n14757), .A2(n14756), .ZN(n14758) );
  NOR2_X2 U17997 ( .A1(n18936), .A2(n19883), .ZN(n18950) );
  OAI22_X1 U17998 ( .A1(n14760), .A2(n18925), .B1(n14759), .B2(n18892), .ZN(
        n14761) );
  AOI211_X1 U17999 ( .C1(n14763), .C2(n18906), .A(n14762), .B(n14761), .ZN(
        n14764) );
  OAI211_X1 U18000 ( .C1(n15255), .C2(n18911), .A(n14765), .B(n14764), .ZN(
        P2_U2828) );
  XOR2_X1 U18001 ( .A(n14767), .B(n15340), .Z(n15337) );
  INV_X1 U18002 ( .A(n15337), .ZN(n14781) );
  INV_X1 U18003 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19799) );
  OAI22_X1 U18004 ( .A1(n14768), .A2(n18892), .B1(n19799), .B2(n18873), .ZN(
        n14775) );
  NOR2_X1 U18005 ( .A1(n14769), .A2(n18934), .ZN(n14773) );
  NAND2_X1 U18006 ( .A1(n18901), .A2(n18915), .ZN(n18839) );
  OR2_X1 U18007 ( .A1(n14770), .A2(n18839), .ZN(n18757) );
  INV_X1 U18008 ( .A(n18757), .ZN(n14772) );
  INV_X1 U18009 ( .A(n14771), .ZN(n15113) );
  MUX2_X1 U18010 ( .A(n14773), .B(n14772), .S(n15113), .Z(n14774) );
  AOI211_X1 U18011 ( .C1(P2_EBX_REG_21__SCAN_IN), .C2(n18935), .A(n14775), .B(
        n14774), .ZN(n14780) );
  NAND2_X1 U18012 ( .A1(n15125), .A2(n14776), .ZN(n14777) );
  NAND2_X1 U18013 ( .A1(n15313), .A2(n14777), .ZN(n15333) );
  INV_X1 U18014 ( .A(n15333), .ZN(n15117) );
  AOI22_X1 U18015 ( .A1(n14778), .A2(n18906), .B1(n15117), .B2(n18944), .ZN(
        n14779) );
  OAI211_X1 U18016 ( .C1(n14781), .C2(n18925), .A(n14780), .B(n14779), .ZN(
        P2_U2834) );
  NAND2_X1 U18017 ( .A1(n14711), .A2(n14792), .ZN(n14782) );
  NOR2_X1 U18018 ( .A1(n18934), .A2(n14782), .ZN(n14797) );
  INV_X1 U18019 ( .A(n14783), .ZN(n15170) );
  NAND2_X1 U18020 ( .A1(n14785), .A2(n14784), .ZN(n14786) );
  NAND2_X1 U18021 ( .A1(n14928), .A2(n14786), .ZN(n18957) );
  INV_X1 U18022 ( .A(n18957), .ZN(n15173) );
  AOI22_X1 U18023 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18950), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n18936), .ZN(n14787) );
  OAI211_X1 U18024 ( .C1(n18909), .C2(n14788), .A(n14787), .B(n18871), .ZN(
        n14789) );
  AOI21_X1 U18025 ( .B1(n15173), .B2(n18944), .A(n14789), .ZN(n14790) );
  OAI21_X1 U18026 ( .B1(n14791), .B2(n18941), .A(n14790), .ZN(n14794) );
  AOI211_X1 U18027 ( .C1(n18915), .C2(n14792), .A(n15170), .B(n18934), .ZN(
        n14793) );
  AOI211_X1 U18028 ( .C1(n14797), .C2(n15170), .A(n14794), .B(n14793), .ZN(
        n14795) );
  OAI21_X1 U18029 ( .B1(n14796), .B2(n18925), .A(n14795), .ZN(P2_U2839) );
  OAI21_X1 U18030 ( .B1(n14798), .B2(n15186), .A(n14797), .ZN(n14801) );
  INV_X1 U18031 ( .A(n15407), .ZN(n14799) );
  AOI22_X1 U18032 ( .A1(n14799), .A2(n18944), .B1(n18935), .B2(
        P2_EBX_REG_15__SCAN_IN), .ZN(n14800) );
  OAI211_X1 U18033 ( .C1(n14802), .C2(n18941), .A(n14801), .B(n14800), .ZN(
        n14806) );
  INV_X1 U18034 ( .A(n18949), .ZN(n14804) );
  AOI22_X1 U18035 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18950), .B1(
        P2_REIP_REG_15__SCAN_IN), .B2(n18936), .ZN(n14803) );
  OAI211_X1 U18036 ( .C1(n15186), .C2(n14804), .A(n14803), .B(n18871), .ZN(
        n14805) );
  NOR2_X1 U18037 ( .A1(n14806), .A2(n14805), .ZN(n14807) );
  OAI21_X1 U18038 ( .B1(n15411), .B2(n18925), .A(n14807), .ZN(P2_U2840) );
  XNOR2_X1 U18039 ( .A(n14809), .B(n14808), .ZN(n18997) );
  NAND2_X1 U18040 ( .A1(n14711), .A2(n18840), .ZN(n14810) );
  XNOR2_X1 U18041 ( .A(n14811), .B(n14810), .ZN(n14812) );
  NAND2_X1 U18042 ( .A1(n14812), .A2(n18901), .ZN(n14822) );
  OR2_X1 U18043 ( .A1(n14814), .A2(n14813), .ZN(n14815) );
  NAND2_X1 U18044 ( .A1(n13514), .A2(n14815), .ZN(n18968) );
  INV_X1 U18045 ( .A(n18968), .ZN(n16143) );
  AOI22_X1 U18046 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(n18935), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18950), .ZN(n14816) );
  OAI211_X1 U18047 ( .C1(n18873), .C2(n14817), .A(n14816), .B(n18871), .ZN(
        n14820) );
  NOR2_X1 U18048 ( .A1(n14818), .A2(n18941), .ZN(n14819) );
  AOI211_X1 U18049 ( .C1(n18944), .C2(n16143), .A(n14820), .B(n14819), .ZN(
        n14821) );
  OAI211_X1 U18050 ( .C1(n18925), .C2(n18997), .A(n14822), .B(n14821), .ZN(
        P2_U2843) );
  XNOR2_X1 U18051 ( .A(n14823), .B(n14824), .ZN(n19000) );
  NAND2_X1 U18052 ( .A1(n14711), .A2(n14825), .ZN(n14826) );
  XNOR2_X1 U18053 ( .A(n14827), .B(n14826), .ZN(n14828) );
  NAND2_X1 U18054 ( .A1(n14828), .A2(n18901), .ZN(n14837) );
  OAI21_X1 U18055 ( .B1(n11970), .B2(n18873), .A(n13051), .ZN(n14834) );
  OR2_X1 U18056 ( .A1(n9711), .A2(n14829), .ZN(n14831) );
  AND2_X1 U18057 ( .A1(n14831), .A2(n14830), .ZN(n16158) );
  INV_X1 U18058 ( .A(n16158), .ZN(n18973) );
  AOI22_X1 U18059 ( .A1(n18935), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18950), .ZN(n14832) );
  OAI21_X1 U18060 ( .B1(n18973), .B2(n18911), .A(n14832), .ZN(n14833) );
  AOI211_X1 U18061 ( .C1(n14835), .C2(n18906), .A(n14834), .B(n14833), .ZN(
        n14836) );
  OAI211_X1 U18062 ( .C1(n18925), .C2(n19000), .A(n14837), .B(n14836), .ZN(
        P2_U2845) );
  NOR2_X1 U18063 ( .A1(n18896), .A2(n14838), .ZN(n14840) );
  XNOR2_X1 U18064 ( .A(n14840), .B(n14839), .ZN(n14852) );
  INV_X1 U18065 ( .A(n18948), .ZN(n18912) );
  NOR2_X1 U18066 ( .A1(n19450), .A2(n18912), .ZN(n14851) );
  NOR2_X1 U18067 ( .A1(n18892), .A2(n14841), .ZN(n14842) );
  AOI21_X1 U18068 ( .B1(n18935), .B2(P2_EBX_REG_3__SCAN_IN), .A(n14842), .ZN(
        n14844) );
  OR2_X1 U18069 ( .A1(n18873), .A2(n13493), .ZN(n14843) );
  OAI211_X1 U18070 ( .C1(n14845), .C2(n18941), .A(n14844), .B(n14843), .ZN(
        n14846) );
  AOI21_X1 U18071 ( .B1(n14847), .B2(n18944), .A(n14846), .ZN(n14848) );
  OAI21_X1 U18072 ( .B1(n14849), .B2(n18925), .A(n14848), .ZN(n14850) );
  AOI211_X1 U18073 ( .C1(n14852), .C2(n18901), .A(n14851), .B(n14850), .ZN(
        n14853) );
  INV_X1 U18074 ( .A(n14853), .ZN(P2_U2852) );
  NAND2_X1 U18075 ( .A1(n14711), .A2(n15538), .ZN(n14854) );
  XNOR2_X1 U18076 ( .A(n14855), .B(n14854), .ZN(n14856) );
  NAND2_X1 U18077 ( .A1(n14856), .A2(n18901), .ZN(n14864) );
  AOI22_X1 U18078 ( .A1(n18935), .A2(P2_EBX_REG_2__SCAN_IN), .B1(n18950), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14857) );
  OAI21_X1 U18079 ( .B1(n19777), .B2(n18873), .A(n14857), .ZN(n14858) );
  AOI21_X1 U18080 ( .B1(n14859), .B2(n18906), .A(n14858), .ZN(n14860) );
  OAI21_X1 U18081 ( .B1(n14861), .B2(n18911), .A(n14860), .ZN(n14862) );
  AOI21_X1 U18082 ( .B1(n19847), .B2(n18937), .A(n14862), .ZN(n14863) );
  OAI211_X1 U18083 ( .C1(n18912), .C2(n19845), .A(n14864), .B(n14863), .ZN(
        P2_U2853) );
  NAND3_X1 U18084 ( .A1(n14933), .A2(n14866), .A3(n18954), .ZN(n14868) );
  NAND2_X1 U18085 ( .A1(n18983), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14867) );
  OAI211_X1 U18086 ( .C1(n18983), .C2(n15032), .A(n14868), .B(n14867), .ZN(
        P2_U2858) );
  NOR2_X1 U18087 ( .A1(n13992), .A2(n14869), .ZN(n14871) );
  XNOR2_X1 U18088 ( .A(n14871), .B(n14870), .ZN(n14949) );
  NOR2_X1 U18089 ( .A1(n14704), .A2(n14872), .ZN(n14873) );
  NOR2_X1 U18090 ( .A1(n16053), .A2(n18983), .ZN(n14874) );
  AOI21_X1 U18091 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n18983), .A(n14874), .ZN(
        n14875) );
  OAI21_X1 U18092 ( .B1(n14949), .B2(n18984), .A(n14875), .ZN(P2_U2859) );
  CLKBUF_X1 U18093 ( .A(n14876), .Z(n14877) );
  OAI21_X1 U18094 ( .B1(n14877), .B2(n14879), .A(n14878), .ZN(n14954) );
  NOR2_X1 U18095 ( .A1(n15255), .A2(n18983), .ZN(n14880) );
  AOI21_X1 U18096 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n18983), .A(n14880), .ZN(
        n14881) );
  OAI21_X1 U18097 ( .B1(n14954), .B2(n18984), .A(n14881), .ZN(P2_U2860) );
  AOI21_X1 U18098 ( .B1(n14882), .B2(n14884), .A(n14883), .ZN(n14885) );
  INV_X1 U18099 ( .A(n14885), .ZN(n14964) );
  NOR2_X1 U18100 ( .A1(n14886), .A2(n14887), .ZN(n14888) );
  OR2_X1 U18101 ( .A1(n14705), .A2(n14888), .ZN(n16056) );
  NOR2_X1 U18102 ( .A1(n16056), .A2(n18983), .ZN(n14889) );
  AOI21_X1 U18103 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n18983), .A(n14889), .ZN(
        n14890) );
  OAI21_X1 U18104 ( .B1(n14964), .B2(n18984), .A(n14890), .ZN(P2_U2861) );
  OAI21_X1 U18105 ( .B1(n14891), .B2(n14893), .A(n14892), .ZN(n14973) );
  NAND2_X1 U18106 ( .A1(n18983), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n14897) );
  AND2_X1 U18107 ( .A1(n14904), .A2(n14894), .ZN(n14895) );
  NOR2_X1 U18108 ( .A1(n14886), .A2(n14895), .ZN(n16067) );
  NAND2_X1 U18109 ( .A1(n16067), .A2(n18988), .ZN(n14896) );
  OAI211_X1 U18110 ( .C1(n14973), .C2(n18984), .A(n14897), .B(n14896), .ZN(
        P2_U2862) );
  OR2_X1 U18111 ( .A1(n14900), .A2(n14899), .ZN(n14974) );
  NAND3_X1 U18112 ( .A1(n14898), .A2(n14974), .A3(n18954), .ZN(n14906) );
  NAND2_X1 U18113 ( .A1(n14901), .A2(n14902), .ZN(n14903) );
  NAND2_X1 U18114 ( .A1(n14904), .A2(n14903), .ZN(n16089) );
  INV_X1 U18115 ( .A(n16089), .ZN(n15291) );
  NAND2_X1 U18116 ( .A1(n15291), .A2(n18988), .ZN(n14905) );
  OAI211_X1 U18117 ( .C1(n18988), .C2(n9809), .A(n14906), .B(n14905), .ZN(
        P2_U2863) );
  OAI21_X1 U18118 ( .B1(n14907), .B2(n14909), .A(n14908), .ZN(n14993) );
  OAI21_X1 U18119 ( .B1(n15315), .B2(n14910), .A(n14901), .ZN(n15294) );
  NOR2_X1 U18120 ( .A1(n15294), .A2(n18983), .ZN(n14911) );
  AOI21_X1 U18121 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n18983), .A(n14911), .ZN(
        n14912) );
  OAI21_X1 U18122 ( .B1(n14993), .B2(n18984), .A(n14912), .ZN(P2_U2864) );
  OR2_X1 U18123 ( .A1(n14914), .A2(n14915), .ZN(n14916) );
  NAND2_X1 U18124 ( .A1(n14913), .A2(n14916), .ZN(n14997) );
  MUX2_X1 U18125 ( .A(n15333), .B(n14917), .S(n18983), .Z(n14918) );
  OAI21_X1 U18126 ( .B1(n14997), .B2(n18984), .A(n14918), .ZN(P2_U2866) );
  OR2_X1 U18127 ( .A1(n15152), .A2(n14919), .ZN(n14920) );
  NAND2_X1 U18128 ( .A1(n15123), .A2(n14920), .ZN(n18775) );
  AOI21_X1 U18129 ( .B1(n14923), .B2(n14921), .A(n14922), .ZN(n20790) );
  NAND2_X1 U18130 ( .A1(n20790), .A2(n18954), .ZN(n14925) );
  NAND2_X1 U18131 ( .A1(n18983), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14924) );
  OAI211_X1 U18132 ( .C1(n18775), .C2(n18983), .A(n14925), .B(n14924), .ZN(
        P2_U2868) );
  AND2_X1 U18133 ( .A1(n14928), .A2(n14927), .ZN(n14929) );
  NOR2_X1 U18134 ( .A1(n14926), .A2(n14929), .ZN(n15387) );
  INV_X1 U18135 ( .A(n15387), .ZN(n18800) );
  NOR2_X1 U18136 ( .A1(n18800), .A2(n18983), .ZN(n14930) );
  AOI21_X1 U18137 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n18983), .A(n14930), .ZN(
        n14931) );
  OAI21_X1 U18138 ( .B1(n14932), .B2(n18984), .A(n14931), .ZN(P2_U2870) );
  NAND3_X1 U18139 ( .A1(n14933), .A2(n14866), .A3(n20791), .ZN(n14939) );
  INV_X1 U18140 ( .A(n19083), .ZN(n14934) );
  AOI22_X1 U18141 ( .A1(n20782), .A2(n14934), .B1(n20780), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n14938) );
  AOI22_X1 U18142 ( .A1(n20784), .A2(BUF2_REG_29__SCAN_IN), .B1(n20783), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14937) );
  INV_X1 U18143 ( .A(n14935), .ZN(n16034) );
  NAND2_X1 U18144 ( .A1(n16034), .A2(n18989), .ZN(n14936) );
  NAND4_X1 U18145 ( .A1(n14939), .A2(n14938), .A3(n14937), .A4(n14936), .ZN(
        P2_U2890) );
  NOR2_X1 U18146 ( .A1(n14941), .A2(n14940), .ZN(n14942) );
  OR2_X1 U18147 ( .A1(n12262), .A2(n14942), .ZN(n16044) );
  AOI22_X1 U18148 ( .A1(n20784), .A2(BUF2_REG_28__SCAN_IN), .B1(n20783), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14946) );
  NAND2_X1 U18149 ( .A1(n19101), .A2(BUF2_REG_12__SCAN_IN), .ZN(n14944) );
  OR2_X1 U18150 ( .A1(n19101), .A2(n16325), .ZN(n14943) );
  NAND2_X1 U18151 ( .A1(n14944), .A2(n14943), .ZN(n19062) );
  AOI22_X1 U18152 ( .A1(n20782), .A2(n19062), .B1(n20780), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n14945) );
  OAI211_X1 U18153 ( .C1(n16044), .C2(n20787), .A(n14946), .B(n14945), .ZN(
        n14947) );
  INV_X1 U18154 ( .A(n14947), .ZN(n14948) );
  OAI21_X1 U18155 ( .B1(n14949), .B2(n14996), .A(n14948), .ZN(P2_U2891) );
  AOI22_X1 U18156 ( .A1(n15251), .A2(n18989), .B1(n20784), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n14953) );
  OAI22_X1 U18157 ( .A1(n14980), .A2(n19078), .B1(n14979), .B2(n14950), .ZN(
        n14951) );
  AOI21_X1 U18158 ( .B1(n20783), .B2(BUF1_REG_27__SCAN_IN), .A(n14951), .ZN(
        n14952) );
  OAI211_X1 U18159 ( .C1(n14954), .C2(n14996), .A(n14953), .B(n14952), .ZN(
        P2_U2892) );
  NAND2_X1 U18160 ( .A1(n14956), .A2(n14955), .ZN(n14957) );
  NAND2_X1 U18161 ( .A1(n14958), .A2(n14957), .ZN(n16055) );
  OAI22_X1 U18162 ( .A1(n20787), .A2(n16055), .B1(n14979), .B2(n12890), .ZN(
        n14962) );
  INV_X1 U18163 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n14960) );
  OAI22_X1 U18164 ( .A1(n14969), .A2(n14960), .B1(n14980), .B2(n14959), .ZN(
        n14961) );
  AOI211_X1 U18165 ( .C1(n20783), .C2(BUF1_REG_26__SCAN_IN), .A(n14962), .B(
        n14961), .ZN(n14963) );
  OAI21_X1 U18166 ( .B1(n14964), .B2(n14996), .A(n14963), .ZN(P2_U2893) );
  XNOR2_X1 U18167 ( .A(n14965), .B(n9710), .ZN(n16066) );
  INV_X1 U18168 ( .A(n16066), .ZN(n14967) );
  OAI22_X1 U18169 ( .A1(n20787), .A2(n14967), .B1(n14979), .B2(n14966), .ZN(
        n14971) );
  OAI22_X1 U18170 ( .A1(n14969), .A2(n19117), .B1(n14980), .B2(n14968), .ZN(
        n14970) );
  AOI211_X1 U18171 ( .C1(n20783), .C2(BUF1_REG_25__SCAN_IN), .A(n14971), .B(
        n14970), .ZN(n14972) );
  OAI21_X1 U18172 ( .B1(n14973), .B2(n14996), .A(n14972), .ZN(P2_U2894) );
  NAND3_X1 U18173 ( .A1(n14898), .A2(n14974), .A3(n20791), .ZN(n14984) );
  OR2_X1 U18174 ( .A1(n14976), .A2(n14975), .ZN(n14977) );
  AND2_X1 U18175 ( .A1(n14965), .A2(n14977), .ZN(n16080) );
  AOI22_X1 U18176 ( .A1(n18989), .A2(n16080), .B1(n20784), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n14983) );
  OAI22_X1 U18177 ( .A1(n14980), .A2(n19076), .B1(n14979), .B2(n14978), .ZN(
        n14981) );
  AOI21_X1 U18178 ( .B1(n20783), .B2(BUF1_REG_24__SCAN_IN), .A(n14981), .ZN(
        n14982) );
  NAND3_X1 U18179 ( .A1(n14984), .A2(n14983), .A3(n14982), .ZN(P2_U2895) );
  INV_X1 U18180 ( .A(n14985), .ZN(n14987) );
  XNOR2_X1 U18181 ( .A(n14987), .B(n14986), .ZN(n16091) );
  AOI22_X1 U18182 ( .A1(n18989), .A2(n16091), .B1(n20784), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n14991) );
  INV_X1 U18183 ( .A(n19161), .ZN(n14988) );
  AOI22_X1 U18184 ( .A1(n20782), .A2(n14988), .B1(n20780), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n14990) );
  NAND2_X1 U18185 ( .A1(n20783), .A2(BUF1_REG_23__SCAN_IN), .ZN(n14989) );
  AND3_X1 U18186 ( .A1(n14991), .A2(n14990), .A3(n14989), .ZN(n14992) );
  OAI21_X1 U18187 ( .B1(n14993), .B2(n14996), .A(n14992), .ZN(P2_U2896) );
  AOI22_X1 U18188 ( .A1(n19103), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19101), .ZN(n19145) );
  INV_X1 U18189 ( .A(n19145), .ZN(n19004) );
  AOI22_X1 U18190 ( .A1(n20782), .A2(n19004), .B1(n20780), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n14995) );
  AOI22_X1 U18191 ( .A1(n20784), .A2(BUF2_REG_21__SCAN_IN), .B1(n20783), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n14994) );
  OAI211_X1 U18192 ( .C1(n14997), .C2(n14996), .A(n14995), .B(n14994), .ZN(
        n14998) );
  AOI21_X1 U18193 ( .B1(n15337), .B2(n18989), .A(n14998), .ZN(n14999) );
  INV_X1 U18194 ( .A(n14999), .ZN(P2_U2898) );
  NOR2_X1 U18195 ( .A1(n15004), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n15005) );
  MUX2_X1 U18196 ( .A(n15006), .B(n15005), .S(n11440), .Z(n16013) );
  NAND2_X1 U18197 ( .A1(n16013), .A2(n11814), .ZN(n15007) );
  XNOR2_X1 U18198 ( .A(n15007), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15008) );
  XNOR2_X1 U18199 ( .A(n15009), .B(n15008), .ZN(n15239) );
  NAND2_X1 U18200 ( .A1(n15013), .A2(n15012), .ZN(n15021) );
  INV_X1 U18201 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19820) );
  NAND2_X1 U18202 ( .A1(n15014), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n15016) );
  NAND2_X1 U18203 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15015) );
  OAI211_X1 U18204 ( .C1(n19820), .C2(n9610), .A(n15016), .B(n15015), .ZN(
        n15018) );
  AOI21_X1 U18205 ( .B1(n15019), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n15018), .ZN(n15020) );
  NOR2_X1 U18206 ( .A1(n18871), .A2(n19820), .ZN(n15234) );
  NOR2_X1 U18207 ( .A1(n16166), .A2(n15022), .ZN(n15023) );
  AOI211_X1 U18208 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n16156), .A(
        n15234), .B(n15023), .ZN(n15024) );
  OAI21_X1 U18209 ( .B1(n16101), .B2(n19102), .A(n15024), .ZN(n15025) );
  AOI21_X1 U18210 ( .B1(n15238), .B2(n19091), .A(n15025), .ZN(n15026) );
  OAI21_X1 U18211 ( .B1(n15239), .B2(n16168), .A(n15026), .ZN(P2_U2983) );
  AOI21_X1 U18212 ( .B1(n15029), .B2(n15046), .A(n15027), .ZN(n16012) );
  OAI21_X1 U18213 ( .B1(n19100), .B2(n15029), .A(n15028), .ZN(n15030) );
  AOI21_X1 U18214 ( .B1(n19089), .B2(n16012), .A(n15030), .ZN(n15031) );
  OAI21_X1 U18215 ( .B1(n15032), .B2(n19102), .A(n15031), .ZN(n15033) );
  AOI21_X1 U18216 ( .B1(n15034), .B2(n19091), .A(n15033), .ZN(n15035) );
  OAI21_X1 U18217 ( .B1(n15036), .B2(n16168), .A(n15035), .ZN(P2_U2985) );
  XNOR2_X1 U18218 ( .A(n15039), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15040) );
  XNOR2_X1 U18219 ( .A(n15041), .B(n15040), .ZN(n15248) );
  XNOR2_X1 U18220 ( .A(n15052), .B(n15042), .ZN(n15246) );
  NOR2_X1 U18221 ( .A1(n16053), .A2(n19102), .ZN(n15049) );
  NAND2_X1 U18222 ( .A1(n15044), .A2(n15043), .ZN(n15045) );
  NAND2_X1 U18223 ( .A1(n15046), .A2(n15045), .ZN(n16050) );
  NAND2_X1 U18224 ( .A1(n19090), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15241) );
  NAND2_X1 U18225 ( .A1(n16156), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15047) );
  OAI211_X1 U18226 ( .C1(n16166), .C2(n16050), .A(n15241), .B(n15047), .ZN(
        n15048) );
  AOI211_X1 U18227 ( .C1(n15246), .C2(n19091), .A(n15049), .B(n15048), .ZN(
        n15050) );
  OAI21_X1 U18228 ( .B1(n15248), .B2(n16168), .A(n15050), .ZN(P2_U2986) );
  XNOR2_X1 U18229 ( .A(n15051), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15259) );
  AOI21_X1 U18230 ( .B1(n15053), .B2(n15063), .A(n15052), .ZN(n15257) );
  NOR2_X1 U18231 ( .A1(n18871), .A2(n19811), .ZN(n15249) );
  NOR2_X1 U18232 ( .A1(n16166), .A2(n15054), .ZN(n15055) );
  AOI211_X1 U18233 ( .C1(n16156), .C2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15249), .B(n15055), .ZN(n15056) );
  OAI21_X1 U18234 ( .B1(n15255), .B2(n19102), .A(n15056), .ZN(n15057) );
  AOI21_X1 U18235 ( .B1(n15257), .B2(n19091), .A(n15057), .ZN(n15058) );
  OAI21_X1 U18236 ( .B1(n15259), .B2(n16168), .A(n15058), .ZN(P2_U2987) );
  AOI21_X1 U18237 ( .B1(n9803), .B2(n15069), .A(n15071), .ZN(n15061) );
  XNOR2_X1 U18238 ( .A(n15061), .B(n15060), .ZN(n15270) );
  OAI21_X1 U18239 ( .B1(n15085), .B2(n15276), .A(n15062), .ZN(n15064) );
  AND2_X1 U18240 ( .A1(n15064), .A2(n15063), .ZN(n15268) );
  INV_X1 U18241 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19808) );
  NOR2_X1 U18242 ( .A1(n18871), .A2(n19808), .ZN(n15261) );
  NOR2_X1 U18243 ( .A1(n16166), .A2(n16060), .ZN(n15065) );
  AOI211_X1 U18244 ( .C1(n16156), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15261), .B(n15065), .ZN(n15066) );
  OAI21_X1 U18245 ( .B1(n16056), .B2(n19102), .A(n15066), .ZN(n15067) );
  AOI21_X1 U18246 ( .B1(n15268), .B2(n19091), .A(n15067), .ZN(n15068) );
  OAI21_X1 U18247 ( .B1(n15270), .B2(n16168), .A(n15068), .ZN(P2_U2988) );
  INV_X1 U18248 ( .A(n15069), .ZN(n15070) );
  NOR2_X1 U18249 ( .A1(n15071), .A2(n15070), .ZN(n15072) );
  XNOR2_X1 U18250 ( .A(n9803), .B(n15072), .ZN(n15282) );
  NAND2_X1 U18251 ( .A1(n19089), .A2(n15073), .ZN(n15074) );
  NAND2_X1 U18252 ( .A1(n19090), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15272) );
  OAI211_X1 U18253 ( .C1(n19100), .C2(n15075), .A(n15074), .B(n15272), .ZN(
        n15077) );
  XNOR2_X1 U18254 ( .A(n15085), .B(n15276), .ZN(n15278) );
  NOR2_X1 U18255 ( .A1(n15278), .A2(n16169), .ZN(n15076) );
  AOI211_X1 U18256 ( .C1(n19094), .C2(n16067), .A(n15077), .B(n15076), .ZN(
        n15078) );
  OAI21_X1 U18257 ( .B1(n15282), .B2(n16168), .A(n15078), .ZN(P2_U2989) );
  INV_X1 U18258 ( .A(n15080), .ZN(n15082) );
  NOR2_X1 U18259 ( .A1(n15082), .A2(n15081), .ZN(n15083) );
  XNOR2_X1 U18260 ( .A(n15079), .B(n15083), .ZN(n15293) );
  NOR2_X1 U18261 ( .A1(n18871), .A2(n19804), .ZN(n15285) );
  AOI21_X1 U18262 ( .B1(n16156), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15285), .ZN(n15084) );
  OAI21_X1 U18263 ( .B1(n16166), .B2(n16086), .A(n15084), .ZN(n15087) );
  OAI21_X1 U18264 ( .B1(n15090), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15085), .ZN(n15288) );
  NOR2_X1 U18265 ( .A1(n15288), .A2(n16169), .ZN(n15086) );
  AOI211_X1 U18266 ( .C1(n19094), .C2(n15291), .A(n15087), .B(n15086), .ZN(
        n15088) );
  OAI21_X1 U18267 ( .B1(n15293), .B2(n16168), .A(n15088), .ZN(P2_U2990) );
  INV_X1 U18268 ( .A(n15305), .ZN(n15089) );
  NAND2_X1 U18269 ( .A1(n15089), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15307) );
  INV_X1 U18270 ( .A(n15307), .ZN(n15091) );
  OAI21_X1 U18271 ( .B1(n15091), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n9834), .ZN(n15304) );
  INV_X1 U18272 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19802) );
  OAI22_X1 U18273 ( .A1(n19100), .A2(n15092), .B1(n19802), .B2(n18871), .ZN(
        n15094) );
  NOR2_X1 U18274 ( .A1(n15294), .A2(n19102), .ZN(n15093) );
  AOI211_X1 U18275 ( .C1(n19089), .C2(n15095), .A(n15094), .B(n15093), .ZN(
        n15100) );
  OR2_X1 U18276 ( .A1(n15097), .A2(n15096), .ZN(n15301) );
  NAND3_X1 U18277 ( .A1(n15301), .A2(n15098), .A3(n19095), .ZN(n15099) );
  OAI211_X1 U18278 ( .C1(n15304), .C2(n16169), .A(n15100), .B(n15099), .ZN(
        P2_U2991) );
  NAND2_X1 U18279 ( .A1(n15102), .A2(n15101), .ZN(n15111) );
  NAND2_X1 U18280 ( .A1(n15183), .A2(n15103), .ZN(n15104) );
  INV_X1 U18281 ( .A(n15167), .ZN(n15106) );
  NAND2_X1 U18282 ( .A1(n15109), .A2(n15108), .ZN(n15161) );
  INV_X1 U18283 ( .A(n15137), .ZN(n15110) );
  OAI211_X1 U18284 ( .C1(n15136), .C2(n15110), .A(n15148), .B(n15138), .ZN(
        n15122) );
  NOR2_X1 U18285 ( .A1(n18871), .A2(n19799), .ZN(n15329) );
  AOI21_X1 U18286 ( .B1(n16156), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15329), .ZN(n15112) );
  OAI21_X1 U18287 ( .B1(n16166), .B2(n15113), .A(n15112), .ZN(n15116) );
  NAND2_X1 U18288 ( .A1(n15131), .A2(n15330), .ZN(n15114) );
  NAND2_X1 U18289 ( .A1(n15305), .A2(n15114), .ZN(n15334) );
  NOR2_X1 U18290 ( .A1(n15334), .A2(n16169), .ZN(n15115) );
  AOI211_X1 U18291 ( .C1(n19094), .C2(n15117), .A(n15116), .B(n15115), .ZN(
        n15118) );
  NAND2_X1 U18292 ( .A1(n15120), .A2(n15119), .ZN(n15121) );
  XNOR2_X1 U18293 ( .A(n15122), .B(n15121), .ZN(n15351) );
  INV_X1 U18294 ( .A(n15123), .ZN(n15127) );
  INV_X1 U18295 ( .A(n15124), .ZN(n15126) );
  OAI21_X1 U18296 ( .B1(n15127), .B2(n15126), .A(n15125), .ZN(n16109) );
  INV_X1 U18297 ( .A(n16109), .ZN(n18762) );
  NOR2_X1 U18298 ( .A1(n18871), .A2(n15128), .ZN(n15343) );
  AOI21_X1 U18299 ( .B1(n16156), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15343), .ZN(n15129) );
  OAI21_X1 U18300 ( .B1(n15130), .B2(n16166), .A(n15129), .ZN(n15134) );
  OAI21_X1 U18301 ( .B1(n9837), .B2(n15357), .A(n15342), .ZN(n15132) );
  NAND2_X1 U18302 ( .A1(n15132), .A2(n15131), .ZN(n15347) );
  NOR2_X1 U18303 ( .A1(n15347), .A2(n16169), .ZN(n15133) );
  AOI211_X1 U18304 ( .C1(n19094), .C2(n18762), .A(n15134), .B(n15133), .ZN(
        n15135) );
  OAI21_X1 U18305 ( .B1(n15351), .B2(n16168), .A(n15135), .ZN(P2_U2994) );
  NAND2_X1 U18306 ( .A1(n15136), .A2(n15148), .ZN(n15140) );
  NAND2_X1 U18307 ( .A1(n15138), .A2(n15137), .ZN(n15139) );
  XNOR2_X1 U18308 ( .A(n15140), .B(n15139), .ZN(n15365) );
  XNOR2_X1 U18309 ( .A(n15150), .B(n15357), .ZN(n15363) );
  INV_X1 U18310 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19796) );
  NOR2_X1 U18311 ( .A1(n18871), .A2(n19796), .ZN(n15356) );
  NOR2_X1 U18312 ( .A1(n15141), .A2(n16166), .ZN(n15142) );
  AOI211_X1 U18313 ( .C1(n16156), .C2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15356), .B(n15142), .ZN(n15143) );
  OAI21_X1 U18314 ( .B1(n19102), .B2(n18775), .A(n15143), .ZN(n15144) );
  AOI21_X1 U18315 ( .B1(n15363), .B2(n19091), .A(n15144), .ZN(n15145) );
  OAI21_X1 U18316 ( .B1(n15365), .B2(n16168), .A(n15145), .ZN(P2_U2995) );
  NAND2_X1 U18317 ( .A1(n15148), .A2(n15147), .ZN(n15149) );
  XNOR2_X1 U18318 ( .A(n15146), .B(n15149), .ZN(n15378) );
  INV_X1 U18319 ( .A(n15421), .ZN(n15175) );
  NOR2_X2 U18320 ( .A1(n15175), .A2(n15385), .ZN(n15380) );
  AOI21_X1 U18321 ( .B1(n15380), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15151) );
  NOR2_X1 U18322 ( .A1(n15151), .A2(n15150), .ZN(n15376) );
  INV_X1 U18323 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19794) );
  NOR2_X1 U18324 ( .A1(n18871), .A2(n19794), .ZN(n15370) );
  INV_X1 U18325 ( .A(n15152), .ZN(n15153) );
  OAI21_X1 U18326 ( .B1(n14926), .B2(n15154), .A(n15153), .ZN(n18792) );
  NOR2_X1 U18327 ( .A1(n18792), .A2(n19102), .ZN(n15155) );
  AOI211_X1 U18328 ( .C1(n16156), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15370), .B(n15155), .ZN(n15156) );
  OAI21_X1 U18329 ( .B1(n16166), .B2(n15157), .A(n15156), .ZN(n15158) );
  AOI21_X1 U18330 ( .B1(n15376), .B2(n19091), .A(n15158), .ZN(n15159) );
  OAI21_X1 U18331 ( .B1(n15378), .B2(n16168), .A(n15159), .ZN(P2_U2996) );
  XOR2_X1 U18332 ( .A(n15161), .B(n15160), .Z(n15393) );
  XNOR2_X1 U18333 ( .A(n15380), .B(n15368), .ZN(n15165) );
  NAND2_X1 U18334 ( .A1(n15387), .A2(n19094), .ZN(n15163) );
  NOR2_X1 U18335 ( .A1(n18871), .A2(n20892), .ZN(n15386) );
  AOI21_X1 U18336 ( .B1(n16156), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15386), .ZN(n15162) );
  OAI211_X1 U18337 ( .C1(n18794), .C2(n16166), .A(n15163), .B(n15162), .ZN(
        n15164) );
  AOI21_X1 U18338 ( .B1(n15165), .B2(n19091), .A(n15164), .ZN(n15166) );
  OAI21_X1 U18339 ( .B1(n15393), .B2(n16168), .A(n15166), .ZN(P2_U2997) );
  XNOR2_X1 U18340 ( .A(n15168), .B(n15167), .ZN(n15399) );
  INV_X1 U18341 ( .A(n15399), .ZN(n15180) );
  NAND2_X1 U18342 ( .A1(n18784), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15394) );
  OAI21_X1 U18343 ( .B1(n19100), .B2(n15169), .A(n15394), .ZN(n15172) );
  NOR2_X1 U18344 ( .A1(n15170), .A2(n16166), .ZN(n15171) );
  AOI211_X1 U18345 ( .C1(n15173), .C2(n19094), .A(n15172), .B(n15171), .ZN(
        n15179) );
  INV_X1 U18346 ( .A(n15380), .ZN(n15177) );
  OAI21_X1 U18347 ( .B1(n15175), .B2(n15404), .A(n15174), .ZN(n15176) );
  NAND3_X1 U18348 ( .A1(n15177), .A2(n19091), .A3(n15176), .ZN(n15178) );
  OAI211_X1 U18349 ( .C1(n15180), .C2(n16168), .A(n15179), .B(n15178), .ZN(
        P2_U2998) );
  NAND2_X1 U18350 ( .A1(n15182), .A2(n15181), .ZN(n15185) );
  NAND2_X1 U18351 ( .A1(n15183), .A2(n15417), .ZN(n15184) );
  XOR2_X1 U18352 ( .A(n15185), .B(n15184), .Z(n15415) );
  XNOR2_X1 U18353 ( .A(n15421), .B(n15404), .ZN(n15413) );
  INV_X1 U18354 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15187) );
  OAI22_X1 U18355 ( .A1(n19100), .A2(n15187), .B1(n16166), .B2(n15186), .ZN(
        n15190) );
  INV_X1 U18356 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n15188) );
  OAI22_X1 U18357 ( .A1(n19102), .A2(n15407), .B1(n15188), .B2(n18871), .ZN(
        n15189) );
  AOI211_X1 U18358 ( .C1(n15413), .C2(n19091), .A(n15190), .B(n15189), .ZN(
        n15191) );
  OAI21_X1 U18359 ( .B1(n15415), .B2(n16168), .A(n15191), .ZN(P2_U2999) );
  NAND2_X1 U18360 ( .A1(n15194), .A2(n15193), .ZN(n15195) );
  XNOR2_X1 U18361 ( .A(n15192), .B(n15195), .ZN(n15450) );
  NAND2_X1 U18362 ( .A1(n15196), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15515) );
  NAND2_X1 U18363 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15461), .ZN(
        n15462) );
  INV_X1 U18364 ( .A(n15461), .ZN(n15474) );
  NOR2_X1 U18365 ( .A1(n15474), .A2(n15433), .ZN(n15420) );
  AOI21_X1 U18366 ( .B1(n15197), .B2(n15462), .A(n15420), .ZN(n15198) );
  INV_X1 U18367 ( .A(n15198), .ZN(n15446) );
  OR2_X1 U18368 ( .A1(n13051), .A2(n15199), .ZN(n15443) );
  OAI21_X1 U18369 ( .B1(n16169), .B2(n15446), .A(n15443), .ZN(n15202) );
  OAI22_X1 U18370 ( .A1(n19100), .A2(n18818), .B1(n16166), .B2(n15200), .ZN(
        n15201) );
  AOI211_X1 U18371 ( .C1(n19094), .C2(n18824), .A(n15202), .B(n15201), .ZN(
        n15203) );
  OAI21_X1 U18372 ( .B1(n15450), .B2(n16168), .A(n15203), .ZN(P2_U3001) );
  XNOR2_X1 U18373 ( .A(n15204), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15205) );
  XNOR2_X1 U18374 ( .A(n15206), .B(n15205), .ZN(n16214) );
  NAND2_X1 U18375 ( .A1(n16178), .A2(n16180), .ZN(n15208) );
  XNOR2_X1 U18376 ( .A(n15207), .B(n15208), .ZN(n16211) );
  INV_X1 U18377 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15209) );
  OAI22_X1 U18378 ( .A1(n19100), .A2(n15209), .B1(n16166), .B2(n18869), .ZN(
        n15212) );
  OAI22_X1 U18379 ( .A1(n19102), .A2(n18874), .B1(n13051), .B2(n15210), .ZN(
        n15211) );
  AOI211_X1 U18380 ( .C1(n16211), .C2(n19095), .A(n15212), .B(n15211), .ZN(
        n15213) );
  OAI21_X1 U18381 ( .B1(n16169), .B2(n16214), .A(n15213), .ZN(P2_U3007) );
  XNOR2_X1 U18382 ( .A(n15214), .B(n16198), .ZN(n15520) );
  INV_X1 U18383 ( .A(n15520), .ZN(n15223) );
  XNOR2_X1 U18384 ( .A(n15216), .B(n15215), .ZN(n15533) );
  NOR2_X1 U18385 ( .A1(n15533), .A2(n16168), .ZN(n15221) );
  NOR2_X1 U18386 ( .A1(n18885), .A2(n19102), .ZN(n15220) );
  OAI22_X1 U18387 ( .A1(n19100), .A2(n15217), .B1(n15526), .B2(n18871), .ZN(
        n15219) );
  AND2_X1 U18388 ( .A1(n19089), .A2(n18884), .ZN(n15218) );
  NOR4_X1 U18389 ( .A1(n15221), .A2(n15220), .A3(n15219), .A4(n15218), .ZN(
        n15222) );
  OAI21_X1 U18390 ( .B1(n15223), .B2(n16169), .A(n15222), .ZN(P2_U3008) );
  AOI22_X1 U18391 ( .A1(n15224), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n12079), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15226) );
  NAND2_X1 U18392 ( .A1(n12119), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n15225) );
  NAND2_X1 U18393 ( .A1(n15226), .A2(n15225), .ZN(n15227) );
  XNOR2_X1 U18394 ( .A(n15228), .B(n15227), .ZN(n18990) );
  NAND2_X1 U18395 ( .A1(n18990), .A2(n16217), .ZN(n15237) );
  OAI21_X1 U18396 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16216), .A(
        n15229), .ZN(n15230) );
  NAND2_X1 U18397 ( .A1(n15230), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15236) );
  NOR4_X1 U18398 ( .A1(n15233), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15232), .A4(n15231), .ZN(n15235) );
  OAI21_X1 U18399 ( .B1(n15239), .B2(n16222), .A(n9632), .ZN(P2_U3015) );
  OAI211_X1 U18400 ( .C1(n16204), .C2(n16044), .A(n15241), .B(n15240), .ZN(
        n15242) );
  AOI21_X1 U18401 ( .B1(n15243), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15242), .ZN(n15244) );
  OAI21_X1 U18402 ( .B1(n16053), .B2(n15521), .A(n15244), .ZN(n15245) );
  AOI21_X1 U18403 ( .B1(n15246), .B2(n16192), .A(n15245), .ZN(n15247) );
  OAI21_X1 U18404 ( .B1(n15248), .B2(n16222), .A(n15247), .ZN(P2_U3018) );
  AOI211_X1 U18405 ( .C1(n16217), .C2(n15251), .A(n15250), .B(n15249), .ZN(
        n15254) );
  NAND2_X1 U18406 ( .A1(n15252), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15253) );
  OAI211_X1 U18407 ( .C1(n15255), .C2(n15521), .A(n15254), .B(n15253), .ZN(
        n15256) );
  AOI21_X1 U18408 ( .B1(n15257), .B2(n16192), .A(n15256), .ZN(n15258) );
  OAI21_X1 U18409 ( .B1(n15259), .B2(n16222), .A(n15258), .ZN(P2_U3019) );
  INV_X1 U18410 ( .A(n16055), .ZN(n15262) );
  OR2_X1 U18411 ( .A1(n15283), .A2(n20927), .ZN(n15264) );
  NOR3_X1 U18412 ( .A1(n15264), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15276), .ZN(n15260) );
  AOI211_X1 U18413 ( .C1(n16217), .C2(n15262), .A(n15261), .B(n15260), .ZN(
        n15266) );
  INV_X1 U18414 ( .A(n15263), .ZN(n16190) );
  AOI21_X1 U18415 ( .B1(n15287), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16190), .ZN(n15271) );
  NOR2_X1 U18416 ( .A1(n15264), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15273) );
  OAI21_X1 U18417 ( .B1(n15271), .B2(n15273), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15265) );
  OAI211_X1 U18418 ( .C1(n16056), .C2(n15521), .A(n15266), .B(n15265), .ZN(
        n15267) );
  AOI21_X1 U18419 ( .B1(n15268), .B2(n16192), .A(n15267), .ZN(n15269) );
  OAI21_X1 U18420 ( .B1(n15270), .B2(n16222), .A(n15269), .ZN(P2_U3020) );
  INV_X1 U18421 ( .A(n15271), .ZN(n15277) );
  INV_X1 U18422 ( .A(n15272), .ZN(n15274) );
  AOI211_X1 U18423 ( .C1(n16217), .C2(n16066), .A(n15274), .B(n15273), .ZN(
        n15275) );
  OAI21_X1 U18424 ( .B1(n15277), .B2(n15276), .A(n15275), .ZN(n15280) );
  NOR2_X1 U18425 ( .A1(n15278), .A2(n16227), .ZN(n15279) );
  AOI211_X1 U18426 ( .C1(n16067), .C2(n16218), .A(n15280), .B(n15279), .ZN(
        n15281) );
  OAI21_X1 U18427 ( .B1(n15282), .B2(n16222), .A(n15281), .ZN(P2_U3021) );
  NOR2_X1 U18428 ( .A1(n15283), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15284) );
  AOI211_X1 U18429 ( .C1(n16217), .C2(n16080), .A(n15285), .B(n15284), .ZN(
        n15286) );
  OAI21_X1 U18430 ( .B1(n15287), .B2(n20927), .A(n15286), .ZN(n15290) );
  NOR2_X1 U18431 ( .A1(n15288), .A2(n16227), .ZN(n15289) );
  AOI211_X1 U18432 ( .C1(n15291), .C2(n16218), .A(n15290), .B(n15289), .ZN(
        n15292) );
  OAI21_X1 U18433 ( .B1(n15293), .B2(n16222), .A(n15292), .ZN(P2_U3022) );
  INV_X1 U18434 ( .A(n15294), .ZN(n16092) );
  NAND2_X1 U18435 ( .A1(n16217), .A2(n16091), .ZN(n15297) );
  INV_X1 U18436 ( .A(n15331), .ZN(n15295) );
  OAI21_X1 U18437 ( .B1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n15295), .A(
        n15327), .ZN(n15318) );
  NAND2_X1 U18438 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n15318), .ZN(
        n15296) );
  OAI211_X1 U18439 ( .C1(n19802), .C2(n18871), .A(n15297), .B(n15296), .ZN(
        n15300) );
  NAND2_X1 U18440 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15331), .ZN(
        n15322) );
  AOI221_X1 U18441 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C1(n15298), .C2(n15321), .A(
        n15322), .ZN(n15299) );
  AOI211_X1 U18442 ( .C1(n16092), .C2(n16218), .A(n15300), .B(n15299), .ZN(
        n15303) );
  INV_X1 U18443 ( .A(n16222), .ZN(n16210) );
  NAND3_X1 U18444 ( .A1(n15301), .A2(n15098), .A3(n16210), .ZN(n15302) );
  OAI211_X1 U18445 ( .C1(n15304), .C2(n16227), .A(n15303), .B(n15302), .ZN(
        P2_U3023) );
  NAND2_X1 U18446 ( .A1(n15305), .A2(n15321), .ZN(n15306) );
  NAND2_X1 U18447 ( .A1(n15307), .A2(n15306), .ZN(n16132) );
  NAND2_X1 U18448 ( .A1(n15310), .A2(n15309), .ZN(n15311) );
  XNOR2_X1 U18449 ( .A(n15308), .B(n15311), .ZN(n16128) );
  NAND2_X1 U18450 ( .A1(n16128), .A2(n16210), .ZN(n15326) );
  AND2_X1 U18451 ( .A1(n15313), .A2(n15312), .ZN(n15314) );
  NOR2_X1 U18452 ( .A1(n15315), .A2(n15314), .ZN(n16129) );
  OAI21_X1 U18453 ( .B1(n15317), .B2(n15316), .A(n14986), .ZN(n15697) );
  NOR2_X1 U18454 ( .A1(n16204), .A2(n15697), .ZN(n15324) );
  INV_X1 U18455 ( .A(n15318), .ZN(n15320) );
  NAND2_X1 U18456 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19090), .ZN(n15319) );
  OAI221_X1 U18457 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15322), 
        .C1(n15321), .C2(n15320), .A(n15319), .ZN(n15323) );
  AOI211_X1 U18458 ( .C1(n16129), .C2(n16218), .A(n15324), .B(n15323), .ZN(
        n15325) );
  OAI211_X1 U18459 ( .C1(n16132), .C2(n16227), .A(n15326), .B(n15325), .ZN(
        P2_U3024) );
  NOR2_X1 U18460 ( .A1(n15327), .A2(n15330), .ZN(n15328) );
  AOI211_X1 U18461 ( .C1(n15331), .C2(n15330), .A(n15329), .B(n15328), .ZN(
        n15332) );
  OAI21_X1 U18462 ( .B1(n15521), .B2(n15333), .A(n15332), .ZN(n15336) );
  NOR2_X1 U18463 ( .A1(n15334), .A2(n16227), .ZN(n15335) );
  AOI211_X1 U18464 ( .C1(n16217), .C2(n15337), .A(n15336), .B(n15335), .ZN(
        n15338) );
  OAI21_X1 U18465 ( .B1(n15339), .B2(n16222), .A(n15338), .ZN(P2_U3025) );
  AOI21_X1 U18466 ( .B1(n15341), .B2(n15355), .A(n15340), .ZN(n18763) );
  XNOR2_X1 U18467 ( .A(n15342), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15344) );
  AOI21_X1 U18468 ( .B1(n15358), .B2(n15344), .A(n15343), .ZN(n15346) );
  NAND2_X1 U18469 ( .A1(n15372), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15345) );
  OAI211_X1 U18470 ( .C1(n16109), .C2(n15521), .A(n15346), .B(n15345), .ZN(
        n15349) );
  NOR2_X1 U18471 ( .A1(n15347), .A2(n16227), .ZN(n15348) );
  AOI211_X1 U18472 ( .C1(n16217), .C2(n18763), .A(n15349), .B(n15348), .ZN(
        n15350) );
  OAI21_X1 U18473 ( .B1(n15351), .B2(n16222), .A(n15350), .ZN(P2_U3026) );
  NAND2_X1 U18474 ( .A1(n15352), .A2(n15353), .ZN(n15354) );
  NAND2_X1 U18475 ( .A1(n15355), .A2(n15354), .ZN(n20788) );
  AOI21_X1 U18476 ( .B1(n15358), .B2(n15357), .A(n15356), .ZN(n15359) );
  OAI21_X1 U18477 ( .B1(n18775), .B2(n15521), .A(n15359), .ZN(n15360) );
  AOI21_X1 U18478 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15372), .A(
        n15360), .ZN(n15361) );
  OAI21_X1 U18479 ( .B1(n20788), .B2(n16204), .A(n15361), .ZN(n15362) );
  AOI21_X1 U18480 ( .B1(n15363), .B2(n16192), .A(n15362), .ZN(n15364) );
  OAI21_X1 U18481 ( .B1(n15365), .B2(n16222), .A(n15364), .ZN(P2_U3027) );
  OR2_X1 U18482 ( .A1(n13697), .A2(n15366), .ZN(n15367) );
  NAND2_X1 U18483 ( .A1(n15352), .A2(n15367), .ZN(n16123) );
  INV_X1 U18484 ( .A(n18792), .ZN(n15371) );
  NOR4_X1 U18485 ( .A1(n15384), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15368), .A4(n15385), .ZN(n15369) );
  AOI211_X1 U18486 ( .C1(n15371), .C2(n16218), .A(n15370), .B(n15369), .ZN(
        n15374) );
  NAND2_X1 U18487 ( .A1(n15372), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15373) );
  OAI211_X1 U18488 ( .C1(n16123), .C2(n16204), .A(n15374), .B(n15373), .ZN(
        n15375) );
  AOI21_X1 U18489 ( .B1(n15376), .B2(n16192), .A(n15375), .ZN(n15377) );
  OAI21_X1 U18490 ( .B1(n15378), .B2(n16222), .A(n15377), .ZN(P2_U3028) );
  INV_X1 U18491 ( .A(n15379), .ZN(n15383) );
  AOI21_X1 U18492 ( .B1(n16227), .B2(n15381), .A(n15380), .ZN(n15382) );
  OAI21_X1 U18493 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n16216), .A(
        n15402), .ZN(n15391) );
  INV_X1 U18494 ( .A(n15384), .ZN(n15405) );
  AOI21_X1 U18495 ( .B1(n15421), .B2(n16192), .A(n15405), .ZN(n15395) );
  NOR3_X1 U18496 ( .A1(n15395), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15385), .ZN(n15390) );
  AOI21_X1 U18497 ( .B1(n15387), .B2(n16218), .A(n15386), .ZN(n15388) );
  OAI21_X1 U18498 ( .B1(n18801), .B2(n16204), .A(n15388), .ZN(n15389) );
  OAI21_X1 U18499 ( .B1(n15393), .B2(n16222), .A(n15392), .ZN(P2_U3029) );
  OAI21_X1 U18500 ( .B1(n18957), .B2(n15521), .A(n15394), .ZN(n15397) );
  NOR3_X1 U18501 ( .A1(n15395), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15404), .ZN(n15396) );
  AOI211_X1 U18502 ( .C1(n16217), .C2(n15398), .A(n15397), .B(n15396), .ZN(
        n15401) );
  NAND2_X1 U18503 ( .A1(n15399), .A2(n16210), .ZN(n15400) );
  OAI211_X1 U18504 ( .C1(n15402), .C2(n15174), .A(n15401), .B(n15400), .ZN(
        P2_U3030) );
  NOR2_X1 U18505 ( .A1(n15188), .A2(n18871), .ZN(n15403) );
  AOI21_X1 U18506 ( .B1(n15405), .B2(n15404), .A(n15403), .ZN(n15406) );
  OAI21_X1 U18507 ( .B1(n15407), .B2(n15521), .A(n15406), .ZN(n15408) );
  AOI21_X1 U18508 ( .B1(n15409), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15408), .ZN(n15410) );
  OAI21_X1 U18509 ( .B1(n15411), .B2(n16204), .A(n15410), .ZN(n15412) );
  AOI21_X1 U18510 ( .B1(n15413), .B2(n16192), .A(n15412), .ZN(n15414) );
  OAI21_X1 U18511 ( .B1(n15415), .B2(n16222), .A(n15414), .ZN(P2_U3031) );
  NAND2_X1 U18512 ( .A1(n15417), .A2(n15416), .ZN(n15418) );
  XNOR2_X1 U18513 ( .A(n15419), .B(n15418), .ZN(n16138) );
  INV_X1 U18514 ( .A(n16138), .ZN(n15440) );
  INV_X1 U18515 ( .A(n15420), .ZN(n15423) );
  AOI21_X1 U18516 ( .B1(n15423), .B2(n15422), .A(n15421), .ZN(n16139) );
  AND2_X1 U18517 ( .A1(n15425), .A2(n15424), .ZN(n15427) );
  OR2_X1 U18518 ( .A1(n15427), .A2(n15426), .ZN(n18962) );
  AOI21_X1 U18519 ( .B1(n15429), .B2(n15428), .A(n13611), .ZN(n18813) );
  INV_X1 U18520 ( .A(n15433), .ZN(n15432) );
  NAND2_X1 U18521 ( .A1(n15430), .A2(n15507), .ZN(n15442) );
  OAI21_X1 U18522 ( .B1(n15430), .B2(n16216), .A(n15514), .ZN(n15457) );
  INV_X1 U18523 ( .A(n15457), .ZN(n15431) );
  OAI21_X1 U18524 ( .B1(n15432), .B2(n15442), .A(n15431), .ZN(n15441) );
  NOR3_X1 U18525 ( .A1(n15433), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n15442), .ZN(n15434) );
  AOI21_X1 U18526 ( .B1(n15441), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15434), .ZN(n15435) );
  OAI21_X1 U18527 ( .B1(n13051), .B2(n11980), .A(n15435), .ZN(n15436) );
  AOI21_X1 U18528 ( .B1(n16217), .B2(n18813), .A(n15436), .ZN(n15437) );
  OAI21_X1 U18529 ( .B1(n15521), .B2(n18962), .A(n15437), .ZN(n15438) );
  AOI21_X1 U18530 ( .B1(n16139), .B2(n16192), .A(n15438), .ZN(n15439) );
  OAI21_X1 U18531 ( .B1(n16222), .B2(n15440), .A(n15439), .ZN(P2_U3032) );
  INV_X1 U18532 ( .A(n15441), .ZN(n15445) );
  INV_X1 U18533 ( .A(n15442), .ZN(n15458) );
  AOI21_X1 U18534 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15458), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15444) );
  OAI21_X1 U18535 ( .B1(n15445), .B2(n15444), .A(n15443), .ZN(n15448) );
  OAI22_X1 U18536 ( .A1(n16204), .A2(n18825), .B1(n16227), .B2(n15446), .ZN(
        n15447) );
  AOI211_X1 U18537 ( .C1(n16218), .C2(n18824), .A(n15448), .B(n15447), .ZN(
        n15449) );
  OAI21_X1 U18538 ( .B1(n15450), .B2(n16222), .A(n15449), .ZN(P2_U3033) );
  INV_X1 U18539 ( .A(n15452), .ZN(n15453) );
  OR2_X1 U18540 ( .A1(n15454), .A2(n15453), .ZN(n15455) );
  XNOR2_X1 U18541 ( .A(n9599), .B(n15455), .ZN(n16142) );
  NOR2_X1 U18542 ( .A1(n14817), .A2(n18871), .ZN(n15456) );
  AOI221_X1 U18543 ( .B1(n15458), .B2(n11772), .C1(n15457), .C2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n15456), .ZN(n15460) );
  NAND2_X1 U18544 ( .A1(n16218), .A2(n16143), .ZN(n15459) );
  OAI211_X1 U18545 ( .C1(n18997), .C2(n16204), .A(n15460), .B(n15459), .ZN(
        n15465) );
  OR2_X1 U18546 ( .A1(n15461), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15463) );
  NAND2_X1 U18547 ( .A1(n15463), .A2(n15462), .ZN(n16146) );
  NOR2_X1 U18548 ( .A1(n16146), .A2(n16227), .ZN(n15464) );
  AOI211_X1 U18549 ( .C1(n16210), .C2(n16142), .A(n15465), .B(n15464), .ZN(
        n15466) );
  INV_X1 U18550 ( .A(n15466), .ZN(P2_U3034) );
  INV_X1 U18551 ( .A(n15467), .ZN(n15468) );
  NAND2_X1 U18552 ( .A1(n15469), .A2(n15468), .ZN(n15473) );
  NOR2_X1 U18553 ( .A1(n15471), .A2(n15470), .ZN(n15472) );
  XNOR2_X1 U18554 ( .A(n15473), .B(n15472), .ZN(n16151) );
  OAI21_X1 U18555 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15496), .A(
        n15474), .ZN(n16152) );
  INV_X1 U18556 ( .A(n16152), .ZN(n15481) );
  OAI21_X1 U18557 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16216), .A(
        n15514), .ZN(n15489) );
  NOR2_X1 U18558 ( .A1(n11973), .A2(n13051), .ZN(n15477) );
  INV_X1 U18559 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15475) );
  NAND2_X1 U18560 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15507), .ZN(
        n15491) );
  AOI221_X1 U18561 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n15475), .C2(n11755), .A(
        n15491), .ZN(n15476) );
  AOI211_X1 U18562 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15489), .A(
        n15477), .B(n15476), .ZN(n15479) );
  NAND2_X1 U18563 ( .A1(n16218), .A2(n18838), .ZN(n15478) );
  OAI211_X1 U18564 ( .C1(n18834), .C2(n16204), .A(n15479), .B(n15478), .ZN(
        n15480) );
  AOI21_X1 U18565 ( .B1(n15481), .B2(n16192), .A(n15480), .ZN(n15482) );
  OAI21_X1 U18566 ( .B1(n16151), .B2(n16222), .A(n15482), .ZN(P2_U3035) );
  INV_X1 U18567 ( .A(n15483), .ZN(n15501) );
  OR2_X1 U18568 ( .A1(n15484), .A2(n15501), .ZN(n15488) );
  NAND2_X1 U18569 ( .A1(n15486), .A2(n15485), .ZN(n15487) );
  XNOR2_X1 U18570 ( .A(n15488), .B(n15487), .ZN(n16157) );
  NOR2_X1 U18571 ( .A1(n11970), .A2(n18871), .ZN(n15493) );
  NAND2_X1 U18572 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15489), .ZN(
        n15490) );
  OAI21_X1 U18573 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n15491), .A(
        n15490), .ZN(n15492) );
  OR2_X1 U18574 ( .A1(n15493), .A2(n15492), .ZN(n15494) );
  AOI21_X1 U18575 ( .B1(n16218), .B2(n16158), .A(n15494), .ZN(n15495) );
  OAI21_X1 U18576 ( .B1(n19000), .B2(n16204), .A(n15495), .ZN(n15499) );
  AND2_X1 U18577 ( .A1(n15515), .A2(n11755), .ZN(n15497) );
  OR2_X1 U18578 ( .A1(n15497), .A2(n15496), .ZN(n16161) );
  NOR2_X1 U18579 ( .A1(n16161), .A2(n16227), .ZN(n15498) );
  AOI211_X1 U18580 ( .C1(n16210), .C2(n16157), .A(n15499), .B(n15498), .ZN(
        n15500) );
  INV_X1 U18581 ( .A(n15500), .ZN(P2_U3036) );
  OR2_X1 U18582 ( .A1(n15502), .A2(n15501), .ZN(n15503) );
  XNOR2_X1 U18583 ( .A(n15504), .B(n15503), .ZN(n16167) );
  OAI21_X1 U18584 ( .B1(n15506), .B2(n15505), .A(n14823), .ZN(n19003) );
  INV_X1 U18585 ( .A(n19003), .ZN(n15518) );
  INV_X1 U18586 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15513) );
  NOR2_X1 U18587 ( .A1(n11967), .A2(n13051), .ZN(n15510) );
  INV_X1 U18588 ( .A(n15507), .ZN(n15508) );
  NOR2_X1 U18589 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15508), .ZN(
        n15509) );
  NOR2_X1 U18590 ( .A1(n15510), .A2(n15509), .ZN(n15512) );
  INV_X1 U18591 ( .A(n18852), .ZN(n16172) );
  NAND2_X1 U18592 ( .A1(n16218), .A2(n16172), .ZN(n15511) );
  OAI211_X1 U18593 ( .C1(n15514), .C2(n15513), .A(n15512), .B(n15511), .ZN(
        n15517) );
  OAI21_X1 U18594 ( .B1(n15196), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15515), .ZN(n16170) );
  NOR2_X1 U18595 ( .A1(n16170), .A2(n16227), .ZN(n15516) );
  AOI211_X1 U18596 ( .C1(n16217), .C2(n15518), .A(n15517), .B(n15516), .ZN(
        n15519) );
  OAI21_X1 U18597 ( .B1(n16222), .B2(n16167), .A(n15519), .ZN(P2_U3037) );
  NAND2_X1 U18598 ( .A1(n15520), .A2(n16192), .ZN(n15532) );
  NOR2_X1 U18599 ( .A1(n18885), .A2(n15521), .ZN(n15529) );
  AOI211_X1 U18600 ( .C1(n15523), .C2(n16197), .A(n15522), .B(n16198), .ZN(
        n16191) );
  AOI21_X1 U18601 ( .B1(n15525), .B2(n15524), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15527) );
  OAI22_X1 U18602 ( .A1(n16191), .A2(n15527), .B1(n13051), .B2(n15526), .ZN(
        n15528) );
  AOI211_X1 U18603 ( .C1(n15530), .C2(n16217), .A(n15529), .B(n15528), .ZN(
        n15531) );
  OAI211_X1 U18604 ( .C1(n16222), .C2(n15533), .A(n15532), .B(n15531), .ZN(
        P2_U3040) );
  INV_X1 U18605 ( .A(n15540), .ZN(n18947) );
  AOI22_X1 U18606 ( .A1(n18896), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18947), .B2(n18915), .ZN(n15542) );
  AOI222_X1 U18607 ( .A1(n15535), .A2(n19833), .B1(n15534), .B2(n10024), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n15542), .ZN(n15537) );
  NAND2_X1 U18608 ( .A1(n15552), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15536) );
  OAI21_X1 U18609 ( .B1(n15537), .B2(n15552), .A(n15536), .ZN(P2_U3601) );
  OAI211_X1 U18610 ( .C1(n15540), .C2(n15539), .A(n18915), .B(n15538), .ZN(
        n18933) );
  OAI21_X1 U18611 ( .B1(n14711), .B2(n15541), .A(n18933), .ZN(n15548) );
  INV_X1 U18612 ( .A(n15548), .ZN(n15543) );
  NOR2_X1 U18613 ( .A1(n15542), .A2(n19757), .ZN(n15547) );
  AOI222_X1 U18614 ( .A1(n15544), .A2(n19833), .B1(n15543), .B2(n15547), .C1(
        n19851), .C2(n10024), .ZN(n15546) );
  NAND2_X1 U18615 ( .A1(n15552), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15545) );
  OAI21_X1 U18616 ( .B1(n15546), .B2(n15552), .A(n15545), .ZN(P2_U3600) );
  AOI222_X1 U18617 ( .A1(n15549), .A2(n19833), .B1(n10024), .B2(n19281), .C1(
        n15548), .C2(n15547), .ZN(n15553) );
  NAND2_X1 U18618 ( .A1(n15552), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15551) );
  OAI21_X1 U18619 ( .B1(n15553), .B2(n15552), .A(n15551), .ZN(P2_U3599) );
  INV_X1 U18620 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16795) );
  INV_X1 U18621 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16518) );
  INV_X1 U18622 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16552) );
  INV_X1 U18623 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16574) );
  INV_X1 U18624 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n15560) );
  INV_X1 U18625 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16638) );
  INV_X1 U18626 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n16730) );
  INV_X1 U18627 ( .A(n9580), .ZN(n15555) );
  NAND3_X1 U18628 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17086) );
  NAND4_X1 U18629 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(P3_EBX_REG_7__SCAN_IN), .ZN(n15559) );
  NAND3_X1 U18630 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .ZN(n16923) );
  NOR4_X2 U18631 ( .A1(n16574), .A2(n15560), .A3(n17005), .A4(n16923), .ZN(
        n16910) );
  NAND2_X1 U18632 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16910), .ZN(n16897) );
  NAND3_X1 U18633 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n16849), .ZN(n16833) );
  NOR2_X2 U18634 ( .A1(n16833), .A2(n16795), .ZN(n16838) );
  NAND2_X1 U18635 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16838), .ZN(n16832) );
  INV_X1 U18636 ( .A(n16832), .ZN(n15640) );
  AOI21_X1 U18637 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17097), .A(n16838), .ZN(
        n15639) );
  AOI22_X1 U18638 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9579), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15564) );
  AOI22_X1 U18639 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15563) );
  AOI22_X1 U18640 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15612), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15562) );
  AOI22_X1 U18641 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15561) );
  NAND4_X1 U18642 ( .A1(n15564), .A2(n15563), .A3(n15562), .A4(n15561), .ZN(
        n15570) );
  AOI22_X1 U18643 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15568) );
  AOI22_X1 U18644 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15627), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15567) );
  AOI22_X1 U18645 ( .A1(n16813), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15615), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15566) );
  AOI22_X1 U18646 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15565) );
  NAND4_X1 U18647 ( .A1(n15568), .A2(n15567), .A3(n15566), .A4(n15565), .ZN(
        n15569) );
  NOR2_X1 U18648 ( .A1(n15570), .A2(n15569), .ZN(n15637) );
  AOI22_X1 U18649 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15612), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15574) );
  AOI22_X1 U18650 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15573) );
  AOI22_X1 U18651 ( .A1(n16813), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15572) );
  AOI22_X1 U18652 ( .A1(n16806), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15571) );
  NAND4_X1 U18653 ( .A1(n15574), .A2(n15573), .A3(n15572), .A4(n15571), .ZN(
        n15580) );
  AOI22_X1 U18654 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15615), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15578) );
  AOI22_X1 U18655 ( .A1(n17065), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15627), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15577) );
  AOI22_X1 U18656 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15576) );
  AOI22_X1 U18657 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9579), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15575) );
  NAND4_X1 U18658 ( .A1(n15578), .A2(n15577), .A3(n15576), .A4(n15575), .ZN(
        n15579) );
  NOR2_X1 U18659 ( .A1(n15580), .A2(n15579), .ZN(n16839) );
  AOI22_X1 U18660 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15612), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15584) );
  AOI22_X1 U18661 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15583) );
  AOI22_X1 U18662 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15582) );
  AOI22_X1 U18663 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15581) );
  NAND4_X1 U18664 ( .A1(n15584), .A2(n15583), .A3(n15582), .A4(n15581), .ZN(
        n15590) );
  AOI22_X1 U18665 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n16806), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15588) );
  AOI22_X1 U18666 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15587) );
  AOI22_X1 U18667 ( .A1(n9579), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15627), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15586) );
  AOI22_X1 U18668 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15615), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15585) );
  NAND4_X1 U18669 ( .A1(n15588), .A2(n15587), .A3(n15586), .A4(n15585), .ZN(
        n15589) );
  NOR2_X1 U18670 ( .A1(n15590), .A2(n15589), .ZN(n16847) );
  AOI22_X1 U18671 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16806), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15601) );
  AOI22_X1 U18672 ( .A1(n16813), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15600) );
  INV_X1 U18673 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18406) );
  AOI22_X1 U18674 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15626), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15591) );
  OAI21_X1 U18675 ( .B1(n15592), .B2(n18406), .A(n15591), .ZN(n15598) );
  AOI22_X1 U18676 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15627), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15596) );
  AOI22_X1 U18677 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15615), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15595) );
  AOI22_X1 U18678 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15612), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15594) );
  AOI22_X1 U18679 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15593) );
  NAND4_X1 U18680 ( .A1(n15596), .A2(n15595), .A3(n15594), .A4(n15593), .ZN(
        n15597) );
  AOI211_X1 U18681 ( .C1(n17035), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n15598), .B(n15597), .ZN(n15599) );
  NAND3_X1 U18682 ( .A1(n15601), .A2(n15600), .A3(n15599), .ZN(n16852) );
  AOI22_X1 U18683 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17055), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15611) );
  AOI22_X1 U18684 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17051), .B1(
        n15626), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15610) );
  INV_X1 U18685 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16951) );
  AOI22_X1 U18686 ( .A1(n17065), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n9608), .ZN(n15602) );
  OAI21_X1 U18687 ( .B1(n12438), .B2(n16951), .A(n15602), .ZN(n15608) );
  AOI22_X1 U18688 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15606) );
  AOI22_X1 U18689 ( .A1(n16813), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n16998), .ZN(n15605) );
  AOI22_X1 U18690 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15615), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15604) );
  AOI22_X1 U18691 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17060), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17036), .ZN(n15603) );
  NAND4_X1 U18692 ( .A1(n15606), .A2(n15605), .A3(n15604), .A4(n15603), .ZN(
        n15607) );
  AOI211_X1 U18693 ( .C1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .C2(n17052), .A(
        n15608), .B(n15607), .ZN(n15609) );
  NAND3_X1 U18694 ( .A1(n15611), .A2(n15610), .A3(n15609), .ZN(n16853) );
  NAND2_X1 U18695 ( .A1(n16852), .A2(n16853), .ZN(n16851) );
  NOR2_X1 U18696 ( .A1(n16847), .A2(n16851), .ZN(n16844) );
  AOI22_X1 U18697 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15626), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15624) );
  AOI22_X1 U18698 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15612), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15623) );
  AOI22_X1 U18699 ( .A1(n17052), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15613) );
  OAI21_X1 U18700 ( .B1(n15614), .B2(n17095), .A(n15613), .ZN(n15621) );
  AOI22_X1 U18701 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15619) );
  AOI22_X1 U18702 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15615), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15618) );
  AOI22_X1 U18703 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15617) );
  AOI22_X1 U18704 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15616) );
  NAND4_X1 U18705 ( .A1(n15619), .A2(n15618), .A3(n15617), .A4(n15616), .ZN(
        n15620) );
  AOI211_X1 U18706 ( .C1(n9579), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n15621), .B(n15620), .ZN(n15622) );
  NAND3_X1 U18707 ( .A1(n15624), .A2(n15623), .A3(n15622), .ZN(n16843) );
  NAND2_X1 U18708 ( .A1(n16844), .A2(n16843), .ZN(n16842) );
  NOR2_X1 U18709 ( .A1(n16839), .A2(n16842), .ZN(n16836) );
  AOI22_X1 U18710 ( .A1(n17034), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15636) );
  AOI22_X1 U18711 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15635) );
  AOI22_X1 U18712 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9579), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15625) );
  OAI21_X1 U18713 ( .B1(n12588), .B2(n20839), .A(n15625), .ZN(n15633) );
  AOI22_X1 U18714 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15626), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15631) );
  AOI22_X1 U18715 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15630) );
  AOI22_X1 U18716 ( .A1(n16965), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15627), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15629) );
  AOI22_X1 U18717 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15628) );
  NAND4_X1 U18718 ( .A1(n15631), .A2(n15630), .A3(n15629), .A4(n15628), .ZN(
        n15632) );
  AOI211_X1 U18719 ( .C1(n17035), .C2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n15633), .B(n15632), .ZN(n15634) );
  NAND3_X1 U18720 ( .A1(n15636), .A2(n15635), .A3(n15634), .ZN(n16835) );
  NAND2_X1 U18721 ( .A1(n16836), .A2(n16835), .ZN(n16834) );
  NOR2_X1 U18722 ( .A1(n15637), .A2(n16834), .ZN(n16830) );
  AOI21_X1 U18723 ( .B1(n15637), .B2(n16834), .A(n16830), .ZN(n17121) );
  INV_X1 U18724 ( .A(n17121), .ZN(n15638) );
  OAI22_X1 U18725 ( .A1(n15640), .A2(n15639), .B1(n17085), .B2(n15638), .ZN(
        P3_U2675) );
  NOR2_X1 U18726 ( .A1(n18667), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18098) );
  NAND3_X1 U18727 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18665)
         );
  INV_X1 U18728 ( .A(n18665), .ZN(n15642) );
  OAI211_X1 U18729 ( .C1(n18672), .C2(n18522), .A(n15641), .B(n18504), .ZN(
        n18053) );
  INV_X1 U18730 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18054) );
  NOR2_X1 U18731 ( .A1(n18054), .A2(n18665), .ZN(n15660) );
  AOI211_X1 U18732 ( .C1(n15642), .C2(n18053), .A(n18300), .B(n15660), .ZN(
        n15643) );
  NOR2_X1 U18733 ( .A1(n18098), .A2(n15643), .ZN(n15645) );
  INV_X1 U18734 ( .A(n18398), .ZN(n18297) );
  INV_X1 U18735 ( .A(n15643), .ZN(n18059) );
  INV_X1 U18736 ( .A(n17632), .ZN(n17687) );
  NAND2_X1 U18737 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18063) );
  OAI21_X1 U18738 ( .B1(n18710), .B2(n17687), .A(n18063), .ZN(n15648) );
  NAND3_X1 U18739 ( .A1(n18534), .A2(n18059), .A3(n15648), .ZN(n15644) );
  OAI221_X1 U18740 ( .B1(n18534), .B2(n15645), .C1(n18534), .C2(n18297), .A(
        n15644), .ZN(P3_U2864) );
  NAND2_X1 U18741 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18227) );
  NOR2_X1 U18742 ( .A1(n18710), .A2(n17687), .ZN(n15647) );
  INV_X1 U18743 ( .A(n15645), .ZN(n15646) );
  AOI221_X1 U18744 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18227), .C1(n15647), 
        .C2(n18227), .A(n15646), .ZN(n18058) );
  OAI221_X1 U18745 ( .B1(n18398), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18398), .C2(n15648), .A(n18059), .ZN(n18056) );
  AOI22_X1 U18746 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18058), .B1(
        n18056), .B2(n20885), .ZN(P3_U2865) );
  NAND2_X1 U18747 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18717) );
  NOR2_X1 U18748 ( .A1(n18578), .A2(n15672), .ZN(n15658) );
  INV_X1 U18749 ( .A(n15649), .ZN(n17307) );
  NAND2_X1 U18750 ( .A1(n18716), .A2(n17307), .ZN(n18555) );
  NAND2_X2 U18751 ( .A1(n18658), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18652) );
  OAI21_X1 U18752 ( .B1(n15653), .B2(n15652), .A(n15651), .ZN(n15655) );
  NAND2_X1 U18753 ( .A1(n15655), .A2(n15654), .ZN(n15673) );
  AOI211_X1 U18754 ( .C1(n15658), .C2(n17252), .A(n15656), .B(n15673), .ZN(
        n15659) );
  INV_X1 U18755 ( .A(n18515), .ZN(n18520) );
  NAND2_X1 U18756 ( .A1(n15659), .A2(n15762), .ZN(n18538) );
  NOR2_X1 U18757 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18667), .ZN(n18061) );
  INV_X1 U18758 ( .A(n18697), .ZN(n18695) );
  INV_X1 U18759 ( .A(n18522), .ZN(n18506) );
  AOI21_X1 U18760 ( .B1(n18506), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15662) );
  INV_X1 U18761 ( .A(n18523), .ZN(n15661) );
  NOR2_X1 U18762 ( .A1(n15662), .A2(n15661), .ZN(n18552) );
  NAND3_X1 U18763 ( .A1(n18695), .A2(n18693), .A3(n18552), .ZN(n15663) );
  OAI21_X1 U18764 ( .B1(n18695), .B2(n18504), .A(n15663), .ZN(P3_U3284) );
  AND4_X1 U18765 ( .A1(n15665), .A2(n19119), .A3(n19833), .A4(n15664), .ZN(
        n15666) );
  NAND2_X1 U18766 ( .A1(n15669), .A2(n15666), .ZN(n15667) );
  OAI21_X1 U18767 ( .B1(n15669), .B2(n15668), .A(n15667), .ZN(P2_U3595) );
  INV_X1 U18768 ( .A(n16252), .ZN(n16251) );
  INV_X1 U18769 ( .A(n18499), .ZN(n15678) );
  OAI21_X1 U18770 ( .B1(n18072), .B2(n16410), .A(n18714), .ZN(n15670) );
  OAI21_X1 U18771 ( .B1(n15671), .B2(n15670), .A(n18717), .ZN(n16391) );
  NOR3_X1 U18772 ( .A1(n15675), .A2(n15672), .A3(n16391), .ZN(n15674) );
  AOI211_X1 U18773 ( .C1(n15675), .C2(n9580), .A(n15674), .B(n15673), .ZN(
        n15677) );
  AOI221_X4 U18774 ( .B1(n15678), .B2(n15677), .C1(n15676), .C2(n15677), .A(
        n18561), .ZN(n18026) );
  NOR2_X1 U18775 ( .A1(n17217), .A2(n18041), .ZN(n17897) );
  INV_X1 U18776 ( .A(n17897), .ZN(n17967) );
  INV_X1 U18777 ( .A(n18519), .ZN(n18017) );
  AOI21_X1 U18778 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17998) );
  NAND3_X1 U18779 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17872) );
  NOR2_X1 U18780 ( .A1(n17998), .A2(n17872), .ZN(n17952) );
  NAND4_X1 U18781 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n17952), .ZN(n17858) );
  NOR2_X1 U18782 ( .A1(n16244), .A2(n17858), .ZN(n15684) );
  INV_X1 U18783 ( .A(n15684), .ZN(n17841) );
  NAND2_X1 U18784 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17997) );
  NOR2_X1 U18785 ( .A1(n17997), .A2(n17872), .ZN(n17954) );
  NAND4_X1 U18786 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n17954), .ZN(n17857) );
  NOR2_X1 U18787 ( .A1(n16244), .A2(n17857), .ZN(n15680) );
  INV_X1 U18788 ( .A(n15680), .ZN(n17840) );
  INV_X1 U18789 ( .A(n18529), .ZN(n17928) );
  AOI21_X1 U18790 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n17928), .A(
        n18532), .ZN(n18018) );
  OAI22_X1 U18791 ( .A1(n18017), .A2(n17841), .B1(n17840), .B2(n18018), .ZN(
        n17766) );
  NAND3_X1 U18792 ( .A1(n18026), .A2(n17749), .A3(n17766), .ZN(n16268) );
  NAND2_X1 U18793 ( .A1(n18494), .A2(n18026), .ZN(n18014) );
  INV_X1 U18794 ( .A(n18014), .ZN(n18045) );
  NAND2_X1 U18795 ( .A1(n16250), .A2(n18045), .ZN(n15679) );
  OAI211_X1 U18796 ( .C1(n17967), .C2(n17745), .A(n16268), .B(n15679), .ZN(
        n15751) );
  NAND2_X1 U18797 ( .A1(n16251), .A2(n15751), .ZN(n15694) );
  NOR2_X1 U18798 ( .A1(n17939), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16284) );
  NAND2_X1 U18799 ( .A1(n17749), .A2(n15680), .ZN(n15683) );
  INV_X1 U18800 ( .A(n17474), .ZN(n17497) );
  NOR2_X1 U18801 ( .A1(n18694), .A2(n17857), .ZN(n17925) );
  NAND2_X1 U18802 ( .A1(n17521), .A2(n17925), .ZN(n17861) );
  NOR2_X1 U18803 ( .A1(n17497), .A2(n17861), .ZN(n17817) );
  NAND4_X1 U18804 ( .A1(n15686), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15681), .A4(n17817), .ZN(n15682) );
  AOI22_X1 U18805 ( .A1(n18532), .A2(n15683), .B1(n17928), .B2(n15682), .ZN(
        n15748) );
  INV_X1 U18806 ( .A(n15748), .ZN(n15688) );
  INV_X2 U18807 ( .A(n18048), .ZN(n18038) );
  NOR2_X2 U18808 ( .A1(n18038), .A2(n18026), .ZN(n18027) );
  INV_X1 U18809 ( .A(n17956), .ZN(n17863) );
  NOR2_X1 U18810 ( .A1(n17863), .A2(n18049), .ZN(n18033) );
  NOR2_X1 U18811 ( .A1(n18027), .A2(n18033), .ZN(n17958) );
  AOI21_X1 U18812 ( .B1(n17474), .B2(n15684), .A(n18017), .ZN(n17801) );
  AOI21_X1 U18813 ( .B1(n18519), .B2(n15685), .A(n17801), .ZN(n17787) );
  OAI21_X1 U18814 ( .B1(n15686), .B2(n18017), .A(n17787), .ZN(n17743) );
  NOR2_X1 U18815 ( .A1(n18027), .A2(n17743), .ZN(n15747) );
  NAND2_X1 U18816 ( .A1(n16267), .A2(n16250), .ZN(n16242) );
  INV_X1 U18817 ( .A(n16243), .ZN(n16253) );
  AOI22_X1 U18818 ( .A1(n18045), .A2(n16242), .B1(n17897), .B2(n16253), .ZN(
        n15749) );
  OAI221_X1 U18819 ( .B1(n17958), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), 
        .C1(n17958), .C2(n15747), .A(n15749), .ZN(n15687) );
  AOI221_X1 U18820 ( .B1(n16284), .B2(n18026), .C1(n15688), .C2(n18026), .A(
        n15687), .ZN(n15693) );
  NOR2_X1 U18821 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17639), .ZN(
        n16282) );
  AOI21_X1 U18822 ( .B1(n16287), .B2(n15690), .A(n16282), .ZN(n15691) );
  XNOR2_X1 U18823 ( .A(n15691), .B(n16265), .ZN(n16263) );
  AOI22_X1 U18824 ( .A1(n18038), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n17936), 
        .B2(n16263), .ZN(n15692) );
  OAI221_X1 U18825 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15694), 
        .C1(n16265), .C2(n15693), .A(n15692), .ZN(P3_U2833) );
  AOI22_X1 U18826 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n18935), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18936), .ZN(n15703) );
  INV_X1 U18827 ( .A(n15695), .ZN(n15696) );
  AOI22_X1 U18828 ( .A1(n15696), .A2(n18906), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18950), .ZN(n15702) );
  INV_X1 U18829 ( .A(n15697), .ZN(n16114) );
  AOI22_X1 U18830 ( .A1(n16129), .A2(n18944), .B1(n16114), .B2(n18937), .ZN(
        n15701) );
  OAI211_X1 U18831 ( .C1(n15699), .C2(n16136), .A(n18901), .B(n15698), .ZN(
        n15700) );
  NAND4_X1 U18832 ( .A1(n15703), .A2(n15702), .A3(n15701), .A4(n15700), .ZN(
        P2_U2833) );
  OAI21_X1 U18833 ( .B1(n20687), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20613), 
        .ZN(n16005) );
  INV_X1 U18834 ( .A(n16005), .ZN(n15736) );
  NAND2_X1 U18835 ( .A1(n20768), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16000) );
  INV_X1 U18836 ( .A(n15704), .ZN(n15730) );
  OAI211_X1 U18837 ( .C1(n9875), .C2(n15706), .A(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15705), .ZN(n15710) );
  INV_X1 U18838 ( .A(n15707), .ZN(n15709) );
  OAI211_X1 U18839 ( .C1(n20505), .C2(n15710), .A(n15709), .B(n15708), .ZN(
        n15712) );
  NAND2_X1 U18840 ( .A1(n20505), .A2(n15710), .ZN(n15711) );
  NAND2_X1 U18841 ( .A1(n15712), .A2(n15711), .ZN(n15714) );
  INV_X1 U18842 ( .A(n15714), .ZN(n15716) );
  AOI21_X1 U18843 ( .B1(n15714), .B2(n20425), .A(n15713), .ZN(n15715) );
  AOI21_X1 U18844 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15716), .A(
        n15715), .ZN(n15718) );
  INV_X1 U18845 ( .A(n15718), .ZN(n15721) );
  INV_X1 U18846 ( .A(n15717), .ZN(n15720) );
  OAI21_X1 U18847 ( .B1(n15718), .B2(n15717), .A(n20473), .ZN(n15719) );
  OAI21_X1 U18848 ( .B1(n15721), .B2(n15720), .A(n15719), .ZN(n15728) );
  OAI21_X1 U18849 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15722), .ZN(n15725) );
  NAND4_X1 U18850 ( .A1(n15725), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n15724), 
        .A4(n15723), .ZN(n15726) );
  AOI211_X1 U18851 ( .C1(n15728), .C2(n20088), .A(n15727), .B(n15726), .ZN(
        n15729) );
  NAND2_X1 U18852 ( .A1(n15730), .A2(n15729), .ZN(n15737) );
  NAND3_X1 U18853 ( .A1(n9616), .A2(n15732), .A3(n15731), .ZN(n15733) );
  AOI21_X1 U18854 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATE2_REG_1__SCAN_IN), .A(n20613), .ZN(n20677) );
  OAI211_X1 U18855 ( .C1(n12753), .C2(n15733), .A(n20677), .B(n16000), .ZN(
        n16007) );
  AOI21_X1 U18856 ( .B1(n15737), .B2(n15734), .A(n16007), .ZN(n16004) );
  AOI211_X1 U18857 ( .C1(n15736), .C2(n16000), .A(n15735), .B(n16004), .ZN(
        n15743) );
  OAI21_X1 U18858 ( .B1(n15738), .B2(n10259), .A(n15737), .ZN(n15742) );
  AOI21_X1 U18859 ( .B1(n15739), .B2(n20772), .A(n16004), .ZN(n15740) );
  INV_X1 U18860 ( .A(n15740), .ZN(n15741) );
  AOI22_X1 U18861 ( .A1(n15743), .A2(n15742), .B1(n10259), .B2(n15741), .ZN(
        P1_U3161) );
  AOI21_X1 U18862 ( .B1(n15745), .B2(n17639), .A(n15744), .ZN(n15746) );
  XOR2_X1 U18863 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n15746), .Z(
        n16249) );
  NAND2_X1 U18864 ( .A1(n15748), .A2(n15747), .ZN(n16283) );
  OAI221_X1 U18865 ( .B1(n16283), .B2(n17956), .C1(n16283), .C2(n15750), .A(
        n18048), .ZN(n16270) );
  NAND2_X1 U18866 ( .A1(n15749), .A2(n16270), .ZN(n15752) );
  NOR2_X1 U18867 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15750), .ZN(
        n16245) );
  AOI22_X1 U18868 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15752), .B1(
        n16245), .B2(n15751), .ZN(n15753) );
  NAND2_X1 U18869 ( .A1(n18038), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16238) );
  OAI211_X1 U18870 ( .C1(n16249), .C2(n17960), .A(n15753), .B(n16238), .ZN(
        P3_U2832) );
  INV_X1 U18871 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20693) );
  INV_X1 U18872 ( .A(HOLD), .ZN(n20683) );
  NOR2_X1 U18873 ( .A1(n20693), .A2(n20683), .ZN(n20680) );
  AOI22_X1 U18874 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15755) );
  INV_X1 U18875 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20686) );
  NOR2_X1 U18876 ( .A1(n20686), .A2(n20768), .ZN(n20684) );
  INV_X1 U18877 ( .A(n20684), .ZN(n20678) );
  OAI211_X1 U18878 ( .C1(n20680), .C2(n15755), .A(n15754), .B(n20678), .ZN(
        P1_U3195) );
  INV_X1 U18879 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16382) );
  NOR2_X1 U18880 ( .A1(n20007), .A2(n16382), .ZN(P1_U2905) );
  INV_X1 U18881 ( .A(n16228), .ZN(n19886) );
  OAI221_X1 U18882 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n19630), .C1(n18737), 
        .C2(n19886), .A(n19491), .ZN(n19756) );
  OAI211_X1 U18883 ( .C1(P2_STATE2_REG_1__SCAN_IN), .C2(
        P2_STATE2_REG_2__SCAN_IN), .A(n15758), .B(n19756), .ZN(n15756) );
  INV_X1 U18884 ( .A(n15756), .ZN(P2_U3178) );
  OAI211_X1 U18885 ( .C1(n19875), .C2(n15758), .A(n15757), .B(n19452), .ZN(
        n19866) );
  NOR2_X1 U18886 ( .A1(n15759), .A2(n19866), .ZN(P2_U3047) );
  NAND2_X1 U18887 ( .A1(n18716), .A2(n18062), .ZN(n15760) );
  NAND2_X1 U18888 ( .A1(n18094), .A2(n17244), .ZN(n17243) );
  INV_X1 U18889 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17334) );
  NAND2_X2 U18890 ( .A1(n17185), .A2(n17244), .ZN(n17221) );
  AOI22_X1 U18891 ( .A1(n17248), .A2(BUF2_REG_0__SCAN_IN), .B1(n17247), .B2(
        n15764), .ZN(n15765) );
  OAI221_X1 U18892 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17243), .C1(n17334), 
        .C2(n17244), .A(n15765), .ZN(P3_U2735) );
  NOR2_X1 U18893 ( .A1(n15785), .A2(n20727), .ZN(n15770) );
  AOI22_X1 U18894 ( .A1(n19982), .A2(P1_EBX_REG_21__SCAN_IN), .B1(n19986), 
        .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15766) );
  OAI21_X1 U18895 ( .B1(n15768), .B2(n15767), .A(n15766), .ZN(n15769) );
  NOR2_X1 U18896 ( .A1(n15770), .A2(n15769), .ZN(n15775) );
  OAI22_X1 U18897 ( .A1(n15772), .A2(n15810), .B1(n19971), .B2(n15771), .ZN(
        n15773) );
  INV_X1 U18898 ( .A(n15773), .ZN(n15774) );
  OAI211_X1 U18899 ( .C1(n15776), .C2(n19981), .A(n15775), .B(n15774), .ZN(
        P1_U2819) );
  AOI21_X1 U18900 ( .B1(n19925), .B2(n15777), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15784) );
  AOI22_X1 U18901 ( .A1(P1_EBX_REG_20__SCAN_IN), .A2(n19982), .B1(n19986), 
        .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15783) );
  OAI22_X1 U18902 ( .A1(n15779), .A2(n15810), .B1(n19971), .B2(n15778), .ZN(
        n15780) );
  AOI21_X1 U18903 ( .B1(n15781), .B2(n19993), .A(n15780), .ZN(n15782) );
  OAI211_X1 U18904 ( .C1(n15785), .C2(n15784), .A(n15783), .B(n15782), .ZN(
        P1_U2820) );
  NOR3_X1 U18905 ( .A1(n15838), .A2(P1_REIP_REG_19__SCAN_IN), .A3(n15786), 
        .ZN(n15791) );
  INV_X1 U18906 ( .A(n15787), .ZN(n15788) );
  NOR3_X1 U18907 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15838), .A3(n15788), 
        .ZN(n15797) );
  OAI21_X1 U18908 ( .B1(n15799), .B2(n15797), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15789) );
  OAI211_X1 U18909 ( .C1(n19928), .C2(n10757), .A(n15789), .B(n19962), .ZN(
        n15790) );
  AOI211_X1 U18910 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n19982), .A(n15791), .B(
        n15790), .ZN(n15794) );
  INV_X1 U18911 ( .A(n15792), .ZN(n15918) );
  AOI22_X1 U18912 ( .A1(n15859), .A2(n19955), .B1(n15918), .B2(n19983), .ZN(
        n15793) );
  OAI211_X1 U18913 ( .C1(n15862), .C2(n19981), .A(n15794), .B(n15793), .ZN(
        P1_U2821) );
  AOI21_X1 U18914 ( .B1(n19982), .B2(P1_EBX_REG_18__SCAN_IN), .A(n19973), .ZN(
        n15795) );
  OAI21_X1 U18915 ( .B1(n15796), .B2(n19928), .A(n15795), .ZN(n15798) );
  AOI211_X1 U18916 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n15799), .A(n15798), 
        .B(n15797), .ZN(n15800) );
  OAI21_X1 U18917 ( .B1(n15801), .B2(n15810), .A(n15800), .ZN(n15802) );
  AOI21_X1 U18918 ( .B1(n15803), .B2(n19993), .A(n15802), .ZN(n15804) );
  OAI21_X1 U18919 ( .B1(n19971), .B2(n15805), .A(n15804), .ZN(P1_U2822) );
  OAI21_X1 U18920 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n15806), .ZN(n15816) );
  AOI22_X1 U18921 ( .A1(n15820), .A2(P1_REIP_REG_16__SCAN_IN), .B1(n19982), 
        .B2(P1_EBX_REG_16__SCAN_IN), .ZN(n15807) );
  OAI211_X1 U18922 ( .C1(n19928), .C2(n15808), .A(n15807), .B(n19962), .ZN(
        n15813) );
  OAI22_X1 U18923 ( .A1(n15811), .A2(n15810), .B1(n19971), .B2(n15809), .ZN(
        n15812) );
  AOI211_X1 U18924 ( .C1(n15814), .C2(n19993), .A(n15813), .B(n15812), .ZN(
        n15815) );
  OAI21_X1 U18925 ( .B1(n15824), .B2(n15816), .A(n15815), .ZN(P1_U2824) );
  AOI22_X1 U18926 ( .A1(n19982), .A2(P1_EBX_REG_15__SCAN_IN), .B1(n19993), 
        .B2(n15880), .ZN(n15817) );
  OAI211_X1 U18927 ( .C1(n19928), .C2(n15818), .A(n15817), .B(n19962), .ZN(
        n15819) );
  AOI21_X1 U18928 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n15820), .A(n15819), 
        .ZN(n15823) );
  INV_X1 U18929 ( .A(n15821), .ZN(n15934) );
  AOI22_X1 U18930 ( .A1(n15881), .A2(n19955), .B1(n19983), .B2(n15934), .ZN(
        n15822) );
  OAI211_X1 U18931 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n15824), .A(n15823), 
        .B(n15822), .ZN(P1_U2825) );
  AOI22_X1 U18932 ( .A1(n19982), .A2(P1_EBX_REG_12__SCAN_IN), .B1(n19986), 
        .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15832) );
  AOI21_X1 U18933 ( .B1(n15951), .B2(n19983), .A(n19973), .ZN(n15831) );
  INV_X1 U18934 ( .A(n15825), .ZN(n15887) );
  AOI22_X1 U18935 ( .A1(n15888), .A2(n19993), .B1(n19955), .B2(n15887), .ZN(
        n15830) );
  INV_X1 U18936 ( .A(n15826), .ZN(n15827) );
  OAI21_X1 U18937 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(n15828), .A(n15827), 
        .ZN(n15829) );
  NAND4_X1 U18938 ( .A1(n15832), .A2(n15831), .A3(n15830), .A4(n15829), .ZN(
        P1_U2828) );
  NAND2_X1 U18939 ( .A1(n15834), .A2(n15833), .ZN(n15853) );
  OAI22_X1 U18940 ( .A1(n15960), .A2(n19971), .B1(n19936), .B2(n15835), .ZN(
        n15836) );
  INV_X1 U18941 ( .A(n15836), .ZN(n15843) );
  NOR2_X1 U18942 ( .A1(n15838), .A2(n15837), .ZN(n15839) );
  AOI22_X1 U18943 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19986), .B1(
        n15839), .B2(n20710), .ZN(n15840) );
  OAI211_X1 U18944 ( .C1(n19981), .C2(n15900), .A(n15840), .B(n19962), .ZN(
        n15841) );
  AOI21_X1 U18945 ( .B1(n19955), .B2(n15897), .A(n15841), .ZN(n15842) );
  OAI211_X1 U18946 ( .C1(n20710), .C2(n15853), .A(n15843), .B(n15842), .ZN(
        P1_U2829) );
  INV_X1 U18947 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20708) );
  NOR2_X1 U18948 ( .A1(n20708), .A2(n15844), .ZN(n19934) );
  NOR2_X1 U18949 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n19934), .ZN(n15854) );
  OAI22_X1 U18950 ( .A1(n15846), .A2(n19971), .B1(n15845), .B2(n19936), .ZN(
        n15847) );
  AOI211_X1 U18951 ( .C1(n19986), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19973), .B(n15847), .ZN(n15852) );
  INV_X1 U18952 ( .A(n15848), .ZN(n15849) );
  AOI22_X1 U18953 ( .A1(n15850), .A2(n19955), .B1(n15849), .B2(n19993), .ZN(
        n15851) );
  OAI211_X1 U18954 ( .C1(n15854), .C2(n15853), .A(n15852), .B(n15851), .ZN(
        P1_U2830) );
  AOI22_X1 U18955 ( .A1(n20025), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20024), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15861) );
  NOR2_X1 U18956 ( .A1(n9581), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15855) );
  MUX2_X1 U18957 ( .A(n9582), .B(n15855), .S(n14453), .Z(n15858) );
  XNOR2_X1 U18958 ( .A(n15858), .B(n15857), .ZN(n15919) );
  AOI22_X1 U18959 ( .A1(n15859), .A2(n20031), .B1(n20032), .B2(n15919), .ZN(
        n15860) );
  OAI211_X1 U18960 ( .C1(n20036), .C2(n15862), .A(n15861), .B(n15860), .ZN(
        P1_U2980) );
  NAND2_X1 U18961 ( .A1(n15892), .A2(n15863), .ZN(n15869) );
  INV_X1 U18962 ( .A(n15864), .ZN(n15866) );
  OAI21_X1 U18963 ( .B1(n15867), .B2(n15866), .A(n15865), .ZN(n15868) );
  MUX2_X1 U18964 ( .A(n15892), .B(n15869), .S(n15868), .Z(n15870) );
  XNOR2_X1 U18965 ( .A(n15870), .B(n11146), .ZN(n15931) );
  AOI22_X1 U18966 ( .A1(n20025), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20024), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15875) );
  INV_X1 U18967 ( .A(n15871), .ZN(n15873) );
  AOI22_X1 U18968 ( .A1(n15873), .A2(n20031), .B1(n15889), .B2(n15872), .ZN(
        n15874) );
  OAI211_X1 U18969 ( .C1(n19908), .C2(n15931), .A(n15875), .B(n15874), .ZN(
        P1_U2982) );
  OAI21_X1 U18970 ( .B1(n15878), .B2(n15877), .A(n15876), .ZN(n15879) );
  INV_X1 U18971 ( .A(n15879), .ZN(n15938) );
  AOI22_X1 U18972 ( .A1(n20025), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20024), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15883) );
  AOI22_X1 U18973 ( .A1(n15881), .A2(n20031), .B1(n15889), .B2(n15880), .ZN(
        n15882) );
  OAI211_X1 U18974 ( .C1(n15938), .C2(n19908), .A(n15883), .B(n15882), .ZN(
        P1_U2984) );
  AOI21_X1 U18975 ( .B1(n15886), .B2(n15885), .A(n15884), .ZN(n15959) );
  AOI22_X1 U18976 ( .A1(n20025), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20024), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15891) );
  AOI22_X1 U18977 ( .A1(n15889), .A2(n15888), .B1(n20031), .B2(n15887), .ZN(
        n15890) );
  OAI211_X1 U18978 ( .C1(n15959), .C2(n19908), .A(n15891), .B(n15890), .ZN(
        P1_U2987) );
  AOI22_X1 U18979 ( .A1(n20025), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20024), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15899) );
  NOR3_X1 U18980 ( .A1(n15893), .A2(n15892), .A3(n11269), .ZN(n15895) );
  NOR2_X1 U18981 ( .A1(n15895), .A2(n15894), .ZN(n15896) );
  XNOR2_X1 U18982 ( .A(n15896), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15963) );
  AOI22_X1 U18983 ( .A1(n20032), .A2(n15963), .B1(n20031), .B2(n15897), .ZN(
        n15898) );
  OAI211_X1 U18984 ( .C1(n20036), .C2(n15900), .A(n15899), .B(n15898), .ZN(
        P1_U2988) );
  AOI22_X1 U18985 ( .A1(n20025), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20024), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15906) );
  NAND2_X1 U18986 ( .A1(n15903), .A2(n15902), .ZN(n15904) );
  XNOR2_X1 U18987 ( .A(n15901), .B(n15904), .ZN(n15990) );
  AOI22_X1 U18988 ( .A1(n15990), .A2(n20032), .B1(n20031), .B2(n19944), .ZN(
        n15905) );
  OAI211_X1 U18989 ( .C1(n20036), .C2(n19947), .A(n15906), .B(n15905), .ZN(
        P1_U2992) );
  AOI22_X1 U18990 ( .A1(n20025), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20024), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15909) );
  AOI22_X1 U18991 ( .A1(n15907), .A2(n20032), .B1(n20031), .B2(n19956), .ZN(
        n15908) );
  OAI211_X1 U18992 ( .C1(n20036), .C2(n19959), .A(n15909), .B(n15908), .ZN(
        P1_U2993) );
  AOI22_X1 U18993 ( .A1(n20025), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20024), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15916) );
  OAI21_X1 U18994 ( .B1(n15912), .B2(n15911), .A(n15910), .ZN(n15913) );
  INV_X1 U18995 ( .A(n15913), .ZN(n15996) );
  INV_X1 U18996 ( .A(n15914), .ZN(n19966) );
  AOI22_X1 U18997 ( .A1(n15996), .A2(n20032), .B1(n20031), .B2(n19966), .ZN(
        n15915) );
  OAI211_X1 U18998 ( .C1(n20036), .C2(n19964), .A(n15916), .B(n15915), .ZN(
        P1_U2994) );
  AOI22_X1 U18999 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15917), .B1(
        n20024), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15921) );
  AOI22_X1 U19000 ( .A1(n15919), .A2(n20062), .B1(n20048), .B2(n15918), .ZN(
        n15920) );
  OAI211_X1 U19001 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15922), .A(
        n15921), .B(n15920), .ZN(P1_U3012) );
  OAI21_X1 U19002 ( .B1(n15923), .B2(n15933), .A(n11146), .ZN(n15928) );
  INV_X1 U19003 ( .A(n15924), .ZN(n15927) );
  INV_X1 U19004 ( .A(n15925), .ZN(n15926) );
  AOI22_X1 U19005 ( .A1(n15928), .A2(n15927), .B1(n20048), .B2(n15926), .ZN(
        n15930) );
  NAND2_X1 U19006 ( .A1(n20024), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15929) );
  OAI211_X1 U19007 ( .C1(n15931), .C2(n20073), .A(n15930), .B(n15929), .ZN(
        P1_U3014) );
  AOI22_X1 U19008 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15932), .B1(
        n20024), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15937) );
  INV_X1 U19009 ( .A(n15933), .ZN(n15935) );
  AOI22_X1 U19010 ( .A1(n15935), .A2(n11145), .B1(n20048), .B2(n15934), .ZN(
        n15936) );
  OAI211_X1 U19011 ( .C1(n15938), .C2(n20073), .A(n15937), .B(n15936), .ZN(
        P1_U3016) );
  AOI22_X1 U19012 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15939), .B1(
        n20024), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n15944) );
  INV_X1 U19013 ( .A(n15940), .ZN(n15942) );
  AOI22_X1 U19014 ( .A1(n15942), .A2(n20062), .B1(n20048), .B2(n15941), .ZN(
        n15943) );
  OAI211_X1 U19015 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n15945), .A(
        n15944), .B(n15943), .ZN(P1_U3018) );
  OAI21_X1 U19016 ( .B1(n15947), .B2(n20057), .A(n15946), .ZN(n15948) );
  AOI21_X1 U19017 ( .B1(n20061), .B2(n15949), .A(n15948), .ZN(n15967) );
  AOI221_X1 U19018 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15967), 
        .C1(n15950), .C2(n15967), .A(n15956), .ZN(n15955) );
  NAND2_X1 U19019 ( .A1(n15951), .A2(n20048), .ZN(n15953) );
  NAND2_X1 U19020 ( .A1(n20024), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15952) );
  NAND2_X1 U19021 ( .A1(n15953), .A2(n15952), .ZN(n15954) );
  NOR2_X1 U19022 ( .A1(n15955), .A2(n15954), .ZN(n15958) );
  NAND3_X1 U19023 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15962), .A3(
        n15956), .ZN(n15957) );
  OAI211_X1 U19024 ( .C1(n15959), .C2(n20073), .A(n15958), .B(n15957), .ZN(
        P1_U3019) );
  OAI22_X1 U19025 ( .A1(n15960), .A2(n20079), .B1(n20065), .B2(n20710), .ZN(
        n15961) );
  INV_X1 U19026 ( .A(n15961), .ZN(n15965) );
  AOI22_X1 U19027 ( .A1(n15963), .A2(n20062), .B1(n15962), .B2(n15966), .ZN(
        n15964) );
  OAI211_X1 U19028 ( .C1(n15967), .C2(n15966), .A(n15965), .B(n15964), .ZN(
        P1_U3020) );
  INV_X1 U19029 ( .A(n15968), .ZN(n15977) );
  NAND2_X1 U19030 ( .A1(n15970), .A2(n15969), .ZN(n15971) );
  AND2_X1 U19031 ( .A1(n15972), .A2(n15971), .ZN(n19998) );
  INV_X1 U19032 ( .A(n19998), .ZN(n15973) );
  OAI22_X1 U19033 ( .A1(n15973), .A2(n20079), .B1(n20708), .B2(n20065), .ZN(
        n15976) );
  NOR2_X1 U19034 ( .A1(n15974), .A2(n20073), .ZN(n15975) );
  AOI211_X1 U19035 ( .C1(n15980), .C2(n15977), .A(n15976), .B(n15975), .ZN(
        n15978) );
  OAI21_X1 U19036 ( .B1(n15980), .B2(n15979), .A(n15978), .ZN(P1_U3022) );
  INV_X1 U19037 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15989) );
  NAND2_X1 U19038 ( .A1(n15982), .A2(n15981), .ZN(n15992) );
  NAND2_X1 U19039 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15983), .ZN(
        n15994) );
  AOI221_X1 U19040 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n15989), .C2(n15993), .A(
        n15994), .ZN(n15986) );
  OAI22_X1 U19041 ( .A1(n15984), .A2(n20079), .B1(n20706), .B2(n20065), .ZN(
        n15985) );
  AOI211_X1 U19042 ( .C1(n15987), .C2(n20062), .A(n15986), .B(n15985), .ZN(
        n15988) );
  OAI21_X1 U19043 ( .B1(n15989), .B2(n15992), .A(n15988), .ZN(P1_U3023) );
  AOI222_X1 U19044 ( .A1(n15990), .A2(n20062), .B1(n20048), .B2(n19935), .C1(
        P1_REIP_REG_7__SCAN_IN), .C2(n20024), .ZN(n15991) );
  OAI221_X1 U19045 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15994), .C1(
        n15993), .C2(n15992), .A(n15991), .ZN(P1_U3024) );
  AOI22_X1 U19046 ( .A1(n20048), .A2(n19960), .B1(n20024), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n15998) );
  AOI22_X1 U19047 ( .A1(n15996), .A2(n20062), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n15995), .ZN(n15997) );
  OAI211_X1 U19048 ( .C1(n20049), .C2(n15999), .A(n15998), .B(n15997), .ZN(
        P1_U3026) );
  INV_X1 U19049 ( .A(n16000), .ZN(n16001) );
  NAND3_X1 U19050 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20613), .A3(n16001), 
        .ZN(n16002) );
  NAND2_X1 U19051 ( .A1(n16003), .A2(n16002), .ZN(n20676) );
  NOR2_X1 U19052 ( .A1(n16004), .A2(n10259), .ZN(n16010) );
  AOI21_X1 U19053 ( .B1(n16010), .B2(n16005), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n16006) );
  AOI221_X1 U19054 ( .B1(n16008), .B2(n16007), .C1(n20676), .C2(n16007), .A(
        n16006), .ZN(P1_U3162) );
  OAI21_X1 U19055 ( .B1(n16010), .B2(n20510), .A(n16009), .ZN(P1_U3466) );
  NAND2_X1 U19056 ( .A1(n18915), .A2(n16011), .ZN(n16049) );
  NAND2_X1 U19057 ( .A1(n16049), .A2(n16050), .ZN(n16048) );
  NAND2_X1 U19058 ( .A1(n18915), .A2(n16048), .ZN(n16037) );
  INV_X1 U19059 ( .A(n16012), .ZN(n16038) );
  NAND2_X1 U19060 ( .A1(n16037), .A2(n16038), .ZN(n16036) );
  NAND2_X1 U19061 ( .A1(n18915), .A2(n16036), .ZN(n16029) );
  NAND2_X1 U19062 ( .A1(n16029), .A2(n16028), .ZN(n16027) );
  INV_X1 U19063 ( .A(n16013), .ZN(n16014) );
  OAI222_X1 U19064 ( .A1(n16015), .A2(n16100), .B1(n18941), .B2(n16014), .C1(
        n19820), .C2(n18873), .ZN(n16016) );
  AOI21_X1 U19065 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n18950), .A(
        n16016), .ZN(n16020) );
  INV_X1 U19066 ( .A(n18990), .ZN(n16017) );
  OAI22_X1 U19067 ( .A1(n16101), .A2(n18911), .B1(n16017), .B2(n18925), .ZN(
        n16018) );
  INV_X1 U19068 ( .A(n16018), .ZN(n16019) );
  OAI211_X1 U19069 ( .C1(n18839), .C2(n16027), .A(n16020), .B(n16019), .ZN(
        P2_U2824) );
  INV_X1 U19070 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n16021) );
  OAI22_X1 U19071 ( .A1(n18909), .A2(n16021), .B1(n12343), .B2(n18873), .ZN(
        n16025) );
  INV_X1 U19072 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16022) );
  OAI22_X1 U19073 ( .A1(n16023), .A2(n18925), .B1(n16022), .B2(n18892), .ZN(
        n16024) );
  AOI211_X1 U19074 ( .C1(n16026), .C2(n18906), .A(n16025), .B(n16024), .ZN(
        n16031) );
  OAI211_X1 U19075 ( .C1(n16029), .C2(n16028), .A(n16027), .B(n18901), .ZN(
        n16030) );
  OAI211_X1 U19076 ( .C1(n18911), .C2(n16032), .A(n16031), .B(n16030), .ZN(
        P2_U2825) );
  AOI22_X1 U19077 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n18935), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n18936), .ZN(n16042) );
  AOI22_X1 U19078 ( .A1(n16033), .A2(n18906), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18950), .ZN(n16041) );
  AOI22_X1 U19079 ( .A1(n16035), .A2(n18944), .B1(n16034), .B2(n18937), .ZN(
        n16040) );
  OAI211_X1 U19080 ( .C1(n16038), .C2(n16037), .A(n18901), .B(n16036), .ZN(
        n16039) );
  NAND4_X1 U19081 ( .A1(n16042), .A2(n16041), .A3(n16040), .A4(n16039), .ZN(
        P2_U2826) );
  INV_X1 U19082 ( .A(n16043), .ZN(n16047) );
  INV_X1 U19083 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19812) );
  OAI22_X1 U19084 ( .A1(n18909), .A2(n11857), .B1(n19812), .B2(n18873), .ZN(
        n16046) );
  OAI22_X1 U19085 ( .A1(n16044), .A2(n18925), .B1(n15043), .B2(n18892), .ZN(
        n16045) );
  AOI211_X1 U19086 ( .C1(n16047), .C2(n18906), .A(n16046), .B(n16045), .ZN(
        n16052) );
  OAI211_X1 U19087 ( .C1(n16050), .C2(n16049), .A(n18901), .B(n16048), .ZN(
        n16051) );
  OAI211_X1 U19088 ( .C1(n18911), .C2(n16053), .A(n16052), .B(n16051), .ZN(
        P2_U2827) );
  AOI22_X1 U19089 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n18935), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n18936), .ZN(n16064) );
  AOI22_X1 U19090 ( .A1(n16054), .A2(n18906), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18950), .ZN(n16063) );
  OAI22_X1 U19091 ( .A1(n16056), .A2(n18911), .B1(n16055), .B2(n18925), .ZN(
        n16057) );
  INV_X1 U19092 ( .A(n16057), .ZN(n16062) );
  OAI211_X1 U19093 ( .C1(n16060), .C2(n16059), .A(n18901), .B(n16058), .ZN(
        n16061) );
  NAND4_X1 U19094 ( .A1(n16064), .A2(n16063), .A3(n16062), .A4(n16061), .ZN(
        P2_U2829) );
  OAI22_X1 U19095 ( .A1(n18909), .A2(n16072), .B1(n19806), .B2(n18873), .ZN(
        n16065) );
  AOI21_X1 U19096 ( .B1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18950), .A(
        n16065), .ZN(n16076) );
  AOI22_X1 U19097 ( .A1(n16067), .A2(n18944), .B1(n18937), .B2(n16066), .ZN(
        n16075) );
  OAI211_X1 U19098 ( .C1(n16070), .C2(n16069), .A(n18901), .B(n16068), .ZN(
        n16074) );
  OAI211_X1 U19099 ( .C1(n9686), .C2(n16072), .A(n16071), .B(n18906), .ZN(
        n16073) );
  NAND4_X1 U19100 ( .A1(n16076), .A2(n16075), .A3(n16074), .A4(n16073), .ZN(
        P2_U2830) );
  OAI22_X1 U19101 ( .A1(n18909), .A2(n9809), .B1(n19804), .B2(n18873), .ZN(
        n16077) );
  INV_X1 U19102 ( .A(n16077), .ZN(n16078) );
  OAI21_X1 U19103 ( .B1(n18892), .B2(n9891), .A(n16078), .ZN(n16079) );
  AOI21_X1 U19104 ( .B1(n18937), .B2(n16080), .A(n16079), .ZN(n16081) );
  OAI21_X1 U19105 ( .B1(n16082), .B2(n18941), .A(n16081), .ZN(n16083) );
  INV_X1 U19106 ( .A(n16083), .ZN(n16088) );
  OAI211_X1 U19107 ( .C1(n16086), .C2(n16085), .A(n18901), .B(n16084), .ZN(
        n16087) );
  OAI211_X1 U19108 ( .C1(n18911), .C2(n16089), .A(n16088), .B(n16087), .ZN(
        P2_U2831) );
  AOI22_X1 U19109 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n18935), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n18936), .ZN(n16099) );
  AOI22_X1 U19110 ( .A1(n16090), .A2(n18906), .B1(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18950), .ZN(n16098) );
  AOI22_X1 U19111 ( .A1(n16092), .A2(n18944), .B1(n18937), .B2(n16091), .ZN(
        n16097) );
  OAI211_X1 U19112 ( .C1(n16095), .C2(n16094), .A(n18901), .B(n16093), .ZN(
        n16096) );
  NAND4_X1 U19113 ( .A1(n16099), .A2(n16098), .A3(n16097), .A4(n16096), .ZN(
        P2_U2832) );
  AOI22_X1 U19114 ( .A1(n18988), .A2(n16101), .B1(n16100), .B2(n18983), .ZN(
        P2_U2856) );
  AOI21_X1 U19115 ( .B1(n16103), .B2(n14913), .A(n16102), .ZN(n16115) );
  AOI22_X1 U19116 ( .A1(n16115), .A2(n18954), .B1(n18988), .B2(n16129), .ZN(
        n16104) );
  OAI21_X1 U19117 ( .B1(n18988), .B2(n16105), .A(n16104), .ZN(P2_U2865) );
  NOR2_X1 U19118 ( .A1(n14922), .A2(n16106), .ZN(n16107) );
  AOI22_X1 U19119 ( .A1(n10028), .A2(n18954), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n18983), .ZN(n16108) );
  OAI21_X1 U19120 ( .B1(n18983), .B2(n16109), .A(n16108), .ZN(P2_U2867) );
  INV_X1 U19121 ( .A(n14921), .ZN(n16110) );
  AOI21_X1 U19122 ( .B1(n16111), .B2(n13791), .A(n16110), .ZN(n16124) );
  AOI22_X1 U19123 ( .A1(n16124), .A2(n18954), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n18983), .ZN(n16112) );
  OAI21_X1 U19124 ( .B1(n18983), .B2(n18792), .A(n16112), .ZN(P2_U2869) );
  INV_X1 U19125 ( .A(n19152), .ZN(n16113) );
  AOI22_X1 U19126 ( .A1(n20782), .A2(n16113), .B1(n20780), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16118) );
  AOI22_X1 U19127 ( .A1(n20783), .A2(BUF1_REG_22__SCAN_IN), .B1(n20784), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16117) );
  AOI22_X1 U19128 ( .A1(n16115), .A2(n20791), .B1(n18989), .B2(n16114), .ZN(
        n16116) );
  NAND3_X1 U19129 ( .A1(n16118), .A2(n16117), .A3(n16116), .ZN(P2_U2897) );
  AOI22_X1 U19130 ( .A1(n20782), .A2(n16119), .B1(n20780), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16122) );
  AOI22_X1 U19131 ( .A1(n20783), .A2(BUF1_REG_20__SCAN_IN), .B1(n20784), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16121) );
  AOI22_X1 U19132 ( .A1(n18763), .A2(n18989), .B1(n20791), .B2(n10028), .ZN(
        n16120) );
  NAND3_X1 U19133 ( .A1(n16122), .A2(n16121), .A3(n16120), .ZN(P2_U2899) );
  AOI22_X1 U19134 ( .A1(n20782), .A2(n19126), .B1(n20780), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16127) );
  AOI22_X1 U19135 ( .A1(n20783), .A2(BUF1_REG_18__SCAN_IN), .B1(n20784), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16126) );
  INV_X1 U19136 ( .A(n16123), .ZN(n18789) );
  AOI22_X1 U19137 ( .A1(n20791), .A2(n16124), .B1(n18789), .B2(n18989), .ZN(
        n16125) );
  NAND3_X1 U19138 ( .A1(n16127), .A2(n16126), .A3(n16125), .ZN(P2_U2901) );
  AOI22_X1 U19139 ( .A1(n16156), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19090), .ZN(n16135) );
  NAND2_X1 U19140 ( .A1(n16128), .A2(n19095), .ZN(n16131) );
  NAND2_X1 U19141 ( .A1(n16129), .A2(n19094), .ZN(n16130) );
  OAI211_X1 U19142 ( .C1(n16169), .C2(n16132), .A(n16131), .B(n16130), .ZN(
        n16133) );
  INV_X1 U19143 ( .A(n16133), .ZN(n16134) );
  OAI211_X1 U19144 ( .C1(n16166), .C2(n16136), .A(n16135), .B(n16134), .ZN(
        P2_U2992) );
  AOI22_X1 U19145 ( .A1(n16156), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19090), .ZN(n16141) );
  INV_X1 U19146 ( .A(n18962), .ZN(n16137) );
  AOI222_X1 U19147 ( .A1(n16139), .A2(n19091), .B1(n19095), .B2(n16138), .C1(
        n19094), .C2(n16137), .ZN(n16140) );
  OAI211_X1 U19148 ( .C1(n16166), .C2(n18808), .A(n16141), .B(n16140), .ZN(
        P2_U3000) );
  AOI22_X1 U19149 ( .A1(n16156), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19090), .ZN(n16149) );
  NAND2_X1 U19150 ( .A1(n16142), .A2(n19095), .ZN(n16145) );
  NAND2_X1 U19151 ( .A1(n19094), .A2(n16143), .ZN(n16144) );
  OAI211_X1 U19152 ( .C1(n16146), .C2(n16169), .A(n16145), .B(n16144), .ZN(
        n16147) );
  INV_X1 U19153 ( .A(n16147), .ZN(n16148) );
  OAI211_X1 U19154 ( .C1(n16166), .C2(n16150), .A(n16149), .B(n16148), .ZN(
        P2_U3002) );
  AOI22_X1 U19155 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19090), .B1(n19089), 
        .B2(n18837), .ZN(n16155) );
  OAI22_X1 U19156 ( .A1(n16152), .A2(n16169), .B1(n16151), .B2(n16168), .ZN(
        n16153) );
  AOI21_X1 U19157 ( .B1(n19094), .B2(n18838), .A(n16153), .ZN(n16154) );
  OAI211_X1 U19158 ( .C1(n19100), .C2(n18831), .A(n16155), .B(n16154), .ZN(
        P2_U3003) );
  AOI22_X1 U19159 ( .A1(n16156), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19090), .ZN(n16164) );
  NAND2_X1 U19160 ( .A1(n16157), .A2(n19095), .ZN(n16160) );
  NAND2_X1 U19161 ( .A1(n19094), .A2(n16158), .ZN(n16159) );
  OAI211_X1 U19162 ( .C1(n16161), .C2(n16169), .A(n16160), .B(n16159), .ZN(
        n16162) );
  INV_X1 U19163 ( .A(n16162), .ZN(n16163) );
  OAI211_X1 U19164 ( .C1(n16166), .C2(n16165), .A(n16164), .B(n16163), .ZN(
        P2_U3004) );
  AOI22_X1 U19165 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19090), .B1(n19089), 
        .B2(n18848), .ZN(n16174) );
  OAI22_X1 U19166 ( .A1(n16170), .A2(n16169), .B1(n16168), .B2(n16167), .ZN(
        n16171) );
  AOI21_X1 U19167 ( .B1(n19094), .B2(n16172), .A(n16171), .ZN(n16173) );
  OAI211_X1 U19168 ( .C1(n19100), .C2(n16175), .A(n16174), .B(n16173), .ZN(
        P2_U3005) );
  AOI22_X1 U19169 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19090), .B1(n19089), 
        .B2(n18862), .ZN(n16188) );
  NAND2_X1 U19170 ( .A1(n16177), .A2(n16176), .ZN(n16182) );
  INV_X1 U19171 ( .A(n16178), .ZN(n16179) );
  AOI21_X1 U19172 ( .B1(n15207), .B2(n16180), .A(n16179), .ZN(n16181) );
  XOR2_X1 U19173 ( .A(n16182), .B(n16181), .Z(n16195) );
  NOR2_X1 U19174 ( .A1(n16183), .A2(n13161), .ZN(n16184) );
  OR2_X1 U19175 ( .A1(n9709), .A2(n16184), .ZN(n18981) );
  INV_X1 U19176 ( .A(n18981), .ZN(n16194) );
  XOR2_X1 U19177 ( .A(n16186), .B(n16185), .Z(n16193) );
  AOI222_X1 U19178 ( .A1(n16195), .A2(n19095), .B1(n19094), .B2(n16194), .C1(
        n16193), .C2(n19091), .ZN(n16187) );
  OAI211_X1 U19179 ( .C1(n19100), .C2(n16189), .A(n16188), .B(n16187), .ZN(
        P2_U3006) );
  NOR2_X1 U19180 ( .A1(n16191), .A2(n16190), .ZN(n16208) );
  AOI22_X1 U19181 ( .A1(n16208), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16217), .B2(n18863), .ZN(n16203) );
  AOI222_X1 U19182 ( .A1(n16195), .A2(n16210), .B1(n16218), .B2(n16194), .C1(
        n16193), .C2(n16192), .ZN(n16202) );
  NAND2_X1 U19183 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19090), .ZN(n16201) );
  NOR3_X1 U19184 ( .A1(n16198), .A2(n16197), .A3(n16196), .ZN(n16207) );
  OAI221_X1 U19185 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16199), .C2(n16206), .A(
        n16207), .ZN(n16200) );
  NAND4_X1 U19186 ( .A1(n16203), .A2(n16202), .A3(n16201), .A4(n16200), .ZN(
        P2_U3038) );
  OAI22_X1 U19187 ( .A1(n18875), .A2(n16204), .B1(n15210), .B2(n18871), .ZN(
        n16205) );
  AOI221_X1 U19188 ( .B1(n16208), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(
        n16207), .C2(n16206), .A(n16205), .ZN(n16213) );
  INV_X1 U19189 ( .A(n18874), .ZN(n16209) );
  AOI22_X1 U19190 ( .A1(n16211), .A2(n16210), .B1(n16218), .B2(n16209), .ZN(
        n16212) );
  OAI211_X1 U19191 ( .C1(n16227), .C2(n16214), .A(n16213), .B(n16212), .ZN(
        P2_U3039) );
  MUX2_X1 U19192 ( .A(n16216), .B(n16215), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n16220) );
  AOI22_X1 U19193 ( .A1(n16218), .A2(n18945), .B1(n16217), .B2(n18938), .ZN(
        n16219) );
  OAI211_X1 U19194 ( .C1(n16222), .C2(n16221), .A(n16220), .B(n16219), .ZN(
        n16223) );
  INV_X1 U19195 ( .A(n16223), .ZN(n16225) );
  OAI211_X1 U19196 ( .C1(n16227), .C2(n16226), .A(n16225), .B(n16224), .ZN(
        P2_U3046) );
  NOR3_X1 U19197 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n18737), .A3(n16228), 
        .ZN(n16230) );
  AOI211_X1 U19198 ( .C1(n16231), .C2(n19875), .A(n16230), .B(n16229), .ZN(
        n16235) );
  INV_X1 U19199 ( .A(n16232), .ZN(n19753) );
  OAI21_X1 U19200 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n10024), .A(n19885), 
        .ZN(n16233) );
  NAND2_X1 U19201 ( .A1(n16232), .A2(n19886), .ZN(n19755) );
  OAI22_X1 U19202 ( .A1(n16232), .A2(n16233), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n19755), .ZN(n16234) );
  OAI211_X1 U19203 ( .C1(n16237), .C2(n16236), .A(n16235), .B(n16234), .ZN(
        P2_U3176) );
  XOR2_X1 U19204 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n16254), .Z(
        n16435) );
  OAI221_X1 U19205 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16240), .C1(
        n9924), .C2(n16239), .A(n16238), .ZN(n16241) );
  AOI21_X1 U19206 ( .B1(n17582), .B2(n16435), .A(n16241), .ZN(n16248) );
  NAND2_X1 U19207 ( .A1(n17727), .A2(n16242), .ZN(n16266) );
  OAI21_X1 U19208 ( .B1(n16243), .B2(n17646), .A(n16266), .ZN(n16246) );
  OAI22_X1 U19209 ( .A1(n17646), .A2(n17920), .B1(n17739), .B2(n17922), .ZN(
        n17599) );
  NOR2_X2 U19210 ( .A1(n17624), .A2(n16244), .ZN(n17533) );
  INV_X1 U19211 ( .A(n17533), .ZN(n17454) );
  INV_X1 U19212 ( .A(n17428), .ZN(n17442) );
  NOR2_X1 U19213 ( .A1(n16280), .A2(n17442), .ZN(n17392) );
  AOI22_X1 U19214 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16246), .B1(
        n16245), .B2(n17392), .ZN(n16247) );
  OAI211_X1 U19215 ( .C1(n16249), .C2(n17642), .A(n16248), .B(n16247), .ZN(
        P3_U2800) );
  NAND2_X1 U19216 ( .A1(n16251), .A2(n16250), .ZN(n16285) );
  NAND2_X1 U19217 ( .A1(n18038), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16261) );
  NOR2_X1 U19218 ( .A1(n17745), .A2(n16252), .ZN(n16291) );
  OAI211_X1 U19219 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16291), .A(
        n17598), .B(n16253), .ZN(n16260) );
  AOI21_X1 U19220 ( .B1(n9923), .B2(n16413), .A(n16254), .ZN(n16443) );
  OAI21_X1 U19221 ( .B1(n16255), .B2(n17582), .A(n16443), .ZN(n16259) );
  OAI221_X1 U19222 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16257), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n18374), .A(n16256), .ZN(
        n16258) );
  NAND4_X1 U19223 ( .A1(n16261), .A2(n16260), .A3(n16259), .A4(n16258), .ZN(
        n16262) );
  AOI21_X1 U19224 ( .B1(n17615), .B2(n16263), .A(n16262), .ZN(n16264) );
  OAI221_X1 U19225 ( .B1(n16266), .B2(n16265), .C1(n16266), .C2(n16285), .A(
        n16264), .ZN(P3_U2801) );
  NAND3_X1 U19226 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16267), .A3(
        n18676), .ZN(n16269) );
  OAI22_X1 U19227 ( .A1(n18676), .A2(n16270), .B1(n16269), .B2(n16268), .ZN(
        n16271) );
  AOI211_X1 U19228 ( .C1(n16273), .C2(n18033), .A(n16272), .B(n16271), .ZN(
        n16277) );
  AOI22_X1 U19229 ( .A1(n16275), .A2(n17897), .B1(n17936), .B2(n16274), .ZN(
        n16276) );
  OAI211_X1 U19230 ( .C1(n16278), .C2(n18014), .A(n16277), .B(n16276), .ZN(
        P3_U2831) );
  INV_X1 U19231 ( .A(n18494), .ZN(n18023) );
  INV_X1 U19232 ( .A(n16288), .ZN(n18500) );
  NOR2_X1 U19233 ( .A1(n17217), .A2(n18500), .ZN(n17921) );
  OAI22_X1 U19234 ( .A1(n18023), .A2(n17922), .B1(n17920), .B2(n17904), .ZN(
        n17901) );
  AOI21_X1 U19235 ( .B1(n17901), .B2(n17521), .A(n17766), .ZN(n17806) );
  NOR2_X1 U19236 ( .A1(n16279), .A2(n17806), .ZN(n17757) );
  INV_X1 U19237 ( .A(n17757), .ZN(n17793) );
  NOR2_X1 U19238 ( .A1(n18049), .A2(n17793), .ZN(n17779) );
  NOR3_X1 U19239 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17752), .A3(
        n16280), .ZN(n17376) );
  AOI22_X1 U19240 ( .A1(n18038), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17779), 
        .B2(n17376), .ZN(n16296) );
  OAI22_X1 U19241 ( .A1(n17639), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n16281), .B2(n17608), .ZN(n17379) );
  OR3_X1 U19242 ( .A1(n16286), .A2(n17960), .A3(n17379), .ZN(n16295) );
  INV_X1 U19243 ( .A(n18041), .ZN(n18047) );
  NAND3_X1 U19244 ( .A1(n17384), .A2(n18047), .A3(n16282), .ZN(n16294) );
  AOI211_X1 U19245 ( .C1(n18494), .C2(n16285), .A(n16284), .B(n16283), .ZN(
        n16290) );
  OAI21_X1 U19246 ( .B1(n17384), .B2(n17639), .A(n16286), .ZN(n17378) );
  NAND2_X1 U19247 ( .A1(n17379), .A2(n17378), .ZN(n17377) );
  NAND4_X1 U19248 ( .A1(n16288), .A2(n17217), .A3(n16287), .A4(n17377), .ZN(
        n16289) );
  OAI211_X1 U19249 ( .C1(n16291), .C2(n17904), .A(n16290), .B(n16289), .ZN(
        n16292) );
  NAND3_X1 U19250 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18048), .A3(
        n16292), .ZN(n16293) );
  NAND4_X1 U19251 ( .A1(n16296), .A2(n16295), .A3(n16294), .A4(n16293), .ZN(
        P3_U2834) );
  NOR3_X1 U19252 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16298) );
  NOR4_X1 U19253 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16297) );
  NAND4_X1 U19254 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16298), .A3(n16297), .A4(
        U215), .ZN(U213) );
  INV_X1 U19255 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19013) );
  NOR2_X1 U19256 ( .A1(n16340), .A2(n16299), .ZN(n16343) );
  OAI222_X1 U19257 ( .A1(U212), .A2(n19013), .B1(n16347), .B2(n16300), .C1(
        U214), .C2(n16382), .ZN(U216) );
  INV_X2 U19258 ( .A(U212), .ZN(n16345) );
  AOI22_X1 U19259 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16345), .ZN(n16301) );
  OAI21_X1 U19260 ( .B1(n14072), .B2(n16347), .A(n16301), .ZN(U217) );
  INV_X1 U19261 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16303) );
  AOI22_X1 U19262 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16345), .ZN(n16302) );
  OAI21_X1 U19263 ( .B1(n16303), .B2(n16347), .A(n16302), .ZN(U218) );
  AOI222_X1 U19264 ( .A1(n16340), .A2(P1_DATAO_REG_28__SCAN_IN), .B1(n16343), 
        .B2(BUF1_REG_28__SCAN_IN), .C1(n16345), .C2(P2_DATAO_REG_28__SCAN_IN), 
        .ZN(n16304) );
  INV_X1 U19265 ( .A(n16304), .ZN(U219) );
  AOI22_X1 U19266 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16345), .ZN(n16305) );
  OAI21_X1 U19267 ( .B1(n16306), .B2(n16347), .A(n16305), .ZN(U220) );
  INV_X1 U19268 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n19124) );
  AOI22_X1 U19269 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16345), .ZN(n16307) );
  OAI21_X1 U19270 ( .B1(n19124), .B2(n16347), .A(n16307), .ZN(U221) );
  AOI22_X1 U19271 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16345), .ZN(n16308) );
  OAI21_X1 U19272 ( .B1(n19118), .B2(n16347), .A(n16308), .ZN(U222) );
  AOI22_X1 U19273 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16345), .ZN(n16309) );
  OAI21_X1 U19274 ( .B1(n14325), .B2(n16347), .A(n16309), .ZN(U223) );
  INV_X1 U19275 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16311) );
  AOI22_X1 U19276 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16345), .ZN(n16310) );
  OAI21_X1 U19277 ( .B1(n16311), .B2(n16347), .A(n16310), .ZN(U224) );
  INV_X1 U19278 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16313) );
  AOI22_X1 U19279 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16345), .ZN(n16312) );
  OAI21_X1 U19280 ( .B1(n16313), .B2(n16347), .A(n16312), .ZN(U225) );
  INV_X1 U19281 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n19143) );
  AOI22_X1 U19282 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16345), .ZN(n16314) );
  OAI21_X1 U19283 ( .B1(n19143), .B2(n16347), .A(n16314), .ZN(U226) );
  INV_X1 U19284 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n19137) );
  AOI22_X1 U19285 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16345), .ZN(n16315) );
  OAI21_X1 U19286 ( .B1(n19137), .B2(n16347), .A(n16315), .ZN(U227) );
  INV_X1 U19287 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n19130) );
  AOI22_X1 U19288 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16345), .ZN(n16316) );
  OAI21_X1 U19289 ( .B1(n19130), .B2(n16347), .A(n16316), .ZN(U228) );
  INV_X1 U19290 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16318) );
  AOI22_X1 U19291 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16345), .ZN(n16317) );
  OAI21_X1 U19292 ( .B1(n16318), .B2(n16347), .A(n16317), .ZN(U229) );
  INV_X1 U19293 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16320) );
  AOI22_X1 U19294 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16345), .ZN(n16319) );
  OAI21_X1 U19295 ( .B1(n16320), .B2(n16347), .A(n16319), .ZN(U230) );
  AOI22_X1 U19296 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16345), .ZN(n16321) );
  OAI21_X1 U19297 ( .B1(n13681), .B2(n16347), .A(n16321), .ZN(U231) );
  AOI22_X1 U19298 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16345), .ZN(n16322) );
  OAI21_X1 U19299 ( .B1(n13394), .B2(n16347), .A(n16322), .ZN(U232) );
  AOI22_X1 U19300 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16345), .ZN(n16323) );
  OAI21_X1 U19301 ( .B1(n12883), .B2(n16347), .A(n16323), .ZN(U233) );
  INV_X1 U19302 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16362) );
  INV_X1 U19303 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n20877) );
  OAI222_X1 U19304 ( .A1(U212), .A2(n16362), .B1(n16347), .B2(n14299), .C1(
        U214), .C2(n20877), .ZN(U234) );
  AOI22_X1 U19305 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16345), .ZN(n16324) );
  OAI21_X1 U19306 ( .B1(n16325), .B2(n16347), .A(n16324), .ZN(U235) );
  AOI22_X1 U19307 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16345), .ZN(n16326) );
  OAI21_X1 U19308 ( .B1(n13429), .B2(n16347), .A(n16326), .ZN(U236) );
  AOI22_X1 U19309 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16345), .ZN(n16327) );
  OAI21_X1 U19310 ( .B1(n16328), .B2(n16347), .A(n16327), .ZN(U237) );
  AOI22_X1 U19311 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16345), .ZN(n16329) );
  OAI21_X1 U19312 ( .B1(n16330), .B2(n16347), .A(n16329), .ZN(U238) );
  INV_X1 U19313 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16332) );
  AOI22_X1 U19314 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16345), .ZN(n16331) );
  OAI21_X1 U19315 ( .B1(n16332), .B2(n16347), .A(n16331), .ZN(U239) );
  INV_X1 U19316 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n20902) );
  AOI22_X1 U19317 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16343), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16345), .ZN(n16333) );
  OAI21_X1 U19318 ( .B1(n20902), .B2(U214), .A(n16333), .ZN(U240) );
  INV_X1 U19319 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16335) );
  AOI22_X1 U19320 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16345), .ZN(n16334) );
  OAI21_X1 U19321 ( .B1(n16335), .B2(n16347), .A(n16334), .ZN(U241) );
  INV_X1 U19322 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16354) );
  AOI22_X1 U19323 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16343), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16340), .ZN(n16336) );
  OAI21_X1 U19324 ( .B1(n16354), .B2(U212), .A(n16336), .ZN(U242) );
  INV_X1 U19325 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16338) );
  AOI22_X1 U19326 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16345), .ZN(n16337) );
  OAI21_X1 U19327 ( .B1(n16338), .B2(n16347), .A(n16337), .ZN(U243) );
  INV_X1 U19328 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16352) );
  AOI22_X1 U19329 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16343), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16340), .ZN(n16339) );
  OAI21_X1 U19330 ( .B1(n16352), .B2(U212), .A(n16339), .ZN(U244) );
  AOI22_X1 U19331 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16345), .ZN(n16341) );
  OAI21_X1 U19332 ( .B1(n16342), .B2(n16347), .A(n16341), .ZN(U245) );
  INV_X1 U19333 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16350) );
  AOI22_X1 U19334 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16343), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16340), .ZN(n16344) );
  OAI21_X1 U19335 ( .B1(n16350), .B2(U212), .A(n16344), .ZN(U246) );
  AOI22_X1 U19336 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16340), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16345), .ZN(n16346) );
  OAI21_X1 U19337 ( .B1(n16348), .B2(n16347), .A(n16346), .ZN(U247) );
  OAI22_X1 U19338 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16381), .ZN(n16349) );
  INV_X1 U19339 ( .A(n16349), .ZN(U251) );
  INV_X1 U19340 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18068) );
  AOI22_X1 U19341 ( .A1(n16381), .A2(n16350), .B1(n18068), .B2(U215), .ZN(U252) );
  INV_X1 U19342 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16351) );
  AOI22_X1 U19343 ( .A1(n16381), .A2(n16351), .B1(n18071), .B2(U215), .ZN(U253) );
  INV_X1 U19344 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18075) );
  AOI22_X1 U19345 ( .A1(n16381), .A2(n16352), .B1(n18075), .B2(U215), .ZN(U254) );
  INV_X1 U19346 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16353) );
  INV_X1 U19347 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18080) );
  AOI22_X1 U19348 ( .A1(n16381), .A2(n16353), .B1(n18080), .B2(U215), .ZN(U255) );
  INV_X1 U19349 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18084) );
  AOI22_X1 U19350 ( .A1(n16381), .A2(n16354), .B1(n18084), .B2(U215), .ZN(U256) );
  INV_X1 U19351 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16355) );
  INV_X1 U19352 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18088) );
  AOI22_X1 U19353 ( .A1(n16376), .A2(n16355), .B1(n18088), .B2(U215), .ZN(U257) );
  OAI22_X1 U19354 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16376), .ZN(n16356) );
  INV_X1 U19355 ( .A(n16356), .ZN(U258) );
  OAI22_X1 U19356 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16376), .ZN(n16357) );
  INV_X1 U19357 ( .A(n16357), .ZN(U259) );
  INV_X1 U19358 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16358) );
  INV_X1 U19359 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17347) );
  AOI22_X1 U19360 ( .A1(n16376), .A2(n16358), .B1(n17347), .B2(U215), .ZN(U260) );
  INV_X1 U19361 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16359) );
  INV_X1 U19362 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17349) );
  AOI22_X1 U19363 ( .A1(n16381), .A2(n16359), .B1(n17349), .B2(U215), .ZN(U261) );
  INV_X1 U19364 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16360) );
  INV_X1 U19365 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17351) );
  AOI22_X1 U19366 ( .A1(n16381), .A2(n16360), .B1(n17351), .B2(U215), .ZN(U262) );
  INV_X1 U19367 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16361) );
  INV_X1 U19368 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U19369 ( .A1(n16381), .A2(n16361), .B1(n17353), .B2(U215), .ZN(U263) );
  INV_X1 U19370 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17358) );
  AOI22_X1 U19371 ( .A1(n16381), .A2(n16362), .B1(n17358), .B2(U215), .ZN(U264) );
  OAI22_X1 U19372 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16381), .ZN(n16363) );
  INV_X1 U19373 ( .A(n16363), .ZN(U265) );
  OAI22_X1 U19374 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16381), .ZN(n16364) );
  INV_X1 U19375 ( .A(n16364), .ZN(U266) );
  OAI22_X1 U19376 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16381), .ZN(n16365) );
  INV_X1 U19377 ( .A(n16365), .ZN(U267) );
  OAI22_X1 U19378 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16381), .ZN(n16366) );
  INV_X1 U19379 ( .A(n16366), .ZN(U268) );
  INV_X1 U19380 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n16367) );
  INV_X1 U19381 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n20907) );
  AOI22_X1 U19382 ( .A1(n16376), .A2(n16367), .B1(n20907), .B2(U215), .ZN(U269) );
  INV_X1 U19383 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n16368) );
  INV_X1 U19384 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n19129) );
  AOI22_X1 U19385 ( .A1(n16381), .A2(n16368), .B1(n19129), .B2(U215), .ZN(U270) );
  INV_X1 U19386 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16369) );
  INV_X1 U19387 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n19136) );
  AOI22_X1 U19388 ( .A1(n16376), .A2(n16369), .B1(n19136), .B2(U215), .ZN(U271) );
  INV_X1 U19389 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16370) );
  INV_X1 U19390 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n19142) );
  AOI22_X1 U19391 ( .A1(n16381), .A2(n16370), .B1(n19142), .B2(U215), .ZN(U272) );
  INV_X1 U19392 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16371) );
  INV_X1 U19393 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n20830) );
  AOI22_X1 U19394 ( .A1(n16376), .A2(n16371), .B1(n20830), .B2(U215), .ZN(U273) );
  OAI22_X1 U19395 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16376), .ZN(n16372) );
  INV_X1 U19396 ( .A(n16372), .ZN(U274) );
  INV_X1 U19397 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16373) );
  INV_X1 U19398 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n19104) );
  AOI22_X1 U19399 ( .A1(n16376), .A2(n16373), .B1(n19104), .B2(U215), .ZN(U275) );
  INV_X1 U19400 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n16374) );
  INV_X1 U19401 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n19117) );
  AOI22_X1 U19402 ( .A1(n16381), .A2(n16374), .B1(n19117), .B2(U215), .ZN(U276) );
  INV_X1 U19403 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n16375) );
  AOI22_X1 U19404 ( .A1(n16381), .A2(n16375), .B1(n14960), .B2(U215), .ZN(U277) );
  OAI22_X1 U19405 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16376), .ZN(n16377) );
  INV_X1 U19406 ( .A(n16377), .ZN(U278) );
  INV_X1 U19407 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n20929) );
  INV_X1 U19408 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18079) );
  AOI22_X1 U19409 ( .A1(n16381), .A2(n20929), .B1(n18079), .B2(U215), .ZN(U279) );
  OAI22_X1 U19410 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16381), .ZN(n16378) );
  INV_X1 U19411 ( .A(n16378), .ZN(U280) );
  INV_X1 U19412 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n16379) );
  INV_X1 U19413 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19149) );
  AOI22_X1 U19414 ( .A1(n16381), .A2(n16379), .B1(n19149), .B2(U215), .ZN(U281) );
  INV_X1 U19415 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n16380) );
  AOI22_X1 U19416 ( .A1(n16381), .A2(n19013), .B1(n16380), .B2(U215), .ZN(U282) );
  INV_X1 U19417 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17253) );
  AOI222_X1 U19418 ( .A1(n16382), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19013), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17253), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16383) );
  INV_X2 U19419 ( .A(n16385), .ZN(n16384) );
  INV_X1 U19420 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18609) );
  AOI22_X1 U19421 ( .A1(n16384), .A2(n18609), .B1(n19786), .B2(n16385), .ZN(
        U347) );
  INV_X1 U19422 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18607) );
  INV_X1 U19423 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19785) );
  AOI22_X1 U19424 ( .A1(n16383), .A2(n18607), .B1(n19785), .B2(n16385), .ZN(
        U348) );
  INV_X1 U19425 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18605) );
  INV_X1 U19426 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19784) );
  AOI22_X1 U19427 ( .A1(n16384), .A2(n18605), .B1(n19784), .B2(n16385), .ZN(
        U349) );
  INV_X1 U19428 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18603) );
  INV_X1 U19429 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19783) );
  AOI22_X1 U19430 ( .A1(n16384), .A2(n18603), .B1(n19783), .B2(n16385), .ZN(
        U350) );
  INV_X1 U19431 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18601) );
  INV_X1 U19432 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19782) );
  AOI22_X1 U19433 ( .A1(n16384), .A2(n18601), .B1(n19782), .B2(n16385), .ZN(
        U351) );
  INV_X1 U19434 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18599) );
  INV_X1 U19435 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19781) );
  AOI22_X1 U19436 ( .A1(n16384), .A2(n18599), .B1(n19781), .B2(n16385), .ZN(
        U352) );
  INV_X1 U19437 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18597) );
  INV_X1 U19438 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19780) );
  AOI22_X1 U19439 ( .A1(n16384), .A2(n18597), .B1(n19780), .B2(n16385), .ZN(
        U353) );
  INV_X1 U19440 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18595) );
  INV_X1 U19441 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19779) );
  AOI22_X1 U19442 ( .A1(n16384), .A2(n18595), .B1(n19779), .B2(n16385), .ZN(
        U354) );
  INV_X1 U19443 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18650) );
  INV_X1 U19444 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19819) );
  AOI22_X1 U19445 ( .A1(n16384), .A2(n18650), .B1(n19819), .B2(n16385), .ZN(
        U355) );
  INV_X1 U19446 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18648) );
  INV_X1 U19447 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19816) );
  AOI22_X1 U19448 ( .A1(n16384), .A2(n18648), .B1(n19816), .B2(n16385), .ZN(
        U356) );
  INV_X1 U19449 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18645) );
  INV_X1 U19450 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19814) );
  AOI22_X1 U19451 ( .A1(n16384), .A2(n18645), .B1(n19814), .B2(n16385), .ZN(
        U357) );
  INV_X1 U19452 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18644) );
  INV_X1 U19453 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19810) );
  AOI22_X1 U19454 ( .A1(n16384), .A2(n18644), .B1(n19810), .B2(n16385), .ZN(
        U358) );
  INV_X1 U19455 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18642) );
  INV_X1 U19456 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19809) );
  AOI22_X1 U19457 ( .A1(n16384), .A2(n18642), .B1(n19809), .B2(n16385), .ZN(
        U359) );
  INV_X1 U19458 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18640) );
  INV_X1 U19459 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19807) );
  AOI22_X1 U19460 ( .A1(n16384), .A2(n18640), .B1(n19807), .B2(n16385), .ZN(
        U360) );
  INV_X1 U19461 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18637) );
  INV_X1 U19462 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19805) );
  AOI22_X1 U19463 ( .A1(n16384), .A2(n18637), .B1(n19805), .B2(n16385), .ZN(
        U361) );
  INV_X1 U19464 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18635) );
  INV_X1 U19465 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19803) );
  AOI22_X1 U19466 ( .A1(n16384), .A2(n18635), .B1(n19803), .B2(n16385), .ZN(
        U362) );
  INV_X1 U19467 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18633) );
  INV_X1 U19468 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19801) );
  AOI22_X1 U19469 ( .A1(n16384), .A2(n18633), .B1(n19801), .B2(n16385), .ZN(
        U363) );
  INV_X1 U19470 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18631) );
  INV_X1 U19471 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19800) );
  AOI22_X1 U19472 ( .A1(n16384), .A2(n18631), .B1(n19800), .B2(n16385), .ZN(
        U364) );
  INV_X1 U19473 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18593) );
  INV_X1 U19474 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19778) );
  AOI22_X1 U19475 ( .A1(n16384), .A2(n18593), .B1(n19778), .B2(n16385), .ZN(
        U365) );
  INV_X1 U19476 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18629) );
  INV_X1 U19477 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19798) );
  AOI22_X1 U19478 ( .A1(n16384), .A2(n18629), .B1(n19798), .B2(n16385), .ZN(
        U366) );
  INV_X1 U19479 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18627) );
  INV_X1 U19480 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19797) );
  AOI22_X1 U19481 ( .A1(n16384), .A2(n18627), .B1(n19797), .B2(n16385), .ZN(
        U367) );
  INV_X1 U19482 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18625) );
  INV_X1 U19483 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19795) );
  AOI22_X1 U19484 ( .A1(n16384), .A2(n18625), .B1(n19795), .B2(n16385), .ZN(
        U368) );
  INV_X1 U19485 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18622) );
  INV_X1 U19486 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19793) );
  AOI22_X1 U19487 ( .A1(n16384), .A2(n18622), .B1(n19793), .B2(n16385), .ZN(
        U369) );
  INV_X1 U19488 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18621) );
  INV_X1 U19489 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19792) );
  AOI22_X1 U19490 ( .A1(n16384), .A2(n18621), .B1(n19792), .B2(n16385), .ZN(
        U370) );
  INV_X1 U19491 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18619) );
  INV_X1 U19492 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19791) );
  AOI22_X1 U19493 ( .A1(n16383), .A2(n18619), .B1(n19791), .B2(n16385), .ZN(
        U371) );
  INV_X1 U19494 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18617) );
  INV_X1 U19495 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19790) );
  AOI22_X1 U19496 ( .A1(n16383), .A2(n18617), .B1(n19790), .B2(n16385), .ZN(
        U372) );
  INV_X1 U19497 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18615) );
  INV_X1 U19498 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19789) );
  AOI22_X1 U19499 ( .A1(n16384), .A2(n18615), .B1(n19789), .B2(n16385), .ZN(
        U373) );
  INV_X1 U19500 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18613) );
  INV_X1 U19501 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19788) );
  AOI22_X1 U19502 ( .A1(n16384), .A2(n18613), .B1(n19788), .B2(n16385), .ZN(
        U374) );
  INV_X1 U19503 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18611) );
  INV_X1 U19504 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19787) );
  AOI22_X1 U19505 ( .A1(n16383), .A2(n18611), .B1(n19787), .B2(n16385), .ZN(
        U375) );
  INV_X1 U19506 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18592) );
  INV_X1 U19507 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19775) );
  AOI22_X1 U19508 ( .A1(n16384), .A2(n18592), .B1(n19775), .B2(n16385), .ZN(
        U376) );
  INV_X1 U19509 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16386) );
  AND2_X1 U19510 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18591), .ZN(n18581) );
  OAI21_X1 U19511 ( .B1(n18589), .B2(n18581), .A(n18725), .ZN(n18660) );
  INV_X1 U19512 ( .A(n18660), .ZN(n18664) );
  OAI21_X1 U19513 ( .B1(n16386), .B2(n18589), .A(n18575), .ZN(P3_U2633) );
  OAI21_X1 U19514 ( .B1(n16387), .B2(n17305), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16388) );
  OAI21_X1 U19515 ( .B1(n16389), .B2(n18566), .A(n16388), .ZN(P3_U2634) );
  AOI21_X1 U19516 ( .B1(n18589), .B2(n18591), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16390) );
  AOI22_X1 U19517 ( .A1(n18658), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16390), 
        .B2(n18725), .ZN(P3_U2635) );
  NOR2_X1 U19518 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18576) );
  OAI21_X1 U19519 ( .B1(n18576), .B2(BS16), .A(n18664), .ZN(n18662) );
  OAI21_X1 U19520 ( .B1(n18664), .B2(n18715), .A(n18662), .ZN(P3_U2636) );
  AND3_X1 U19521 ( .A1(n18498), .A2(n16392), .A3(n16391), .ZN(n18501) );
  NOR2_X1 U19522 ( .A1(n18501), .A2(n18561), .ZN(n18708) );
  OAI21_X1 U19523 ( .B1(n18708), .B2(n18054), .A(n16393), .ZN(P3_U2637) );
  NOR4_X1 U19524 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16397) );
  NOR4_X1 U19525 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16396) );
  NOR4_X1 U19526 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16395) );
  NOR4_X1 U19527 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16394) );
  NAND4_X1 U19528 ( .A1(n16397), .A2(n16396), .A3(n16395), .A4(n16394), .ZN(
        n16403) );
  NOR4_X1 U19529 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16401) );
  AOI211_X1 U19530 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16400) );
  NOR4_X1 U19531 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16399) );
  NOR4_X1 U19532 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16398) );
  NAND4_X1 U19533 ( .A1(n16401), .A2(n16400), .A3(n16399), .A4(n16398), .ZN(
        n16402) );
  NOR2_X1 U19534 ( .A1(n16403), .A2(n16402), .ZN(n18702) );
  INV_X1 U19535 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20862) );
  NOR3_X1 U19536 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16405) );
  OAI21_X1 U19537 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16405), .A(n18702), .ZN(
        n16404) );
  OAI21_X1 U19538 ( .B1(n18702), .B2(n20862), .A(n16404), .ZN(P3_U2638) );
  INV_X1 U19539 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18698) );
  INV_X1 U19540 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18663) );
  AOI21_X1 U19541 ( .B1(n18698), .B2(n18663), .A(n16405), .ZN(n16406) );
  INV_X1 U19542 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18654) );
  INV_X1 U19543 ( .A(n18702), .ZN(n18705) );
  AOI22_X1 U19544 ( .A1(n18702), .A2(n16406), .B1(n18654), .B2(n18705), .ZN(
        P3_U2639) );
  NOR4_X4 U19545 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n18675), .ZN(n16739) );
  NOR2_X1 U19546 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18667), .ZN(n18564) );
  OR2_X1 U19547 ( .A1(n18566), .A2(n18433), .ZN(n18559) );
  AOI211_X1 U19548 ( .C1(n18716), .C2(n18714), .A(n18578), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16408) );
  AOI211_X4 U19549 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n16410), .A(n16408), .B(
        n16412), .ZN(n16768) );
  INV_X1 U19550 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18651) );
  INV_X1 U19551 ( .A(n16408), .ZN(n18554) );
  INV_X1 U19552 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18636) );
  INV_X1 U19553 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18632) );
  INV_X1 U19554 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18630) );
  INV_X1 U19555 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18623) );
  INV_X1 U19556 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18620) );
  INV_X1 U19557 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18616) );
  INV_X1 U19558 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18614) );
  INV_X1 U19559 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18610) );
  INV_X1 U19560 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18606) );
  INV_X1 U19561 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18602) );
  INV_X1 U19562 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18598) );
  INV_X1 U19563 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18594) );
  NAND2_X1 U19564 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n16764) );
  NOR2_X1 U19565 ( .A1(n18594), .A2(n16764), .ZN(n16727) );
  NAND2_X1 U19566 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16727), .ZN(n16713) );
  NOR2_X1 U19567 ( .A1(n18598), .A2(n16713), .ZN(n16686) );
  NAND2_X1 U19568 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16686), .ZN(n16692) );
  NOR2_X1 U19569 ( .A1(n18602), .A2(n16692), .ZN(n16672) );
  NAND2_X1 U19570 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16672), .ZN(n16651) );
  NOR2_X1 U19571 ( .A1(n18606), .A2(n16651), .ZN(n16650) );
  NAND2_X1 U19572 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n16650), .ZN(n16637) );
  NOR2_X1 U19573 ( .A1(n18610), .A2(n16637), .ZN(n16626) );
  NAND2_X1 U19574 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16626), .ZN(n16600) );
  NOR3_X1 U19575 ( .A1(n18616), .A2(n18614), .A3(n16600), .ZN(n16580) );
  NAND2_X1 U19576 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16580), .ZN(n16564) );
  NOR3_X1 U19577 ( .A1(n18623), .A2(n18620), .A3(n16564), .ZN(n16546) );
  NAND4_X1 U19578 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16546), .A3(
        P3_REIP_REG_19__SCAN_IN), .A4(P3_REIP_REG_18__SCAN_IN), .ZN(n16517) );
  NOR3_X1 U19579 ( .A1(n18632), .A2(n18630), .A3(n16517), .ZN(n16503) );
  NAND2_X1 U19580 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16503), .ZN(n16499) );
  NOR2_X1 U19581 ( .A1(n18636), .A2(n16499), .ZN(n16471) );
  NAND3_X1 U19582 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n16471), .ZN(n16425) );
  NAND4_X1 U19583 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16466), .ZN(n16427) );
  NOR3_X1 U19584 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18651), .A3(n16427), 
        .ZN(n16409) );
  AOI21_X1 U19585 ( .B1(n16768), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16409), .ZN(
        n16432) );
  NAND2_X1 U19586 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n16410), .ZN(n16411) );
  AOI211_X4 U19587 ( .C1(n18715), .C2(n18717), .A(n16412), .B(n16411), .ZN(
        n16748) );
  NOR3_X1 U19588 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16755) );
  NAND2_X1 U19589 ( .A1(n16755), .A2(n16749), .ZN(n16747) );
  NOR2_X1 U19590 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16747), .ZN(n16728) );
  INV_X1 U19591 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16721) );
  NAND2_X1 U19592 ( .A1(n16728), .A2(n16721), .ZN(n16714) );
  NAND2_X1 U19593 ( .A1(n16705), .A2(n17007), .ZN(n16696) );
  NAND2_X1 U19594 ( .A1(n16671), .A2(n17031), .ZN(n16667) );
  NAND2_X1 U19595 ( .A1(n16647), .A2(n16638), .ZN(n16641) );
  INV_X1 U19596 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16990) );
  NAND2_X1 U19597 ( .A1(n16623), .A2(n16990), .ZN(n16612) );
  INV_X1 U19598 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20894) );
  NAND2_X1 U19599 ( .A1(n16599), .A2(n20894), .ZN(n16589) );
  NAND2_X1 U19600 ( .A1(n16577), .A2(n16574), .ZN(n16573) );
  NAND2_X1 U19601 ( .A1(n16557), .A2(n16552), .ZN(n16551) );
  INV_X1 U19602 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20835) );
  NAND2_X1 U19603 ( .A1(n16533), .A2(n20835), .ZN(n16529) );
  INV_X1 U19604 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16509) );
  NAND2_X1 U19605 ( .A1(n16514), .A2(n16509), .ZN(n16508) );
  INV_X1 U19606 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16487) );
  NAND2_X1 U19607 ( .A1(n16491), .A2(n16487), .ZN(n16486) );
  NOR2_X1 U19608 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16486), .ZN(n16474) );
  NAND2_X1 U19609 ( .A1(n16474), .A2(n16795), .ZN(n16467) );
  NOR2_X1 U19610 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16467), .ZN(n16452) );
  INV_X1 U19611 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n20915) );
  NAND2_X1 U19612 ( .A1(n16452), .A2(n20915), .ZN(n16433) );
  NOR2_X1 U19613 ( .A1(n16784), .A2(n16433), .ZN(n16438) );
  INV_X1 U19614 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16800) );
  NOR2_X1 U19615 ( .A1(n17728), .A2(n17366), .ZN(n16414) );
  OAI21_X1 U19616 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16414), .A(
        n16413), .ZN(n17373) );
  INV_X1 U19617 ( .A(n17373), .ZN(n16455) );
  INV_X1 U19618 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17367) );
  NOR2_X1 U19619 ( .A1(n17728), .A2(n9917), .ZN(n16419) );
  NAND3_X1 U19620 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(n16419), .ZN(n17370) );
  NOR2_X1 U19621 ( .A1(n17396), .A2(n17370), .ZN(n16416) );
  INV_X1 U19622 ( .A(n16416), .ZN(n16415) );
  AOI21_X1 U19623 ( .B1(n17367), .B2(n16415), .A(n16414), .ZN(n17386) );
  AOI21_X1 U19624 ( .B1(n17396), .B2(n17370), .A(n16416), .ZN(n17399) );
  INV_X1 U19625 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17421) );
  INV_X1 U19626 ( .A(n16419), .ZN(n16418) );
  NOR2_X1 U19627 ( .A1(n17421), .A2(n16418), .ZN(n16417) );
  OAI21_X1 U19628 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16417), .A(
        n17370), .ZN(n17409) );
  INV_X1 U19629 ( .A(n17409), .ZN(n16482) );
  AOI21_X1 U19630 ( .B1(n17421), .B2(n16418), .A(n16417), .ZN(n17419) );
  NAND2_X1 U19631 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9705), .ZN(
        n17407) );
  AOI21_X1 U19632 ( .B1(n17437), .B2(n17407), .A(n16419), .ZN(n17434) );
  INV_X1 U19633 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17460) );
  INV_X1 U19634 ( .A(n16420), .ZN(n17481) );
  NAND2_X1 U19635 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17481), .ZN(
        n17443) );
  NOR2_X1 U19636 ( .A1(n17445), .A2(n17443), .ZN(n16423) );
  NAND2_X1 U19637 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16423), .ZN(
        n16422) );
  INV_X1 U19638 ( .A(n17407), .ZN(n16421) );
  AOI21_X1 U19639 ( .B1(n17460), .B2(n16422), .A(n16421), .ZN(n17449) );
  INV_X1 U19640 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17462) );
  XNOR2_X1 U19641 ( .A(n17462), .B(n16423), .ZN(n17465) );
  AOI21_X1 U19642 ( .B1(n17445), .B2(n17443), .A(n16423), .ZN(n17483) );
  INV_X1 U19643 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17542) );
  INV_X1 U19644 ( .A(n16424), .ZN(n17526) );
  NOR2_X1 U19645 ( .A1(n17728), .A2(n17526), .ZN(n17524) );
  INV_X1 U19646 ( .A(n17524), .ZN(n16544) );
  NOR2_X1 U19647 ( .A1(n17542), .A2(n16544), .ZN(n16567) );
  INV_X1 U19648 ( .A(n16567), .ZN(n16588) );
  NOR2_X1 U19649 ( .A1(n17465), .A2(n16525), .ZN(n16524) );
  NOR2_X1 U19650 ( .A1(n16524), .A2(n16738), .ZN(n16516) );
  NOR2_X1 U19651 ( .A1(n17449), .A2(n16516), .ZN(n16515) );
  NOR2_X1 U19652 ( .A1(n16515), .A2(n16738), .ZN(n16502) );
  NOR2_X1 U19653 ( .A1(n17434), .A2(n16502), .ZN(n16501) );
  NOR2_X1 U19654 ( .A1(n16481), .A2(n16738), .ZN(n16473) );
  NOR2_X1 U19655 ( .A1(n17399), .A2(n16473), .ZN(n16472) );
  NOR2_X1 U19656 ( .A1(n16472), .A2(n16738), .ZN(n16463) );
  NOR2_X1 U19657 ( .A1(n17386), .A2(n16463), .ZN(n16462) );
  NOR2_X1 U19658 ( .A1(n16462), .A2(n16738), .ZN(n16454) );
  NOR2_X1 U19659 ( .A1(n16455), .A2(n16454), .ZN(n16453) );
  NOR2_X1 U19660 ( .A1(n16453), .A2(n16738), .ZN(n16442) );
  NAND2_X1 U19661 ( .A1(n16723), .A2(n16739), .ZN(n16775) );
  NOR3_X1 U19662 ( .A1(n16435), .A2(n16434), .A3(n16775), .ZN(n16430) );
  NAND3_X1 U19663 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16426) );
  INV_X1 U19664 ( .A(n16782), .ZN(n16787) );
  AOI21_X1 U19665 ( .B1(n16425), .B2(n16763), .A(n16787), .ZN(n16470) );
  INV_X1 U19666 ( .A(n16470), .ZN(n16478) );
  AOI21_X1 U19667 ( .B1(n16763), .B2(n16426), .A(n16478), .ZN(n16451) );
  NOR2_X1 U19668 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16427), .ZN(n16437) );
  INV_X1 U19669 ( .A(n16437), .ZN(n16428) );
  AOI21_X1 U19670 ( .B1(n16451), .B2(n16428), .A(n18649), .ZN(n16429) );
  OAI211_X1 U19671 ( .C1(n12693), .C2(n16774), .A(n16432), .B(n16431), .ZN(
        P3_U2640) );
  NAND2_X1 U19672 ( .A1(n16748), .A2(n16433), .ZN(n16447) );
  OAI22_X1 U19673 ( .A1(n16451), .A2(n18651), .B1(n9924), .B2(n16774), .ZN(
        n16436) );
  OAI21_X1 U19674 ( .B1(n16768), .B2(n16438), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16439) );
  OAI211_X1 U19675 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16447), .A(n16440), .B(
        n16439), .ZN(P3_U2641) );
  INV_X1 U19676 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18647) );
  AOI211_X1 U19677 ( .C1(n16443), .C2(n16442), .A(n16441), .B(n18569), .ZN(
        n16446) );
  NAND3_X1 U19678 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16466), .ZN(n16444) );
  OAI22_X1 U19679 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16444), .B1(n9923), 
        .B2(n16774), .ZN(n16445) );
  AOI211_X1 U19680 ( .C1(n16768), .C2(P3_EBX_REG_29__SCAN_IN), .A(n16446), .B(
        n16445), .ZN(n16450) );
  INV_X1 U19681 ( .A(n16447), .ZN(n16448) );
  OAI21_X1 U19682 ( .B1(n16452), .B2(n20915), .A(n16448), .ZN(n16449) );
  OAI211_X1 U19683 ( .C1(n16451), .C2(n18647), .A(n16450), .B(n16449), .ZN(
        P3_U2642) );
  AOI22_X1 U19684 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16759), .B1(
        n16768), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16461) );
  AOI211_X1 U19685 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16467), .A(n16452), .B(
        n16784), .ZN(n16457) );
  AOI211_X1 U19686 ( .C1(n16455), .C2(n16454), .A(n16453), .B(n18569), .ZN(
        n16456) );
  AOI211_X1 U19687 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16478), .A(n16457), 
        .B(n16456), .ZN(n16460) );
  NAND2_X1 U19688 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16458) );
  OAI211_X1 U19689 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16466), .B(n16458), .ZN(n16459) );
  NAND3_X1 U19690 ( .A1(n16461), .A2(n16460), .A3(n16459), .ZN(P3_U2643) );
  INV_X1 U19691 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18643) );
  AOI211_X1 U19692 ( .C1(n17386), .C2(n16463), .A(n16462), .B(n18569), .ZN(
        n16465) );
  OAI22_X1 U19693 ( .A1(n17367), .A2(n16774), .B1(n16785), .B2(n16795), .ZN(
        n16464) );
  AOI211_X1 U19694 ( .C1(n16466), .C2(n18643), .A(n16465), .B(n16464), .ZN(
        n16469) );
  OAI211_X1 U19695 ( .C1(n16474), .C2(n16795), .A(n16748), .B(n16467), .ZN(
        n16468) );
  OAI211_X1 U19696 ( .C1(n16470), .C2(n18643), .A(n16469), .B(n16468), .ZN(
        P3_U2644) );
  AOI22_X1 U19697 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16759), .B1(
        n16768), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16480) );
  INV_X1 U19698 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18639) );
  NAND2_X1 U19699 ( .A1(n16763), .A2(n16471), .ZN(n16483) );
  INV_X1 U19700 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18641) );
  OAI21_X1 U19701 ( .B1(n18639), .B2(n16483), .A(n18641), .ZN(n16477) );
  AOI211_X1 U19702 ( .C1(n17399), .C2(n16473), .A(n16472), .B(n18569), .ZN(
        n16476) );
  AOI211_X1 U19703 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16486), .A(n16474), .B(
        n16784), .ZN(n16475) );
  AOI211_X1 U19704 ( .C1(n16478), .C2(n16477), .A(n16476), .B(n16475), .ZN(
        n16479) );
  NAND2_X1 U19705 ( .A1(n16480), .A2(n16479), .ZN(P3_U2645) );
  NAND2_X1 U19706 ( .A1(n16763), .A2(n16499), .ZN(n16504) );
  NAND2_X1 U19707 ( .A1(n16782), .A2(n16504), .ZN(n16500) );
  AOI21_X1 U19708 ( .B1(n16763), .B2(n18636), .A(n16500), .ZN(n16490) );
  AOI211_X1 U19709 ( .C1(n16482), .C2(n9707), .A(n16481), .B(n18569), .ZN(
        n16485) );
  OAI22_X1 U19710 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16483), .B1(n16487), 
        .B2(n16785), .ZN(n16484) );
  AOI211_X1 U19711 ( .C1(n16759), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16485), .B(n16484), .ZN(n16489) );
  OAI211_X1 U19712 ( .C1(n16491), .C2(n16487), .A(n16748), .B(n16486), .ZN(
        n16488) );
  OAI211_X1 U19713 ( .C1(n16490), .C2(n18639), .A(n16489), .B(n16488), .ZN(
        P3_U2646) );
  NAND2_X1 U19714 ( .A1(n16763), .A2(n18636), .ZN(n16498) );
  AOI22_X1 U19715 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16759), .B1(
        n16768), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n16497) );
  AOI211_X1 U19716 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16508), .A(n16491), .B(
        n16784), .ZN(n16495) );
  AOI211_X1 U19717 ( .C1(n17419), .C2(n16493), .A(n16492), .B(n18569), .ZN(
        n16494) );
  AOI211_X1 U19718 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16500), .A(n16495), 
        .B(n16494), .ZN(n16496) );
  OAI211_X1 U19719 ( .C1(n16499), .C2(n16498), .A(n16497), .B(n16496), .ZN(
        P3_U2647) );
  INV_X1 U19720 ( .A(n16500), .ZN(n16512) );
  INV_X1 U19721 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18634) );
  AOI211_X1 U19722 ( .C1(n17434), .C2(n16502), .A(n16501), .B(n18569), .ZN(
        n16507) );
  INV_X1 U19723 ( .A(n16503), .ZN(n16505) );
  OAI22_X1 U19724 ( .A1(n16785), .A2(n16509), .B1(n16505), .B2(n16504), .ZN(
        n16506) );
  AOI211_X1 U19725 ( .C1(n16759), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16507), .B(n16506), .ZN(n16511) );
  OAI211_X1 U19726 ( .C1(n16514), .C2(n16509), .A(n16748), .B(n16508), .ZN(
        n16510) );
  OAI211_X1 U19727 ( .C1(n16512), .C2(n18634), .A(n16511), .B(n16510), .ZN(
        P3_U2648) );
  AOI21_X1 U19728 ( .B1(n16763), .B2(n16517), .A(n16787), .ZN(n16541) );
  NOR2_X1 U19729 ( .A1(n16781), .A2(n16517), .ZN(n16513) );
  NAND2_X1 U19730 ( .A1(n16513), .A2(n18630), .ZN(n16531) );
  AOI211_X1 U19731 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16529), .A(n16514), .B(
        n16784), .ZN(n16522) );
  AOI211_X1 U19732 ( .C1(n17449), .C2(n16516), .A(n16515), .B(n18569), .ZN(
        n16521) );
  NOR4_X1 U19733 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16781), .A3(n18630), 
        .A4(n16517), .ZN(n16520) );
  OAI22_X1 U19734 ( .A1(n17460), .A2(n16774), .B1(n16785), .B2(n16518), .ZN(
        n16519) );
  NOR4_X1 U19735 ( .A1(n16522), .A2(n16521), .A3(n16520), .A4(n16519), .ZN(
        n16523) );
  OAI221_X1 U19736 ( .B1(n18632), .B2(n16541), .C1(n18632), .C2(n16531), .A(
        n16523), .ZN(P3_U2649) );
  INV_X1 U19737 ( .A(n16541), .ZN(n16528) );
  AOI211_X1 U19738 ( .C1(n17465), .C2(n16525), .A(n16524), .B(n18569), .ZN(
        n16527) );
  OAI22_X1 U19739 ( .A1(n17462), .A2(n16774), .B1(n20835), .B2(n16785), .ZN(
        n16526) );
  AOI211_X1 U19740 ( .C1(n16528), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16527), 
        .B(n16526), .ZN(n16532) );
  OAI211_X1 U19741 ( .C1(n16533), .C2(n20835), .A(n16748), .B(n16529), .ZN(
        n16530) );
  NAND3_X1 U19742 ( .A1(n16532), .A2(n16531), .A3(n16530), .ZN(P3_U2650) );
  INV_X1 U19743 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18628) );
  AOI211_X1 U19744 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16551), .A(n16533), .B(
        n16784), .ZN(n16534) );
  AOI21_X1 U19745 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16768), .A(n16534), .ZN(
        n16540) );
  AOI211_X1 U19746 ( .C1(n17483), .C2(n16536), .A(n16535), .B(n18569), .ZN(
        n16538) );
  NAND2_X1 U19747 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16542) );
  NAND2_X1 U19748 ( .A1(n16763), .A2(n16546), .ZN(n16558) );
  NOR3_X1 U19749 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16542), .A3(n16558), 
        .ZN(n16537) );
  AOI211_X1 U19750 ( .C1(n16759), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16538), .B(n16537), .ZN(n16539) );
  OAI211_X1 U19751 ( .C1(n18628), .C2(n16541), .A(n16540), .B(n16539), .ZN(
        P3_U2651) );
  INV_X1 U19752 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17491) );
  OAI21_X1 U19753 ( .B1(P3_REIP_REG_19__SCAN_IN), .B2(P3_REIP_REG_18__SCAN_IN), 
        .A(n16542), .ZN(n16543) );
  OAI22_X1 U19754 ( .A1(n16785), .A2(n16552), .B1(n16558), .B2(n16543), .ZN(
        n16550) );
  INV_X1 U19755 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17502) );
  OR2_X1 U19756 ( .A1(n17528), .A2(n16544), .ZN(n16566) );
  NOR2_X1 U19757 ( .A1(n17511), .A2(n16566), .ZN(n16565) );
  INV_X1 U19758 ( .A(n16565), .ZN(n17488) );
  NOR2_X1 U19759 ( .A1(n17502), .A2(n17488), .ZN(n16555) );
  AOI21_X1 U19760 ( .B1(n16786), .B2(n16555), .A(n16738), .ZN(n16545) );
  OAI21_X1 U19761 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16555), .A(
        n17443), .ZN(n17490) );
  XOR2_X1 U19762 ( .A(n16545), .B(n17490), .Z(n16548) );
  INV_X1 U19763 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18626) );
  INV_X1 U19764 ( .A(n16546), .ZN(n16547) );
  AOI21_X1 U19765 ( .B1(n16763), .B2(n16547), .A(n16787), .ZN(n16570) );
  OAI22_X1 U19766 ( .A1(n18569), .A2(n16548), .B1(n18626), .B2(n16570), .ZN(
        n16549) );
  NOR3_X1 U19767 ( .A1(n18038), .A2(n16550), .A3(n16549), .ZN(n16554) );
  OAI211_X1 U19768 ( .C1(n16557), .C2(n16552), .A(n16748), .B(n16551), .ZN(
        n16553) );
  OAI211_X1 U19769 ( .C1(n16774), .C2(n17491), .A(n16554), .B(n16553), .ZN(
        P3_U2652) );
  INV_X1 U19770 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18624) );
  AOI22_X1 U19771 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16759), .B1(
        n16768), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n16563) );
  AOI21_X1 U19772 ( .B1(n17502), .B2(n17488), .A(n16555), .ZN(n17505) );
  NOR2_X1 U19773 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17728), .ZN(
        n16673) );
  AOI21_X1 U19774 ( .B1(n17487), .B2(n16673), .A(n16738), .ZN(n16556) );
  XOR2_X1 U19775 ( .A(n17505), .B(n16556), .Z(n16561) );
  AOI211_X1 U19776 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16573), .A(n16557), .B(
        n16784), .ZN(n16560) );
  OAI21_X1 U19777 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16558), .A(n18048), 
        .ZN(n16559) );
  AOI211_X1 U19778 ( .C1(n16561), .C2(n16739), .A(n16560), .B(n16559), .ZN(
        n16562) );
  OAI211_X1 U19779 ( .C1(n18624), .C2(n16570), .A(n16563), .B(n16562), .ZN(
        P3_U2653) );
  NOR2_X1 U19780 ( .A1(n16781), .A2(n16564), .ZN(n16579) );
  AOI21_X1 U19781 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n16579), .A(
        P3_REIP_REG_17__SCAN_IN), .ZN(n16571) );
  AOI21_X1 U19782 ( .B1(n17511), .B2(n16566), .A(n16565), .ZN(n17516) );
  OAI21_X1 U19783 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16567), .A(
        n16566), .ZN(n16581) );
  INV_X1 U19784 ( .A(n16581), .ZN(n17525) );
  OAI21_X1 U19785 ( .B1(n16595), .B2(n17525), .A(n16723), .ZN(n16568) );
  XOR2_X1 U19786 ( .A(n17516), .B(n16568), .Z(n16569) );
  OAI22_X1 U19787 ( .A1(n16571), .A2(n16570), .B1(n18569), .B2(n16569), .ZN(
        n16572) );
  AOI211_X1 U19788 ( .C1(n16768), .C2(P3_EBX_REG_17__SCAN_IN), .A(n18038), .B(
        n16572), .ZN(n16576) );
  OAI211_X1 U19789 ( .C1(n16577), .C2(n16574), .A(n16748), .B(n16573), .ZN(
        n16575) );
  OAI211_X1 U19790 ( .C1(n16774), .C2(n17511), .A(n16576), .B(n16575), .ZN(
        P3_U2654) );
  AOI22_X1 U19791 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16759), .B1(
        n16768), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n16586) );
  AOI211_X1 U19792 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16589), .A(n16577), .B(
        n16784), .ZN(n16578) );
  AOI211_X1 U19793 ( .C1(n16579), .C2(n18620), .A(n18038), .B(n16578), .ZN(
        n16585) );
  OAI21_X1 U19794 ( .B1(n16580), .B2(n16781), .A(n16782), .ZN(n16591) );
  INV_X1 U19795 ( .A(n16580), .ZN(n16601) );
  NOR3_X1 U19796 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16781), .A3(n16601), 
        .ZN(n16594) );
  OAI21_X1 U19797 ( .B1(n16591), .B2(n16594), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n16584) );
  OAI221_X1 U19798 ( .B1(n16595), .B2(n17525), .C1(n16582), .C2(n16581), .A(
        n16739), .ZN(n16583) );
  NAND4_X1 U19799 ( .A1(n16586), .A2(n16585), .A3(n16584), .A4(n16583), .ZN(
        P3_U2655) );
  NOR2_X1 U19800 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18569), .ZN(
        n16587) );
  NOR2_X1 U19801 ( .A1(n16723), .A2(n18569), .ZN(n16754) );
  AOI21_X1 U19802 ( .B1(n16587), .B2(n17542), .A(n16754), .ZN(n16598) );
  OAI21_X1 U19803 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17524), .A(
        n16588), .ZN(n17539) );
  OAI211_X1 U19804 ( .C1(n16599), .C2(n20894), .A(n16748), .B(n16589), .ZN(
        n16590) );
  OAI211_X1 U19805 ( .C1(n20894), .C2(n16785), .A(n18048), .B(n16590), .ZN(
        n16593) );
  INV_X1 U19806 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18618) );
  INV_X1 U19807 ( .A(n16591), .ZN(n16609) );
  OAI22_X1 U19808 ( .A1(n17542), .A2(n16774), .B1(n18618), .B2(n16609), .ZN(
        n16592) );
  NOR3_X1 U19809 ( .A1(n16594), .A2(n16593), .A3(n16592), .ZN(n16597) );
  NAND3_X1 U19810 ( .A1(n16595), .A2(n16739), .A3(n17539), .ZN(n16596) );
  OAI211_X1 U19811 ( .C1(n16598), .C2(n17539), .A(n16597), .B(n16596), .ZN(
        P3_U2656) );
  AOI211_X1 U19812 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16612), .A(n16599), .B(
        n16784), .ZN(n16604) );
  NOR2_X1 U19813 ( .A1(n16781), .A2(n16600), .ZN(n16618) );
  NAND3_X1 U19814 ( .A1(n16601), .A2(n16618), .A3(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n16602) );
  OAI211_X1 U19815 ( .C1(n17551), .C2(n16774), .A(n18048), .B(n16602), .ZN(
        n16603) );
  AOI211_X1 U19816 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16768), .A(n16604), .B(
        n16603), .ZN(n16608) );
  NOR3_X1 U19817 ( .A1(n17728), .A2(n16634), .A3(n17596), .ZN(n17565) );
  NAND3_X1 U19818 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A3(n17565), .ZN(n16610) );
  AOI21_X1 U19819 ( .B1(n17551), .B2(n16610), .A(n17524), .ZN(n17554) );
  INV_X1 U19820 ( .A(n16673), .ZN(n16761) );
  OAI21_X1 U19821 ( .B1(n17552), .B2(n16761), .A(n16723), .ZN(n16605) );
  INV_X1 U19822 ( .A(n16605), .ZN(n16619) );
  INV_X1 U19823 ( .A(n17554), .ZN(n16606) );
  OAI221_X1 U19824 ( .B1(n17554), .B2(n16619), .C1(n16606), .C2(n16605), .A(
        n16739), .ZN(n16607) );
  OAI211_X1 U19825 ( .C1(n16609), .C2(n18616), .A(n16608), .B(n16607), .ZN(
        P3_U2657) );
  INV_X1 U19826 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16628) );
  INV_X1 U19827 ( .A(n17565), .ZN(n16635) );
  NOR2_X1 U19828 ( .A1(n16628), .A2(n16635), .ZN(n16627) );
  OAI21_X1 U19829 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16627), .A(
        n16610), .ZN(n17567) );
  AOI21_X1 U19830 ( .B1(n16723), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18569), .ZN(n16777) );
  OAI21_X1 U19831 ( .B1(n16627), .B2(n16754), .A(n16777), .ZN(n16622) );
  OAI21_X1 U19832 ( .B1(n16626), .B2(n16781), .A(n16782), .ZN(n16643) );
  INV_X1 U19833 ( .A(n16643), .ZN(n16611) );
  OAI21_X1 U19834 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n16781), .A(n16611), 
        .ZN(n16617) );
  INV_X1 U19835 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16615) );
  AOI21_X1 U19836 ( .B1(n16768), .B2(P3_EBX_REG_13__SCAN_IN), .A(n18038), .ZN(
        n16614) );
  OAI211_X1 U19837 ( .C1(n16623), .C2(n16990), .A(n16748), .B(n16612), .ZN(
        n16613) );
  OAI211_X1 U19838 ( .C1(n16774), .C2(n16615), .A(n16614), .B(n16613), .ZN(
        n16616) );
  AOI221_X1 U19839 ( .B1(n16618), .B2(n18614), .C1(n16617), .C2(
        P3_REIP_REG_13__SCAN_IN), .A(n16616), .ZN(n16621) );
  NAND3_X1 U19840 ( .A1(n16739), .A2(n16619), .A3(n17567), .ZN(n16620) );
  OAI211_X1 U19841 ( .C1(n17567), .C2(n16622), .A(n16621), .B(n16620), .ZN(
        P3_U2658) );
  AOI211_X1 U19842 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16641), .A(n16623), .B(
        n16784), .ZN(n16624) );
  AOI21_X1 U19843 ( .B1(n16759), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16624), .ZN(n16633) );
  NOR2_X1 U19844 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16781), .ZN(n16625) );
  AOI22_X1 U19845 ( .A1(n16768), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n16626), 
        .B2(n16625), .ZN(n16632) );
  AOI21_X1 U19846 ( .B1(n16628), .B2(n16635), .A(n16627), .ZN(n17581) );
  OAI21_X1 U19847 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16635), .A(
        n16723), .ZN(n16629) );
  XNOR2_X1 U19848 ( .A(n17581), .B(n16629), .ZN(n16630) );
  AOI22_X1 U19849 ( .A1(n16739), .A2(n16630), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n16643), .ZN(n16631) );
  NAND4_X1 U19850 ( .A1(n16633), .A2(n16632), .A3(n16631), .A4(n18048), .ZN(
        P3_U2659) );
  INV_X1 U19851 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17604) );
  NAND2_X1 U19852 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17633), .ZN(
        n16701) );
  OAI21_X1 U19853 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16701), .A(
        n16723), .ZN(n16688) );
  OAI21_X1 U19854 ( .B1(n17593), .B2(n16738), .A(n16688), .ZN(n16654) );
  AOI21_X1 U19855 ( .B1(n16723), .B2(n17604), .A(n16654), .ZN(n16636) );
  NOR2_X1 U19856 ( .A1(n17728), .A2(n16634), .ZN(n16652) );
  OAI21_X1 U19857 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16652), .A(
        n16635), .ZN(n17594) );
  XNOR2_X1 U19858 ( .A(n16636), .B(n17594), .ZN(n16646) );
  AOI21_X1 U19859 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16759), .A(
        n18038), .ZN(n16645) );
  OAI21_X1 U19860 ( .B1(n16781), .B2(n16637), .A(n18610), .ZN(n16642) );
  NOR2_X1 U19861 ( .A1(n16647), .A2(n16638), .ZN(n16639) );
  OAI22_X1 U19862 ( .A1(n16784), .A2(n16639), .B1(n16785), .B2(n16638), .ZN(
        n16640) );
  AOI22_X1 U19863 ( .A1(n16643), .A2(n16642), .B1(n16641), .B2(n16640), .ZN(
        n16644) );
  OAI211_X1 U19864 ( .C1(n18569), .C2(n16646), .A(n16645), .B(n16644), .ZN(
        P3_U2660) );
  AOI22_X1 U19865 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16759), .B1(
        n16768), .B2(P3_EBX_REG_10__SCAN_IN), .ZN(n16658) );
  NOR2_X1 U19866 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n16781), .ZN(n16649) );
  AOI211_X1 U19867 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16667), .A(n16647), .B(
        n16784), .ZN(n16648) );
  AOI211_X1 U19868 ( .C1(n16650), .C2(n16649), .A(n18038), .B(n16648), .ZN(
        n16657) );
  AOI21_X1 U19869 ( .B1(n16651), .B2(n16763), .A(n16787), .ZN(n16679) );
  INV_X1 U19870 ( .A(n16679), .ZN(n16665) );
  NOR3_X1 U19871 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16781), .A3(n16651), .ZN(
        n16666) );
  OAI21_X1 U19872 ( .B1(n16665), .B2(n16666), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n16656) );
  NOR2_X1 U19873 ( .A1(n17634), .A2(n16701), .ZN(n16675) );
  NAND2_X1 U19874 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16675), .ZN(
        n16659) );
  AOI21_X1 U19875 ( .B1(n17604), .B2(n16659), .A(n16652), .ZN(n17607) );
  INV_X1 U19876 ( .A(n17607), .ZN(n16653) );
  INV_X1 U19877 ( .A(n16654), .ZN(n16660) );
  OAI221_X1 U19878 ( .B1(n17607), .B2(n16654), .C1(n16653), .C2(n16660), .A(
        n16739), .ZN(n16655) );
  NAND4_X1 U19879 ( .A1(n16658), .A2(n16657), .A3(n16656), .A4(n16655), .ZN(
        P3_U2661) );
  OAI21_X1 U19880 ( .B1(n16675), .B2(n16754), .A(n16777), .ZN(n16662) );
  OAI21_X1 U19881 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16675), .A(
        n16659), .ZN(n17622) );
  NAND2_X1 U19882 ( .A1(n16739), .A2(n17622), .ZN(n16661) );
  AOI22_X1 U19883 ( .A1(n16662), .A2(n16661), .B1(n16660), .B2(n17622), .ZN(
        n16664) );
  OAI22_X1 U19884 ( .A1(n17621), .A2(n16774), .B1(n16785), .B2(n17031), .ZN(
        n16663) );
  AOI211_X1 U19885 ( .C1(n16665), .C2(P3_REIP_REG_9__SCAN_IN), .A(n16664), .B(
        n16663), .ZN(n16670) );
  INV_X1 U19886 ( .A(n16666), .ZN(n16669) );
  OAI211_X1 U19887 ( .C1(n16671), .C2(n17031), .A(n16748), .B(n16667), .ZN(
        n16668) );
  NAND4_X1 U19888 ( .A1(n16670), .A2(n18048), .A3(n16669), .A4(n16668), .ZN(
        P3_U2662) );
  INV_X1 U19889 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n16684) );
  AOI211_X1 U19890 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16696), .A(n16671), .B(
        n16784), .ZN(n16682) );
  AOI21_X1 U19891 ( .B1(n16763), .B2(n16672), .A(P3_REIP_REG_8__SCAN_IN), .ZN(
        n16680) );
  NAND2_X1 U19892 ( .A1(n17633), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16674) );
  INV_X1 U19893 ( .A(n16674), .ZN(n17635) );
  AOI21_X1 U19894 ( .B1(n17635), .B2(n16673), .A(n16738), .ZN(n16677) );
  NOR2_X1 U19895 ( .A1(n17728), .A2(n16674), .ZN(n16687) );
  INV_X1 U19896 ( .A(n16675), .ZN(n16676) );
  OAI21_X1 U19897 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16687), .A(
        n16676), .ZN(n17637) );
  XOR2_X1 U19898 ( .A(n16677), .B(n17637), .Z(n16678) );
  OAI22_X1 U19899 ( .A1(n16680), .A2(n16679), .B1(n18569), .B2(n16678), .ZN(
        n16681) );
  AOI211_X1 U19900 ( .C1(n16759), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16682), .B(n16681), .ZN(n16683) );
  OAI211_X1 U19901 ( .C1(n16785), .C2(n16684), .A(n16683), .B(n18048), .ZN(
        P3_U2663) );
  OAI21_X1 U19902 ( .B1(n16781), .B2(n16686), .A(n16782), .ZN(n16685) );
  INV_X1 U19903 ( .A(n16685), .ZN(n16712) );
  INV_X1 U19904 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18600) );
  NAND3_X1 U19905 ( .A1(n18600), .A2(n16763), .A3(n16686), .ZN(n16699) );
  AOI21_X1 U19906 ( .B1(n16712), .B2(n16699), .A(n18602), .ZN(n16695) );
  INV_X1 U19907 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17651) );
  AOI21_X1 U19908 ( .B1(n17651), .B2(n16701), .A(n16687), .ZN(n17657) );
  INV_X1 U19909 ( .A(n16688), .ZN(n16690) );
  INV_X1 U19910 ( .A(n17657), .ZN(n16689) );
  AOI221_X1 U19911 ( .B1(n17657), .B2(n16690), .C1(n16689), .C2(n16688), .A(
        n18569), .ZN(n16694) );
  NAND2_X1 U19912 ( .A1(n16763), .A2(n18602), .ZN(n16691) );
  OAI22_X1 U19913 ( .A1(n17651), .A2(n16774), .B1(n16692), .B2(n16691), .ZN(
        n16693) );
  NOR4_X1 U19914 ( .A1(n18038), .A2(n16695), .A3(n16694), .A4(n16693), .ZN(
        n16698) );
  OAI211_X1 U19915 ( .C1(n16705), .C2(n17007), .A(n16748), .B(n16696), .ZN(
        n16697) );
  OAI211_X1 U19916 ( .C1(n17007), .C2(n16785), .A(n16698), .B(n16697), .ZN(
        P3_U2664) );
  INV_X1 U19917 ( .A(n16699), .ZN(n16700) );
  AOI211_X1 U19918 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16768), .A(n18038), .B(
        n16700), .ZN(n16709) );
  NOR2_X1 U19919 ( .A1(n17728), .A2(n17662), .ZN(n16710) );
  OAI21_X1 U19920 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16710), .A(
        n16701), .ZN(n17669) );
  INV_X1 U19921 ( .A(n17669), .ZN(n16704) );
  OAI21_X1 U19922 ( .B1(n16754), .B2(n17663), .A(n16777), .ZN(n16703) );
  NOR2_X1 U19923 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16701), .ZN(
        n16702) );
  AOI221_X1 U19924 ( .B1(n16704), .B2(n16703), .C1(n17669), .C2(n16775), .A(
        n16702), .ZN(n16707) );
  AOI211_X1 U19925 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16714), .A(n16705), .B(
        n16784), .ZN(n16706) );
  AOI211_X1 U19926 ( .C1(n16759), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16707), .B(n16706), .ZN(n16708) );
  OAI211_X1 U19927 ( .C1(n18600), .C2(n16712), .A(n16709), .B(n16708), .ZN(
        P3_U2665) );
  INV_X1 U19928 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16716) );
  NAND2_X1 U19929 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17683), .ZN(
        n16722) );
  AOI21_X1 U19930 ( .B1(n16716), .B2(n16722), .A(n16710), .ZN(n17681) );
  INV_X1 U19931 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16786) );
  INV_X1 U19932 ( .A(n16722), .ZN(n16711) );
  AOI21_X1 U19933 ( .B1(n16786), .B2(n16711), .A(n16738), .ZN(n16725) );
  XOR2_X1 U19934 ( .A(n17681), .B(n16725), .Z(n16719) );
  AOI221_X1 U19935 ( .B1(n16781), .B2(n18598), .C1(n16713), .C2(n18598), .A(
        n16712), .ZN(n16718) );
  OAI211_X1 U19936 ( .C1(n16728), .C2(n16721), .A(n16748), .B(n16714), .ZN(
        n16715) );
  OAI21_X1 U19937 ( .B1(n16774), .B2(n16716), .A(n16715), .ZN(n16717) );
  AOI211_X1 U19938 ( .C1(n16739), .C2(n16719), .A(n16718), .B(n16717), .ZN(
        n16720) );
  OAI211_X1 U19939 ( .C1(n16785), .C2(n16721), .A(n16720), .B(n18048), .ZN(
        P3_U2666) );
  NOR2_X1 U19940 ( .A1(n17728), .A2(n17686), .ZN(n16737) );
  OAI21_X1 U19941 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16737), .A(
        n16722), .ZN(n17696) );
  OR2_X1 U19942 ( .A1(n17686), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17692) );
  OAI22_X1 U19943 ( .A1(n16723), .A2(n17696), .B1(n16761), .B2(n17692), .ZN(
        n16724) );
  AOI21_X1 U19944 ( .B1(n16725), .B2(n17696), .A(n16724), .ZN(n16735) );
  NOR2_X1 U19945 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16781), .ZN(n16726) );
  AOI22_X1 U19946 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16759), .B1(
        n16727), .B2(n16726), .ZN(n16734) );
  OAI21_X1 U19947 ( .B1(n16727), .B2(n16781), .A(n16782), .ZN(n16746) );
  AOI211_X1 U19948 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16747), .A(n16728), .B(
        n16784), .ZN(n16732) );
  NAND2_X1 U19949 ( .A1(n18062), .A2(n18731), .ZN(n16792) );
  INV_X1 U19950 ( .A(n16792), .ZN(n18732) );
  OAI21_X1 U19951 ( .B1(n16998), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n18732), .ZN(n16729) );
  OAI211_X1 U19952 ( .C1(n16785), .C2(n16730), .A(n18048), .B(n16729), .ZN(
        n16731) );
  AOI211_X1 U19953 ( .C1(P3_REIP_REG_4__SCAN_IN), .C2(n16746), .A(n16732), .B(
        n16731), .ZN(n16733) );
  OAI211_X1 U19954 ( .C1(n16735), .C2(n18569), .A(n16734), .B(n16733), .ZN(
        P3_U2667) );
  NOR2_X1 U19955 ( .A1(n16736), .A2(n18522), .ZN(n18512) );
  OAI21_X1 U19956 ( .B1(n18672), .B2(n18512), .A(n10014), .ZN(n18668) );
  INV_X1 U19957 ( .A(n18668), .ZN(n16752) );
  OAI21_X1 U19958 ( .B1(n16781), .B2(n16764), .A(n18594), .ZN(n16745) );
  INV_X1 U19959 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16742) );
  NAND2_X1 U19960 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16753) );
  AOI21_X1 U19961 ( .B1(n16742), .B2(n16753), .A(n16737), .ZN(n17710) );
  NOR2_X1 U19962 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16753), .ZN(
        n16760) );
  NOR2_X1 U19963 ( .A1(n16760), .A2(n16738), .ZN(n16741) );
  OAI21_X1 U19964 ( .B1(n17710), .B2(n16741), .A(n16739), .ZN(n16740) );
  AOI21_X1 U19965 ( .B1(n17710), .B2(n16741), .A(n16740), .ZN(n16744) );
  OAI22_X1 U19966 ( .A1(n16742), .A2(n16774), .B1(n16785), .B2(n16749), .ZN(
        n16743) );
  AOI211_X1 U19967 ( .C1(n16746), .C2(n16745), .A(n16744), .B(n16743), .ZN(
        n16751) );
  OAI211_X1 U19968 ( .C1(n16755), .C2(n16749), .A(n16748), .B(n16747), .ZN(
        n16750) );
  OAI211_X1 U19969 ( .C1(n16752), .C2(n16792), .A(n16751), .B(n16750), .ZN(
        P3_U2668) );
  OAI21_X1 U19970 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16753), .ZN(n17718) );
  INV_X1 U19971 ( .A(n16754), .ZN(n16771) );
  INV_X1 U19972 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n16783) );
  INV_X1 U19973 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17100) );
  NAND2_X1 U19974 ( .A1(n16783), .A2(n17100), .ZN(n16756) );
  AOI211_X1 U19975 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16756), .A(n16755), .B(
        n16784), .ZN(n16758) );
  INV_X1 U19976 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20923) );
  NAND2_X1 U19977 ( .A1(n18682), .A2(n18517), .ZN(n18511) );
  OAI21_X1 U19978 ( .B1(n18522), .B2(n16736), .A(n18511), .ZN(n18678) );
  OAI22_X1 U19979 ( .A1(n20923), .A2(n16782), .B1(n18678), .B2(n16792), .ZN(
        n16757) );
  AOI211_X1 U19980 ( .C1(n16759), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n16758), .B(n16757), .ZN(n16770) );
  INV_X1 U19981 ( .A(n17718), .ZN(n16762) );
  AOI211_X1 U19982 ( .C1(n16762), .C2(n16761), .A(n16760), .B(n16775), .ZN(
        n16767) );
  OAI211_X1 U19983 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n16764), .B(n16763), .ZN(n16765) );
  INV_X1 U19984 ( .A(n16765), .ZN(n16766) );
  AOI211_X1 U19985 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16768), .A(n16767), .B(
        n16766), .ZN(n16769) );
  OAI211_X1 U19986 ( .C1(n17718), .C2(n16771), .A(n16770), .B(n16769), .ZN(
        P3_U2669) );
  NOR2_X1 U19987 ( .A1(n16783), .A2(n17100), .ZN(n17093) );
  INV_X1 U19988 ( .A(n17093), .ZN(n16772) );
  OAI21_X1 U19989 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n16772), .ZN(n17101) );
  AND2_X1 U19990 ( .A1(n18517), .A2(n16773), .ZN(n18687) );
  AOI22_X1 U19991 ( .A1(n16787), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18687), 
        .B2(n18732), .ZN(n16780) );
  OAI21_X1 U19992 ( .B1(n16786), .B2(n16775), .A(n16774), .ZN(n16778) );
  OAI22_X1 U19993 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16781), .B1(n16785), 
        .B2(n17100), .ZN(n16776) );
  AOI221_X1 U19994 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16778), .C1(
        n17728), .C2(n16777), .A(n16776), .ZN(n16779) );
  OAI211_X1 U19995 ( .C1(n16784), .C2(n17101), .A(n16780), .B(n16779), .ZN(
        P3_U2670) );
  NAND2_X1 U19996 ( .A1(n16782), .A2(n16781), .ZN(n16790) );
  AOI21_X1 U19997 ( .B1(n16785), .B2(n16784), .A(n16783), .ZN(n16789) );
  NOR3_X1 U19998 ( .A1(n18693), .A2(n16787), .A3(n16786), .ZN(n16788) );
  AOI211_X1 U19999 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(n16790), .A(n16789), .B(
        n16788), .ZN(n16791) );
  OAI21_X1 U20000 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16792), .A(
        n16791), .ZN(P3_U2671) );
  INV_X1 U20001 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16794) );
  NAND2_X1 U20002 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16909), .ZN(n16879) );
  NAND4_X1 U20003 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(P3_EBX_REG_29__SCAN_IN), 
        .A3(P3_EBX_REG_23__SCAN_IN), .A4(P3_EBX_REG_22__SCAN_IN), .ZN(n16793)
         );
  NOR4_X1 U20004 ( .A1(n16795), .A2(n16794), .A3(n16879), .A4(n16793), .ZN(
        n16796) );
  NAND4_X1 U20005 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(P3_EBX_REG_25__SCAN_IN), .A4(n16796), .ZN(n16799) );
  NOR2_X1 U20006 ( .A1(n16800), .A2(n16799), .ZN(n16827) );
  NAND2_X1 U20007 ( .A1(n17097), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16798) );
  NAND2_X1 U20008 ( .A1(n16827), .A2(n18094), .ZN(n16797) );
  OAI22_X1 U20009 ( .A1(n16827), .A2(n16798), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16797), .ZN(P3_U2672) );
  NAND2_X1 U20010 ( .A1(n16800), .A2(n16799), .ZN(n16801) );
  NAND2_X1 U20011 ( .A1(n16801), .A2(n17097), .ZN(n16826) );
  AOI22_X1 U20012 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n16998), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16805) );
  AOI22_X1 U20013 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17060), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n17064), .ZN(n16804) );
  AOI22_X1 U20014 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n9608), .ZN(n16803) );
  AOI22_X1 U20015 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16802) );
  NAND4_X1 U20016 ( .A1(n16805), .A2(n16804), .A3(n16803), .A4(n16802), .ZN(
        n16812) );
  AOI22_X1 U20017 ( .A1(n17065), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17062), .ZN(n16810) );
  AOI22_X1 U20018 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n16806), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16809) );
  AOI22_X1 U20019 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17051), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16808) );
  AOI22_X1 U20020 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n17036), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17052), .ZN(n16807) );
  NAND4_X1 U20021 ( .A1(n16810), .A2(n16809), .A3(n16808), .A4(n16807), .ZN(
        n16811) );
  NOR2_X1 U20022 ( .A1(n16812), .A2(n16811), .ZN(n16825) );
  AOI22_X1 U20023 ( .A1(n16813), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16824) );
  AOI22_X1 U20024 ( .A1(n17065), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16823) );
  AOI22_X1 U20025 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16814) );
  OAI21_X1 U20026 ( .B1(n16815), .B2(n20820), .A(n16814), .ZN(n16821) );
  AOI22_X1 U20027 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16819) );
  AOI22_X1 U20028 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16818) );
  AOI22_X1 U20029 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16817) );
  AOI22_X1 U20030 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16816) );
  NAND4_X1 U20031 ( .A1(n16819), .A2(n16818), .A3(n16817), .A4(n16816), .ZN(
        n16820) );
  AOI211_X1 U20032 ( .C1(n17064), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n16821), .B(n16820), .ZN(n16822) );
  NAND3_X1 U20033 ( .A1(n16824), .A2(n16823), .A3(n16822), .ZN(n16829) );
  NAND2_X1 U20034 ( .A1(n16830), .A2(n16829), .ZN(n16828) );
  XNOR2_X1 U20035 ( .A(n16825), .B(n16828), .ZN(n17116) );
  OAI22_X1 U20036 ( .A1(n16827), .A2(n16826), .B1(n17116), .B2(n17097), .ZN(
        P3_U2673) );
  OAI21_X1 U20037 ( .B1(n16830), .B2(n16829), .A(n16828), .ZN(n17120) );
  NAND3_X1 U20038 ( .A1(n16832), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n17097), 
        .ZN(n16831) );
  OAI221_X1 U20039 ( .B1(n16832), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n17085), 
        .C2(n17120), .A(n16831), .ZN(P3_U2674) );
  INV_X1 U20040 ( .A(n16833), .ZN(n16841) );
  AOI21_X1 U20041 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17097), .A(n16841), .ZN(
        n16837) );
  OAI21_X1 U20042 ( .B1(n16836), .B2(n16835), .A(n16834), .ZN(n17129) );
  OAI22_X1 U20043 ( .A1(n16838), .A2(n16837), .B1(n17097), .B2(n17129), .ZN(
        P3_U2676) );
  AOI22_X1 U20044 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17097), .B1(
        P3_EBX_REG_25__SCAN_IN), .B2(n16849), .ZN(n16840) );
  XNOR2_X1 U20045 ( .A(n16839), .B(n16842), .ZN(n17133) );
  OAI22_X1 U20046 ( .A1(n16841), .A2(n16840), .B1(n17085), .B2(n17133), .ZN(
        P3_U2677) );
  OAI21_X1 U20047 ( .B1(n16844), .B2(n16843), .A(n16842), .ZN(n17138) );
  NAND3_X1 U20048 ( .A1(n16846), .A2(P3_EBX_REG_25__SCAN_IN), .A3(n17097), 
        .ZN(n16845) );
  OAI221_X1 U20049 ( .B1(n16846), .B2(P3_EBX_REG_25__SCAN_IN), .C1(n17085), 
        .C2(n17138), .A(n16845), .ZN(P3_U2678) );
  AOI21_X1 U20050 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17097), .A(n16855), .ZN(
        n16848) );
  XNOR2_X1 U20051 ( .A(n16847), .B(n16851), .ZN(n17143) );
  OAI22_X1 U20052 ( .A1(n16849), .A2(n16848), .B1(n17085), .B2(n17143), .ZN(
        P3_U2679) );
  AOI21_X1 U20053 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17097), .A(n16850), .ZN(
        n16854) );
  OAI21_X1 U20054 ( .B1(n16853), .B2(n16852), .A(n16851), .ZN(n17148) );
  OAI22_X1 U20055 ( .A1(n16855), .A2(n16854), .B1(n17097), .B2(n17148), .ZN(
        P3_U2680) );
  AOI22_X1 U20056 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16865) );
  AOI22_X1 U20057 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16864) );
  AOI22_X1 U20058 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16856) );
  OAI21_X1 U20059 ( .B1(n10014), .B2(n20820), .A(n16856), .ZN(n16862) );
  AOI22_X1 U20060 ( .A1(n17034), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17064), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16860) );
  AOI22_X1 U20061 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16859) );
  AOI22_X1 U20062 ( .A1(n17065), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9579), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16858) );
  AOI22_X1 U20063 ( .A1(n16965), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16857) );
  NAND4_X1 U20064 ( .A1(n16860), .A2(n16859), .A3(n16858), .A4(n16857), .ZN(
        n16861) );
  AOI211_X1 U20065 ( .C1(n17061), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n16862), .B(n16861), .ZN(n16863) );
  NAND3_X1 U20066 ( .A1(n16865), .A2(n16864), .A3(n16863), .ZN(n17149) );
  INV_X1 U20067 ( .A(n17149), .ZN(n16867) );
  NAND3_X1 U20068 ( .A1(n16868), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17097), 
        .ZN(n16866) );
  OAI221_X1 U20069 ( .B1(n16868), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17085), 
        .C2(n16867), .A(n16866), .ZN(P3_U2681) );
  AOI22_X1 U20070 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16872) );
  AOI22_X1 U20071 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16871) );
  AOI22_X1 U20072 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16870) );
  AOI22_X1 U20073 ( .A1(n16965), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16869) );
  NAND4_X1 U20074 ( .A1(n16872), .A2(n16871), .A3(n16870), .A4(n16869), .ZN(
        n16878) );
  AOI22_X1 U20075 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16876) );
  AOI22_X1 U20076 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16875) );
  AOI22_X1 U20077 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16874) );
  AOI22_X1 U20078 ( .A1(n17065), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17064), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16873) );
  NAND4_X1 U20079 ( .A1(n16876), .A2(n16875), .A3(n16874), .A4(n16873), .ZN(
        n16877) );
  NOR2_X1 U20080 ( .A1(n16878), .A2(n16877), .ZN(n17157) );
  AND2_X1 U20081 ( .A1(n17085), .A2(n16879), .ZN(n16893) );
  AOI22_X1 U20082 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16893), .B1(n16880), 
        .B2(n20835), .ZN(n16881) );
  OAI21_X1 U20083 ( .B1(n17157), .B2(n17085), .A(n16881), .ZN(P3_U2682) );
  AOI22_X1 U20084 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16892) );
  AOI22_X1 U20085 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17064), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16891) );
  AOI22_X1 U20086 ( .A1(n17034), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16882) );
  OAI21_X1 U20087 ( .B1(n16883), .B2(n20839), .A(n16882), .ZN(n16889) );
  AOI22_X1 U20088 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16887) );
  AOI22_X1 U20089 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16886) );
  AOI22_X1 U20090 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16885) );
  AOI22_X1 U20091 ( .A1(n16965), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16884) );
  NAND4_X1 U20092 ( .A1(n16887), .A2(n16886), .A3(n16885), .A4(n16884), .ZN(
        n16888) );
  AOI211_X1 U20093 ( .C1(n17061), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n16889), .B(n16888), .ZN(n16890) );
  NAND3_X1 U20094 ( .A1(n16892), .A2(n16891), .A3(n16890), .ZN(n17158) );
  INV_X1 U20095 ( .A(n17158), .ZN(n16896) );
  OAI21_X1 U20096 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16894), .A(n16893), .ZN(
        n16895) );
  OAI21_X1 U20097 ( .B1(n16896), .B2(n17097), .A(n16895), .ZN(P3_U2683) );
  INV_X1 U20098 ( .A(n16897), .ZN(n16922) );
  OAI21_X1 U20099 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n16922), .A(n17097), .ZN(
        n16908) );
  AOI22_X1 U20100 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16901) );
  AOI22_X1 U20101 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16900) );
  AOI22_X1 U20102 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16899) );
  AOI22_X1 U20103 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16898) );
  NAND4_X1 U20104 ( .A1(n16901), .A2(n16900), .A3(n16899), .A4(n16898), .ZN(
        n16907) );
  AOI22_X1 U20105 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16905) );
  AOI22_X1 U20106 ( .A1(n17034), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16904) );
  AOI22_X1 U20107 ( .A1(n16965), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16903) );
  AOI22_X1 U20108 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16902) );
  NAND4_X1 U20109 ( .A1(n16905), .A2(n16904), .A3(n16903), .A4(n16902), .ZN(
        n16906) );
  NOR2_X1 U20110 ( .A1(n16907), .A2(n16906), .ZN(n17167) );
  OAI22_X1 U20111 ( .A1(n16909), .A2(n16908), .B1(n17167), .B2(n17097), .ZN(
        P3_U2684) );
  AOI22_X1 U20112 ( .A1(n18094), .A2(n16910), .B1(P3_EBX_REG_18__SCAN_IN), 
        .B2(n17085), .ZN(n16921) );
  AOI22_X1 U20113 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16914) );
  AOI22_X1 U20114 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16913) );
  AOI22_X1 U20115 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16912) );
  AOI22_X1 U20116 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16911) );
  NAND4_X1 U20117 ( .A1(n16914), .A2(n16913), .A3(n16912), .A4(n16911), .ZN(
        n16920) );
  AOI22_X1 U20118 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16918) );
  AOI22_X1 U20119 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16917) );
  AOI22_X1 U20120 ( .A1(n17034), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16916) );
  AOI22_X1 U20121 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16915) );
  NAND4_X1 U20122 ( .A1(n16918), .A2(n16917), .A3(n16916), .A4(n16915), .ZN(
        n16919) );
  NOR2_X1 U20123 ( .A1(n16920), .A2(n16919), .ZN(n17172) );
  OAI22_X1 U20124 ( .A1(n16922), .A2(n16921), .B1(n17172), .B2(n17097), .ZN(
        P3_U2685) );
  NOR3_X1 U20125 ( .A1(n17185), .A2(n17005), .A3(n16923), .ZN(n16963) );
  NAND2_X1 U20126 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16963), .ZN(n16945) );
  AOI22_X1 U20127 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16927) );
  AOI22_X1 U20128 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17064), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16926) );
  AOI22_X1 U20129 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16925) );
  AOI22_X1 U20130 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16924) );
  NAND4_X1 U20131 ( .A1(n16927), .A2(n16926), .A3(n16925), .A4(n16924), .ZN(
        n16933) );
  AOI22_X1 U20132 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16931) );
  AOI22_X1 U20133 ( .A1(n17034), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16930) );
  AOI22_X1 U20134 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16929) );
  AOI22_X1 U20135 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16928) );
  NAND4_X1 U20136 ( .A1(n16931), .A2(n16930), .A3(n16929), .A4(n16928), .ZN(
        n16932) );
  NOR2_X1 U20137 ( .A1(n16933), .A2(n16932), .ZN(n17177) );
  NAND3_X1 U20138 ( .A1(n16945), .A2(P3_EBX_REG_17__SCAN_IN), .A3(n17097), 
        .ZN(n16934) );
  OAI221_X1 U20139 ( .B1(n16945), .B2(P3_EBX_REG_17__SCAN_IN), .C1(n17085), 
        .C2(n17177), .A(n16934), .ZN(P3_U2686) );
  AOI22_X1 U20140 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16938) );
  AOI22_X1 U20141 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16937) );
  AOI22_X1 U20142 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16936) );
  AOI22_X1 U20143 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16935) );
  NAND4_X1 U20144 ( .A1(n16938), .A2(n16937), .A3(n16936), .A4(n16935), .ZN(
        n16944) );
  AOI22_X1 U20145 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16942) );
  AOI22_X1 U20146 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16983), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16941) );
  AOI22_X1 U20147 ( .A1(n9579), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16940) );
  AOI22_X1 U20148 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16939) );
  NAND4_X1 U20149 ( .A1(n16942), .A2(n16941), .A3(n16940), .A4(n16939), .ZN(
        n16943) );
  NOR2_X1 U20150 ( .A1(n16944), .A2(n16943), .ZN(n17184) );
  INV_X1 U20151 ( .A(n16945), .ZN(n16947) );
  AOI21_X1 U20152 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17097), .A(n16963), .ZN(
        n16946) );
  OAI22_X1 U20153 ( .A1(n17184), .A2(n17097), .B1(n16947), .B2(n16946), .ZN(
        P3_U2687) );
  INV_X1 U20154 ( .A(n17005), .ZN(n16949) );
  INV_X1 U20155 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16975) );
  NOR2_X1 U20156 ( .A1(n16975), .A2(n16990), .ZN(n16948) );
  OAI221_X1 U20157 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n16949), .C1(
        P3_EBX_REG_15__SCAN_IN), .C2(n16948), .A(n17097), .ZN(n16962) );
  AOI22_X1 U20158 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16960) );
  AOI22_X1 U20159 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17054), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n9608), .ZN(n16959) );
  AOI22_X1 U20160 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17036), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n16965), .ZN(n16950) );
  OAI21_X1 U20161 ( .B1(n10022), .B2(n16951), .A(n16950), .ZN(n16957) );
  AOI22_X1 U20162 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17060), .ZN(n16955) );
  AOI22_X1 U20163 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17012), .ZN(n16954) );
  AOI22_X1 U20164 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n17052), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16953) );
  AOI22_X1 U20165 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16952) );
  NAND4_X1 U20166 ( .A1(n16955), .A2(n16954), .A3(n16953), .A4(n16952), .ZN(
        n16956) );
  AOI211_X1 U20167 ( .C1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .C2(n17034), .A(
        n16957), .B(n16956), .ZN(n16958) );
  NAND3_X1 U20168 ( .A1(n16960), .A2(n16959), .A3(n16958), .ZN(n17187) );
  INV_X1 U20169 ( .A(n17187), .ZN(n16961) );
  OAI22_X1 U20170 ( .A1(n16963), .A2(n16962), .B1(n16961), .B2(n17097), .ZN(
        P3_U2688) );
  AOI22_X1 U20171 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16974) );
  AOI22_X1 U20172 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17064), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16973) );
  AOI22_X1 U20173 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16983), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16964) );
  OAI21_X1 U20174 ( .B1(n12588), .B2(n20820), .A(n16964), .ZN(n16971) );
  AOI22_X1 U20175 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16969) );
  AOI22_X1 U20176 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16968) );
  AOI22_X1 U20177 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16967) );
  AOI22_X1 U20178 ( .A1(n16965), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16966) );
  NAND4_X1 U20179 ( .A1(n16969), .A2(n16968), .A3(n16967), .A4(n16966), .ZN(
        n16970) );
  AOI211_X1 U20180 ( .C1(n17061), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n16971), .B(n16970), .ZN(n16972) );
  NAND3_X1 U20181 ( .A1(n16974), .A2(n16973), .A3(n16972), .ZN(n17190) );
  INV_X1 U20182 ( .A(n17190), .ZN(n16978) );
  OAI211_X1 U20183 ( .C1(n16990), .C2(n17005), .A(P3_EBX_REG_14__SCAN_IN), .B(
        n17097), .ZN(n16977) );
  NOR2_X1 U20184 ( .A1(n17185), .A2(n17005), .ZN(n16991) );
  NAND3_X1 U20185 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16991), .A3(n16975), 
        .ZN(n16976) );
  OAI211_X1 U20186 ( .C1(n16978), .C2(n17085), .A(n16977), .B(n16976), .ZN(
        P3_U2689) );
  AOI22_X1 U20187 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16982) );
  AOI22_X1 U20188 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17064), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16981) );
  AOI22_X1 U20189 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16980) );
  AOI22_X1 U20190 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16979) );
  NAND4_X1 U20191 ( .A1(n16982), .A2(n16981), .A3(n16980), .A4(n16979), .ZN(
        n16989) );
  AOI22_X1 U20192 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16987) );
  AOI22_X1 U20193 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16986) );
  AOI22_X1 U20194 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16985) );
  AOI22_X1 U20195 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16984) );
  NAND4_X1 U20196 ( .A1(n16987), .A2(n16986), .A3(n16985), .A4(n16984), .ZN(
        n16988) );
  NOR2_X1 U20197 ( .A1(n16989), .A2(n16988), .ZN(n17194) );
  AOI21_X1 U20198 ( .B1(n17097), .B2(n17005), .A(n16990), .ZN(n16993) );
  NOR2_X1 U20199 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16991), .ZN(n16992) );
  OAI22_X1 U20200 ( .A1(n17194), .A2(n17097), .B1(n16993), .B2(n16992), .ZN(
        P3_U2690) );
  AOI22_X1 U20201 ( .A1(n17034), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16997) );
  AOI22_X1 U20202 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16996) );
  AOI22_X1 U20203 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16995) );
  AOI22_X1 U20204 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16994) );
  NAND4_X1 U20205 ( .A1(n16997), .A2(n16996), .A3(n16995), .A4(n16994), .ZN(
        n17004) );
  AOI22_X1 U20206 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17064), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17002) );
  AOI22_X1 U20207 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17001) );
  AOI22_X1 U20208 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17000) );
  AOI22_X1 U20209 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16999) );
  NAND4_X1 U20210 ( .A1(n17002), .A2(n17001), .A3(n17000), .A4(n16999), .ZN(
        n17003) );
  NOR2_X1 U20211 ( .A1(n17004), .A2(n17003), .ZN(n17198) );
  OAI211_X1 U20212 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17020), .A(n17005), .B(
        n17097), .ZN(n17006) );
  OAI21_X1 U20213 ( .B1(n17198), .B2(n17097), .A(n17006), .ZN(P3_U2691) );
  NOR2_X1 U20214 ( .A1(n17007), .A2(n17075), .ZN(n17079) );
  NAND2_X1 U20215 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17079), .ZN(n17073) );
  INV_X1 U20216 ( .A(n17073), .ZN(n17048) );
  AND3_X1 U20217 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(n17048), .ZN(n17033) );
  OAI21_X1 U20218 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17033), .A(n17097), .ZN(
        n17019) );
  AOI22_X1 U20219 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17064), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17011) );
  AOI22_X1 U20220 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U20221 ( .A1(n17052), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17009) );
  AOI22_X1 U20222 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17008) );
  NAND4_X1 U20223 ( .A1(n17011), .A2(n17010), .A3(n17009), .A4(n17008), .ZN(
        n17018) );
  AOI22_X1 U20224 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17016) );
  AOI22_X1 U20225 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17015) );
  AOI22_X1 U20226 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17014) );
  AOI22_X1 U20227 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17013) );
  NAND4_X1 U20228 ( .A1(n17016), .A2(n17015), .A3(n17014), .A4(n17013), .ZN(
        n17017) );
  NOR2_X1 U20229 ( .A1(n17018), .A2(n17017), .ZN(n17201) );
  OAI22_X1 U20230 ( .A1(n17020), .A2(n17019), .B1(n17201), .B2(n17097), .ZN(
        P3_U2692) );
  AOI22_X1 U20231 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17024) );
  AOI22_X1 U20232 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17023) );
  AOI22_X1 U20233 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17064), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17022) );
  AOI22_X1 U20234 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17021) );
  NAND4_X1 U20235 ( .A1(n17024), .A2(n17023), .A3(n17022), .A4(n17021), .ZN(
        n17030) );
  AOI22_X1 U20236 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20237 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17027) );
  AOI22_X1 U20238 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17026) );
  AOI22_X1 U20239 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17025) );
  NAND4_X1 U20240 ( .A1(n17028), .A2(n17027), .A3(n17026), .A4(n17025), .ZN(
        n17029) );
  NOR2_X1 U20241 ( .A1(n17030), .A2(n17029), .ZN(n17207) );
  NOR2_X1 U20242 ( .A1(n17031), .A2(n17073), .ZN(n17050) );
  OAI21_X1 U20243 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17050), .A(n17097), .ZN(
        n17032) );
  OAI22_X1 U20244 ( .A1(n17207), .A2(n17097), .B1(n17033), .B2(n17032), .ZN(
        P3_U2693) );
  AOI22_X1 U20245 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17040) );
  AOI22_X1 U20246 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20247 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20248 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17037) );
  NAND4_X1 U20249 ( .A1(n17040), .A2(n17039), .A3(n17038), .A4(n17037), .ZN(
        n17047) );
  AOI22_X1 U20250 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17045) );
  AOI22_X1 U20251 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U20252 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9579), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U20253 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17042) );
  NAND4_X1 U20254 ( .A1(n17045), .A2(n17044), .A3(n17043), .A4(n17042), .ZN(
        n17046) );
  NOR2_X1 U20255 ( .A1(n17047), .A2(n17046), .ZN(n17209) );
  OAI21_X1 U20256 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17048), .A(n17097), .ZN(
        n17049) );
  OAI22_X1 U20257 ( .A1(n17209), .A2(n17097), .B1(n17050), .B2(n17049), .ZN(
        P3_U2694) );
  AOI22_X1 U20258 ( .A1(n17034), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17059) );
  AOI22_X1 U20259 ( .A1(n9608), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17058) );
  AOI22_X1 U20260 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U20261 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17056) );
  NAND4_X1 U20262 ( .A1(n17059), .A2(n17058), .A3(n17057), .A4(n17056), .ZN(
        n17072) );
  AOI22_X1 U20263 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U20264 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17069) );
  AOI22_X1 U20265 ( .A1(n17065), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17064), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U20266 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17067) );
  NAND4_X1 U20267 ( .A1(n17070), .A2(n17069), .A3(n17068), .A4(n17067), .ZN(
        n17071) );
  NOR2_X1 U20268 ( .A1(n17072), .A2(n17071), .ZN(n17216) );
  OAI211_X1 U20269 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17079), .A(n17073), .B(
        n17097), .ZN(n17074) );
  OAI21_X1 U20270 ( .B1(n17216), .B2(n17097), .A(n17074), .ZN(P3_U2695) );
  INV_X1 U20271 ( .A(n17075), .ZN(n17076) );
  AOI22_X1 U20272 ( .A1(n18094), .A2(n17076), .B1(P3_EBX_REG_7__SCAN_IN), .B2(
        n17085), .ZN(n17078) );
  INV_X1 U20273 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17077) );
  OAI22_X1 U20274 ( .A1(n17079), .A2(n17078), .B1(n17077), .B2(n17097), .ZN(
        P3_U2696) );
  NAND3_X1 U20275 ( .A1(n18094), .A2(P3_EBX_REG_5__SCAN_IN), .A3(n17089), .ZN(
        n17082) );
  INV_X1 U20276 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17081) );
  NAND3_X1 U20277 ( .A1(n17082), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n17097), .ZN(
        n17080) );
  OAI221_X1 U20278 ( .B1(n17082), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n17085), 
        .C2(n17081), .A(n17080), .ZN(P3_U2697) );
  INV_X1 U20279 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17084) );
  OAI211_X1 U20280 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17089), .A(n17082), .B(
        n17097), .ZN(n17083) );
  OAI21_X1 U20281 ( .B1(n17085), .B2(n17084), .A(n17083), .ZN(P3_U2698) );
  NAND2_X1 U20282 ( .A1(n18094), .A2(n17099), .ZN(n17105) );
  NOR2_X1 U20283 ( .A1(n17086), .A2(n17105), .ZN(n17094) );
  AND2_X1 U20284 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17094), .ZN(n17092) );
  AOI21_X1 U20285 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17097), .A(n17092), .ZN(
        n17088) );
  INV_X1 U20286 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17087) );
  OAI22_X1 U20287 ( .A1(n17089), .A2(n17088), .B1(n17087), .B2(n17097), .ZN(
        P3_U2699) );
  AOI21_X1 U20288 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17097), .A(n17094), .ZN(
        n17091) );
  INV_X1 U20289 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17090) );
  OAI22_X1 U20290 ( .A1(n17092), .A2(n17091), .B1(n17090), .B2(n17097), .ZN(
        P3_U2700) );
  AOI21_X1 U20291 ( .B1(n17099), .B2(n17093), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17096) );
  AOI221_X1 U20292 ( .B1(n17096), .B2(n17097), .C1(n17095), .C2(n17103), .A(
        n17094), .ZN(P3_U2701) );
  INV_X1 U20293 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17098) );
  OAI222_X1 U20294 ( .A1(n17105), .A2(n17101), .B1(n17100), .B2(n17099), .C1(
        n17098), .C2(n17097), .ZN(P3_U2702) );
  AOI22_X1 U20295 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17103), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17102), .ZN(n17104) );
  OAI21_X1 U20296 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17105), .A(n17104), .ZN(
        P3_U2703) );
  INV_X1 U20297 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17258) );
  INV_X1 U20298 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17326) );
  INV_X1 U20299 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n20819) );
  INV_X1 U20300 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17365) );
  NAND4_X1 U20301 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .A4(P3_EAX_REG_1__SCAN_IN), .ZN(n17106) );
  NAND2_X1 U20302 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17224), .ZN(n17218) );
  NAND4_X1 U20303 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n17107)
         );
  NAND4_X1 U20304 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_8__SCAN_IN), .A4(n17108), .ZN(n17186) );
  INV_X1 U20305 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17320) );
  NAND2_X1 U20306 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17134), .ZN(n17130) );
  NAND2_X1 U20307 ( .A1(n17113), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17112) );
  NOR2_X2 U20308 ( .A1(n18089), .A2(n17221), .ZN(n17178) );
  OAI22_X1 U20309 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17243), .B1(n17213), 
        .B2(n17113), .ZN(n17109) );
  AOI22_X1 U20310 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17178), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17109), .ZN(n17110) );
  OAI21_X1 U20311 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17112), .A(n17110), .ZN(
        P3_U2704) );
  NOR2_X2 U20312 ( .A1(n17111), .A2(n17221), .ZN(n17179) );
  AOI22_X1 U20313 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17179), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17178), .ZN(n17115) );
  OAI211_X1 U20314 ( .C1(n17113), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17221), .B(
        n17112), .ZN(n17114) );
  OAI211_X1 U20315 ( .C1(n17116), .C2(n17239), .A(n17115), .B(n17114), .ZN(
        P3_U2705) );
  AOI22_X1 U20316 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17179), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17178), .ZN(n17119) );
  OAI211_X1 U20317 ( .C1(n9658), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17221), .B(
        n17117), .ZN(n17118) );
  OAI211_X1 U20318 ( .C1(n17120), .C2(n17239), .A(n17119), .B(n17118), .ZN(
        P3_U2706) );
  INV_X1 U20319 ( .A(n17179), .ZN(n17162) );
  AOI22_X1 U20320 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n17178), .B1(n17247), .B2(
        n17121), .ZN(n17124) );
  AOI211_X1 U20321 ( .C1(n17258), .C2(n17125), .A(n9658), .B(n17213), .ZN(
        n17122) );
  INV_X1 U20322 ( .A(n17122), .ZN(n17123) );
  OAI211_X1 U20323 ( .C1(n17162), .C2(n17353), .A(n17124), .B(n17123), .ZN(
        P3_U2707) );
  AOI22_X1 U20324 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17179), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17178), .ZN(n17128) );
  OAI211_X1 U20325 ( .C1(n17126), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17221), .B(
        n17125), .ZN(n17127) );
  OAI211_X1 U20326 ( .C1(n17129), .C2(n17239), .A(n17128), .B(n17127), .ZN(
        P3_U2708) );
  AOI22_X1 U20327 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17179), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17178), .ZN(n17132) );
  OAI211_X1 U20328 ( .C1(n17134), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17221), .B(
        n17130), .ZN(n17131) );
  OAI211_X1 U20329 ( .C1(n17133), .C2(n17239), .A(n17132), .B(n17131), .ZN(
        P3_U2709) );
  AOI22_X1 U20330 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17179), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17178), .ZN(n17137) );
  AOI211_X1 U20331 ( .C1(n17326), .C2(n17139), .A(n17134), .B(n17213), .ZN(
        n17135) );
  INV_X1 U20332 ( .A(n17135), .ZN(n17136) );
  OAI211_X1 U20333 ( .C1(n17138), .C2(n17239), .A(n17137), .B(n17136), .ZN(
        P3_U2710) );
  AOI22_X1 U20334 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17179), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17178), .ZN(n17142) );
  OAI211_X1 U20335 ( .C1(n17140), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17221), .B(
        n17139), .ZN(n17141) );
  OAI211_X1 U20336 ( .C1(n17143), .C2(n17239), .A(n17142), .B(n17141), .ZN(
        P3_U2711) );
  AOI22_X1 U20337 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17179), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17178), .ZN(n17147) );
  OAI211_X1 U20338 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17145), .A(n17221), .B(
        n17144), .ZN(n17146) );
  OAI211_X1 U20339 ( .C1(n17148), .C2(n17239), .A(n17147), .B(n17146), .ZN(
        P3_U2712) );
  AOI22_X1 U20340 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17178), .B1(n17247), .B2(
        n17149), .ZN(n17152) );
  INV_X1 U20341 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17315) );
  NOR2_X1 U20342 ( .A1(n17185), .A2(n17180), .ZN(n17174) );
  NAND2_X1 U20343 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17174), .ZN(n17173) );
  NAND2_X1 U20344 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17163), .ZN(n17159) );
  NAND2_X1 U20345 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17154), .ZN(n17153) );
  OAI21_X1 U20346 ( .B1(n17320), .B2(n17213), .A(n17153), .ZN(n17150) );
  OAI21_X1 U20347 ( .B1(n17320), .B2(n17153), .A(n17150), .ZN(n17151) );
  OAI211_X1 U20348 ( .C1(n18088), .C2(n17162), .A(n17152), .B(n17151), .ZN(
        P3_U2713) );
  AOI22_X1 U20349 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17179), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17178), .ZN(n17156) );
  OAI211_X1 U20350 ( .C1(n17154), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17221), .B(
        n17153), .ZN(n17155) );
  OAI211_X1 U20351 ( .C1(n17157), .C2(n17239), .A(n17156), .B(n17155), .ZN(
        P3_U2714) );
  AOI22_X1 U20352 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17178), .B1(n17247), .B2(
        n17158), .ZN(n17161) );
  OAI211_X1 U20353 ( .C1(n17163), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17221), .B(
        n17159), .ZN(n17160) );
  OAI211_X1 U20354 ( .C1(n17162), .C2(n18080), .A(n17161), .B(n17160), .ZN(
        P3_U2715) );
  AOI22_X1 U20355 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17179), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17178), .ZN(n17166) );
  AOI211_X1 U20356 ( .C1(n17315), .C2(n17168), .A(n17163), .B(n17213), .ZN(
        n17164) );
  INV_X1 U20357 ( .A(n17164), .ZN(n17165) );
  OAI211_X1 U20358 ( .C1(n17167), .C2(n17239), .A(n17166), .B(n17165), .ZN(
        P3_U2716) );
  AOI22_X1 U20359 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17178), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n17179), .ZN(n17171) );
  OAI211_X1 U20360 ( .C1(n17169), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17221), .B(
        n17168), .ZN(n17170) );
  OAI211_X1 U20361 ( .C1(n17172), .C2(n17239), .A(n17171), .B(n17170), .ZN(
        P3_U2717) );
  AOI22_X1 U20362 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17179), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17178), .ZN(n17176) );
  OAI211_X1 U20363 ( .C1(n17174), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17221), .B(
        n17173), .ZN(n17175) );
  OAI211_X1 U20364 ( .C1(n17177), .C2(n17239), .A(n17176), .B(n17175), .ZN(
        P3_U2718) );
  AOI22_X1 U20365 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17179), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17178), .ZN(n17183) );
  OAI211_X1 U20366 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17181), .A(n17221), .B(
        n17180), .ZN(n17182) );
  OAI211_X1 U20367 ( .C1(n17184), .C2(n17239), .A(n17183), .B(n17182), .ZN(
        P3_U2719) );
  OR2_X1 U20368 ( .A1(n17185), .A2(n17186), .ZN(n17189) );
  NAND2_X1 U20369 ( .A1(n17221), .A2(n17186), .ZN(n17192) );
  AOI22_X1 U20370 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17248), .B1(n17247), .B2(
        n17187), .ZN(n17188) );
  OAI221_X1 U20371 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n17189), .C1(n17365), 
        .C2(n17192), .A(n17188), .ZN(P3_U2720) );
  INV_X1 U20372 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17281) );
  INV_X1 U20373 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17285) );
  AND4_X1 U20374 ( .A1(n18094), .A2(P3_EAX_REG_7__SCAN_IN), .A3(n17224), .A4(
        P3_EAX_REG_8__SCAN_IN), .ZN(n17212) );
  NAND2_X1 U20375 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17212), .ZN(n17208) );
  NOR2_X1 U20376 ( .A1(n17285), .A2(n17208), .ZN(n17204) );
  NAND2_X1 U20377 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17204), .ZN(n17197) );
  NOR2_X1 U20378 ( .A1(n17281), .A2(n17197), .ZN(n17200) );
  NAND2_X1 U20379 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17200), .ZN(n17193) );
  INV_X1 U20380 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17360) );
  AOI22_X1 U20381 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17248), .B1(n17247), .B2(
        n17190), .ZN(n17191) );
  OAI221_X1 U20382 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17193), .C1(n17360), 
        .C2(n17192), .A(n17191), .ZN(P3_U2721) );
  INV_X1 U20383 ( .A(n17193), .ZN(n17196) );
  AOI21_X1 U20384 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17221), .A(n17200), .ZN(
        n17195) );
  OAI222_X1 U20385 ( .A1(n17242), .A2(n17358), .B1(n17196), .B2(n17195), .C1(
        n17239), .C2(n17194), .ZN(P3_U2722) );
  INV_X1 U20386 ( .A(n17197), .ZN(n17203) );
  AOI21_X1 U20387 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17221), .A(n17203), .ZN(
        n17199) );
  OAI222_X1 U20388 ( .A1(n17242), .A2(n17353), .B1(n17200), .B2(n17199), .C1(
        n17239), .C2(n17198), .ZN(P3_U2723) );
  AOI21_X1 U20389 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17221), .A(n17204), .ZN(
        n17202) );
  OAI222_X1 U20390 ( .A1(n17242), .A2(n17351), .B1(n17203), .B2(n17202), .C1(
        n17239), .C2(n17201), .ZN(P3_U2724) );
  AOI211_X1 U20391 ( .C1(n17285), .C2(n17208), .A(n17213), .B(n17204), .ZN(
        n17205) );
  AOI21_X1 U20392 ( .B1(n17248), .B2(BUF2_REG_10__SCAN_IN), .A(n17205), .ZN(
        n17206) );
  OAI21_X1 U20393 ( .B1(n17207), .B2(n17239), .A(n17206), .ZN(P3_U2725) );
  INV_X1 U20394 ( .A(n17208), .ZN(n17211) );
  AOI21_X1 U20395 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17221), .A(n17212), .ZN(
        n17210) );
  OAI222_X1 U20396 ( .A1(n17242), .A2(n17347), .B1(n17211), .B2(n17210), .C1(
        n17239), .C2(n17209), .ZN(P3_U2726) );
  INV_X1 U20397 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17345) );
  AOI211_X1 U20398 ( .C1(n17218), .C2(n17345), .A(n17213), .B(n17212), .ZN(
        n17214) );
  AOI21_X1 U20399 ( .B1(n17248), .B2(BUF2_REG_8__SCAN_IN), .A(n17214), .ZN(
        n17215) );
  OAI21_X1 U20400 ( .B1(n17216), .B2(n17239), .A(n17215), .ZN(P3_U2727) );
  AOI22_X1 U20401 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17248), .B1(n17247), .B2(
        n17217), .ZN(n17220) );
  OAI211_X1 U20402 ( .C1(P3_EAX_REG_7__SCAN_IN), .C2(n17224), .A(n17221), .B(
        n17218), .ZN(n17219) );
  NAND2_X1 U20403 ( .A1(n17220), .A2(n17219), .ZN(P3_U2728) );
  INV_X1 U20404 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17293) );
  INV_X1 U20405 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17297) );
  INV_X1 U20406 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17336) );
  NOR3_X1 U20407 ( .A1(n17336), .A2(n17334), .A3(n17243), .ZN(n17236) );
  NAND2_X1 U20408 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17236), .ZN(n17232) );
  NOR2_X1 U20409 ( .A1(n17297), .A2(n17232), .ZN(n17235) );
  NAND2_X1 U20410 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17235), .ZN(n17225) );
  NOR2_X1 U20411 ( .A1(n17293), .A2(n17225), .ZN(n17228) );
  AOI21_X1 U20412 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17221), .A(n17228), .ZN(
        n17223) );
  OAI222_X1 U20413 ( .A1(n18088), .A2(n17242), .B1(n17224), .B2(n17223), .C1(
        n17239), .C2(n17222), .ZN(P3_U2729) );
  INV_X1 U20414 ( .A(n17225), .ZN(n17231) );
  AOI21_X1 U20415 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17221), .A(n17231), .ZN(
        n17227) );
  OAI222_X1 U20416 ( .A1(n18084), .A2(n17242), .B1(n17228), .B2(n17227), .C1(
        n17239), .C2(n17226), .ZN(P3_U2730) );
  AOI21_X1 U20417 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17221), .A(n17235), .ZN(
        n17230) );
  OAI222_X1 U20418 ( .A1(n18080), .A2(n17242), .B1(n17231), .B2(n17230), .C1(
        n17239), .C2(n17229), .ZN(P3_U2731) );
  INV_X1 U20419 ( .A(n17232), .ZN(n17241) );
  AOI21_X1 U20420 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17221), .A(n17241), .ZN(
        n17234) );
  OAI222_X1 U20421 ( .A1(n18075), .A2(n17242), .B1(n17235), .B2(n17234), .C1(
        n17239), .C2(n17233), .ZN(P3_U2732) );
  AOI21_X1 U20422 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17221), .A(n17236), .ZN(
        n17240) );
  INV_X1 U20423 ( .A(n17237), .ZN(n17238) );
  OAI222_X1 U20424 ( .A1(n18071), .A2(n17242), .B1(n17241), .B2(n17240), .C1(
        n17239), .C2(n17238), .ZN(P3_U2733) );
  OR2_X1 U20425 ( .A1(n17334), .A2(n17243), .ZN(n17251) );
  INV_X1 U20426 ( .A(n17244), .ZN(n17245) );
  AOI21_X1 U20427 ( .B1(n18094), .B2(n17334), .A(n17245), .ZN(n17250) );
  AOI22_X1 U20428 ( .A1(n17248), .A2(BUF2_REG_1__SCAN_IN), .B1(n17247), .B2(
        n17246), .ZN(n17249) );
  OAI221_X1 U20429 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17251), .C1(n17336), 
        .C2(n17250), .A(n17249), .ZN(P3_U2734) );
  INV_X1 U20430 ( .A(n17489), .ZN(n18574) );
  NOR2_X1 U20431 ( .A1(n18675), .A2(n18574), .ZN(n18713) );
  INV_X1 U20432 ( .A(n17305), .ZN(n17306) );
  NOR2_X1 U20433 ( .A1(n17276), .A2(n17253), .ZN(P3_U2736) );
  INV_X1 U20434 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17332) );
  NOR2_X1 U20435 ( .A1(n17304), .A2(n18062), .ZN(n17261) );
  AOI22_X1 U20436 ( .A1(n18713), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17254) );
  OAI21_X1 U20437 ( .B1(n17332), .B2(n17273), .A(n17254), .ZN(P3_U2737) );
  INV_X1 U20438 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17256) );
  AOI22_X1 U20439 ( .A1(n18713), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17255) );
  OAI21_X1 U20440 ( .B1(n17256), .B2(n17273), .A(n17255), .ZN(P3_U2738) );
  AOI22_X1 U20441 ( .A1(n18713), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17257) );
  OAI21_X1 U20442 ( .B1(n17258), .B2(n17273), .A(n17257), .ZN(P3_U2739) );
  INV_X1 U20443 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17260) );
  AOI22_X1 U20444 ( .A1(n18713), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17259) );
  OAI21_X1 U20445 ( .B1(n17260), .B2(n17273), .A(n17259), .ZN(P3_U2740) );
  INV_X1 U20446 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n20910) );
  AOI22_X1 U20447 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17261), .B1(n18713), 
        .B2(P3_UWORD_REG_10__SCAN_IN), .ZN(n17262) );
  OAI21_X1 U20448 ( .B1(n20910), .B2(n17276), .A(n17262), .ZN(P3_U2741) );
  CLKBUF_X1 U20449 ( .A(n18713), .Z(n17302) );
  AOI22_X1 U20450 ( .A1(n17302), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17263) );
  OAI21_X1 U20451 ( .B1(n17326), .B2(n17273), .A(n17263), .ZN(P3_U2742) );
  INV_X1 U20452 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17324) );
  AOI22_X1 U20453 ( .A1(n18713), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17264) );
  OAI21_X1 U20454 ( .B1(n17324), .B2(n17273), .A(n17264), .ZN(P3_U2743) );
  INV_X1 U20455 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17322) );
  AOI22_X1 U20456 ( .A1(n17302), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17265) );
  OAI21_X1 U20457 ( .B1(n17322), .B2(n17273), .A(n17265), .ZN(P3_U2744) );
  AOI22_X1 U20458 ( .A1(n17302), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17266) );
  OAI21_X1 U20459 ( .B1(n17320), .B2(n17273), .A(n17266), .ZN(P3_U2745) );
  AOI22_X1 U20460 ( .A1(n17302), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17267) );
  OAI21_X1 U20461 ( .B1(n20819), .B2(n17273), .A(n17267), .ZN(P3_U2746) );
  INV_X1 U20462 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17317) );
  AOI22_X1 U20463 ( .A1(n17302), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17268) );
  OAI21_X1 U20464 ( .B1(n17317), .B2(n17273), .A(n17268), .ZN(P3_U2747) );
  AOI22_X1 U20465 ( .A1(n17302), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17269) );
  OAI21_X1 U20466 ( .B1(n17315), .B2(n17273), .A(n17269), .ZN(P3_U2748) );
  INV_X1 U20467 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17313) );
  AOI22_X1 U20468 ( .A1(n17302), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17270) );
  OAI21_X1 U20469 ( .B1(n17313), .B2(n17273), .A(n17270), .ZN(P3_U2749) );
  INV_X1 U20470 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17311) );
  INV_X2 U20471 ( .A(n17276), .ZN(n17301) );
  AOI22_X1 U20472 ( .A1(n17302), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17271) );
  OAI21_X1 U20473 ( .B1(n17311), .B2(n17273), .A(n17271), .ZN(P3_U2750) );
  INV_X1 U20474 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17309) );
  AOI22_X1 U20475 ( .A1(n17302), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17272) );
  OAI21_X1 U20476 ( .B1(n17309), .B2(n17273), .A(n17272), .ZN(P3_U2751) );
  INV_X1 U20477 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n20881) );
  AOI22_X1 U20478 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n17274), .B1(n18713), 
        .B2(P3_LWORD_REG_15__SCAN_IN), .ZN(n17275) );
  OAI21_X1 U20479 ( .B1(n20881), .B2(n17276), .A(n17275), .ZN(P3_U2752) );
  AOI22_X1 U20480 ( .A1(n17302), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17277) );
  OAI21_X1 U20481 ( .B1(n17360), .B2(n17304), .A(n17277), .ZN(P3_U2753) );
  INV_X1 U20482 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17279) );
  AOI22_X1 U20483 ( .A1(n17302), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17278) );
  OAI21_X1 U20484 ( .B1(n17279), .B2(n17304), .A(n17278), .ZN(P3_U2754) );
  AOI22_X1 U20485 ( .A1(n17302), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17280) );
  OAI21_X1 U20486 ( .B1(n17281), .B2(n17304), .A(n17280), .ZN(P3_U2755) );
  INV_X1 U20487 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17283) );
  AOI22_X1 U20488 ( .A1(n17302), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17282) );
  OAI21_X1 U20489 ( .B1(n17283), .B2(n17304), .A(n17282), .ZN(P3_U2756) );
  AOI22_X1 U20490 ( .A1(n17302), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17284) );
  OAI21_X1 U20491 ( .B1(n17285), .B2(n17304), .A(n17284), .ZN(P3_U2757) );
  INV_X1 U20492 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U20493 ( .A1(n17302), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17286) );
  OAI21_X1 U20494 ( .B1(n17287), .B2(n17304), .A(n17286), .ZN(P3_U2758) );
  AOI22_X1 U20495 ( .A1(n17302), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17288) );
  OAI21_X1 U20496 ( .B1(n17345), .B2(n17304), .A(n17288), .ZN(P3_U2759) );
  INV_X1 U20497 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17343) );
  AOI22_X1 U20498 ( .A1(n17302), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17289) );
  OAI21_X1 U20499 ( .B1(n17343), .B2(n17304), .A(n17289), .ZN(P3_U2760) );
  INV_X1 U20500 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17291) );
  AOI22_X1 U20501 ( .A1(n17302), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17290) );
  OAI21_X1 U20502 ( .B1(n17291), .B2(n17304), .A(n17290), .ZN(P3_U2761) );
  AOI22_X1 U20503 ( .A1(n17302), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17292) );
  OAI21_X1 U20504 ( .B1(n17293), .B2(n17304), .A(n17292), .ZN(P3_U2762) );
  INV_X1 U20505 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17295) );
  AOI22_X1 U20506 ( .A1(n17302), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17294) );
  OAI21_X1 U20507 ( .B1(n17295), .B2(n17304), .A(n17294), .ZN(P3_U2763) );
  AOI22_X1 U20508 ( .A1(n17302), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17296) );
  OAI21_X1 U20509 ( .B1(n17297), .B2(n17304), .A(n17296), .ZN(P3_U2764) );
  INV_X1 U20510 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17299) );
  AOI22_X1 U20511 ( .A1(n17302), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17298) );
  OAI21_X1 U20512 ( .B1(n17299), .B2(n17304), .A(n17298), .ZN(P3_U2765) );
  AOI22_X1 U20513 ( .A1(n17302), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17300) );
  OAI21_X1 U20514 ( .B1(n17336), .B2(n17304), .A(n17300), .ZN(P3_U2766) );
  AOI22_X1 U20515 ( .A1(n17302), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17301), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17303) );
  OAI21_X1 U20516 ( .B1(n17334), .B2(n17304), .A(n17303), .ZN(P3_U2767) );
  NOR2_X2 U20517 ( .A1(n17305), .A2(n18555), .ZN(n17355) );
  NOR2_X2 U20518 ( .A1(n18716), .A2(n17354), .ZN(n17362) );
  AOI22_X1 U20519 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17354), .ZN(n17308) );
  OAI21_X1 U20520 ( .B1(n17309), .B2(n17364), .A(n17308), .ZN(P3_U2768) );
  AOI22_X1 U20521 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17354), .ZN(n17310) );
  OAI21_X1 U20522 ( .B1(n17311), .B2(n17364), .A(n17310), .ZN(P3_U2769) );
  AOI22_X1 U20523 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17354), .ZN(n17312) );
  OAI21_X1 U20524 ( .B1(n17313), .B2(n17364), .A(n17312), .ZN(P3_U2770) );
  AOI22_X1 U20525 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17354), .ZN(n17314) );
  OAI21_X1 U20526 ( .B1(n17315), .B2(n17364), .A(n17314), .ZN(P3_U2771) );
  AOI22_X1 U20527 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17354), .ZN(n17316) );
  OAI21_X1 U20528 ( .B1(n17317), .B2(n17364), .A(n17316), .ZN(P3_U2772) );
  AOI22_X1 U20529 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17354), .ZN(n17318) );
  OAI21_X1 U20530 ( .B1(n20819), .B2(n17364), .A(n17318), .ZN(P3_U2773) );
  AOI22_X1 U20531 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17354), .ZN(n17319) );
  OAI21_X1 U20532 ( .B1(n17320), .B2(n17364), .A(n17319), .ZN(P3_U2774) );
  AOI22_X1 U20533 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17354), .ZN(n17321) );
  OAI21_X1 U20534 ( .B1(n17322), .B2(n17364), .A(n17321), .ZN(P3_U2775) );
  AOI22_X1 U20535 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17354), .ZN(n17323) );
  OAI21_X1 U20536 ( .B1(n17324), .B2(n17364), .A(n17323), .ZN(P3_U2776) );
  AOI22_X1 U20537 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17354), .ZN(n17325) );
  OAI21_X1 U20538 ( .B1(n17326), .B2(n17364), .A(n17325), .ZN(P3_U2777) );
  AOI22_X1 U20539 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17355), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17354), .ZN(n17327) );
  OAI21_X1 U20540 ( .B1(n17349), .B2(n17357), .A(n17327), .ZN(P3_U2778) );
  AOI22_X1 U20541 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17355), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17354), .ZN(n17328) );
  OAI21_X1 U20542 ( .B1(n17351), .B2(n17357), .A(n17328), .ZN(P3_U2779) );
  AOI22_X1 U20543 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17355), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17354), .ZN(n17329) );
  OAI21_X1 U20544 ( .B1(n17353), .B2(n17357), .A(n17329), .ZN(P3_U2780) );
  AOI22_X1 U20545 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17355), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17354), .ZN(n17330) );
  OAI21_X1 U20546 ( .B1(n17358), .B2(n17357), .A(n17330), .ZN(P3_U2781) );
  AOI22_X1 U20547 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17354), .ZN(n17331) );
  OAI21_X1 U20548 ( .B1(n17332), .B2(n17364), .A(n17331), .ZN(P3_U2782) );
  AOI22_X1 U20549 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17362), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17354), .ZN(n17333) );
  OAI21_X1 U20550 ( .B1(n17334), .B2(n17364), .A(n17333), .ZN(P3_U2783) );
  AOI22_X1 U20551 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17362), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17354), .ZN(n17335) );
  OAI21_X1 U20552 ( .B1(n17336), .B2(n17364), .A(n17335), .ZN(P3_U2784) );
  AOI22_X1 U20553 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17355), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17354), .ZN(n17337) );
  OAI21_X1 U20554 ( .B1(n18071), .B2(n17357), .A(n17337), .ZN(P3_U2785) );
  AOI22_X1 U20555 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17355), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17354), .ZN(n17338) );
  OAI21_X1 U20556 ( .B1(n18075), .B2(n17357), .A(n17338), .ZN(P3_U2786) );
  AOI22_X1 U20557 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17355), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17361), .ZN(n17339) );
  OAI21_X1 U20558 ( .B1(n18080), .B2(n17357), .A(n17339), .ZN(P3_U2787) );
  AOI22_X1 U20559 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17355), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17361), .ZN(n17340) );
  OAI21_X1 U20560 ( .B1(n18084), .B2(n17357), .A(n17340), .ZN(P3_U2788) );
  AOI22_X1 U20561 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17355), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17361), .ZN(n17341) );
  OAI21_X1 U20562 ( .B1(n18088), .B2(n17357), .A(n17341), .ZN(P3_U2789) );
  AOI22_X1 U20563 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17362), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17361), .ZN(n17342) );
  OAI21_X1 U20564 ( .B1(n17343), .B2(n17364), .A(n17342), .ZN(P3_U2790) );
  AOI22_X1 U20565 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17362), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17361), .ZN(n17344) );
  OAI21_X1 U20566 ( .B1(n17345), .B2(n17364), .A(n17344), .ZN(P3_U2791) );
  AOI22_X1 U20567 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17355), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17361), .ZN(n17346) );
  OAI21_X1 U20568 ( .B1(n17347), .B2(n17357), .A(n17346), .ZN(P3_U2792) );
  AOI22_X1 U20569 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17355), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17361), .ZN(n17348) );
  OAI21_X1 U20570 ( .B1(n17349), .B2(n17357), .A(n17348), .ZN(P3_U2793) );
  AOI22_X1 U20571 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17355), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17361), .ZN(n17350) );
  OAI21_X1 U20572 ( .B1(n17351), .B2(n17357), .A(n17350), .ZN(P3_U2794) );
  AOI22_X1 U20573 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17355), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17354), .ZN(n17352) );
  OAI21_X1 U20574 ( .B1(n17353), .B2(n17357), .A(n17352), .ZN(P3_U2795) );
  AOI22_X1 U20575 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17355), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17354), .ZN(n17356) );
  OAI21_X1 U20576 ( .B1(n17358), .B2(n17357), .A(n17356), .ZN(P3_U2796) );
  AOI22_X1 U20577 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17362), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17361), .ZN(n17359) );
  OAI21_X1 U20578 ( .B1(n17360), .B2(n17364), .A(n17359), .ZN(P3_U2797) );
  AOI22_X1 U20579 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17362), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17361), .ZN(n17363) );
  OAI21_X1 U20580 ( .B1(n17365), .B2(n17364), .A(n17363), .ZN(P3_U2798) );
  NOR3_X1 U20581 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17527), .A3(
        n17366), .ZN(n17375) );
  AND3_X1 U20582 ( .A1(n17367), .A2(n17579), .A3(n17368), .ZN(n17389) );
  OAI21_X1 U20583 ( .B1(n17368), .B2(n17632), .A(n17735), .ZN(n17369) );
  AOI21_X1 U20584 ( .B1(n17489), .B2(n17370), .A(n17369), .ZN(n17395) );
  OAI21_X1 U20585 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17482), .A(
        n17395), .ZN(n17390) );
  OAI21_X1 U20586 ( .B1(n17389), .B2(n17390), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17372) );
  NAND2_X1 U20587 ( .A1(n18038), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17371) );
  OAI211_X1 U20588 ( .C1(n17566), .C2(n17373), .A(n17372), .B(n17371), .ZN(
        n17374) );
  AOI211_X1 U20589 ( .C1(n17376), .C2(n17428), .A(n17375), .B(n17374), .ZN(
        n17382) );
  NAND2_X1 U20590 ( .A1(n17646), .A2(n17739), .ZN(n17475) );
  AOI22_X1 U20591 ( .A1(n17598), .A2(n17745), .B1(n17727), .B2(n17746), .ZN(
        n17405) );
  NAND2_X1 U20592 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17405), .ZN(
        n17391) );
  NAND3_X1 U20593 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17475), .A3(
        n17391), .ZN(n17381) );
  OAI211_X1 U20594 ( .C1(n17379), .C2(n17378), .A(n17615), .B(n17377), .ZN(
        n17380) );
  NAND3_X1 U20595 ( .A1(n17382), .A2(n17381), .A3(n17380), .ZN(P3_U2802) );
  NOR2_X1 U20596 ( .A1(n17384), .A2(n17383), .ZN(n17385) );
  XNOR2_X1 U20597 ( .A(n17385), .B(n17639), .ZN(n17755) );
  INV_X1 U20598 ( .A(n17386), .ZN(n17387) );
  OAI22_X1 U20599 ( .A1(n18048), .A2(n18643), .B1(n17566), .B2(n17387), .ZN(
        n17388) );
  AOI211_X1 U20600 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17390), .A(
        n17389), .B(n17388), .ZN(n17394) );
  OAI21_X1 U20601 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17392), .A(
        n17391), .ZN(n17393) );
  OAI211_X1 U20602 ( .C1(n17755), .C2(n17642), .A(n17394), .B(n17393), .ZN(
        P3_U2803) );
  NAND2_X1 U20603 ( .A1(n17566), .A2(n17482), .ZN(n17729) );
  NOR2_X1 U20604 ( .A1(n18048), .A2(n18641), .ZN(n17760) );
  AOI221_X1 U20605 ( .B1(n17397), .B2(n17396), .C1(n18204), .C2(n17396), .A(
        n17395), .ZN(n17398) );
  AOI211_X1 U20606 ( .C1(n17399), .C2(n17729), .A(n17760), .B(n17398), .ZN(
        n17403) );
  OAI21_X1 U20607 ( .B1(n17401), .B2(n17404), .A(n17400), .ZN(n17759) );
  NOR3_X1 U20608 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17764), .A3(
        n17742), .ZN(n17756) );
  AOI22_X1 U20609 ( .A1(n17615), .A2(n17759), .B1(n17428), .B2(n17756), .ZN(
        n17402) );
  OAI211_X1 U20610 ( .C1(n17405), .C2(n17404), .A(n17403), .B(n17402), .ZN(
        P3_U2804) );
  NAND2_X1 U20611 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17423), .ZN(
        n17765) );
  INV_X1 U20612 ( .A(n17765), .ZN(n17767) );
  NAND2_X1 U20613 ( .A1(n17767), .A2(n17871), .ZN(n17406) );
  XNOR2_X1 U20614 ( .A(n17406), .B(n17764), .ZN(n17777) );
  INV_X1 U20615 ( .A(n17735), .ZN(n17722) );
  NOR2_X1 U20616 ( .A1(n17408), .A2(n18204), .ZN(n17435) );
  AOI211_X1 U20617 ( .C1(n17489), .C2(n17407), .A(n17722), .B(n17435), .ZN(
        n17438) );
  OAI21_X1 U20618 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17482), .A(
        n17438), .ZN(n17420) );
  NOR2_X1 U20619 ( .A1(n18048), .A2(n18639), .ZN(n17772) );
  AND2_X1 U20620 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17411) );
  OAI211_X1 U20621 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17408), .B(n17579), .ZN(n17410) );
  OAI22_X1 U20622 ( .A1(n17411), .A2(n17410), .B1(n17409), .B2(n17566), .ZN(
        n17412) );
  AOI211_X1 U20623 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17420), .A(
        n17772), .B(n17412), .ZN(n17418) );
  AND2_X1 U20624 ( .A1(n17870), .A2(n17767), .ZN(n17413) );
  XNOR2_X1 U20625 ( .A(n17413), .B(n17764), .ZN(n17774) );
  AOI21_X1 U20626 ( .B1(n17608), .B2(n17415), .A(n17414), .ZN(n17416) );
  XNOR2_X1 U20627 ( .A(n17416), .B(n17764), .ZN(n17773) );
  AOI22_X1 U20628 ( .A1(n17727), .A2(n17774), .B1(n17615), .B2(n17773), .ZN(
        n17417) );
  OAI211_X1 U20629 ( .C1(n17646), .C2(n17777), .A(n17418), .B(n17417), .ZN(
        P3_U2805) );
  NOR2_X1 U20630 ( .A1(n17527), .A2(n9917), .ZN(n17422) );
  NOR2_X1 U20631 ( .A1(n18048), .A2(n18636), .ZN(n17778) );
  AOI221_X1 U20632 ( .B1(n17422), .B2(n17421), .C1(n17420), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17778), .ZN(n17430) );
  NOR2_X1 U20633 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17792), .ZN(
        n17780) );
  NAND2_X1 U20634 ( .A1(n17871), .A2(n17423), .ZN(n17781) );
  NAND2_X1 U20635 ( .A1(n17870), .A2(n17423), .ZN(n17783) );
  AOI22_X1 U20636 ( .A1(n17598), .A2(n17781), .B1(n17727), .B2(n17783), .ZN(
        n17441) );
  INV_X1 U20637 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17426) );
  AOI21_X1 U20638 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17425), .A(
        n17424), .ZN(n17791) );
  OAI22_X1 U20639 ( .A1(n17441), .A2(n17426), .B1(n17791), .B2(n17642), .ZN(
        n17427) );
  AOI21_X1 U20640 ( .B1(n17428), .B2(n17780), .A(n17427), .ZN(n17429) );
  OAI211_X1 U20641 ( .C1(n17566), .C2(n9911), .A(n17430), .B(n17429), .ZN(
        P3_U2806) );
  AOI22_X1 U20642 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17639), .B1(
        n17452), .B2(n17431), .ZN(n17432) );
  NAND2_X1 U20643 ( .A1(n17476), .A2(n17432), .ZN(n17433) );
  XNOR2_X1 U20644 ( .A(n17433), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17796) );
  AOI22_X1 U20645 ( .A1(n9705), .A2(n17435), .B1(n17434), .B2(n17729), .ZN(
        n17436) );
  NAND2_X1 U20646 ( .A1(n18038), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17797) );
  OAI211_X1 U20647 ( .C1(n17438), .C2(n17437), .A(n17436), .B(n17797), .ZN(
        n17439) );
  AOI21_X1 U20648 ( .B1(n17615), .B2(n17796), .A(n17439), .ZN(n17440) );
  OAI221_X1 U20649 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17442), 
        .C1(n17792), .C2(n17441), .A(n17440), .ZN(P3_U2807) );
  INV_X1 U20650 ( .A(n17482), .ZN(n17446) );
  AOI21_X1 U20651 ( .B1(n17489), .B2(n17443), .A(n17722), .ZN(n17444) );
  OAI21_X1 U20652 ( .B1(n17447), .B2(n17632), .A(n17444), .ZN(n17480) );
  AOI21_X1 U20653 ( .B1(n17446), .B2(n17445), .A(n17480), .ZN(n17461) );
  NOR2_X1 U20654 ( .A1(n18048), .A2(n18632), .ZN(n17799) );
  NAND2_X1 U20655 ( .A1(n17447), .A2(n17579), .ZN(n17463) );
  AOI221_X1 U20656 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n17462), .C2(n17460), .A(
        n17463), .ZN(n17448) );
  AOI211_X1 U20657 ( .C1(n17449), .C2(n17582), .A(n17799), .B(n17448), .ZN(
        n17459) );
  INV_X1 U20658 ( .A(n17450), .ZN(n17522) );
  OR2_X1 U20659 ( .A1(n17469), .A2(n17472), .ZN(n17805) );
  INV_X1 U20660 ( .A(n17476), .ZN(n17451) );
  AOI221_X1 U20661 ( .B1(n17522), .B2(n17452), .C1(n17805), .C2(n17452), .A(
        n17451), .ZN(n17453) );
  XNOR2_X1 U20662 ( .A(n17453), .B(n17811), .ZN(n17800) );
  NOR2_X1 U20663 ( .A1(n17454), .A2(n17805), .ZN(n17456) );
  OAI22_X1 U20664 ( .A1(n17871), .A2(n17646), .B1(n17870), .B2(n17739), .ZN(
        n17532) );
  AOI21_X1 U20665 ( .B1(n17475), .B2(n17805), .A(n17532), .ZN(n17473) );
  INV_X1 U20666 ( .A(n17473), .ZN(n17455) );
  MUX2_X1 U20667 ( .A(n17456), .B(n17455), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17457) );
  AOI21_X1 U20668 ( .B1(n17615), .B2(n17800), .A(n17457), .ZN(n17458) );
  OAI211_X1 U20669 ( .C1(n17461), .C2(n17460), .A(n17459), .B(n17458), .ZN(
        P3_U2808) );
  NAND2_X1 U20670 ( .A1(n18038), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n17820) );
  OAI221_X1 U20671 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17463), .C1(
        n17462), .C2(n17461), .A(n17820), .ZN(n17464) );
  AOI21_X1 U20672 ( .B1(n17582), .B2(n17465), .A(n17464), .ZN(n17471) );
  NOR3_X1 U20673 ( .A1(n17639), .A2(n17850), .A3(n17466), .ZN(n17494) );
  INV_X1 U20674 ( .A(n17507), .ZN(n17495) );
  AOI22_X1 U20675 ( .A1(n17815), .A2(n17494), .B1(n17467), .B2(n17495), .ZN(
        n17468) );
  XNOR2_X1 U20676 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17468), .ZN(
        n17813) );
  NOR2_X1 U20677 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17469), .ZN(
        n17812) );
  AOI22_X1 U20678 ( .A1(n17615), .A2(n17813), .B1(n17533), .B2(n17812), .ZN(
        n17470) );
  OAI211_X1 U20679 ( .C1(n17473), .C2(n17472), .A(n17471), .B(n17470), .ZN(
        P3_U2809) );
  NAND2_X1 U20680 ( .A1(n17474), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17824) );
  NOR2_X1 U20681 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17824), .ZN(
        n17829) );
  AOI21_X1 U20682 ( .B1(n17475), .B2(n17824), .A(n17532), .ZN(n17500) );
  OAI221_X1 U20683 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17506), 
        .C1(n17839), .C2(n17494), .A(n17476), .ZN(n17477) );
  XNOR2_X1 U20684 ( .A(n17478), .B(n17477), .ZN(n17833) );
  OAI22_X1 U20685 ( .A1(n17500), .A2(n17478), .B1(n17642), .B2(n17833), .ZN(
        n17479) );
  AOI21_X1 U20686 ( .B1(n17533), .B2(n17829), .A(n17479), .ZN(n17486) );
  NAND2_X1 U20687 ( .A1(n18038), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17831) );
  OAI221_X1 U20688 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17481), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n18374), .A(n17480), .ZN(
        n17485) );
  OAI21_X1 U20689 ( .B1(n17582), .B2(n17446), .A(n17483), .ZN(n17484) );
  NAND4_X1 U20690 ( .A1(n17486), .A2(n17831), .A3(n17485), .A4(n17484), .ZN(
        P3_U2810) );
  NAND2_X1 U20691 ( .A1(n17487), .A2(n17579), .ZN(n17503) );
  AOI221_X1 U20692 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C1(n17502), .C2(n17491), .A(
        n17503), .ZN(n17493) );
  OAI21_X1 U20693 ( .B1(n17487), .B2(n17632), .A(n17735), .ZN(n17514) );
  AOI21_X1 U20694 ( .B1(n17489), .B2(n17488), .A(n17514), .ZN(n17501) );
  OAI22_X1 U20695 ( .A1(n17501), .A2(n17491), .B1(n17566), .B2(n17490), .ZN(
        n17492) );
  AOI211_X1 U20696 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n18038), .A(n17493), 
        .B(n17492), .ZN(n17499) );
  AOI21_X1 U20697 ( .B1(n17495), .B2(n17506), .A(n17494), .ZN(n17496) );
  XNOR2_X1 U20698 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n17496), .ZN(
        n17835) );
  NOR2_X1 U20699 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17497), .ZN(
        n17834) );
  AOI22_X1 U20700 ( .A1(n17615), .A2(n17835), .B1(n17533), .B2(n17834), .ZN(
        n17498) );
  OAI211_X1 U20701 ( .C1(n17500), .C2(n17839), .A(n17499), .B(n17498), .ZN(
        P3_U2811) );
  AOI21_X1 U20702 ( .B1(n17533), .B2(n17842), .A(n17532), .ZN(n17520) );
  NAND2_X1 U20703 ( .A1(n18038), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17847) );
  OAI221_X1 U20704 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17503), .C1(
        n17502), .C2(n17501), .A(n17847), .ZN(n17504) );
  AOI21_X1 U20705 ( .B1(n17582), .B2(n17505), .A(n17504), .ZN(n17510) );
  AOI21_X1 U20706 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17608), .A(
        n17506), .ZN(n17508) );
  XNOR2_X1 U20707 ( .A(n17508), .B(n17507), .ZN(n17846) );
  NOR2_X1 U20708 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17842), .ZN(
        n17845) );
  AOI22_X1 U20709 ( .A1(n17615), .A2(n17846), .B1(n17533), .B2(n17845), .ZN(
        n17509) );
  OAI211_X1 U20710 ( .C1(n17520), .C2(n17850), .A(n17510), .B(n17509), .ZN(
        P3_U2812) );
  AOI21_X1 U20711 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17533), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17519) );
  OAI21_X1 U20712 ( .B1(n17512), .B2(n18204), .A(n17511), .ZN(n17513) );
  AOI22_X1 U20713 ( .A1(n18038), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n17514), 
        .B2(n17513), .ZN(n17518) );
  OAI21_X1 U20714 ( .B1(n9704), .B2(n17853), .A(n17515), .ZN(n17851) );
  AOI22_X1 U20715 ( .A1(n17615), .A2(n17851), .B1(n17516), .B2(n17729), .ZN(
        n17517) );
  OAI211_X1 U20716 ( .C1(n17520), .C2(n17519), .A(n17518), .B(n17517), .ZN(
        P3_U2813) );
  AOI22_X1 U20717 ( .A1(n17639), .A2(n17522), .B1(n17618), .B2(n17521), .ZN(
        n17523) );
  XNOR2_X1 U20718 ( .A(n17865), .B(n17523), .ZN(n17869) );
  AOI21_X1 U20719 ( .B1(n17687), .B2(n17526), .A(n17722), .ZN(n17550) );
  OAI21_X1 U20720 ( .B1(n17524), .B2(n18574), .A(n17550), .ZN(n17541) );
  AOI22_X1 U20721 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17541), .B1(
        n17582), .B2(n17525), .ZN(n17530) );
  NOR2_X1 U20722 ( .A1(n17527), .A2(n17526), .ZN(n17543) );
  OAI211_X1 U20723 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17543), .B(n17528), .ZN(n17529) );
  OAI211_X1 U20724 ( .C1(n18620), .C2(n18048), .A(n17530), .B(n17529), .ZN(
        n17531) );
  AOI221_X1 U20725 ( .B1(n17533), .B2(n17865), .C1(n17532), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n17531), .ZN(n17534) );
  OAI21_X1 U20726 ( .B1(n17869), .B2(n17642), .A(n17534), .ZN(P3_U2814) );
  NAND3_X1 U20727 ( .A1(n17929), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n17535), .ZN(n17537) );
  NOR2_X1 U20728 ( .A1(n17608), .A2(n12542), .ZN(n17619) );
  NAND3_X1 U20729 ( .A1(n17612), .A2(n17619), .A3(n17591), .ZN(n17576) );
  INV_X1 U20730 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17892) );
  INV_X1 U20731 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17588) );
  AOI22_X1 U20732 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17608), .B1(
        n17892), .B2(n17588), .ZN(n17536) );
  AOI221_X1 U20733 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n17537), 
        .C1(n17573), .C2(n17576), .A(n17536), .ZN(n17538) );
  XNOR2_X1 U20734 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17538), .ZN(
        n17878) );
  OAI22_X1 U20735 ( .A1(n18048), .A2(n18618), .B1(n17566), .B2(n17539), .ZN(
        n17540) );
  AOI221_X1 U20736 ( .B1(n17543), .B2(n17542), .C1(n17541), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17540), .ZN(n17547) );
  NOR2_X1 U20737 ( .A1(n17870), .A2(n17739), .ZN(n17545) );
  NOR2_X1 U20738 ( .A1(n17563), .A2(n17922), .ZN(n17571) );
  INV_X1 U20739 ( .A(n17571), .ZN(n17908) );
  NOR2_X1 U20740 ( .A1(n17573), .A2(n17908), .ZN(n17549) );
  NAND2_X1 U20741 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17549), .ZN(
        n17548) );
  NAND2_X1 U20742 ( .A1(n17885), .A2(n17548), .ZN(n17881) );
  NOR2_X1 U20743 ( .A1(n17871), .A2(n17646), .ZN(n17544) );
  OAI21_X1 U20744 ( .B1(n17555), .B2(n17920), .A(n17885), .ZN(n17876) );
  AOI22_X1 U20745 ( .A1(n17545), .A2(n17881), .B1(n17544), .B2(n17876), .ZN(
        n17546) );
  OAI211_X1 U20746 ( .C1(n17642), .C2(n17878), .A(n17547), .B(n17546), .ZN(
        P3_U2815) );
  OAI21_X1 U20747 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17549), .A(
        n17548), .ZN(n17900) );
  AOI221_X1 U20748 ( .B1(n17552), .B2(n17551), .C1(n18204), .C2(n17551), .A(
        n17550), .ZN(n17553) );
  NOR2_X1 U20749 ( .A1(n18048), .A2(n18616), .ZN(n17894) );
  AOI211_X1 U20750 ( .C1(n17554), .C2(n17729), .A(n17553), .B(n17894), .ZN(
        n17562) );
  INV_X1 U20751 ( .A(n17555), .ZN(n17859) );
  INV_X1 U20752 ( .A(n17920), .ZN(n17557) );
  NOR2_X1 U20753 ( .A1(n17920), .A2(n17563), .ZN(n17905) );
  AOI21_X1 U20754 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n17905), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17556) );
  AOI21_X1 U20755 ( .B1(n17859), .B2(n17557), .A(n17556), .ZN(n17896) );
  INV_X1 U20756 ( .A(n17576), .ZN(n17558) );
  AOI22_X1 U20757 ( .A1(n17887), .A2(n17618), .B1(n17559), .B2(n17558), .ZN(
        n17560) );
  XNOR2_X1 U20758 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17560), .ZN(
        n17895) );
  AOI22_X1 U20759 ( .A1(n17598), .A2(n17896), .B1(n17615), .B2(n17895), .ZN(
        n17561) );
  OAI211_X1 U20760 ( .C1(n17739), .C2(n17900), .A(n17562), .B(n17561), .ZN(
        P3_U2816) );
  INV_X1 U20761 ( .A(n17563), .ZN(n17886) );
  NAND2_X1 U20762 ( .A1(n17886), .A2(n17573), .ZN(n17912) );
  OR2_X1 U20763 ( .A1(n17632), .A2(n17580), .ZN(n17564) );
  OAI211_X1 U20764 ( .C1(n17565), .C2(n18574), .A(n17564), .B(n17735), .ZN(
        n17583) );
  NOR2_X1 U20765 ( .A1(n18048), .A2(n18614), .ZN(n17570) );
  OAI211_X1 U20766 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17580), .B(n17579), .ZN(n17568) );
  OAI22_X1 U20767 ( .A1(n10031), .A2(n17568), .B1(n17567), .B2(n17566), .ZN(
        n17569) );
  AOI211_X1 U20768 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17583), .A(
        n17570), .B(n17569), .ZN(n17575) );
  OAI22_X1 U20769 ( .A1(n17571), .A2(n17739), .B1(n17905), .B2(n17646), .ZN(
        n17587) );
  NAND2_X1 U20770 ( .A1(n17929), .A2(n17618), .ZN(n17577) );
  AOI22_X1 U20771 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17577), .B1(
        n17576), .B2(n17588), .ZN(n17572) );
  XNOR2_X1 U20772 ( .A(n17573), .B(n17572), .ZN(n17903) );
  AOI22_X1 U20773 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17587), .B1(
        n17615), .B2(n17903), .ZN(n17574) );
  OAI211_X1 U20774 ( .C1(n17624), .C2(n17912), .A(n17575), .B(n17574), .ZN(
        P3_U2817) );
  NAND2_X1 U20775 ( .A1(n17577), .A2(n17576), .ZN(n17578) );
  XNOR2_X1 U20776 ( .A(n17578), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17918) );
  AND2_X1 U20777 ( .A1(n17599), .A2(n17929), .ZN(n17589) );
  NAND2_X1 U20778 ( .A1(n17580), .A2(n17579), .ZN(n17585) );
  AOI22_X1 U20779 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17583), .B1(
        n17582), .B2(n17581), .ZN(n17584) );
  NAND2_X1 U20780 ( .A1(n18038), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n17916) );
  OAI211_X1 U20781 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17585), .A(
        n17584), .B(n17916), .ZN(n17586) );
  AOI221_X1 U20782 ( .B1(n17589), .B2(n17588), .C1(n17587), .C2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17586), .ZN(n17590) );
  OAI21_X1 U20783 ( .B1(n17918), .B2(n17642), .A(n17590), .ZN(P3_U2818) );
  INV_X1 U20784 ( .A(n17926), .ZN(n17611) );
  AOI22_X1 U20785 ( .A1(n17611), .A2(n17618), .B1(n17612), .B2(n17619), .ZN(
        n17592) );
  XNOR2_X1 U20786 ( .A(n17592), .B(n17591), .ZN(n17933) );
  NAND3_X1 U20787 ( .A1(n17633), .A2(n17593), .A3(n18374), .ZN(n17629) );
  NOR2_X1 U20788 ( .A1(n17604), .A2(n17629), .ZN(n17603) );
  NOR2_X1 U20789 ( .A1(n17596), .A2(n17603), .ZN(n17597) );
  OAI22_X1 U20790 ( .A1(n17719), .A2(n17594), .B1(n18048), .B2(n18610), .ZN(
        n17595) );
  AOI221_X1 U20791 ( .B1(n17730), .B2(n17597), .C1(n17596), .C2(n17603), .A(
        n17595), .ZN(n17602) );
  AOI22_X1 U20792 ( .A1(n17598), .A2(n17920), .B1(n17727), .B2(n17922), .ZN(
        n17625) );
  OAI21_X1 U20793 ( .B1(n17611), .B2(n17624), .A(n17625), .ZN(n17600) );
  NOR2_X1 U20794 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17926), .ZN(
        n17919) );
  AOI22_X1 U20795 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17600), .B1(
        n17919), .B2(n17599), .ZN(n17601) );
  OAI211_X1 U20796 ( .C1(n17933), .C2(n17642), .A(n17602), .B(n17601), .ZN(
        P3_U2819) );
  INV_X1 U20797 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17934) );
  INV_X1 U20798 ( .A(n17730), .ZN(n17665) );
  AOI211_X1 U20799 ( .C1(n17629), .C2(n17604), .A(n17665), .B(n17603), .ZN(
        n17606) );
  INV_X1 U20800 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18608) );
  NOR2_X1 U20801 ( .A1(n18048), .A2(n18608), .ZN(n17605) );
  AOI211_X1 U20802 ( .C1(n17607), .C2(n17729), .A(n17606), .B(n17605), .ZN(
        n17617) );
  NOR4_X1 U20803 ( .A1(n17608), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17535), .A4(n17934), .ZN(n17610) );
  INV_X1 U20804 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17623) );
  AOI221_X1 U20805 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17618), .C1(
        n17623), .C2(n17619), .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17609) );
  AOI211_X1 U20806 ( .C1(n17618), .C2(n17611), .A(n17610), .B(n17609), .ZN(
        n17935) );
  NOR2_X1 U20807 ( .A1(n17611), .A2(n17624), .ZN(n17614) );
  INV_X1 U20808 ( .A(n17612), .ZN(n17613) );
  AOI22_X1 U20809 ( .A1(n17615), .A2(n17935), .B1(n17614), .B2(n17613), .ZN(
        n17616) );
  OAI211_X1 U20810 ( .C1(n17625), .C2(n17934), .A(n17617), .B(n17616), .ZN(
        P3_U2820) );
  NOR2_X1 U20811 ( .A1(n17619), .A2(n17618), .ZN(n17620) );
  XNOR2_X1 U20812 ( .A(n17620), .B(n17623), .ZN(n17950) );
  NAND2_X1 U20813 ( .A1(n17633), .A2(n18374), .ZN(n17649) );
  OAI22_X1 U20814 ( .A1(n17665), .A2(n17621), .B1(n17634), .B2(n17649), .ZN(
        n17628) );
  NAND2_X1 U20815 ( .A1(n18038), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n17948) );
  OAI21_X1 U20816 ( .B1(n17719), .B2(n17622), .A(n17948), .ZN(n17627) );
  AOI22_X1 U20817 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17625), .B1(
        n17624), .B2(n17623), .ZN(n17626) );
  AOI211_X1 U20818 ( .C1(n17629), .C2(n17628), .A(n17627), .B(n17626), .ZN(
        n17630) );
  OAI21_X1 U20819 ( .B1(n17950), .B2(n17642), .A(n17630), .ZN(P3_U2821) );
  OAI21_X1 U20820 ( .B1(n17633), .B2(n17632), .A(n17735), .ZN(n17650) );
  OAI211_X1 U20821 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17635), .A(
        n18374), .B(n17634), .ZN(n17636) );
  NAND2_X1 U20822 ( .A1(n18038), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n17951) );
  OAI211_X1 U20823 ( .C1(n17719), .C2(n17637), .A(n17636), .B(n17951), .ZN(
        n17644) );
  AOI21_X1 U20824 ( .B1(n17639), .B2(n17631), .A(n17638), .ZN(n17961) );
  OAI21_X1 U20825 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17641), .A(
        n17640), .ZN(n17959) );
  OAI22_X1 U20826 ( .A1(n17961), .A2(n17642), .B1(n17739), .B2(n17959), .ZN(
        n17643) );
  AOI211_X1 U20827 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17650), .A(
        n17644), .B(n17643), .ZN(n17645) );
  OAI21_X1 U20828 ( .B1(n17646), .B2(n17631), .A(n17645), .ZN(P3_U2822) );
  OAI21_X1 U20829 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17648), .A(
        n17647), .ZN(n17976) );
  INV_X1 U20830 ( .A(n17649), .ZN(n17652) );
  NOR2_X1 U20831 ( .A1(n18048), .A2(n18602), .ZN(n17972) );
  AOI221_X1 U20832 ( .B1(n17652), .B2(n17651), .C1(n17650), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n17972), .ZN(n17659) );
  AOI21_X1 U20833 ( .B1(n17655), .B2(n17654), .A(n17653), .ZN(n17656) );
  XNOR2_X1 U20834 ( .A(n17656), .B(n17970), .ZN(n17973) );
  AOI22_X1 U20835 ( .A1(n17727), .A2(n17973), .B1(n17657), .B2(n17729), .ZN(
        n17658) );
  OAI211_X1 U20836 ( .C1(n17738), .C2(n17976), .A(n17659), .B(n17658), .ZN(
        P3_U2823) );
  OAI21_X1 U20837 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17661), .A(
        n17660), .ZN(n17979) );
  NOR2_X1 U20838 ( .A1(n17662), .A2(n18204), .ZN(n17664) );
  AOI22_X1 U20839 ( .A1(n18038), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n17664), 
        .B2(n17663), .ZN(n17672) );
  NOR2_X1 U20840 ( .A1(n17665), .A2(n17664), .ZN(n17682) );
  OAI21_X1 U20841 ( .B1(n17668), .B2(n17667), .A(n17666), .ZN(n17978) );
  OAI22_X1 U20842 ( .A1(n17719), .A2(n17669), .B1(n17738), .B2(n17978), .ZN(
        n17670) );
  AOI21_X1 U20843 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17682), .A(
        n17670), .ZN(n17671) );
  OAI211_X1 U20844 ( .C1(n17739), .C2(n17979), .A(n17672), .B(n17671), .ZN(
        P3_U2824) );
  OAI21_X1 U20845 ( .B1(n17675), .B2(n17674), .A(n17673), .ZN(n17676) );
  XNOR2_X1 U20846 ( .A(n17676), .B(n17988), .ZN(n17986) );
  OAI21_X1 U20847 ( .B1(n17679), .B2(n17678), .A(n17677), .ZN(n17993) );
  OAI22_X1 U20848 ( .A1(n17739), .A2(n17993), .B1(n18048), .B2(n18598), .ZN(
        n17680) );
  AOI21_X1 U20849 ( .B1(n17681), .B2(n17729), .A(n17680), .ZN(n17685) );
  OAI221_X1 U20850 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17683), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n17735), .A(n17682), .ZN(n17684) );
  OAI211_X1 U20851 ( .C1(n17738), .C2(n17986), .A(n17685), .B(n17684), .ZN(
        P3_U2825) );
  AOI21_X1 U20852 ( .B1(n17687), .B2(n17686), .A(n17722), .ZN(n17708) );
  OAI21_X1 U20853 ( .B1(n17690), .B2(n17689), .A(n17688), .ZN(n17691) );
  XNOR2_X1 U20854 ( .A(n17691), .B(n12529), .ZN(n18005) );
  OAI22_X1 U20855 ( .A1(n17739), .A2(n18005), .B1(n18204), .B2(n17692), .ZN(
        n17698) );
  OAI21_X1 U20856 ( .B1(n17695), .B2(n17694), .A(n17693), .ZN(n17999) );
  OAI22_X1 U20857 ( .A1(n17719), .A2(n17696), .B1(n17738), .B2(n17999), .ZN(
        n17697) );
  AOI211_X1 U20858 ( .C1(n18038), .C2(P3_REIP_REG_4__SCAN_IN), .A(n17698), .B(
        n17697), .ZN(n17699) );
  OAI21_X1 U20859 ( .B1(n17708), .B2(n17700), .A(n17699), .ZN(P3_U2826) );
  OAI21_X1 U20860 ( .B1(n17703), .B2(n17702), .A(n17701), .ZN(n18013) );
  AOI21_X1 U20861 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17735), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17707) );
  OAI21_X1 U20862 ( .B1(n17706), .B2(n17705), .A(n17704), .ZN(n18010) );
  OAI22_X1 U20863 ( .A1(n17708), .A2(n17707), .B1(n17738), .B2(n18010), .ZN(
        n17709) );
  AOI21_X1 U20864 ( .B1(n17710), .B2(n17729), .A(n17709), .ZN(n17711) );
  NAND2_X1 U20865 ( .A1(n18038), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18009) );
  OAI211_X1 U20866 ( .C1(n17739), .C2(n18013), .A(n17711), .B(n18009), .ZN(
        P3_U2827) );
  OAI21_X1 U20867 ( .B1(n17714), .B2(n17713), .A(n17712), .ZN(n18024) );
  INV_X1 U20868 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17721) );
  OAI21_X1 U20869 ( .B1(n17717), .B2(n17716), .A(n17715), .ZN(n18030) );
  OAI22_X1 U20870 ( .A1(n17719), .A2(n17718), .B1(n17738), .B2(n18030), .ZN(
        n17720) );
  AOI221_X1 U20871 ( .B1(n17722), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18374), .C2(n17721), .A(n17720), .ZN(n17723) );
  NAND2_X1 U20872 ( .A1(n18038), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18028) );
  OAI211_X1 U20873 ( .C1(n17739), .C2(n18024), .A(n17723), .B(n18028), .ZN(
        P3_U2828) );
  OAI21_X1 U20874 ( .B1(n17733), .B2(n17725), .A(n17724), .ZN(n18042) );
  NAND2_X1 U20875 ( .A1(n18694), .A2(n17734), .ZN(n17726) );
  XNOR2_X1 U20876 ( .A(n17726), .B(n17725), .ZN(n18037) );
  AOI22_X1 U20877 ( .A1(n17727), .A2(n18037), .B1(n18038), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17732) );
  AOI22_X1 U20878 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17730), .B1(
        n17729), .B2(n17728), .ZN(n17731) );
  OAI211_X1 U20879 ( .C1(n17738), .C2(n18042), .A(n17732), .B(n17731), .ZN(
        P3_U2829) );
  AOI21_X1 U20880 ( .B1(n17734), .B2(n18694), .A(n17733), .ZN(n18046) );
  INV_X1 U20881 ( .A(n18046), .ZN(n18044) );
  NAND3_X1 U20882 ( .A1(n18675), .A2(n18574), .A3(n17735), .ZN(n17736) );
  AOI22_X1 U20883 ( .A1(n18038), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17736), .ZN(n17737) );
  OAI221_X1 U20884 ( .B1(n18046), .B2(n17739), .C1(n18044), .C2(n17738), .A(
        n17737), .ZN(P3_U2830) );
  AOI22_X1 U20885 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18027), .B1(
        n18038), .B2(P3_REIP_REG_27__SCAN_IN), .ZN(n17754) );
  INV_X1 U20886 ( .A(n18532), .ZN(n18505) );
  NAND2_X1 U20887 ( .A1(n18505), .A2(n18529), .ZN(n17996) );
  NOR2_X1 U20888 ( .A1(n17840), .A2(n17805), .ZN(n17741) );
  INV_X1 U20889 ( .A(n17741), .ZN(n17740) );
  AOI221_X1 U20890 ( .B1(n18694), .B2(n17928), .C1(n17740), .C2(n17928), .A(
        n17811), .ZN(n17803) );
  INV_X1 U20891 ( .A(n17996), .ZN(n17953) );
  AOI21_X1 U20892 ( .B1(n17741), .B2(n17803), .A(n17953), .ZN(n17782) );
  AOI21_X1 U20893 ( .B1(n17742), .B2(n17996), .A(n17782), .ZN(n17770) );
  AOI21_X1 U20894 ( .B1(n17744), .B2(n17996), .A(n17743), .ZN(n17748) );
  AOI22_X1 U20895 ( .A1(n18494), .A2(n17746), .B1(n17921), .B2(n17745), .ZN(
        n17747) );
  NAND3_X1 U20896 ( .A1(n17770), .A2(n17748), .A3(n17747), .ZN(n17758) );
  NOR2_X1 U20897 ( .A1(n18049), .A2(n17806), .ZN(n17866) );
  AOI22_X1 U20898 ( .A1(n17749), .A2(n17866), .B1(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18026), .ZN(n17750) );
  INV_X1 U20899 ( .A(n17750), .ZN(n17751) );
  OAI21_X1 U20900 ( .B1(n17752), .B2(n17758), .A(n17751), .ZN(n17753) );
  OAI211_X1 U20901 ( .C1(n17755), .C2(n17960), .A(n17754), .B(n17753), .ZN(
        P3_U2835) );
  AOI22_X1 U20902 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17758), .B1(
        n17757), .B2(n17756), .ZN(n17763) );
  AOI22_X1 U20903 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18027), .B1(
        n17936), .B2(n17759), .ZN(n17762) );
  INV_X1 U20904 ( .A(n17760), .ZN(n17761) );
  OAI211_X1 U20905 ( .C1(n17763), .C2(n18049), .A(n17762), .B(n17761), .ZN(
        P3_U2836) );
  AOI221_X1 U20906 ( .B1(n17841), .B2(n18519), .C1(n17765), .C2(n18519), .A(
        n17764), .ZN(n17769) );
  AOI21_X1 U20907 ( .B1(n17767), .B2(n17766), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17768) );
  AOI211_X1 U20908 ( .C1(n17770), .C2(n17769), .A(n17768), .B(n18049), .ZN(
        n17771) );
  AOI211_X1 U20909 ( .C1(n18027), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17772), .B(n17771), .ZN(n17776) );
  AOI22_X1 U20910 ( .A1(n18045), .A2(n17774), .B1(n17936), .B2(n17773), .ZN(
        n17775) );
  OAI211_X1 U20911 ( .C1(n17967), .C2(n17777), .A(n17776), .B(n17775), .ZN(
        P3_U2837) );
  AOI21_X1 U20912 ( .B1(n17780), .B2(n17779), .A(n17778), .ZN(n17790) );
  INV_X1 U20913 ( .A(n17781), .ZN(n17785) );
  AOI211_X1 U20914 ( .C1(n18494), .C2(n17783), .A(n17782), .B(n18027), .ZN(
        n17784) );
  OAI21_X1 U20915 ( .B1(n17785), .B2(n17904), .A(n17784), .ZN(n17788) );
  NOR2_X1 U20916 ( .A1(n17792), .A2(n17788), .ZN(n17786) );
  AOI21_X1 U20917 ( .B1(n17787), .B2(n17786), .A(n18038), .ZN(n17795) );
  OAI211_X1 U20918 ( .C1(n17956), .C2(n17788), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17795), .ZN(n17789) );
  OAI211_X1 U20919 ( .C1(n17791), .C2(n17960), .A(n17790), .B(n17789), .ZN(
        P3_U2838) );
  OAI21_X1 U20920 ( .B1(n18027), .B2(n17793), .A(n17792), .ZN(n17794) );
  AOI22_X1 U20921 ( .A1(n17936), .A2(n17796), .B1(n17795), .B2(n17794), .ZN(
        n17798) );
  NAND2_X1 U20922 ( .A1(n17798), .A2(n17797), .ZN(P3_U2839) );
  INV_X1 U20923 ( .A(n18027), .ZN(n18032) );
  AOI21_X1 U20924 ( .B1(n17800), .B2(n17936), .A(n17799), .ZN(n17810) );
  OAI22_X1 U20925 ( .A1(n17871), .A2(n17904), .B1(n17870), .B2(n18023), .ZN(
        n17816) );
  AND2_X1 U20926 ( .A1(n17815), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n17804) );
  NAND2_X1 U20927 ( .A1(n18023), .A2(n17904), .ZN(n17927) );
  AOI221_X1 U20928 ( .B1(n17840), .B2(n18532), .C1(n17824), .C2(n18532), .A(
        n17801), .ZN(n17822) );
  OAI21_X1 U20929 ( .B1(n18505), .B2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n17822), .ZN(n17802) );
  AOI21_X1 U20930 ( .B1(n17805), .B2(n17927), .A(n17802), .ZN(n17814) );
  OAI211_X1 U20931 ( .C1(n17939), .C2(n17804), .A(n17803), .B(n17814), .ZN(
        n17808) );
  OAI21_X1 U20932 ( .B1(n17806), .B2(n17805), .A(n17811), .ZN(n17807) );
  OAI211_X1 U20933 ( .C1(n17816), .C2(n17808), .A(n18026), .B(n17807), .ZN(
        n17809) );
  OAI211_X1 U20934 ( .C1(n18032), .C2(n17811), .A(n17810), .B(n17809), .ZN(
        P3_U2840) );
  AOI22_X1 U20935 ( .A1(n17936), .A2(n17813), .B1(n17866), .B2(n17812), .ZN(
        n17821) );
  NOR2_X1 U20936 ( .A1(n18519), .A2(n17928), .ZN(n18031) );
  OAI21_X1 U20937 ( .B1(n17815), .B2(n18031), .A(n17814), .ZN(n17818) );
  NOR2_X1 U20938 ( .A1(n18049), .A2(n17816), .ZN(n17862) );
  OAI21_X1 U20939 ( .B1(n18529), .B2(n17817), .A(n17862), .ZN(n17827) );
  OAI211_X1 U20940 ( .C1(n17818), .C2(n17827), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18048), .ZN(n17819) );
  NAND3_X1 U20941 ( .A1(n17821), .A2(n17820), .A3(n17819), .ZN(P3_U2841) );
  NAND2_X1 U20942 ( .A1(n17839), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17828) );
  INV_X1 U20943 ( .A(n17822), .ZN(n17823) );
  AOI21_X1 U20944 ( .B1(n17824), .B2(n17927), .A(n17823), .ZN(n17825) );
  INV_X1 U20945 ( .A(n17825), .ZN(n17826) );
  OAI21_X1 U20946 ( .B1(n17827), .B2(n17826), .A(n18048), .ZN(n17838) );
  OAI21_X1 U20947 ( .B1(n18031), .B2(n17828), .A(n17838), .ZN(n17830) );
  AOI22_X1 U20948 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17830), .B1(
        n17866), .B2(n17829), .ZN(n17832) );
  OAI211_X1 U20949 ( .C1(n17833), .C2(n17960), .A(n17832), .B(n17831), .ZN(
        P3_U2842) );
  AOI22_X1 U20950 ( .A1(n17936), .A2(n17835), .B1(n17866), .B2(n17834), .ZN(
        n17837) );
  NAND2_X1 U20951 ( .A1(n18038), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17836) );
  OAI211_X1 U20952 ( .C1(n17839), .C2(n17838), .A(n17837), .B(n17836), .ZN(
        P3_U2843) );
  NOR2_X1 U20953 ( .A1(n18529), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17995) );
  NOR3_X1 U20954 ( .A1(n17995), .A2(n17840), .A3(n17865), .ZN(n17844) );
  AOI222_X1 U20955 ( .A1(n18519), .A2(n17842), .B1(n18519), .B2(n17841), .C1(
        n17842), .C2(n17927), .ZN(n17843) );
  OAI211_X1 U20956 ( .C1(n17953), .C2(n17844), .A(n17862), .B(n17843), .ZN(
        n17852) );
  OAI221_X1 U20957 ( .B1(n17852), .B2(n17853), .C1(n17852), .C2(n17996), .A(
        n18048), .ZN(n17849) );
  AOI22_X1 U20958 ( .A1(n17936), .A2(n17846), .B1(n17845), .B2(n17866), .ZN(
        n17848) );
  OAI211_X1 U20959 ( .C1(n17850), .C2(n17849), .A(n17848), .B(n17847), .ZN(
        P3_U2844) );
  AOI22_X1 U20960 ( .A1(n18038), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n17936), 
        .B2(n17851), .ZN(n17856) );
  NAND3_X1 U20961 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18048), .A3(
        n17852), .ZN(n17855) );
  NAND3_X1 U20962 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17866), .A3(
        n17853), .ZN(n17854) );
  NAND3_X1 U20963 ( .A1(n17856), .A2(n17855), .A3(n17854), .ZN(P3_U2845) );
  AOI22_X1 U20964 ( .A1(n18519), .A2(n17858), .B1(n18532), .B2(n17857), .ZN(
        n17924) );
  OAI21_X1 U20965 ( .B1(n17939), .B2(n17859), .A(n17924), .ZN(n17860) );
  AOI211_X1 U20966 ( .C1(n17861), .C2(n17928), .A(n17860), .B(n17885), .ZN(
        n17874) );
  AOI221_X1 U20967 ( .B1(n17863), .B2(n17862), .C1(n17874), .C2(n17862), .A(
        n18038), .ZN(n17867) );
  NOR2_X1 U20968 ( .A1(n18048), .A2(n18620), .ZN(n17864) );
  AOI221_X1 U20969 ( .B1(n17867), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), 
        .C1(n17866), .C2(n17865), .A(n17864), .ZN(n17868) );
  OAI21_X1 U20970 ( .B1(n17869), .B2(n17960), .A(n17868), .ZN(P3_U2846) );
  NOR2_X1 U20971 ( .A1(n17870), .A2(n18014), .ZN(n17882) );
  NOR2_X1 U20972 ( .A1(n17871), .A2(n17904), .ZN(n17877) );
  INV_X1 U20973 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17957) );
  INV_X1 U20974 ( .A(n17872), .ZN(n17981) );
  OAI22_X1 U20975 ( .A1(n17998), .A2(n18017), .B1(n17997), .B2(n18018), .ZN(
        n18007) );
  NAND3_X1 U20976 ( .A1(n17981), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n18007), .ZN(n17969) );
  NOR3_X1 U20977 ( .A1(n17970), .A2(n17957), .A3(n17969), .ZN(n17902) );
  NAND2_X1 U20978 ( .A1(n17887), .A2(n17902), .ZN(n17891) );
  AOI211_X1 U20979 ( .C1(n17885), .C2(n17891), .A(n17874), .B(n17873), .ZN(
        n17875) );
  AOI21_X1 U20980 ( .B1(n17877), .B2(n17876), .A(n17875), .ZN(n17879) );
  OAI22_X1 U20981 ( .A1(n17879), .A2(n18049), .B1(n17960), .B2(n17878), .ZN(
        n17880) );
  AOI21_X1 U20982 ( .B1(n17882), .B2(n17881), .A(n17880), .ZN(n17884) );
  NAND2_X1 U20983 ( .A1(n18038), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17883) );
  OAI211_X1 U20984 ( .C1(n18032), .C2(n17885), .A(n17884), .B(n17883), .ZN(
        P3_U2847) );
  OAI221_X1 U20985 ( .B1(n18529), .B2(n17886), .C1(n18529), .C2(n17925), .A(
        n17924), .ZN(n17907) );
  OAI21_X1 U20986 ( .B1(n17886), .B2(n18017), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17889) );
  OAI22_X1 U20987 ( .A1(n18505), .A2(n17887), .B1(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n18031), .ZN(n17888) );
  NOR3_X1 U20988 ( .A1(n17907), .A2(n17889), .A3(n17888), .ZN(n17890) );
  AOI211_X1 U20989 ( .C1(n17892), .C2(n17891), .A(n17890), .B(n18049), .ZN(
        n17893) );
  AOI211_X1 U20990 ( .C1(n18027), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17894), .B(n17893), .ZN(n17899) );
  AOI22_X1 U20991 ( .A1(n17897), .A2(n17896), .B1(n17936), .B2(n17895), .ZN(
        n17898) );
  OAI211_X1 U20992 ( .C1(n18014), .C2(n17900), .A(n17899), .B(n17898), .ZN(
        P3_U2848) );
  OAI21_X1 U20993 ( .B1(n17902), .B2(n17901), .A(n18026), .ZN(n17943) );
  AOI22_X1 U20994 ( .A1(n18038), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n17936), 
        .B2(n17903), .ZN(n17911) );
  OAI22_X1 U20995 ( .A1(n17939), .A2(n17929), .B1(n17905), .B2(n17904), .ZN(
        n17906) );
  AOI211_X1 U20996 ( .C1(n18494), .C2(n17908), .A(n17907), .B(n17906), .ZN(
        n17914) );
  OAI211_X1 U20997 ( .C1(n17939), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18026), .B(n17914), .ZN(n17909) );
  NAND3_X1 U20998 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18048), .A3(
        n17909), .ZN(n17910) );
  OAI211_X1 U20999 ( .C1(n17912), .C2(n17943), .A(n17911), .B(n17910), .ZN(
        P3_U2849) );
  INV_X1 U21000 ( .A(n17943), .ZN(n17947) );
  AOI22_X1 U21001 ( .A1(n17929), .A2(n17947), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18026), .ZN(n17913) );
  AOI21_X1 U21002 ( .B1(n17914), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17913), .ZN(n17915) );
  AOI21_X1 U21003 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18027), .A(
        n17915), .ZN(n17917) );
  OAI211_X1 U21004 ( .C1(n17918), .C2(n17960), .A(n17917), .B(n17916), .ZN(
        P3_U2850) );
  AOI22_X1 U21005 ( .A1(n18038), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17947), 
        .B2(n17919), .ZN(n17932) );
  AOI22_X1 U21006 ( .A1(n18494), .A2(n17922), .B1(n17921), .B2(n17920), .ZN(
        n17923) );
  OAI211_X1 U21007 ( .C1(n18529), .C2(n17925), .A(n17924), .B(n17923), .ZN(
        n17937) );
  OAI21_X1 U21008 ( .B1(n17928), .B2(n17927), .A(n17926), .ZN(n17938) );
  OAI211_X1 U21009 ( .C1(n17939), .C2(n17929), .A(n17938), .B(n18032), .ZN(
        n17930) );
  OAI211_X1 U21010 ( .C1(n17937), .C2(n17930), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18048), .ZN(n17931) );
  OAI211_X1 U21011 ( .C1(n17933), .C2(n17960), .A(n17932), .B(n17931), .ZN(
        P3_U2851) );
  NAND2_X1 U21012 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17934), .ZN(
        n17944) );
  AOI22_X1 U21013 ( .A1(n18038), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17936), 
        .B2(n17935), .ZN(n17942) );
  NOR2_X1 U21014 ( .A1(n18049), .A2(n17937), .ZN(n17945) );
  OAI211_X1 U21015 ( .C1(n17939), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17945), .B(n17938), .ZN(n17940) );
  NAND3_X1 U21016 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18048), .A3(
        n17940), .ZN(n17941) );
  OAI211_X1 U21017 ( .C1(n17944), .C2(n17943), .A(n17942), .B(n17941), .ZN(
        P3_U2852) );
  OAI21_X1 U21018 ( .B1(n18038), .B2(n17945), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17946) );
  OAI21_X1 U21019 ( .B1(n17947), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17946), .ZN(n17949) );
  OAI211_X1 U21020 ( .C1(n17950), .C2(n17960), .A(n17949), .B(n17948), .ZN(
        P3_U2853) );
  INV_X1 U21021 ( .A(n17951), .ZN(n17965) );
  OAI22_X1 U21022 ( .A1(n17954), .A2(n17953), .B1(n17952), .B2(n18017), .ZN(
        n17955) );
  OR2_X1 U21023 ( .A1(n17995), .A2(n17955), .ZN(n17977) );
  AOI211_X1 U21024 ( .C1(n17956), .C2(n17985), .A(n17970), .B(n17977), .ZN(
        n17968) );
  AOI211_X1 U21025 ( .C1(n17968), .C2(n18032), .A(n17958), .B(n17957), .ZN(
        n17964) );
  NOR4_X1 U21026 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17970), .A3(
        n18049), .A4(n17969), .ZN(n17963) );
  OAI22_X1 U21027 ( .A1(n17961), .A2(n17960), .B1(n18014), .B2(n17959), .ZN(
        n17962) );
  NOR4_X1 U21028 ( .A1(n17965), .A2(n17964), .A3(n17963), .A4(n17962), .ZN(
        n17966) );
  OAI21_X1 U21029 ( .B1(n17631), .B2(n17967), .A(n17966), .ZN(P3_U2854) );
  AOI211_X1 U21030 ( .C1(n17970), .C2(n17969), .A(n17968), .B(n18049), .ZN(
        n17971) );
  AOI211_X1 U21031 ( .C1(n18027), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17972), .B(n17971), .ZN(n17975) );
  NAND2_X1 U21032 ( .A1(n18045), .A2(n17973), .ZN(n17974) );
  OAI211_X1 U21033 ( .C1(n17976), .C2(n18041), .A(n17975), .B(n17974), .ZN(
        P3_U2855) );
  OAI21_X1 U21034 ( .B1(n18049), .B2(n17977), .A(n18048), .ZN(n17987) );
  NAND2_X1 U21035 ( .A1(n18026), .A2(n18007), .ZN(n17994) );
  NOR2_X1 U21036 ( .A1(n17994), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17982) );
  OAI22_X1 U21037 ( .A1(n18014), .A2(n17979), .B1(n18041), .B2(n17978), .ZN(
        n17980) );
  AOI21_X1 U21038 ( .B1(n17982), .B2(n17981), .A(n17980), .ZN(n17984) );
  NAND2_X1 U21039 ( .A1(n18038), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n17983) );
  OAI211_X1 U21040 ( .C1(n17985), .C2(n17987), .A(n17984), .B(n17983), .ZN(
        P3_U2856) );
  NOR4_X1 U21041 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12525), .A3(
        n12529), .A4(n17994), .ZN(n17990) );
  OAI22_X1 U21042 ( .A1(n17988), .A2(n17987), .B1(n18041), .B2(n17986), .ZN(
        n17989) );
  NOR2_X1 U21043 ( .A1(n17990), .A2(n17989), .ZN(n17992) );
  NAND2_X1 U21044 ( .A1(n18038), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n17991) );
  OAI211_X1 U21045 ( .C1(n18014), .C2(n17993), .A(n17992), .B(n17991), .ZN(
        P3_U2857) );
  NOR2_X1 U21046 ( .A1(n12525), .A2(n17994), .ZN(n18002) );
  AOI21_X1 U21047 ( .B1(n17997), .B2(n17996), .A(n17995), .ZN(n18015) );
  NAND2_X1 U21048 ( .A1(n18519), .A2(n17998), .ZN(n18021) );
  NAND3_X1 U21049 ( .A1(n18015), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18021), .ZN(n18006) );
  AOI21_X1 U21050 ( .B1(n18033), .B2(n18006), .A(n18027), .ZN(n18000) );
  OAI22_X1 U21051 ( .A1(n18000), .A2(n12529), .B1(n18041), .B2(n17999), .ZN(
        n18001) );
  AOI21_X1 U21052 ( .B1(n18002), .B2(n12529), .A(n18001), .ZN(n18004) );
  NAND2_X1 U21053 ( .A1(n18038), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n18003) );
  OAI211_X1 U21054 ( .C1(n18014), .C2(n18005), .A(n18004), .B(n18003), .ZN(
        P3_U2858) );
  OAI211_X1 U21055 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18007), .A(
        n18026), .B(n18006), .ZN(n18008) );
  OAI211_X1 U21056 ( .C1(n18010), .C2(n18041), .A(n18009), .B(n18008), .ZN(
        n18011) );
  AOI21_X1 U21057 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18027), .A(
        n18011), .ZN(n18012) );
  OAI21_X1 U21058 ( .B1(n18014), .B2(n18013), .A(n18012), .ZN(P3_U2859) );
  NAND2_X1 U21059 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18016) );
  OAI21_X1 U21060 ( .B1(n18017), .B2(n18016), .A(n18015), .ZN(n18020) );
  NOR2_X1 U21061 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18018), .ZN(
        n18019) );
  AOI22_X1 U21062 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18020), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18019), .ZN(n18022) );
  OAI211_X1 U21063 ( .C1(n18024), .C2(n18023), .A(n18022), .B(n18021), .ZN(
        n18025) );
  AOI22_X1 U21064 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18027), .B1(
        n18026), .B2(n18025), .ZN(n18029) );
  OAI211_X1 U21065 ( .C1(n18030), .C2(n18041), .A(n18029), .B(n18028), .ZN(
        P3_U2860) );
  OR3_X1 U21066 ( .A1(n18049), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n18031), .ZN(n18051) );
  INV_X1 U21067 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18677) );
  AOI21_X1 U21068 ( .B1(n18032), .B2(n18051), .A(n18677), .ZN(n18036) );
  OAI211_X1 U21069 ( .C1(n18532), .C2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18677), .B(n18033), .ZN(n18034) );
  INV_X1 U21070 ( .A(n18034), .ZN(n18035) );
  AOI211_X1 U21071 ( .C1(n18045), .C2(n18037), .A(n18036), .B(n18035), .ZN(
        n18040) );
  NAND2_X1 U21072 ( .A1(n18038), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18039) );
  OAI211_X1 U21073 ( .C1(n18042), .C2(n18041), .A(n18040), .B(n18039), .ZN(
        P3_U2861) );
  INV_X1 U21074 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18704) );
  NOR2_X1 U21075 ( .A1(n18048), .A2(n18704), .ZN(n18043) );
  AOI221_X1 U21076 ( .B1(n18047), .B2(n18046), .C1(n18045), .C2(n18044), .A(
        n18043), .ZN(n18052) );
  OAI211_X1 U21077 ( .C1(n18532), .C2(n18049), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18048), .ZN(n18050) );
  NAND3_X1 U21078 ( .A1(n18052), .A2(n18051), .A3(n18050), .ZN(P3_U2862) );
  AOI211_X1 U21079 ( .C1(n18054), .C2(n18053), .A(n18563), .B(n18675), .ZN(
        n18556) );
  OAI21_X1 U21080 ( .B1(n18556), .B2(n18098), .A(n18059), .ZN(n18055) );
  OAI221_X1 U21081 ( .B1(n18533), .B2(n18710), .C1(n18533), .C2(n18059), .A(
        n18055), .ZN(P3_U2863) );
  INV_X1 U21082 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18544) );
  NOR2_X1 U21083 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20885), .ZN(
        n18228) );
  NAND2_X1 U21084 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20885), .ZN(
        n18321) );
  NOR2_X1 U21085 ( .A1(n18297), .A2(n18321), .ZN(n18349) );
  NOR2_X1 U21086 ( .A1(n18228), .A2(n18349), .ZN(n18057) );
  OAI22_X1 U21087 ( .A1(n18058), .A2(n18544), .B1(n18057), .B2(n18056), .ZN(
        P3_U2866) );
  NOR2_X1 U21088 ( .A1(n18545), .A2(n18059), .ZN(P3_U2867) );
  NAND2_X1 U21089 ( .A1(n18061), .A2(n18060), .ZN(n18093) );
  NOR2_X1 U21090 ( .A1(n18062), .A2(n18093), .ZN(n18403) );
  NOR2_X1 U21091 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18537) );
  NOR2_X1 U21092 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18139) );
  NAND2_X1 U21093 ( .A1(n18537), .A2(n18139), .ZN(n18159) );
  NOR2_X1 U21094 ( .A1(n20885), .A2(n18544), .ZN(n18065) );
  NOR2_X1 U21095 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18534), .ZN(
        n18296) );
  NAND2_X1 U21096 ( .A1(n18065), .A2(n18296), .ZN(n18401) );
  INV_X1 U21097 ( .A(n18401), .ZN(n18428) );
  AND2_X1 U21098 ( .A1(n18374), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18435) );
  AND2_X1 U21099 ( .A1(n18300), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18434) );
  NOR2_X1 U21100 ( .A1(n18544), .A2(n18227), .ZN(n18437) );
  NAND2_X1 U21101 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18437), .ZN(
        n18448) );
  AOI21_X1 U21102 ( .B1(n18448), .B2(n18159), .A(n18564), .ZN(n18092) );
  AOI22_X1 U21103 ( .A1(n18428), .A2(n18435), .B1(n18434), .B2(n18092), .ZN(
        n18067) );
  NOR2_X1 U21104 ( .A1(n18533), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18272) );
  OR2_X1 U21105 ( .A1(n18296), .A2(n18272), .ZN(n18348) );
  NAND2_X1 U21106 ( .A1(n18065), .A2(n18348), .ZN(n18402) );
  INV_X1 U21107 ( .A(n18402), .ZN(n18064) );
  AOI21_X1 U21108 ( .B1(n18448), .B2(n18159), .A(n18399), .ZN(n18117) );
  AOI22_X1 U21109 ( .A1(n18374), .A2(n18064), .B1(n18117), .B2(n18063), .ZN(
        n18095) );
  NAND2_X1 U21110 ( .A1(n18065), .A2(n18534), .ZN(n18372) );
  NOR2_X1 U21111 ( .A1(n18533), .A2(n18372), .ZN(n18472) );
  NOR2_X2 U21112 ( .A1(n19104), .A2(n18204), .ZN(n18439) );
  AOI22_X1 U21113 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18095), .B1(
        n18472), .B2(n18439), .ZN(n18066) );
  OAI211_X1 U21114 ( .C1(n18442), .C2(n18159), .A(n18067), .B(n18066), .ZN(
        P3_U2868) );
  NOR2_X1 U21115 ( .A1(n18716), .A2(n18093), .ZN(n18408) );
  INV_X1 U21116 ( .A(n18408), .ZN(n18449) );
  NAND2_X1 U21117 ( .A1(n18374), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18411) );
  INV_X1 U21118 ( .A(n18411), .ZN(n18444) );
  NOR2_X2 U21119 ( .A1(n18399), .A2(n18068), .ZN(n18443) );
  AOI22_X1 U21120 ( .A1(n18428), .A2(n18444), .B1(n18443), .B2(n18092), .ZN(
        n18070) );
  NOR2_X2 U21121 ( .A1(n19117), .A2(n18204), .ZN(n18445) );
  AOI22_X1 U21122 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18095), .B1(
        n18472), .B2(n18445), .ZN(n18069) );
  OAI211_X1 U21123 ( .C1(n18449), .C2(n18159), .A(n18070), .B(n18069), .ZN(
        P3_U2869) );
  NAND2_X1 U21124 ( .A1(n18374), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18455) );
  CLKBUF_X1 U21125 ( .A(n18472), .Z(n18486) );
  NOR2_X1 U21126 ( .A1(n14960), .A2(n18204), .ZN(n18451) );
  NOR2_X2 U21127 ( .A1(n18399), .A2(n18071), .ZN(n18450) );
  AOI22_X1 U21128 ( .A1(n18486), .A2(n18451), .B1(n18450), .B2(n18092), .ZN(
        n18074) );
  NOR2_X2 U21129 ( .A1(n18072), .A2(n18093), .ZN(n18452) );
  AOI22_X1 U21130 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18095), .B1(
        n18452), .B2(n18150), .ZN(n18073) );
  OAI211_X1 U21131 ( .C1(n18401), .C2(n18455), .A(n18074), .B(n18073), .ZN(
        P3_U2870) );
  NAND2_X1 U21132 ( .A1(n18374), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18461) );
  NAND2_X1 U21133 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18374), .ZN(n18332) );
  INV_X1 U21134 ( .A(n18332), .ZN(n18457) );
  NOR2_X2 U21135 ( .A1(n18399), .A2(n18075), .ZN(n18456) );
  AOI22_X1 U21136 ( .A1(n18486), .A2(n18457), .B1(n18456), .B2(n18092), .ZN(
        n18078) );
  NOR2_X2 U21137 ( .A1(n18076), .A2(n18093), .ZN(n18458) );
  AOI22_X1 U21138 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18095), .B1(
        n18458), .B2(n18150), .ZN(n18077) );
  OAI211_X1 U21139 ( .C1(n18401), .C2(n18461), .A(n18078), .B(n18077), .ZN(
        P3_U2871) );
  NAND2_X1 U21140 ( .A1(n18374), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18468) );
  NOR2_X1 U21141 ( .A1(n18079), .A2(n18204), .ZN(n18463) );
  NOR2_X2 U21142 ( .A1(n18399), .A2(n18080), .ZN(n18462) );
  AOI22_X1 U21143 ( .A1(n18472), .A2(n18463), .B1(n18462), .B2(n18092), .ZN(
        n18083) );
  NOR2_X2 U21144 ( .A1(n18081), .A2(n18093), .ZN(n18465) );
  AOI22_X1 U21145 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18095), .B1(
        n18465), .B2(n18150), .ZN(n18082) );
  OAI211_X1 U21146 ( .C1(n18401), .C2(n18468), .A(n18083), .B(n18082), .ZN(
        P3_U2872) );
  NAND2_X1 U21147 ( .A1(n18374), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18421) );
  NAND2_X1 U21148 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18374), .ZN(n18476) );
  INV_X1 U21149 ( .A(n18476), .ZN(n18418) );
  NOR2_X2 U21150 ( .A1(n18399), .A2(n18084), .ZN(n18470) );
  AOI22_X1 U21151 ( .A1(n18472), .A2(n18418), .B1(n18470), .B2(n18092), .ZN(
        n18087) );
  NOR2_X2 U21152 ( .A1(n18085), .A2(n18093), .ZN(n18473) );
  AOI22_X1 U21153 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18095), .B1(
        n18473), .B2(n18150), .ZN(n18086) );
  OAI211_X1 U21154 ( .C1(n18401), .C2(n18421), .A(n18087), .B(n18086), .ZN(
        P3_U2873) );
  INV_X1 U21155 ( .A(n18472), .ZN(n18469) );
  NAND2_X1 U21156 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18374), .ZN(n18482) );
  NOR2_X1 U21157 ( .A1(n18204), .A2(n20830), .ZN(n18478) );
  NOR2_X2 U21158 ( .A1(n18399), .A2(n18088), .ZN(n18477) );
  AOI22_X1 U21159 ( .A1(n18428), .A2(n18478), .B1(n18477), .B2(n18092), .ZN(
        n18091) );
  NOR2_X2 U21160 ( .A1(n18089), .A2(n18093), .ZN(n18479) );
  AOI22_X1 U21161 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18095), .B1(
        n18479), .B2(n18150), .ZN(n18090) );
  OAI211_X1 U21162 ( .C1(n18469), .C2(n18482), .A(n18091), .B(n18090), .ZN(
        P3_U2874) );
  NAND2_X1 U21163 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18374), .ZN(n18432) );
  NAND2_X1 U21164 ( .A1(n18374), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18492) );
  INV_X1 U21165 ( .A(n18492), .ZN(n18426) );
  AND2_X1 U21166 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18300), .ZN(n18484) );
  AOI22_X1 U21167 ( .A1(n18486), .A2(n18426), .B1(n18484), .B2(n18092), .ZN(
        n18097) );
  NOR2_X2 U21168 ( .A1(n18094), .A2(n18093), .ZN(n18488) );
  AOI22_X1 U21169 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18095), .B1(
        n18488), .B2(n18150), .ZN(n18096) );
  OAI211_X1 U21170 ( .C1(n18401), .C2(n18432), .A(n18097), .B(n18096), .ZN(
        P3_U2875) );
  NAND2_X1 U21171 ( .A1(n18272), .A2(n18139), .ZN(n18181) );
  INV_X1 U21172 ( .A(n18139), .ZN(n18138) );
  NAND2_X1 U21173 ( .A1(n18534), .A2(n18433), .ZN(n18273) );
  NOR2_X1 U21174 ( .A1(n18138), .A2(n18273), .ZN(n18113) );
  AOI22_X1 U21175 ( .A1(n18428), .A2(n18439), .B1(n18434), .B2(n18113), .ZN(
        n18100) );
  NOR2_X1 U21176 ( .A1(n18399), .A2(n18098), .ZN(n18436) );
  AND2_X1 U21177 ( .A1(n18534), .A2(n18436), .ZN(n18274) );
  AOI22_X1 U21178 ( .A1(n18374), .A2(n18437), .B1(n18139), .B2(n18274), .ZN(
        n18114) );
  INV_X1 U21179 ( .A(n18448), .ZN(n18487) );
  AOI22_X1 U21180 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18114), .B1(
        n18435), .B2(n18487), .ZN(n18099) );
  OAI211_X1 U21181 ( .C1(n18442), .C2(n18181), .A(n18100), .B(n18099), .ZN(
        P3_U2876) );
  AOI22_X1 U21182 ( .A1(n18428), .A2(n18445), .B1(n18443), .B2(n18113), .ZN(
        n18102) );
  AOI22_X1 U21183 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18114), .B1(
        n18444), .B2(n18487), .ZN(n18101) );
  OAI211_X1 U21184 ( .C1(n18449), .C2(n18181), .A(n18102), .B(n18101), .ZN(
        P3_U2877) );
  AOI22_X1 U21185 ( .A1(n18428), .A2(n18451), .B1(n18450), .B2(n18113), .ZN(
        n18104) );
  AOI22_X1 U21186 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18114), .B1(
        n18452), .B2(n18174), .ZN(n18103) );
  OAI211_X1 U21187 ( .C1(n18455), .C2(n18448), .A(n18104), .B(n18103), .ZN(
        P3_U2878) );
  AOI22_X1 U21188 ( .A1(n18428), .A2(n18457), .B1(n18456), .B2(n18113), .ZN(
        n18106) );
  AOI22_X1 U21189 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18114), .B1(
        n18458), .B2(n18174), .ZN(n18105) );
  OAI211_X1 U21190 ( .C1(n18461), .C2(n18448), .A(n18106), .B(n18105), .ZN(
        P3_U2879) );
  INV_X1 U21191 ( .A(n18463), .ZN(n18336) );
  INV_X1 U21192 ( .A(n18468), .ZN(n18333) );
  AOI22_X1 U21193 ( .A1(n18333), .A2(n18487), .B1(n18462), .B2(n18113), .ZN(
        n18108) );
  AOI22_X1 U21194 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18114), .B1(
        n18465), .B2(n18174), .ZN(n18107) );
  OAI211_X1 U21195 ( .C1(n18401), .C2(n18336), .A(n18108), .B(n18107), .ZN(
        P3_U2880) );
  INV_X1 U21196 ( .A(n18421), .ZN(n18471) );
  AOI22_X1 U21197 ( .A1(n18471), .A2(n18487), .B1(n18470), .B2(n18113), .ZN(
        n18110) );
  AOI22_X1 U21198 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18114), .B1(
        n18473), .B2(n18174), .ZN(n18109) );
  OAI211_X1 U21199 ( .C1(n18401), .C2(n18476), .A(n18110), .B(n18109), .ZN(
        P3_U2881) );
  INV_X1 U21200 ( .A(n18478), .ZN(n18366) );
  INV_X1 U21201 ( .A(n18482), .ZN(n18363) );
  AOI22_X1 U21202 ( .A1(n18428), .A2(n18363), .B1(n18477), .B2(n18113), .ZN(
        n18112) );
  AOI22_X1 U21203 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18114), .B1(
        n18479), .B2(n18174), .ZN(n18111) );
  OAI211_X1 U21204 ( .C1(n18366), .C2(n18448), .A(n18112), .B(n18111), .ZN(
        P3_U2882) );
  INV_X1 U21205 ( .A(n18432), .ZN(n18485) );
  AOI22_X1 U21206 ( .A1(n18485), .A2(n18487), .B1(n18484), .B2(n18113), .ZN(
        n18116) );
  AOI22_X1 U21207 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18114), .B1(
        n18488), .B2(n18174), .ZN(n18115) );
  OAI211_X1 U21208 ( .C1(n18401), .C2(n18492), .A(n18116), .B(n18115), .ZN(
        P3_U2883) );
  NAND2_X1 U21209 ( .A1(n18296), .A2(n18139), .ZN(n18203) );
  INV_X1 U21210 ( .A(n18203), .ZN(n18194) );
  NOR2_X1 U21211 ( .A1(n18174), .A2(n18194), .ZN(n18160) );
  NOR2_X1 U21212 ( .A1(n18564), .A2(n18160), .ZN(n18134) );
  AOI22_X1 U21213 ( .A1(n18434), .A2(n18134), .B1(n18435), .B2(n18150), .ZN(
        n18121) );
  INV_X1 U21214 ( .A(n18117), .ZN(n18118) );
  OAI22_X1 U21215 ( .A1(n18160), .A2(n18399), .B1(n18297), .B2(n18118), .ZN(
        n18119) );
  OAI21_X1 U21216 ( .B1(n18194), .B2(n18667), .A(n18119), .ZN(n18135) );
  AOI22_X1 U21217 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18135), .B1(
        n18439), .B2(n18487), .ZN(n18120) );
  OAI211_X1 U21218 ( .C1(n18442), .C2(n18203), .A(n18121), .B(n18120), .ZN(
        P3_U2884) );
  AOI22_X1 U21219 ( .A1(n18443), .A2(n18134), .B1(n18445), .B2(n18487), .ZN(
        n18123) );
  AOI22_X1 U21220 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18135), .B1(
        n18408), .B2(n18194), .ZN(n18122) );
  OAI211_X1 U21221 ( .C1(n18411), .C2(n18159), .A(n18123), .B(n18122), .ZN(
        P3_U2885) );
  INV_X1 U21222 ( .A(n18451), .ZN(n18382) );
  INV_X1 U21223 ( .A(n18455), .ZN(n18379) );
  AOI22_X1 U21224 ( .A1(n18379), .A2(n18150), .B1(n18450), .B2(n18134), .ZN(
        n18125) );
  AOI22_X1 U21225 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18135), .B1(
        n18452), .B2(n18194), .ZN(n18124) );
  OAI211_X1 U21226 ( .C1(n18382), .C2(n18448), .A(n18125), .B(n18124), .ZN(
        P3_U2886) );
  INV_X1 U21227 ( .A(n18461), .ZN(n18329) );
  AOI22_X1 U21228 ( .A1(n18329), .A2(n18150), .B1(n18456), .B2(n18134), .ZN(
        n18127) );
  AOI22_X1 U21229 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18135), .B1(
        n18458), .B2(n18194), .ZN(n18126) );
  OAI211_X1 U21230 ( .C1(n18332), .C2(n18448), .A(n18127), .B(n18126), .ZN(
        P3_U2887) );
  AOI22_X1 U21231 ( .A1(n18333), .A2(n18150), .B1(n18462), .B2(n18134), .ZN(
        n18129) );
  AOI22_X1 U21232 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18135), .B1(
        n18465), .B2(n18194), .ZN(n18128) );
  OAI211_X1 U21233 ( .C1(n18336), .C2(n18448), .A(n18129), .B(n18128), .ZN(
        P3_U2888) );
  AOI22_X1 U21234 ( .A1(n18471), .A2(n18150), .B1(n18470), .B2(n18134), .ZN(
        n18131) );
  AOI22_X1 U21235 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18135), .B1(
        n18473), .B2(n18194), .ZN(n18130) );
  OAI211_X1 U21236 ( .C1(n18476), .C2(n18448), .A(n18131), .B(n18130), .ZN(
        P3_U2889) );
  AOI22_X1 U21237 ( .A1(n18477), .A2(n18134), .B1(n18478), .B2(n18150), .ZN(
        n18133) );
  AOI22_X1 U21238 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18135), .B1(
        n18479), .B2(n18194), .ZN(n18132) );
  OAI211_X1 U21239 ( .C1(n18482), .C2(n18448), .A(n18133), .B(n18132), .ZN(
        P3_U2890) );
  AOI22_X1 U21240 ( .A1(n18485), .A2(n18150), .B1(n18484), .B2(n18134), .ZN(
        n18137) );
  AOI22_X1 U21241 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18135), .B1(
        n18488), .B2(n18194), .ZN(n18136) );
  OAI211_X1 U21242 ( .C1(n18492), .C2(n18448), .A(n18137), .B(n18136), .ZN(
        P3_U2891) );
  NOR2_X1 U21243 ( .A1(n18534), .A2(n18138), .ZN(n18183) );
  NAND2_X1 U21244 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18183), .ZN(
        n18215) );
  AOI21_X1 U21245 ( .B1(n18534), .B2(n18297), .A(n18399), .ZN(n18229) );
  OAI211_X1 U21246 ( .C1(n18223), .C2(n18667), .A(n18139), .B(n18229), .ZN(
        n18156) );
  AND2_X1 U21247 ( .A1(n18433), .A2(n18183), .ZN(n18155) );
  AOI22_X1 U21248 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18156), .B1(
        n18434), .B2(n18155), .ZN(n18141) );
  AOI22_X1 U21249 ( .A1(n18439), .A2(n18150), .B1(n18435), .B2(n18174), .ZN(
        n18140) );
  OAI211_X1 U21250 ( .C1(n18442), .C2(n18215), .A(n18141), .B(n18140), .ZN(
        P3_U2892) );
  AOI22_X1 U21251 ( .A1(n18443), .A2(n18155), .B1(n18445), .B2(n18150), .ZN(
        n18143) );
  AOI22_X1 U21252 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18156), .B1(
        n18408), .B2(n18223), .ZN(n18142) );
  OAI211_X1 U21253 ( .C1(n18411), .C2(n18181), .A(n18143), .B(n18142), .ZN(
        P3_U2893) );
  AOI22_X1 U21254 ( .A1(n18451), .A2(n18150), .B1(n18450), .B2(n18155), .ZN(
        n18145) );
  AOI22_X1 U21255 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18156), .B1(
        n18452), .B2(n18223), .ZN(n18144) );
  OAI211_X1 U21256 ( .C1(n18455), .C2(n18181), .A(n18145), .B(n18144), .ZN(
        P3_U2894) );
  AOI22_X1 U21257 ( .A1(n18329), .A2(n18174), .B1(n18456), .B2(n18155), .ZN(
        n18147) );
  AOI22_X1 U21258 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18156), .B1(
        n18458), .B2(n18223), .ZN(n18146) );
  OAI211_X1 U21259 ( .C1(n18332), .C2(n18159), .A(n18147), .B(n18146), .ZN(
        P3_U2895) );
  AOI22_X1 U21260 ( .A1(n18463), .A2(n18150), .B1(n18462), .B2(n18155), .ZN(
        n18149) );
  AOI22_X1 U21261 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18156), .B1(
        n18465), .B2(n18223), .ZN(n18148) );
  OAI211_X1 U21262 ( .C1(n18468), .C2(n18181), .A(n18149), .B(n18148), .ZN(
        P3_U2896) );
  AOI22_X1 U21263 ( .A1(n18418), .A2(n18150), .B1(n18470), .B2(n18155), .ZN(
        n18152) );
  AOI22_X1 U21264 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18156), .B1(
        n18473), .B2(n18223), .ZN(n18151) );
  OAI211_X1 U21265 ( .C1(n18421), .C2(n18181), .A(n18152), .B(n18151), .ZN(
        P3_U2897) );
  AOI22_X1 U21266 ( .A1(n18477), .A2(n18155), .B1(n18478), .B2(n18174), .ZN(
        n18154) );
  AOI22_X1 U21267 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18156), .B1(
        n18479), .B2(n18223), .ZN(n18153) );
  OAI211_X1 U21268 ( .C1(n18482), .C2(n18159), .A(n18154), .B(n18153), .ZN(
        P3_U2898) );
  AOI22_X1 U21269 ( .A1(n18485), .A2(n18174), .B1(n18484), .B2(n18155), .ZN(
        n18158) );
  AOI22_X1 U21270 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18156), .B1(
        n18488), .B2(n18223), .ZN(n18157) );
  OAI211_X1 U21271 ( .C1(n18492), .C2(n18159), .A(n18158), .B(n18157), .ZN(
        P3_U2899) );
  NAND2_X1 U21272 ( .A1(n18537), .A2(n18228), .ZN(n18249) );
  AOI21_X1 U21273 ( .B1(n18215), .B2(n18249), .A(n18564), .ZN(n18177) );
  AOI22_X1 U21274 ( .A1(n18434), .A2(n18177), .B1(n18435), .B2(n18194), .ZN(
        n18163) );
  INV_X1 U21275 ( .A(n18249), .ZN(n18242) );
  AOI221_X1 U21276 ( .B1(n18160), .B2(n18215), .C1(n18297), .C2(n18215), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18161) );
  OAI21_X1 U21277 ( .B1(n18242), .B2(n18161), .A(n18300), .ZN(n18178) );
  AOI22_X1 U21278 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18178), .B1(
        n18439), .B2(n18174), .ZN(n18162) );
  OAI211_X1 U21279 ( .C1(n18442), .C2(n18249), .A(n18163), .B(n18162), .ZN(
        P3_U2900) );
  AOI22_X1 U21280 ( .A1(n18444), .A2(n18194), .B1(n18443), .B2(n18177), .ZN(
        n18165) );
  AOI22_X1 U21281 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18178), .B1(
        n18445), .B2(n18174), .ZN(n18164) );
  OAI211_X1 U21282 ( .C1(n18449), .C2(n18249), .A(n18165), .B(n18164), .ZN(
        P3_U2901) );
  AOI22_X1 U21283 ( .A1(n18451), .A2(n18174), .B1(n18450), .B2(n18177), .ZN(
        n18167) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18178), .B1(
        n18452), .B2(n18242), .ZN(n18166) );
  OAI211_X1 U21285 ( .C1(n18455), .C2(n18203), .A(n18167), .B(n18166), .ZN(
        P3_U2902) );
  AOI22_X1 U21286 ( .A1(n18457), .A2(n18174), .B1(n18456), .B2(n18177), .ZN(
        n18169) );
  AOI22_X1 U21287 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18178), .B1(
        n18458), .B2(n18242), .ZN(n18168) );
  OAI211_X1 U21288 ( .C1(n18461), .C2(n18203), .A(n18169), .B(n18168), .ZN(
        P3_U2903) );
  AOI22_X1 U21289 ( .A1(n18333), .A2(n18194), .B1(n18462), .B2(n18177), .ZN(
        n18171) );
  AOI22_X1 U21290 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18178), .B1(
        n18465), .B2(n18242), .ZN(n18170) );
  OAI211_X1 U21291 ( .C1(n18336), .C2(n18181), .A(n18171), .B(n18170), .ZN(
        P3_U2904) );
  AOI22_X1 U21292 ( .A1(n18418), .A2(n18174), .B1(n18470), .B2(n18177), .ZN(
        n18173) );
  AOI22_X1 U21293 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18178), .B1(
        n18473), .B2(n18242), .ZN(n18172) );
  OAI211_X1 U21294 ( .C1(n18421), .C2(n18203), .A(n18173), .B(n18172), .ZN(
        P3_U2905) );
  AOI22_X1 U21295 ( .A1(n18363), .A2(n18174), .B1(n18477), .B2(n18177), .ZN(
        n18176) );
  AOI22_X1 U21296 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18178), .B1(
        n18479), .B2(n18242), .ZN(n18175) );
  OAI211_X1 U21297 ( .C1(n18366), .C2(n18203), .A(n18176), .B(n18175), .ZN(
        P3_U2906) );
  AOI22_X1 U21298 ( .A1(n18485), .A2(n18194), .B1(n18484), .B2(n18177), .ZN(
        n18180) );
  AOI22_X1 U21299 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18178), .B1(
        n18488), .B2(n18242), .ZN(n18179) );
  OAI211_X1 U21300 ( .C1(n18492), .C2(n18181), .A(n18180), .B(n18179), .ZN(
        P3_U2907) );
  NAND2_X1 U21301 ( .A1(n18272), .A2(n18228), .ZN(n18266) );
  INV_X1 U21302 ( .A(n18228), .ZN(n18182) );
  NOR2_X1 U21303 ( .A1(n18273), .A2(n18182), .ZN(n18199) );
  AOI22_X1 U21304 ( .A1(n18439), .A2(n18194), .B1(n18434), .B2(n18199), .ZN(
        n18185) );
  AOI22_X1 U21305 ( .A1(n18374), .A2(n18183), .B1(n18274), .B2(n18228), .ZN(
        n18200) );
  AOI22_X1 U21306 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18200), .B1(
        n18435), .B2(n18223), .ZN(n18184) );
  OAI211_X1 U21307 ( .C1(n18442), .C2(n18266), .A(n18185), .B(n18184), .ZN(
        P3_U2908) );
  AOI22_X1 U21308 ( .A1(n18444), .A2(n18223), .B1(n18443), .B2(n18199), .ZN(
        n18187) );
  AOI22_X1 U21309 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18200), .B1(
        n18445), .B2(n18194), .ZN(n18186) );
  OAI211_X1 U21310 ( .C1(n18449), .C2(n18266), .A(n18187), .B(n18186), .ZN(
        P3_U2909) );
  AOI22_X1 U21311 ( .A1(n18451), .A2(n18194), .B1(n18450), .B2(n18199), .ZN(
        n18189) );
  AOI22_X1 U21312 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18200), .B1(
        n18452), .B2(n18268), .ZN(n18188) );
  OAI211_X1 U21313 ( .C1(n18455), .C2(n18215), .A(n18189), .B(n18188), .ZN(
        P3_U2910) );
  AOI22_X1 U21314 ( .A1(n18329), .A2(n18223), .B1(n18456), .B2(n18199), .ZN(
        n18191) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18200), .B1(
        n18458), .B2(n18268), .ZN(n18190) );
  OAI211_X1 U21316 ( .C1(n18332), .C2(n18203), .A(n18191), .B(n18190), .ZN(
        P3_U2911) );
  AOI22_X1 U21317 ( .A1(n18333), .A2(n18223), .B1(n18462), .B2(n18199), .ZN(
        n18193) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18200), .B1(
        n18465), .B2(n18268), .ZN(n18192) );
  OAI211_X1 U21319 ( .C1(n18336), .C2(n18203), .A(n18193), .B(n18192), .ZN(
        P3_U2912) );
  AOI22_X1 U21320 ( .A1(n18418), .A2(n18194), .B1(n18470), .B2(n18199), .ZN(
        n18196) );
  AOI22_X1 U21321 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18200), .B1(
        n18473), .B2(n18268), .ZN(n18195) );
  OAI211_X1 U21322 ( .C1(n18421), .C2(n18215), .A(n18196), .B(n18195), .ZN(
        P3_U2913) );
  AOI22_X1 U21323 ( .A1(n18477), .A2(n18199), .B1(n18478), .B2(n18223), .ZN(
        n18198) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18200), .B1(
        n18479), .B2(n18268), .ZN(n18197) );
  OAI211_X1 U21325 ( .C1(n18482), .C2(n18203), .A(n18198), .B(n18197), .ZN(
        P3_U2914) );
  AOI22_X1 U21326 ( .A1(n18485), .A2(n18223), .B1(n18484), .B2(n18199), .ZN(
        n18202) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18200), .B1(
        n18488), .B2(n18268), .ZN(n18201) );
  OAI211_X1 U21328 ( .C1(n18492), .C2(n18203), .A(n18202), .B(n18201), .ZN(
        P3_U2915) );
  NAND2_X1 U21329 ( .A1(n18296), .A2(n18228), .ZN(n18295) );
  NOR2_X1 U21330 ( .A1(n18268), .A2(n18288), .ZN(n18250) );
  NOR2_X1 U21331 ( .A1(n18564), .A2(n18250), .ZN(n18222) );
  AOI22_X1 U21332 ( .A1(n18439), .A2(n18223), .B1(n18434), .B2(n18222), .ZN(
        n18208) );
  NOR2_X1 U21333 ( .A1(n18223), .A2(n18242), .ZN(n18205) );
  OAI22_X1 U21334 ( .A1(n18205), .A2(n18204), .B1(n18250), .B2(n18399), .ZN(
        n18206) );
  OAI21_X1 U21335 ( .B1(n18288), .B2(n18667), .A(n18206), .ZN(n18224) );
  AOI22_X1 U21336 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18224), .B1(
        n18435), .B2(n18242), .ZN(n18207) );
  OAI211_X1 U21337 ( .C1(n18442), .C2(n18295), .A(n18208), .B(n18207), .ZN(
        P3_U2916) );
  AOI22_X1 U21338 ( .A1(n18443), .A2(n18222), .B1(n18445), .B2(n18223), .ZN(
        n18210) );
  AOI22_X1 U21339 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18224), .B1(
        n18408), .B2(n18288), .ZN(n18209) );
  OAI211_X1 U21340 ( .C1(n18411), .C2(n18249), .A(n18210), .B(n18209), .ZN(
        P3_U2917) );
  AOI22_X1 U21341 ( .A1(n18451), .A2(n18223), .B1(n18450), .B2(n18222), .ZN(
        n18212) );
  AOI22_X1 U21342 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18224), .B1(
        n18452), .B2(n18288), .ZN(n18211) );
  OAI211_X1 U21343 ( .C1(n18455), .C2(n18249), .A(n18212), .B(n18211), .ZN(
        P3_U2918) );
  AOI22_X1 U21344 ( .A1(n18329), .A2(n18242), .B1(n18456), .B2(n18222), .ZN(
        n18214) );
  AOI22_X1 U21345 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18224), .B1(
        n18458), .B2(n18288), .ZN(n18213) );
  OAI211_X1 U21346 ( .C1(n18332), .C2(n18215), .A(n18214), .B(n18213), .ZN(
        P3_U2919) );
  AOI22_X1 U21347 ( .A1(n18463), .A2(n18223), .B1(n18462), .B2(n18222), .ZN(
        n18217) );
  AOI22_X1 U21348 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18224), .B1(
        n18465), .B2(n18288), .ZN(n18216) );
  OAI211_X1 U21349 ( .C1(n18468), .C2(n18249), .A(n18217), .B(n18216), .ZN(
        P3_U2920) );
  AOI22_X1 U21350 ( .A1(n18418), .A2(n18223), .B1(n18470), .B2(n18222), .ZN(
        n18219) );
  AOI22_X1 U21351 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18224), .B1(
        n18473), .B2(n18288), .ZN(n18218) );
  OAI211_X1 U21352 ( .C1(n18421), .C2(n18249), .A(n18219), .B(n18218), .ZN(
        P3_U2921) );
  AOI22_X1 U21353 ( .A1(n18363), .A2(n18223), .B1(n18477), .B2(n18222), .ZN(
        n18221) );
  AOI22_X1 U21354 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18224), .B1(
        n18479), .B2(n18288), .ZN(n18220) );
  OAI211_X1 U21355 ( .C1(n18366), .C2(n18249), .A(n18221), .B(n18220), .ZN(
        P3_U2922) );
  AOI22_X1 U21356 ( .A1(n18426), .A2(n18223), .B1(n18484), .B2(n18222), .ZN(
        n18226) );
  AOI22_X1 U21357 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18224), .B1(
        n18488), .B2(n18288), .ZN(n18225) );
  OAI211_X1 U21358 ( .C1(n18432), .C2(n18249), .A(n18226), .B(n18225), .ZN(
        P3_U2923) );
  NOR2_X1 U21359 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18227), .ZN(
        n18275) );
  NAND2_X1 U21360 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18275), .ZN(
        n18320) );
  AOI22_X1 U21361 ( .A1(n18434), .A2(n18245), .B1(n18435), .B2(n18268), .ZN(
        n18231) );
  INV_X1 U21362 ( .A(n18320), .ZN(n18311) );
  OAI211_X1 U21363 ( .C1(n18311), .C2(n18667), .A(n18229), .B(n18228), .ZN(
        n18246) );
  AOI22_X1 U21364 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18246), .B1(
        n18439), .B2(n18242), .ZN(n18230) );
  OAI211_X1 U21365 ( .C1(n18442), .C2(n18320), .A(n18231), .B(n18230), .ZN(
        P3_U2924) );
  AOI22_X1 U21366 ( .A1(n18444), .A2(n18268), .B1(n18443), .B2(n18245), .ZN(
        n18233) );
  AOI22_X1 U21367 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18246), .B1(
        n18445), .B2(n18242), .ZN(n18232) );
  OAI211_X1 U21368 ( .C1(n18449), .C2(n18320), .A(n18233), .B(n18232), .ZN(
        P3_U2925) );
  AOI22_X1 U21369 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18246), .B1(
        n18450), .B2(n18245), .ZN(n18235) );
  AOI22_X1 U21370 ( .A1(n18379), .A2(n18268), .B1(n18452), .B2(n18311), .ZN(
        n18234) );
  OAI211_X1 U21371 ( .C1(n18382), .C2(n18249), .A(n18235), .B(n18234), .ZN(
        P3_U2926) );
  AOI22_X1 U21372 ( .A1(n18329), .A2(n18268), .B1(n18456), .B2(n18245), .ZN(
        n18237) );
  AOI22_X1 U21373 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18246), .B1(
        n18458), .B2(n18311), .ZN(n18236) );
  OAI211_X1 U21374 ( .C1(n18332), .C2(n18249), .A(n18237), .B(n18236), .ZN(
        P3_U2927) );
  AOI22_X1 U21375 ( .A1(n18463), .A2(n18242), .B1(n18462), .B2(n18245), .ZN(
        n18239) );
  AOI22_X1 U21376 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18246), .B1(
        n18465), .B2(n18311), .ZN(n18238) );
  OAI211_X1 U21377 ( .C1(n18468), .C2(n18266), .A(n18239), .B(n18238), .ZN(
        P3_U2928) );
  AOI22_X1 U21378 ( .A1(n18418), .A2(n18242), .B1(n18470), .B2(n18245), .ZN(
        n18241) );
  AOI22_X1 U21379 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18246), .B1(
        n18473), .B2(n18311), .ZN(n18240) );
  OAI211_X1 U21380 ( .C1(n18421), .C2(n18266), .A(n18241), .B(n18240), .ZN(
        P3_U2929) );
  AOI22_X1 U21381 ( .A1(n18363), .A2(n18242), .B1(n18477), .B2(n18245), .ZN(
        n18244) );
  AOI22_X1 U21382 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18246), .B1(
        n18479), .B2(n18311), .ZN(n18243) );
  OAI211_X1 U21383 ( .C1(n18366), .C2(n18266), .A(n18244), .B(n18243), .ZN(
        P3_U2930) );
  AOI22_X1 U21384 ( .A1(n18485), .A2(n18268), .B1(n18484), .B2(n18245), .ZN(
        n18248) );
  AOI22_X1 U21385 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18246), .B1(
        n18488), .B2(n18311), .ZN(n18247) );
  OAI211_X1 U21386 ( .C1(n18492), .C2(n18249), .A(n18248), .B(n18247), .ZN(
        P3_U2931) );
  INV_X1 U21387 ( .A(n18321), .ZN(n18322) );
  NAND2_X1 U21388 ( .A1(n18537), .A2(n18322), .ZN(n18346) );
  AOI21_X1 U21389 ( .B1(n18320), .B2(n18346), .A(n18564), .ZN(n18267) );
  AOI22_X1 U21390 ( .A1(n18434), .A2(n18267), .B1(n18435), .B2(n18288), .ZN(
        n18253) );
  AOI221_X1 U21391 ( .B1(n18250), .B2(n18320), .C1(n18297), .C2(n18320), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18251) );
  OAI21_X1 U21392 ( .B1(n18339), .B2(n18251), .A(n18300), .ZN(n18269) );
  AOI22_X1 U21393 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18269), .B1(
        n18439), .B2(n18268), .ZN(n18252) );
  OAI211_X1 U21394 ( .C1(n18442), .C2(n18346), .A(n18253), .B(n18252), .ZN(
        P3_U2932) );
  AOI22_X1 U21395 ( .A1(n18443), .A2(n18267), .B1(n18445), .B2(n18268), .ZN(
        n18255) );
  AOI22_X1 U21396 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18269), .B1(
        n18408), .B2(n18339), .ZN(n18254) );
  OAI211_X1 U21397 ( .C1(n18411), .C2(n18295), .A(n18255), .B(n18254), .ZN(
        P3_U2933) );
  AOI22_X1 U21398 ( .A1(n18451), .A2(n18268), .B1(n18450), .B2(n18267), .ZN(
        n18257) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18269), .B1(
        n18452), .B2(n18339), .ZN(n18256) );
  OAI211_X1 U21400 ( .C1(n18455), .C2(n18295), .A(n18257), .B(n18256), .ZN(
        P3_U2934) );
  AOI22_X1 U21401 ( .A1(n18457), .A2(n18268), .B1(n18456), .B2(n18267), .ZN(
        n18259) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18269), .B1(
        n18458), .B2(n18339), .ZN(n18258) );
  OAI211_X1 U21403 ( .C1(n18461), .C2(n18295), .A(n18259), .B(n18258), .ZN(
        P3_U2935) );
  AOI22_X1 U21404 ( .A1(n18463), .A2(n18268), .B1(n18462), .B2(n18267), .ZN(
        n18261) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18269), .B1(
        n18465), .B2(n18339), .ZN(n18260) );
  OAI211_X1 U21406 ( .C1(n18468), .C2(n18295), .A(n18261), .B(n18260), .ZN(
        P3_U2936) );
  AOI22_X1 U21407 ( .A1(n18418), .A2(n18268), .B1(n18470), .B2(n18267), .ZN(
        n18263) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18269), .B1(
        n18473), .B2(n18339), .ZN(n18262) );
  OAI211_X1 U21409 ( .C1(n18421), .C2(n18295), .A(n18263), .B(n18262), .ZN(
        P3_U2937) );
  AOI22_X1 U21410 ( .A1(n18477), .A2(n18267), .B1(n18478), .B2(n18288), .ZN(
        n18265) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18269), .B1(
        n18479), .B2(n18339), .ZN(n18264) );
  OAI211_X1 U21412 ( .C1(n18482), .C2(n18266), .A(n18265), .B(n18264), .ZN(
        P3_U2938) );
  AOI22_X1 U21413 ( .A1(n18426), .A2(n18268), .B1(n18484), .B2(n18267), .ZN(
        n18271) );
  AOI22_X1 U21414 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18269), .B1(
        n18488), .B2(n18339), .ZN(n18270) );
  OAI211_X1 U21415 ( .C1(n18432), .C2(n18295), .A(n18271), .B(n18270), .ZN(
        P3_U2939) );
  NAND2_X1 U21416 ( .A1(n18322), .A2(n18272), .ZN(n18362) );
  NOR2_X1 U21417 ( .A1(n18321), .A2(n18273), .ZN(n18291) );
  AOI22_X1 U21418 ( .A1(n18434), .A2(n18291), .B1(n18435), .B2(n18311), .ZN(
        n18277) );
  AOI22_X1 U21419 ( .A1(n18374), .A2(n18275), .B1(n18322), .B2(n18274), .ZN(
        n18292) );
  AOI22_X1 U21420 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18292), .B1(
        n18439), .B2(n18288), .ZN(n18276) );
  OAI211_X1 U21421 ( .C1(n18442), .C2(n18362), .A(n18277), .B(n18276), .ZN(
        P3_U2940) );
  AOI22_X1 U21422 ( .A1(n18444), .A2(n18311), .B1(n18443), .B2(n18291), .ZN(
        n18279) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18292), .B1(
        n18445), .B2(n18288), .ZN(n18278) );
  OAI211_X1 U21424 ( .C1(n18449), .C2(n18362), .A(n18279), .B(n18278), .ZN(
        P3_U2941) );
  AOI22_X1 U21425 ( .A1(n18451), .A2(n18288), .B1(n18450), .B2(n18291), .ZN(
        n18281) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18292), .B1(
        n18452), .B2(n18369), .ZN(n18280) );
  OAI211_X1 U21427 ( .C1(n18455), .C2(n18320), .A(n18281), .B(n18280), .ZN(
        P3_U2942) );
  AOI22_X1 U21428 ( .A1(n18457), .A2(n18288), .B1(n18456), .B2(n18291), .ZN(
        n18283) );
  AOI22_X1 U21429 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18292), .B1(
        n18458), .B2(n18369), .ZN(n18282) );
  OAI211_X1 U21430 ( .C1(n18461), .C2(n18320), .A(n18283), .B(n18282), .ZN(
        P3_U2943) );
  AOI22_X1 U21431 ( .A1(n18463), .A2(n18288), .B1(n18462), .B2(n18291), .ZN(
        n18285) );
  AOI22_X1 U21432 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18292), .B1(
        n18465), .B2(n18369), .ZN(n18284) );
  OAI211_X1 U21433 ( .C1(n18468), .C2(n18320), .A(n18285), .B(n18284), .ZN(
        P3_U2944) );
  AOI22_X1 U21434 ( .A1(n18471), .A2(n18311), .B1(n18470), .B2(n18291), .ZN(
        n18287) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18292), .B1(
        n18473), .B2(n18369), .ZN(n18286) );
  OAI211_X1 U21436 ( .C1(n18476), .C2(n18295), .A(n18287), .B(n18286), .ZN(
        P3_U2945) );
  AOI22_X1 U21437 ( .A1(n18363), .A2(n18288), .B1(n18477), .B2(n18291), .ZN(
        n18290) );
  AOI22_X1 U21438 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18292), .B1(
        n18479), .B2(n18369), .ZN(n18289) );
  OAI211_X1 U21439 ( .C1(n18366), .C2(n18320), .A(n18290), .B(n18289), .ZN(
        P3_U2946) );
  AOI22_X1 U21440 ( .A1(n18485), .A2(n18311), .B1(n18484), .B2(n18291), .ZN(
        n18294) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18292), .B1(
        n18488), .B2(n18369), .ZN(n18293) );
  OAI211_X1 U21442 ( .C1(n18492), .C2(n18295), .A(n18294), .B(n18293), .ZN(
        P3_U2947) );
  NAND2_X1 U21443 ( .A1(n18296), .A2(n18322), .ZN(n18396) );
  AOI21_X1 U21444 ( .B1(n18362), .B2(n18396), .A(n18564), .ZN(n18316) );
  AOI22_X1 U21445 ( .A1(n18439), .A2(n18311), .B1(n18434), .B2(n18316), .ZN(
        n18302) );
  NOR2_X1 U21446 ( .A1(n18311), .A2(n18339), .ZN(n18298) );
  OAI211_X1 U21447 ( .C1(n18298), .C2(n18297), .A(n18362), .B(n18396), .ZN(
        n18299) );
  OAI211_X1 U21448 ( .C1(n18387), .C2(n18667), .A(n18300), .B(n18299), .ZN(
        n18317) );
  AOI22_X1 U21449 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18317), .B1(
        n18435), .B2(n18339), .ZN(n18301) );
  OAI211_X1 U21450 ( .C1(n18442), .C2(n18396), .A(n18302), .B(n18301), .ZN(
        P3_U2948) );
  AOI22_X1 U21451 ( .A1(n18443), .A2(n18316), .B1(n18445), .B2(n18311), .ZN(
        n18304) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18317), .B1(
        n18408), .B2(n18387), .ZN(n18303) );
  OAI211_X1 U21453 ( .C1(n18411), .C2(n18346), .A(n18304), .B(n18303), .ZN(
        P3_U2949) );
  AOI22_X1 U21454 ( .A1(n18379), .A2(n18339), .B1(n18450), .B2(n18316), .ZN(
        n18306) );
  AOI22_X1 U21455 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18317), .B1(
        n18452), .B2(n18387), .ZN(n18305) );
  OAI211_X1 U21456 ( .C1(n18382), .C2(n18320), .A(n18306), .B(n18305), .ZN(
        P3_U2950) );
  AOI22_X1 U21457 ( .A1(n18457), .A2(n18311), .B1(n18456), .B2(n18316), .ZN(
        n18308) );
  AOI22_X1 U21458 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18317), .B1(
        n18458), .B2(n18387), .ZN(n18307) );
  OAI211_X1 U21459 ( .C1(n18461), .C2(n18346), .A(n18308), .B(n18307), .ZN(
        P3_U2951) );
  AOI22_X1 U21460 ( .A1(n18333), .A2(n18339), .B1(n18462), .B2(n18316), .ZN(
        n18310) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18317), .B1(
        n18465), .B2(n18387), .ZN(n18309) );
  OAI211_X1 U21462 ( .C1(n18336), .C2(n18320), .A(n18310), .B(n18309), .ZN(
        P3_U2952) );
  AOI22_X1 U21463 ( .A1(n18418), .A2(n18311), .B1(n18470), .B2(n18316), .ZN(
        n18313) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18317), .B1(
        n18473), .B2(n18387), .ZN(n18312) );
  OAI211_X1 U21465 ( .C1(n18421), .C2(n18346), .A(n18313), .B(n18312), .ZN(
        P3_U2953) );
  AOI22_X1 U21466 ( .A1(n18477), .A2(n18316), .B1(n18478), .B2(n18339), .ZN(
        n18315) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18317), .B1(
        n18479), .B2(n18387), .ZN(n18314) );
  OAI211_X1 U21468 ( .C1(n18482), .C2(n18320), .A(n18315), .B(n18314), .ZN(
        P3_U2954) );
  AOI22_X1 U21469 ( .A1(n18485), .A2(n18339), .B1(n18484), .B2(n18316), .ZN(
        n18319) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18317), .B1(
        n18488), .B2(n18387), .ZN(n18318) );
  OAI211_X1 U21471 ( .C1(n18492), .C2(n18320), .A(n18319), .B(n18318), .ZN(
        P3_U2955) );
  NOR2_X1 U21472 ( .A1(n18534), .A2(n18321), .ZN(n18373) );
  NAND2_X1 U21473 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18373), .ZN(
        n18424) );
  AND2_X1 U21474 ( .A1(n18433), .A2(n18373), .ZN(n18342) );
  AOI22_X1 U21475 ( .A1(n18439), .A2(n18339), .B1(n18434), .B2(n18342), .ZN(
        n18324) );
  AOI22_X1 U21476 ( .A1(n18374), .A2(n18322), .B1(n18373), .B2(n18436), .ZN(
        n18343) );
  AOI22_X1 U21477 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18343), .B1(
        n18435), .B2(n18369), .ZN(n18323) );
  OAI211_X1 U21478 ( .C1(n18424), .C2(n18442), .A(n18324), .B(n18323), .ZN(
        P3_U2956) );
  AOI22_X1 U21479 ( .A1(n18444), .A2(n18369), .B1(n18443), .B2(n18342), .ZN(
        n18326) );
  AOI22_X1 U21480 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18343), .B1(
        n18445), .B2(n18339), .ZN(n18325) );
  OAI211_X1 U21481 ( .C1(n18424), .C2(n18449), .A(n18326), .B(n18325), .ZN(
        P3_U2957) );
  AOI22_X1 U21482 ( .A1(n18379), .A2(n18369), .B1(n18450), .B2(n18342), .ZN(
        n18328) );
  AOI22_X1 U21483 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18343), .B1(
        n18427), .B2(n18452), .ZN(n18327) );
  OAI211_X1 U21484 ( .C1(n18382), .C2(n18346), .A(n18328), .B(n18327), .ZN(
        P3_U2958) );
  AOI22_X1 U21485 ( .A1(n18329), .A2(n18369), .B1(n18456), .B2(n18342), .ZN(
        n18331) );
  AOI22_X1 U21486 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18343), .B1(
        n18427), .B2(n18458), .ZN(n18330) );
  OAI211_X1 U21487 ( .C1(n18332), .C2(n18346), .A(n18331), .B(n18330), .ZN(
        P3_U2959) );
  AOI22_X1 U21488 ( .A1(n18333), .A2(n18369), .B1(n18462), .B2(n18342), .ZN(
        n18335) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18343), .B1(
        n18427), .B2(n18465), .ZN(n18334) );
  OAI211_X1 U21490 ( .C1(n18336), .C2(n18346), .A(n18335), .B(n18334), .ZN(
        P3_U2960) );
  AOI22_X1 U21491 ( .A1(n18418), .A2(n18339), .B1(n18470), .B2(n18342), .ZN(
        n18338) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18343), .B1(
        n18427), .B2(n18473), .ZN(n18337) );
  OAI211_X1 U21493 ( .C1(n18421), .C2(n18362), .A(n18338), .B(n18337), .ZN(
        P3_U2961) );
  AOI22_X1 U21494 ( .A1(n18363), .A2(n18339), .B1(n18477), .B2(n18342), .ZN(
        n18341) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18343), .B1(
        n18427), .B2(n18479), .ZN(n18340) );
  OAI211_X1 U21496 ( .C1(n18366), .C2(n18362), .A(n18341), .B(n18340), .ZN(
        P3_U2962) );
  AOI22_X1 U21497 ( .A1(n18485), .A2(n18369), .B1(n18484), .B2(n18342), .ZN(
        n18345) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18343), .B1(
        n18427), .B2(n18488), .ZN(n18344) );
  OAI211_X1 U21499 ( .C1(n18492), .C2(n18346), .A(n18345), .B(n18344), .ZN(
        P3_U2963) );
  INV_X1 U21500 ( .A(n18372), .ZN(n18438) );
  NAND2_X1 U21501 ( .A1(n18438), .A2(n18533), .ZN(n18493) );
  NAND2_X1 U21502 ( .A1(n18493), .A2(n18424), .ZN(n18397) );
  AOI21_X1 U21503 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18493), .A(n18399), 
        .ZN(n18347) );
  OAI221_X1 U21504 ( .B1(n18397), .B2(n18349), .C1(n18397), .C2(n18348), .A(
        n18347), .ZN(n18368) );
  AND2_X1 U21505 ( .A1(n18433), .A2(n18397), .ZN(n18367) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18368), .B1(
        n18434), .B2(n18367), .ZN(n18351) );
  AOI22_X1 U21507 ( .A1(n18439), .A2(n18369), .B1(n18435), .B2(n18387), .ZN(
        n18350) );
  OAI211_X1 U21508 ( .C1(n18493), .C2(n18442), .A(n18351), .B(n18350), .ZN(
        P3_U2964) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18368), .B1(
        n18443), .B2(n18367), .ZN(n18353) );
  INV_X1 U21510 ( .A(n18493), .ZN(n18464) );
  AOI22_X1 U21511 ( .A1(n18464), .A2(n18408), .B1(n18445), .B2(n18369), .ZN(
        n18352) );
  OAI211_X1 U21512 ( .C1(n18411), .C2(n18396), .A(n18353), .B(n18352), .ZN(
        P3_U2965) );
  AOI22_X1 U21513 ( .A1(n18379), .A2(n18387), .B1(n18450), .B2(n18367), .ZN(
        n18355) );
  AOI22_X1 U21514 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18368), .B1(
        n18464), .B2(n18452), .ZN(n18354) );
  OAI211_X1 U21515 ( .C1(n18382), .C2(n18362), .A(n18355), .B(n18354), .ZN(
        P3_U2966) );
  AOI22_X1 U21516 ( .A1(n18457), .A2(n18369), .B1(n18456), .B2(n18367), .ZN(
        n18357) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18368), .B1(
        n18464), .B2(n18458), .ZN(n18356) );
  OAI211_X1 U21518 ( .C1(n18461), .C2(n18396), .A(n18357), .B(n18356), .ZN(
        P3_U2967) );
  AOI22_X1 U21519 ( .A1(n18463), .A2(n18369), .B1(n18462), .B2(n18367), .ZN(
        n18359) );
  AOI22_X1 U21520 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18368), .B1(
        n18464), .B2(n18465), .ZN(n18358) );
  OAI211_X1 U21521 ( .C1(n18468), .C2(n18396), .A(n18359), .B(n18358), .ZN(
        P3_U2968) );
  AOI22_X1 U21522 ( .A1(n18471), .A2(n18387), .B1(n18470), .B2(n18367), .ZN(
        n18361) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18368), .B1(
        n18464), .B2(n18473), .ZN(n18360) );
  OAI211_X1 U21524 ( .C1(n18476), .C2(n18362), .A(n18361), .B(n18360), .ZN(
        P3_U2969) );
  AOI22_X1 U21525 ( .A1(n18363), .A2(n18369), .B1(n18477), .B2(n18367), .ZN(
        n18365) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18368), .B1(
        n18464), .B2(n18479), .ZN(n18364) );
  OAI211_X1 U21527 ( .C1(n18366), .C2(n18396), .A(n18365), .B(n18364), .ZN(
        P3_U2970) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18368), .B1(
        n18484), .B2(n18367), .ZN(n18371) );
  AOI22_X1 U21529 ( .A1(n18464), .A2(n18488), .B1(n18426), .B2(n18369), .ZN(
        n18370) );
  OAI211_X1 U21530 ( .C1(n18432), .C2(n18396), .A(n18371), .B(n18370), .ZN(
        P3_U2971) );
  NOR2_X1 U21531 ( .A1(n18564), .A2(n18372), .ZN(n18392) );
  AOI22_X1 U21532 ( .A1(n18439), .A2(n18387), .B1(n18434), .B2(n18392), .ZN(
        n18376) );
  AOI22_X1 U21533 ( .A1(n18374), .A2(n18373), .B1(n18438), .B2(n18436), .ZN(
        n18393) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18393), .B1(
        n18427), .B2(n18435), .ZN(n18375) );
  OAI211_X1 U21535 ( .C1(n18469), .C2(n18442), .A(n18376), .B(n18375), .ZN(
        P3_U2972) );
  AOI22_X1 U21536 ( .A1(n18443), .A2(n18392), .B1(n18445), .B2(n18387), .ZN(
        n18378) );
  AOI22_X1 U21537 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18393), .B1(
        n18486), .B2(n18408), .ZN(n18377) );
  OAI211_X1 U21538 ( .C1(n18424), .C2(n18411), .A(n18378), .B(n18377), .ZN(
        P3_U2973) );
  AOI22_X1 U21539 ( .A1(n18427), .A2(n18379), .B1(n18450), .B2(n18392), .ZN(
        n18381) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18393), .B1(
        n18486), .B2(n18452), .ZN(n18380) );
  OAI211_X1 U21541 ( .C1(n18382), .C2(n18396), .A(n18381), .B(n18380), .ZN(
        P3_U2974) );
  AOI22_X1 U21542 ( .A1(n18457), .A2(n18387), .B1(n18456), .B2(n18392), .ZN(
        n18384) );
  AOI22_X1 U21543 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18393), .B1(
        n18472), .B2(n18458), .ZN(n18383) );
  OAI211_X1 U21544 ( .C1(n18424), .C2(n18461), .A(n18384), .B(n18383), .ZN(
        P3_U2975) );
  AOI22_X1 U21545 ( .A1(n18463), .A2(n18387), .B1(n18462), .B2(n18392), .ZN(
        n18386) );
  AOI22_X1 U21546 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18393), .B1(
        n18472), .B2(n18465), .ZN(n18385) );
  OAI211_X1 U21547 ( .C1(n18424), .C2(n18468), .A(n18386), .B(n18385), .ZN(
        P3_U2976) );
  AOI22_X1 U21548 ( .A1(n18418), .A2(n18387), .B1(n18470), .B2(n18392), .ZN(
        n18389) );
  AOI22_X1 U21549 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18393), .B1(
        n18486), .B2(n18473), .ZN(n18388) );
  OAI211_X1 U21550 ( .C1(n18424), .C2(n18421), .A(n18389), .B(n18388), .ZN(
        P3_U2977) );
  AOI22_X1 U21551 ( .A1(n18427), .A2(n18478), .B1(n18477), .B2(n18392), .ZN(
        n18391) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18393), .B1(
        n18486), .B2(n18479), .ZN(n18390) );
  OAI211_X1 U21553 ( .C1(n18482), .C2(n18396), .A(n18391), .B(n18390), .ZN(
        P3_U2978) );
  AOI22_X1 U21554 ( .A1(n18427), .A2(n18485), .B1(n18484), .B2(n18392), .ZN(
        n18395) );
  AOI22_X1 U21555 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18393), .B1(
        n18472), .B2(n18488), .ZN(n18394) );
  OAI211_X1 U21556 ( .C1(n18492), .C2(n18396), .A(n18395), .B(n18394), .ZN(
        P3_U2979) );
  OAI221_X1 U21557 ( .B1(n18486), .B2(n18398), .C1(n18486), .C2(n18397), .A(
        n18667), .ZN(n18400) );
  AOI21_X1 U21558 ( .B1(n18401), .B2(n18400), .A(n18399), .ZN(n18407) );
  NOR2_X1 U21559 ( .A1(n18564), .A2(n18402), .ZN(n18425) );
  AOI22_X1 U21560 ( .A1(n18464), .A2(n18435), .B1(n18434), .B2(n18425), .ZN(
        n18405) );
  AOI22_X1 U21561 ( .A1(n18428), .A2(n18403), .B1(n18427), .B2(n18439), .ZN(
        n18404) );
  OAI211_X1 U21562 ( .C1(n18407), .C2(n18406), .A(n18405), .B(n18404), .ZN(
        P3_U2980) );
  AOI22_X1 U21563 ( .A1(n18427), .A2(n18445), .B1(n18425), .B2(n18443), .ZN(
        n18410) );
  INV_X1 U21564 ( .A(n18407), .ZN(n18429) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18429), .B1(
        n18428), .B2(n18408), .ZN(n18409) );
  OAI211_X1 U21566 ( .C1(n18493), .C2(n18411), .A(n18410), .B(n18409), .ZN(
        P3_U2981) );
  AOI22_X1 U21567 ( .A1(n18427), .A2(n18451), .B1(n18425), .B2(n18450), .ZN(
        n18413) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18429), .B1(
        n18428), .B2(n18452), .ZN(n18412) );
  OAI211_X1 U21569 ( .C1(n18493), .C2(n18455), .A(n18413), .B(n18412), .ZN(
        P3_U2982) );
  AOI22_X1 U21570 ( .A1(n18427), .A2(n18457), .B1(n18425), .B2(n18456), .ZN(
        n18415) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18429), .B1(
        n18428), .B2(n18458), .ZN(n18414) );
  OAI211_X1 U21572 ( .C1(n18493), .C2(n18461), .A(n18415), .B(n18414), .ZN(
        P3_U2983) );
  AOI22_X1 U21573 ( .A1(n18427), .A2(n18463), .B1(n18425), .B2(n18462), .ZN(
        n18417) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18429), .B1(
        n18428), .B2(n18465), .ZN(n18416) );
  OAI211_X1 U21575 ( .C1(n18493), .C2(n18468), .A(n18417), .B(n18416), .ZN(
        P3_U2984) );
  AOI22_X1 U21576 ( .A1(n18427), .A2(n18418), .B1(n18425), .B2(n18470), .ZN(
        n18420) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18429), .B1(
        n18428), .B2(n18473), .ZN(n18419) );
  OAI211_X1 U21578 ( .C1(n18493), .C2(n18421), .A(n18420), .B(n18419), .ZN(
        P3_U2985) );
  AOI22_X1 U21579 ( .A1(n18464), .A2(n18478), .B1(n18425), .B2(n18477), .ZN(
        n18423) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18429), .B1(
        n18428), .B2(n18479), .ZN(n18422) );
  OAI211_X1 U21581 ( .C1(n18424), .C2(n18482), .A(n18423), .B(n18422), .ZN(
        P3_U2986) );
  AOI22_X1 U21582 ( .A1(n18427), .A2(n18426), .B1(n18425), .B2(n18484), .ZN(
        n18431) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18429), .B1(
        n18428), .B2(n18488), .ZN(n18430) );
  OAI211_X1 U21584 ( .C1(n18493), .C2(n18432), .A(n18431), .B(n18430), .ZN(
        P3_U2987) );
  AND2_X1 U21585 ( .A1(n18433), .A2(n18437), .ZN(n18483) );
  AOI22_X1 U21586 ( .A1(n18486), .A2(n18435), .B1(n18434), .B2(n18483), .ZN(
        n18441) );
  AOI22_X1 U21587 ( .A1(n18374), .A2(n18438), .B1(n18437), .B2(n18436), .ZN(
        n18489) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18489), .B1(
        n18464), .B2(n18439), .ZN(n18440) );
  OAI211_X1 U21589 ( .C1(n18442), .C2(n18448), .A(n18441), .B(n18440), .ZN(
        P3_U2988) );
  AOI22_X1 U21590 ( .A1(n18472), .A2(n18444), .B1(n18443), .B2(n18483), .ZN(
        n18447) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18489), .B1(
        n18464), .B2(n18445), .ZN(n18446) );
  OAI211_X1 U21592 ( .C1(n18449), .C2(n18448), .A(n18447), .B(n18446), .ZN(
        P3_U2989) );
  AOI22_X1 U21593 ( .A1(n18464), .A2(n18451), .B1(n18450), .B2(n18483), .ZN(
        n18454) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18489), .B1(
        n18452), .B2(n18487), .ZN(n18453) );
  OAI211_X1 U21595 ( .C1(n18469), .C2(n18455), .A(n18454), .B(n18453), .ZN(
        P3_U2990) );
  AOI22_X1 U21596 ( .A1(n18464), .A2(n18457), .B1(n18456), .B2(n18483), .ZN(
        n18460) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18489), .B1(
        n18458), .B2(n18487), .ZN(n18459) );
  OAI211_X1 U21598 ( .C1(n18469), .C2(n18461), .A(n18460), .B(n18459), .ZN(
        P3_U2991) );
  AOI22_X1 U21599 ( .A1(n18464), .A2(n18463), .B1(n18462), .B2(n18483), .ZN(
        n18467) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18489), .B1(
        n18465), .B2(n18487), .ZN(n18466) );
  OAI211_X1 U21601 ( .C1(n18469), .C2(n18468), .A(n18467), .B(n18466), .ZN(
        P3_U2992) );
  AOI22_X1 U21602 ( .A1(n18472), .A2(n18471), .B1(n18470), .B2(n18483), .ZN(
        n18475) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18489), .B1(
        n18473), .B2(n18487), .ZN(n18474) );
  OAI211_X1 U21604 ( .C1(n18493), .C2(n18476), .A(n18475), .B(n18474), .ZN(
        P3_U2993) );
  AOI22_X1 U21605 ( .A1(n18486), .A2(n18478), .B1(n18477), .B2(n18483), .ZN(
        n18481) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18489), .B1(
        n18479), .B2(n18487), .ZN(n18480) );
  OAI211_X1 U21607 ( .C1(n18493), .C2(n18482), .A(n18481), .B(n18480), .ZN(
        P3_U2994) );
  AOI22_X1 U21608 ( .A1(n18486), .A2(n18485), .B1(n18484), .B2(n18483), .ZN(
        n18491) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18489), .B1(
        n18488), .B2(n18487), .ZN(n18490) );
  OAI211_X1 U21610 ( .C1(n18493), .C2(n18492), .A(n18491), .B(n18490), .ZN(
        P3_U2995) );
  NOR2_X1 U21611 ( .A1(n18519), .A2(n18494), .ZN(n18496) );
  OAI222_X1 U21612 ( .A1(n18500), .A2(n18499), .B1(n18498), .B2(n18497), .C1(
        n18496), .C2(n9580), .ZN(n18709) );
  OAI21_X1 U21613 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18501), .ZN(n18502) );
  OAI211_X1 U21614 ( .C1(n18504), .C2(n18538), .A(n18503), .B(n18502), .ZN(
        n18551) );
  NAND2_X1 U21615 ( .A1(n18505), .A2(n16736), .ZN(n18530) );
  AOI22_X1 U21616 ( .A1(n18506), .A2(n18530), .B1(n18519), .B2(n18511), .ZN(
        n18507) );
  NOR2_X1 U21617 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18507), .ZN(
        n18669) );
  AOI21_X1 U21618 ( .B1(n18510), .B2(n18509), .A(n18508), .ZN(n18516) );
  OAI21_X1 U21619 ( .B1(n18516), .B2(n18512), .A(n18511), .ZN(n18513) );
  AOI21_X1 U21620 ( .B1(n18522), .B2(n18532), .A(n18513), .ZN(n18670) );
  AOI21_X1 U21621 ( .B1(n18670), .B2(n18538), .A(n18672), .ZN(n18514) );
  AOI21_X1 U21622 ( .B1(n18538), .B2(n18669), .A(n18514), .ZN(n18549) );
  INV_X1 U21623 ( .A(n18538), .ZN(n18527) );
  AOI221_X1 U21624 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18516), 
        .C1(n18515), .C2(n18516), .A(n18682), .ZN(n18518) );
  AOI22_X1 U21625 ( .A1(n18519), .A2(n18678), .B1(n18518), .B2(n18517), .ZN(
        n18526) );
  NOR2_X1 U21626 ( .A1(n18529), .A2(n16736), .ZN(n18521) );
  OAI211_X1 U21627 ( .C1(n18521), .C2(n18520), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n18682), .ZN(n18525) );
  OAI211_X1 U21628 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18523), .B(n18522), .ZN(
        n18524) );
  NAND3_X1 U21629 ( .A1(n18526), .A2(n18525), .A3(n18524), .ZN(n18680) );
  AOI22_X1 U21630 ( .A1(n18527), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18680), .B2(n18538), .ZN(n18541) );
  NAND2_X1 U21631 ( .A1(n18529), .A2(n18528), .ZN(n18531) );
  AOI22_X1 U21632 ( .A1(n18687), .A2(n18531), .B1(n18690), .B2(n18530), .ZN(
        n18683) );
  AOI22_X1 U21633 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18532), .B1(
        n18531), .B2(n16736), .ZN(n18535) );
  INV_X1 U21634 ( .A(n18535), .ZN(n18692) );
  NOR3_X1 U21635 ( .A1(n18534), .A2(n18533), .A3(n18692), .ZN(n18536) );
  OAI22_X1 U21636 ( .A1(n18683), .A2(n18536), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18535), .ZN(n18539) );
  AOI21_X1 U21637 ( .B1(n18539), .B2(n18538), .A(n18537), .ZN(n18540) );
  AOI21_X1 U21638 ( .B1(n18541), .B2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n18540), .ZN(n18542) );
  INV_X1 U21639 ( .A(n18541), .ZN(n18543) );
  AOI221_X1 U21640 ( .B1(n18542), .B2(n18545), .C1(n18544), .C2(n18545), .A(
        n18543), .ZN(n18548) );
  AOI21_X1 U21641 ( .B1(n20885), .B2(n18543), .A(n18542), .ZN(n18547) );
  NAND2_X1 U21642 ( .A1(n18545), .A2(n18544), .ZN(n18546) );
  OAI22_X1 U21643 ( .A1(n18549), .A2(n18548), .B1(n18547), .B2(n18546), .ZN(
        n18550) );
  NOR4_X1 U21644 ( .A1(n18552), .A2(n18709), .A3(n18551), .A4(n18550), .ZN(
        n18562) );
  AOI22_X1 U21645 ( .A1(n18691), .A2(n18720), .B1(n18578), .B2(n18713), .ZN(
        n18553) );
  INV_X1 U21646 ( .A(n18553), .ZN(n18558) );
  OAI211_X1 U21647 ( .C1(n18555), .C2(n18554), .A(n18711), .B(n18562), .ZN(
        n18666) );
  OAI21_X1 U21648 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18717), .A(n18666), 
        .ZN(n18565) );
  NOR2_X1 U21649 ( .A1(n18556), .A2(n18565), .ZN(n18557) );
  MUX2_X1 U21650 ( .A(n18558), .B(n18557), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18560) );
  OAI211_X1 U21651 ( .C1(n18562), .C2(n18561), .A(n18560), .B(n18559), .ZN(
        P3_U2996) );
  NAND2_X1 U21652 ( .A1(n18578), .A2(n18713), .ZN(n18568) );
  NAND4_X1 U21653 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18578), .A4(n18563), .ZN(n18571) );
  OR3_X1 U21654 ( .A1(n18566), .A2(n18565), .A3(n18564), .ZN(n18567) );
  NAND4_X1 U21655 ( .A1(n18569), .A2(n18568), .A3(n18571), .A4(n18567), .ZN(
        P3_U2997) );
  OAI21_X1 U21656 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18570), .ZN(n18573) );
  INV_X1 U21657 ( .A(n18571), .ZN(n18572) );
  AOI21_X1 U21658 ( .B1(n18574), .B2(n18573), .A(n18572), .ZN(P3_U2998) );
  AND2_X1 U21659 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18660), .ZN(
        P3_U2999) );
  AND2_X1 U21660 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18660), .ZN(
        P3_U3000) );
  AND2_X1 U21661 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18575), .ZN(
        P3_U3001) );
  AND2_X1 U21662 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18575), .ZN(
        P3_U3002) );
  AND2_X1 U21663 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18575), .ZN(
        P3_U3003) );
  AND2_X1 U21664 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18575), .ZN(
        P3_U3004) );
  AND2_X1 U21665 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18575), .ZN(
        P3_U3005) );
  AND2_X1 U21666 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18575), .ZN(
        P3_U3006) );
  AND2_X1 U21667 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18575), .ZN(
        P3_U3007) );
  AND2_X1 U21668 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18575), .ZN(
        P3_U3008) );
  AND2_X1 U21669 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18575), .ZN(
        P3_U3009) );
  AND2_X1 U21670 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18575), .ZN(
        P3_U3010) );
  AND2_X1 U21671 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18575), .ZN(
        P3_U3011) );
  AND2_X1 U21672 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18575), .ZN(
        P3_U3012) );
  AND2_X1 U21673 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18575), .ZN(
        P3_U3013) );
  AND2_X1 U21674 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18575), .ZN(
        P3_U3014) );
  AND2_X1 U21675 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18575), .ZN(
        P3_U3015) );
  AND2_X1 U21676 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18575), .ZN(
        P3_U3016) );
  AND2_X1 U21677 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18575), .ZN(
        P3_U3017) );
  AND2_X1 U21678 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18575), .ZN(
        P3_U3018) );
  AND2_X1 U21679 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18660), .ZN(
        P3_U3019) );
  AND2_X1 U21680 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18660), .ZN(
        P3_U3020) );
  AND2_X1 U21681 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18575), .ZN(P3_U3021) );
  AND2_X1 U21682 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18660), .ZN(P3_U3022) );
  AND2_X1 U21683 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18660), .ZN(P3_U3023) );
  AND2_X1 U21684 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18660), .ZN(P3_U3024) );
  AND2_X1 U21685 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18660), .ZN(P3_U3025) );
  AND2_X1 U21686 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18660), .ZN(P3_U3026) );
  AND2_X1 U21687 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18660), .ZN(P3_U3027) );
  AND2_X1 U21688 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18660), .ZN(P3_U3028) );
  OAI21_X1 U21689 ( .B1(n18576), .B2(n20683), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18577) );
  AOI21_X1 U21690 ( .B1(NA), .B2(n18589), .A(n18577), .ZN(n18580) );
  NAND2_X1 U21691 ( .A1(n18578), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18584) );
  NAND2_X1 U21692 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18584), .ZN(n18587) );
  INV_X1 U21693 ( .A(n18587), .ZN(n18579) );
  OAI22_X1 U21694 ( .A1(n18658), .A2(n18580), .B1(P3_STATE_REG_2__SCAN_IN), 
        .B2(n18579), .ZN(P3_U3029) );
  NOR2_X1 U21695 ( .A1(n18591), .A2(n20683), .ZN(n18586) );
  INV_X1 U21696 ( .A(n18586), .ZN(n18582) );
  AOI22_X1 U21697 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n18582), .B1(HOLD), 
        .B2(n18581), .ZN(n18583) );
  OAI211_X1 U21698 ( .C1(n18583), .C2(n18589), .A(n18584), .B(n18714), .ZN(
        P3_U3030) );
  OAI22_X1 U21699 ( .A1(NA), .A2(n18584), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18585) );
  OAI22_X1 U21700 ( .A1(n18586), .A2(n18585), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18590) );
  INV_X1 U21701 ( .A(NA), .ZN(n20689) );
  OAI211_X1 U21702 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(n20689), .A(
        P3_STATE_REG_2__SCAN_IN), .B(n18587), .ZN(n18588) );
  OAI21_X1 U21703 ( .B1(n18590), .B2(n18589), .A(n18588), .ZN(P3_U3031) );
  OAI222_X1 U21704 ( .A1(n18638), .A2(n20923), .B1(n18592), .B2(n18658), .C1(
        n18698), .C2(n18652), .ZN(P3_U3032) );
  OAI222_X1 U21705 ( .A1(n20923), .A2(n18652), .B1(n18593), .B2(n18658), .C1(
        n18594), .C2(n18638), .ZN(P3_U3033) );
  INV_X1 U21706 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18596) );
  OAI222_X1 U21707 ( .A1(n18638), .A2(n18596), .B1(n18595), .B2(n18658), .C1(
        n18594), .C2(n18652), .ZN(P3_U3034) );
  OAI222_X1 U21708 ( .A1(n18638), .A2(n18598), .B1(n18597), .B2(n18658), .C1(
        n18596), .C2(n18652), .ZN(P3_U3035) );
  OAI222_X1 U21709 ( .A1(n18638), .A2(n18600), .B1(n18599), .B2(n18658), .C1(
        n18598), .C2(n18652), .ZN(P3_U3036) );
  OAI222_X1 U21710 ( .A1(n18638), .A2(n18602), .B1(n18601), .B2(n18658), .C1(
        n18600), .C2(n18652), .ZN(P3_U3037) );
  INV_X1 U21711 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18604) );
  OAI222_X1 U21712 ( .A1(n18638), .A2(n18604), .B1(n18603), .B2(n18658), .C1(
        n18602), .C2(n18652), .ZN(P3_U3038) );
  OAI222_X1 U21713 ( .A1(n18638), .A2(n18606), .B1(n18605), .B2(n18658), .C1(
        n18604), .C2(n18652), .ZN(P3_U3039) );
  OAI222_X1 U21714 ( .A1(n18638), .A2(n18608), .B1(n18607), .B2(n18658), .C1(
        n18606), .C2(n18652), .ZN(P3_U3040) );
  OAI222_X1 U21715 ( .A1(n18638), .A2(n18610), .B1(n18609), .B2(n18658), .C1(
        n18608), .C2(n18652), .ZN(P3_U3041) );
  INV_X1 U21716 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18612) );
  OAI222_X1 U21717 ( .A1(n18638), .A2(n18612), .B1(n18611), .B2(n18658), .C1(
        n18610), .C2(n18652), .ZN(P3_U3042) );
  OAI222_X1 U21718 ( .A1(n18638), .A2(n18614), .B1(n18613), .B2(n18658), .C1(
        n18612), .C2(n18652), .ZN(P3_U3043) );
  OAI222_X1 U21719 ( .A1(n18638), .A2(n18616), .B1(n18615), .B2(n18658), .C1(
        n18614), .C2(n18652), .ZN(P3_U3044) );
  OAI222_X1 U21720 ( .A1(n18638), .A2(n18618), .B1(n18617), .B2(n18658), .C1(
        n18616), .C2(n18652), .ZN(P3_U3045) );
  OAI222_X1 U21721 ( .A1(n18638), .A2(n18620), .B1(n18619), .B2(n18658), .C1(
        n18618), .C2(n18652), .ZN(P3_U3046) );
  OAI222_X1 U21722 ( .A1(n18638), .A2(n18623), .B1(n18621), .B2(n18658), .C1(
        n18620), .C2(n18652), .ZN(P3_U3047) );
  OAI222_X1 U21723 ( .A1(n18623), .A2(n18652), .B1(n18622), .B2(n18658), .C1(
        n18624), .C2(n18638), .ZN(P3_U3048) );
  OAI222_X1 U21724 ( .A1(n18638), .A2(n18626), .B1(n18625), .B2(n18658), .C1(
        n18624), .C2(n18652), .ZN(P3_U3049) );
  OAI222_X1 U21725 ( .A1(n18638), .A2(n18628), .B1(n18627), .B2(n18658), .C1(
        n18626), .C2(n18652), .ZN(P3_U3050) );
  OAI222_X1 U21726 ( .A1(n18638), .A2(n18630), .B1(n18629), .B2(n18658), .C1(
        n18628), .C2(n18652), .ZN(P3_U3051) );
  OAI222_X1 U21727 ( .A1(n18638), .A2(n18632), .B1(n18631), .B2(n18658), .C1(
        n18630), .C2(n18652), .ZN(P3_U3052) );
  OAI222_X1 U21728 ( .A1(n18638), .A2(n18634), .B1(n18633), .B2(n18658), .C1(
        n18632), .C2(n18652), .ZN(P3_U3053) );
  OAI222_X1 U21729 ( .A1(n18638), .A2(n18636), .B1(n18635), .B2(n18658), .C1(
        n18634), .C2(n18652), .ZN(P3_U3054) );
  OAI222_X1 U21730 ( .A1(n18638), .A2(n18639), .B1(n18637), .B2(n18658), .C1(
        n18636), .C2(n18652), .ZN(P3_U3055) );
  OAI222_X1 U21731 ( .A1(n18638), .A2(n18641), .B1(n18640), .B2(n18658), .C1(
        n18639), .C2(n18652), .ZN(P3_U3056) );
  OAI222_X1 U21732 ( .A1(n18638), .A2(n18643), .B1(n18642), .B2(n18658), .C1(
        n18641), .C2(n18652), .ZN(P3_U3057) );
  INV_X1 U21733 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18646) );
  OAI222_X1 U21734 ( .A1(n18638), .A2(n18646), .B1(n18644), .B2(n18658), .C1(
        n18643), .C2(n18652), .ZN(P3_U3058) );
  OAI222_X1 U21735 ( .A1(n18646), .A2(n18652), .B1(n18645), .B2(n18658), .C1(
        n18647), .C2(n18638), .ZN(P3_U3059) );
  OAI222_X1 U21736 ( .A1(n18638), .A2(n18651), .B1(n18648), .B2(n18658), .C1(
        n18647), .C2(n18652), .ZN(P3_U3060) );
  OAI222_X1 U21737 ( .A1(n18652), .A2(n18651), .B1(n18650), .B2(n18658), .C1(
        n18649), .C2(n18638), .ZN(P3_U3061) );
  INV_X1 U21738 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18653) );
  AOI22_X1 U21739 ( .A1(n18658), .A2(n18654), .B1(n18653), .B2(n18725), .ZN(
        P3_U3274) );
  INV_X1 U21740 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18700) );
  INV_X1 U21741 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18655) );
  AOI22_X1 U21742 ( .A1(n18658), .A2(n18700), .B1(n18655), .B2(n18725), .ZN(
        P3_U3275) );
  INV_X1 U21743 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18656) );
  AOI22_X1 U21744 ( .A1(n18658), .A2(n20862), .B1(n18656), .B2(n18725), .ZN(
        P3_U3276) );
  INV_X1 U21745 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18706) );
  INV_X1 U21746 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18657) );
  AOI22_X1 U21747 ( .A1(n18658), .A2(n18706), .B1(n18657), .B2(n18725), .ZN(
        P3_U3277) );
  INV_X1 U21748 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18661) );
  INV_X1 U21749 ( .A(n18662), .ZN(n18659) );
  AOI21_X1 U21750 ( .B1(n18661), .B2(n18660), .A(n18659), .ZN(P3_U3280) );
  OAI21_X1 U21751 ( .B1(n18664), .B2(n18663), .A(n18662), .ZN(P3_U3281) );
  OAI221_X1 U21752 ( .B1(n18667), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18667), 
        .C2(n18666), .A(n18665), .ZN(P3_U3282) );
  AOI22_X1 U21753 ( .A1(n18693), .A2(n18669), .B1(n18691), .B2(n18668), .ZN(
        n18674) );
  INV_X1 U21754 ( .A(n18670), .ZN(n18671) );
  AOI21_X1 U21755 ( .B1(n18693), .B2(n18671), .A(n18697), .ZN(n18673) );
  OAI22_X1 U21756 ( .A1(n18697), .A2(n18674), .B1(n18673), .B2(n18672), .ZN(
        P3_U3285) );
  NOR2_X1 U21757 ( .A1(n18675), .A2(n18694), .ZN(n18685) );
  AOI22_X1 U21758 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18677), .B2(n18676), .ZN(
        n18684) );
  INV_X1 U21759 ( .A(n18678), .ZN(n18679) );
  AOI222_X1 U21760 ( .A1(n18680), .A2(n18693), .B1(n18685), .B2(n18684), .C1(
        n18691), .C2(n18679), .ZN(n18681) );
  AOI22_X1 U21761 ( .A1(n18697), .A2(n18682), .B1(n18681), .B2(n18695), .ZN(
        P3_U3288) );
  INV_X1 U21762 ( .A(n18683), .ZN(n18688) );
  INV_X1 U21763 ( .A(n18684), .ZN(n18686) );
  AOI222_X1 U21764 ( .A1(n18688), .A2(n18693), .B1(n18691), .B2(n18687), .C1(
        n18686), .C2(n18685), .ZN(n18689) );
  AOI22_X1 U21765 ( .A1(n18697), .A2(n18690), .B1(n18689), .B2(n18695), .ZN(
        P3_U3289) );
  AOI222_X1 U21766 ( .A1(n18694), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18693), 
        .B2(n18692), .C1(n16736), .C2(n18691), .ZN(n18696) );
  AOI22_X1 U21767 ( .A1(n18697), .A2(n16736), .B1(n18696), .B2(n18695), .ZN(
        P3_U3290) );
  AOI21_X1 U21768 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18699) );
  AOI22_X1 U21769 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18699), .B2(n18698), .ZN(n18701) );
  AOI22_X1 U21770 ( .A1(n18702), .A2(n18701), .B1(n18700), .B2(n18705), .ZN(
        P3_U3292) );
  NOR2_X1 U21771 ( .A1(n18705), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18703) );
  AOI22_X1 U21772 ( .A1(n18706), .A2(n18705), .B1(n18704), .B2(n18703), .ZN(
        P3_U3293) );
  INV_X1 U21773 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18707) );
  AOI22_X1 U21774 ( .A1(n18658), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18707), 
        .B2(n18725), .ZN(P3_U3294) );
  MUX2_X1 U21775 ( .A(P3_MORE_REG_SCAN_IN), .B(n18709), .S(n18708), .Z(
        P3_U3295) );
  OAI21_X1 U21776 ( .B1(n18711), .B2(n18710), .A(n18729), .ZN(n18712) );
  AOI21_X1 U21777 ( .B1(n18713), .B2(n18717), .A(n18712), .ZN(n18724) );
  INV_X1 U21778 ( .A(n18728), .ZN(n18719) );
  AOI21_X1 U21779 ( .B1(n18716), .B2(n18715), .A(n18714), .ZN(n18718) );
  OAI211_X1 U21780 ( .C1(n18719), .C2(n18718), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18717), .ZN(n18721) );
  AOI21_X1 U21781 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18721), .A(n18720), 
        .ZN(n18723) );
  NAND2_X1 U21782 ( .A1(n18724), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18722) );
  OAI21_X1 U21783 ( .B1(n18724), .B2(n18723), .A(n18722), .ZN(P3_U3296) );
  INV_X1 U21784 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n20867) );
  INV_X1 U21785 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18726) );
  AOI22_X1 U21786 ( .A1(n18658), .A2(n20867), .B1(n18726), .B2(n18725), .ZN(
        P3_U3297) );
  OAI21_X1 U21787 ( .B1(n18730), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n18729), 
        .ZN(n18727) );
  OAI21_X1 U21788 ( .B1(n18729), .B2(n18728), .A(n18727), .ZN(P3_U3298) );
  NOR3_X1 U21789 ( .A1(n18731), .A2(n18730), .A3(P3_MEMORYFETCH_REG_SCAN_IN), 
        .ZN(n18733) );
  NOR2_X1 U21790 ( .A1(n18733), .A2(n18732), .ZN(P3_U3299) );
  INV_X1 U21791 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18735) );
  NAND2_X1 U21792 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19774), .ZN(n19767) );
  NAND2_X1 U21793 ( .A1(n19763), .A2(n18734), .ZN(n19764) );
  OAI21_X1 U21794 ( .B1(n19763), .B2(n19767), .A(n19764), .ZN(n19831) );
  OAI21_X1 U21795 ( .B1(n19763), .B2(n18735), .A(n19758), .ZN(P2_U2815) );
  INV_X1 U21796 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18738) );
  OAI22_X1 U21797 ( .A1(n19878), .A2(n18738), .B1(n18737), .B2(n18736), .ZN(
        P2_U2816) );
  AOI21_X1 U21798 ( .B1(n19763), .B2(n19774), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18739) );
  AOI22_X1 U21799 ( .A1(n19813), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18739), 
        .B2(n19897), .ZN(P2_U2817) );
  INV_X1 U21800 ( .A(n19768), .ZN(n18740) );
  OAI21_X1 U21801 ( .B1(n18740), .B2(BS16), .A(n19831), .ZN(n19829) );
  OAI21_X1 U21802 ( .B1(n19831), .B2(n19630), .A(n19829), .ZN(P2_U2818) );
  INV_X1 U21803 ( .A(P2_DATAWIDTH_REG_12__SCAN_IN), .ZN(n20836) );
  INV_X1 U21804 ( .A(P2_DATAWIDTH_REG_29__SCAN_IN), .ZN(n20859) );
  NAND2_X1 U21805 ( .A1(n20836), .A2(n20859), .ZN(n20800) );
  INV_X1 U21806 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20822) );
  INV_X1 U21807 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19830) );
  INV_X1 U21808 ( .A(P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20845) );
  INV_X1 U21809 ( .A(P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(n20878) );
  OAI211_X1 U21810 ( .C1(n20822), .C2(n19830), .A(n20845), .B(n20878), .ZN(
        n18741) );
  NOR4_X1 U21811 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(n20800), .A4(n18741), .ZN(n18749)
         );
  NOR4_X1 U21812 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18748) );
  NOR4_X1 U21813 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18747) );
  NOR4_X1 U21814 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_19__SCAN_IN), .A3(P2_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_21__SCAN_IN), .ZN(n18745) );
  NOR4_X1 U21815 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_14__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_16__SCAN_IN), .ZN(n18744) );
  NOR4_X1 U21816 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18743) );
  NOR4_X1 U21817 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_23__SCAN_IN), .A3(P2_DATAWIDTH_REG_24__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_25__SCAN_IN), .ZN(n18742) );
  AND4_X1 U21818 ( .A1(n18745), .A2(n18744), .A3(n18743), .A4(n18742), .ZN(
        n18746) );
  NAND4_X1 U21819 ( .A1(n18749), .A2(n18748), .A3(n18747), .A4(n18746), .ZN(
        n18755) );
  NOR2_X1 U21820 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18755), .ZN(n18750) );
  INV_X1 U21821 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19827) );
  AOI22_X1 U21822 ( .A1(n18750), .A2(n20815), .B1(n18755), .B2(n19827), .ZN(
        P2_U2820) );
  NAND3_X1 U21823 ( .A1(n20815), .A2(n20822), .A3(n19830), .ZN(n18754) );
  INV_X1 U21824 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19825) );
  AOI22_X1 U21825 ( .A1(n18750), .A2(n18754), .B1(n18755), .B2(n19825), .ZN(
        P2_U2821) );
  NAND2_X1 U21826 ( .A1(n18750), .A2(n19830), .ZN(n18753) );
  INV_X1 U21827 ( .A(n18755), .ZN(n18756) );
  OAI21_X1 U21828 ( .B1(n20815), .B2(n19776), .A(n18756), .ZN(n18751) );
  OAI21_X1 U21829 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18756), .A(n18751), 
        .ZN(n18752) );
  OAI221_X1 U21830 ( .B1(n18753), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18753), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18752), .ZN(P2_U2822) );
  INV_X1 U21831 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19823) );
  OAI221_X1 U21832 ( .B1(n18756), .B2(n19823), .C1(n18755), .C2(n18754), .A(
        n18753), .ZN(P2_U2823) );
  AOI21_X1 U21833 ( .B1(n18761), .B2(n18758), .A(n18757), .ZN(n18759) );
  AOI21_X1 U21834 ( .B1(n18906), .B2(n18760), .A(n18759), .ZN(n18767) );
  AOI22_X1 U21835 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18950), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18936), .ZN(n18766) );
  AOI22_X1 U21836 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n18935), .B1(n18761), 
        .B2(n18949), .ZN(n18765) );
  AOI22_X1 U21837 ( .A1(n18763), .A2(n18937), .B1(n18762), .B2(n18944), .ZN(
        n18764) );
  NAND4_X1 U21838 ( .A1(n18767), .A2(n18766), .A3(n18765), .A4(n18764), .ZN(
        P2_U2835) );
  NOR2_X1 U21839 ( .A1(n18896), .A2(n18768), .ZN(n18769) );
  XNOR2_X1 U21840 ( .A(n18770), .B(n18769), .ZN(n18779) );
  OAI21_X1 U21841 ( .B1(n19796), .B2(n18873), .A(n13051), .ZN(n18774) );
  INV_X1 U21842 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18771) );
  OAI22_X1 U21843 ( .A1(n18772), .A2(n18941), .B1(n18771), .B2(n18892), .ZN(
        n18773) );
  AOI211_X1 U21844 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n18935), .A(n18774), .B(
        n18773), .ZN(n18778) );
  OAI22_X1 U21845 ( .A1(n20788), .A2(n18925), .B1(n18775), .B2(n18911), .ZN(
        n18776) );
  INV_X1 U21846 ( .A(n18776), .ZN(n18777) );
  OAI211_X1 U21847 ( .C1(n18934), .C2(n18779), .A(n18778), .B(n18777), .ZN(
        P2_U2836) );
  INV_X1 U21848 ( .A(n18780), .ZN(n18782) );
  AOI22_X1 U21849 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18950), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n18935), .ZN(n18781) );
  OAI21_X1 U21850 ( .B1(n18782), .B2(n18941), .A(n18781), .ZN(n18783) );
  AOI211_X1 U21851 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n18936), .A(n18784), 
        .B(n18783), .ZN(n18791) );
  NAND2_X1 U21852 ( .A1(n18915), .A2(n18785), .ZN(n18787) );
  XNOR2_X1 U21853 ( .A(n18787), .B(n18786), .ZN(n18788) );
  AOI22_X1 U21854 ( .A1(n18789), .A2(n18937), .B1(n18901), .B2(n18788), .ZN(
        n18790) );
  OAI211_X1 U21855 ( .C1(n18792), .C2(n18911), .A(n18791), .B(n18790), .ZN(
        P2_U2837) );
  NOR2_X1 U21856 ( .A1(n18896), .A2(n18793), .ZN(n18795) );
  XOR2_X1 U21857 ( .A(n18795), .B(n18794), .Z(n18805) );
  OAI21_X1 U21858 ( .B1(n20892), .B2(n18873), .A(n13051), .ZN(n18799) );
  INV_X1 U21859 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18796) );
  OAI22_X1 U21860 ( .A1(n18797), .A2(n18941), .B1(n18796), .B2(n18892), .ZN(
        n18798) );
  AOI211_X1 U21861 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n18935), .A(n18799), .B(
        n18798), .ZN(n18804) );
  OAI22_X1 U21862 ( .A1(n18801), .A2(n18925), .B1(n18800), .B2(n18911), .ZN(
        n18802) );
  INV_X1 U21863 ( .A(n18802), .ZN(n18803) );
  OAI211_X1 U21864 ( .C1(n18934), .C2(n18805), .A(n18804), .B(n18803), .ZN(
        P2_U2838) );
  NAND2_X1 U21865 ( .A1(n18915), .A2(n18806), .ZN(n18807) );
  XNOR2_X1 U21866 ( .A(n18808), .B(n18807), .ZN(n18817) );
  INV_X1 U21867 ( .A(n18809), .ZN(n18811) );
  AOI22_X1 U21868 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18950), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n18935), .ZN(n18810) );
  OAI21_X1 U21869 ( .B1(n18811), .B2(n18941), .A(n18810), .ZN(n18812) );
  AOI211_X1 U21870 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n18936), .A(n19090), 
        .B(n18812), .ZN(n18816) );
  INV_X1 U21871 ( .A(n18813), .ZN(n18995) );
  OAI22_X1 U21872 ( .A1(n18962), .A2(n18911), .B1(n18995), .B2(n18925), .ZN(
        n18814) );
  INV_X1 U21873 ( .A(n18814), .ZN(n18815) );
  OAI211_X1 U21874 ( .C1(n18934), .C2(n18817), .A(n18816), .B(n18815), .ZN(
        P2_U2841) );
  OAI22_X1 U21875 ( .A1(n18819), .A2(n18941), .B1(n18818), .B2(n18892), .ZN(
        n18820) );
  AOI211_X1 U21876 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n18936), .A(n19090), 
        .B(n18820), .ZN(n18830) );
  NOR2_X1 U21877 ( .A1(n18896), .A2(n18821), .ZN(n18822) );
  XOR2_X1 U21878 ( .A(n18823), .B(n18822), .Z(n18828) );
  INV_X1 U21879 ( .A(n18824), .ZN(n18826) );
  OAI22_X1 U21880 ( .A1(n18826), .A2(n18911), .B1(n18825), .B2(n18925), .ZN(
        n18827) );
  AOI21_X1 U21881 ( .B1(n18828), .B2(n18901), .A(n18827), .ZN(n18829) );
  OAI211_X1 U21882 ( .C1(n18909), .C2(n11774), .A(n18830), .B(n18829), .ZN(
        P2_U2842) );
  OAI22_X1 U21883 ( .A1(n18831), .A2(n18892), .B1(n11973), .B2(n18873), .ZN(
        n18832) );
  NOR2_X1 U21884 ( .A1(n18832), .A2(n19090), .ZN(n18833) );
  OAI21_X1 U21885 ( .B1(n18834), .B2(n18925), .A(n18833), .ZN(n18835) );
  INV_X1 U21886 ( .A(n18835), .ZN(n18846) );
  AOI22_X1 U21887 ( .A1(n18836), .A2(n18906), .B1(P2_EBX_REG_11__SCAN_IN), 
        .B2(n18935), .ZN(n18845) );
  AOI22_X1 U21888 ( .A1(n18838), .A2(n18944), .B1(n18837), .B2(n18949), .ZN(
        n18844) );
  INV_X1 U21889 ( .A(n18839), .ZN(n18946) );
  OAI211_X1 U21890 ( .C1(n18842), .C2(n18841), .A(n18946), .B(n18840), .ZN(
        n18843) );
  NAND4_X1 U21891 ( .A1(n18846), .A2(n18845), .A3(n18844), .A4(n18843), .ZN(
        P2_U2844) );
  NOR2_X1 U21892 ( .A1(n18896), .A2(n18847), .ZN(n18849) );
  XNOR2_X1 U21893 ( .A(n18849), .B(n18848), .ZN(n18856) );
  AOI22_X1 U21894 ( .A1(n18850), .A2(n18906), .B1(n18950), .B2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18851) );
  OAI211_X1 U21895 ( .C1(n11967), .C2(n18873), .A(n18851), .B(n18871), .ZN(
        n18854) );
  OAI22_X1 U21896 ( .A1(n19003), .A2(n18925), .B1(n18911), .B2(n18852), .ZN(
        n18853) );
  AOI211_X1 U21897 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n18935), .A(n18854), .B(
        n18853), .ZN(n18855) );
  OAI21_X1 U21898 ( .B1(n18934), .B2(n18856), .A(n18855), .ZN(P2_U2846) );
  AOI22_X1 U21899 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(n18935), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18950), .ZN(n18857) );
  OAI21_X1 U21900 ( .B1(n18858), .B2(n18941), .A(n18857), .ZN(n18859) );
  AOI211_X1 U21901 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n18936), .A(n19090), .B(
        n18859), .ZN(n18866) );
  NAND2_X1 U21902 ( .A1(n14711), .A2(n18860), .ZN(n18861) );
  XNOR2_X1 U21903 ( .A(n18862), .B(n18861), .ZN(n18864) );
  AOI22_X1 U21904 ( .A1(n18864), .A2(n18901), .B1(n18937), .B2(n18863), .ZN(
        n18865) );
  OAI211_X1 U21905 ( .C1(n18911), .C2(n18981), .A(n18866), .B(n18865), .ZN(
        P2_U2847) );
  NOR2_X1 U21906 ( .A1(n18896), .A2(n18867), .ZN(n18868) );
  XOR2_X1 U21907 ( .A(n18869), .B(n18868), .Z(n18879) );
  AOI22_X1 U21908 ( .A1(n18870), .A2(n18906), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n18935), .ZN(n18872) );
  OAI211_X1 U21909 ( .C1(n15210), .C2(n18873), .A(n18872), .B(n18871), .ZN(
        n18877) );
  OAI22_X1 U21910 ( .A1(n18875), .A2(n18925), .B1(n18874), .B2(n18911), .ZN(
        n18876) );
  AOI211_X1 U21911 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n18950), .A(
        n18877), .B(n18876), .ZN(n18878) );
  OAI21_X1 U21912 ( .B1(n18934), .B2(n18879), .A(n18878), .ZN(P2_U2848) );
  OAI22_X1 U21913 ( .A1(n18880), .A2(n18941), .B1(n15217), .B2(n18892), .ZN(
        n18881) );
  AOI211_X1 U21914 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n18936), .A(n19090), .B(
        n18881), .ZN(n18890) );
  NAND2_X1 U21915 ( .A1(n14711), .A2(n18882), .ZN(n18883) );
  XNOR2_X1 U21916 ( .A(n18884), .B(n18883), .ZN(n18888) );
  OAI22_X1 U21917 ( .A1(n18886), .A2(n18925), .B1(n18911), .B2(n18885), .ZN(
        n18887) );
  AOI21_X1 U21918 ( .B1(n18901), .B2(n18888), .A(n18887), .ZN(n18889) );
  OAI211_X1 U21919 ( .C1(n18909), .C2(n18891), .A(n18890), .B(n18889), .ZN(
        P2_U2849) );
  OAI22_X1 U21920 ( .A1(n18893), .A2(n18941), .B1(n9898), .B2(n18892), .ZN(
        n18894) );
  AOI211_X1 U21921 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18936), .A(n19090), .B(
        n18894), .ZN(n18904) );
  NOR2_X1 U21922 ( .A1(n18896), .A2(n18895), .ZN(n18897) );
  XNOR2_X1 U21923 ( .A(n18898), .B(n18897), .ZN(n18902) );
  OAI22_X1 U21924 ( .A1(n19011), .A2(n18925), .B1(n18911), .B2(n18899), .ZN(
        n18900) );
  AOI21_X1 U21925 ( .B1(n18902), .B2(n18901), .A(n18900), .ZN(n18903) );
  OAI211_X1 U21926 ( .C1(n18909), .C2(n18905), .A(n18904), .B(n18903), .ZN(
        P2_U2850) );
  AOI22_X1 U21927 ( .A1(n18907), .A2(n18906), .B1(n18950), .B2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18921) );
  OAI22_X1 U21928 ( .A1(n18909), .A2(n18987), .B1(n18925), .B2(n18908), .ZN(
        n18910) );
  AOI211_X1 U21929 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n18936), .A(n19090), .B(
        n18910), .ZN(n18920) );
  OAI22_X1 U21930 ( .A1(n19006), .A2(n18912), .B1(n18911), .B2(n18982), .ZN(
        n18913) );
  INV_X1 U21931 ( .A(n18913), .ZN(n18919) );
  AND2_X1 U21932 ( .A1(n18915), .A2(n18914), .ZN(n18917) );
  AOI21_X1 U21933 ( .B1(n19088), .B2(n18917), .A(n18934), .ZN(n18916) );
  OAI21_X1 U21934 ( .B1(n19088), .B2(n18917), .A(n18916), .ZN(n18918) );
  NAND4_X1 U21935 ( .A1(n18921), .A2(n18920), .A3(n18919), .A4(n18918), .ZN(
        P2_U2851) );
  AOI22_X1 U21936 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18950), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n18936), .ZN(n18923) );
  NAND2_X1 U21937 ( .A1(n18935), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n18922) );
  OAI211_X1 U21938 ( .C1(n18941), .C2(n18924), .A(n18923), .B(n18922), .ZN(
        n18928) );
  NOR2_X1 U21939 ( .A1(n18926), .A2(n18925), .ZN(n18927) );
  AOI211_X1 U21940 ( .C1(n18944), .C2(n18929), .A(n18928), .B(n18927), .ZN(
        n18932) );
  AOI22_X1 U21941 ( .A1(n18949), .A2(n18930), .B1(n18948), .B2(n19851), .ZN(
        n18931) );
  OAI211_X1 U21942 ( .C1(n18934), .C2(n18933), .A(n18932), .B(n18931), .ZN(
        P2_U2854) );
  AOI22_X1 U21943 ( .A1(n18936), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n18935), 
        .B2(P2_EBX_REG_0__SCAN_IN), .ZN(n18940) );
  NAND2_X1 U21944 ( .A1(n18938), .A2(n18937), .ZN(n18939) );
  OAI211_X1 U21945 ( .C1(n18942), .C2(n18941), .A(n18940), .B(n18939), .ZN(
        n18943) );
  AOI21_X1 U21946 ( .B1(n18945), .B2(n18944), .A(n18943), .ZN(n18953) );
  AOI22_X1 U21947 ( .A1(n19413), .A2(n18948), .B1(n18947), .B2(n18946), .ZN(
        n18952) );
  OAI21_X1 U21948 ( .B1(n18950), .B2(n18949), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18951) );
  NAND3_X1 U21949 ( .A1(n18953), .A2(n18952), .A3(n18951), .ZN(P2_U2855) );
  AOI22_X1 U21950 ( .A1(n18955), .A2(n18954), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n18983), .ZN(n18956) );
  OAI21_X1 U21951 ( .B1(n18983), .B2(n18957), .A(n18956), .ZN(P2_U2871) );
  AOI21_X1 U21952 ( .B1(n13671), .B2(n18958), .A(n18984), .ZN(n18960) );
  AOI22_X1 U21953 ( .A1(n18960), .A2(n18959), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n18983), .ZN(n18961) );
  OAI21_X1 U21954 ( .B1(n18962), .B2(n18983), .A(n18961), .ZN(P2_U2873) );
  AOI21_X1 U21955 ( .B1(n13511), .B2(n18964), .A(n18963), .ZN(n18965) );
  NOR3_X1 U21956 ( .A1(n18965), .A2(n13512), .A3(n18984), .ZN(n18966) );
  AOI21_X1 U21957 ( .B1(P2_EBX_REG_12__SCAN_IN), .B2(n18983), .A(n18966), .ZN(
        n18967) );
  OAI21_X1 U21958 ( .B1(n18968), .B2(n18983), .A(n18967), .ZN(P2_U2875) );
  AOI21_X1 U21959 ( .B1(n18977), .B2(n18970), .A(n18969), .ZN(n18971) );
  OR3_X1 U21960 ( .A1(n18971), .A2(n13511), .A3(n18984), .ZN(n18972) );
  OAI21_X1 U21961 ( .B1(n18973), .B2(n18983), .A(n18972), .ZN(n18974) );
  INV_X1 U21962 ( .A(n18974), .ZN(n18975) );
  OAI21_X1 U21963 ( .B1(n18988), .B2(n9816), .A(n18975), .ZN(P2_U2877) );
  AOI211_X1 U21964 ( .C1(n18978), .C2(n18976), .A(n18984), .B(n18977), .ZN(
        n18979) );
  AOI21_X1 U21965 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n18983), .A(n18979), .ZN(
        n18980) );
  OAI21_X1 U21966 ( .B1(n18981), .B2(n18983), .A(n18980), .ZN(P2_U2879) );
  OAI22_X1 U21967 ( .A1(n19006), .A2(n18984), .B1(n18983), .B2(n18982), .ZN(
        n18985) );
  INV_X1 U21968 ( .A(n18985), .ZN(n18986) );
  OAI21_X1 U21969 ( .B1(n18988), .B2(n18987), .A(n18986), .ZN(P2_U2883) );
  AOI22_X1 U21970 ( .A1(n18990), .A2(n18989), .B1(n20784), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n18992) );
  AOI22_X1 U21971 ( .A1(n20783), .A2(BUF1_REG_31__SCAN_IN), .B1(n20780), .B2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n18991) );
  NAND2_X1 U21972 ( .A1(n18992), .A2(n18991), .ZN(P2_U2888) );
  AOI22_X1 U21973 ( .A1(n19005), .A2(n18993), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n20780), .ZN(n18994) );
  OAI21_X1 U21974 ( .B1(n19012), .B2(n18995), .A(n18994), .ZN(P2_U2905) );
  AOI22_X1 U21975 ( .A1(n19005), .A2(n19062), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n20780), .ZN(n18996) );
  OAI21_X1 U21976 ( .B1(n19012), .B2(n18997), .A(n18996), .ZN(P2_U2907) );
  AOI22_X1 U21977 ( .A1(n19005), .A2(n18998), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n20780), .ZN(n18999) );
  OAI21_X1 U21978 ( .B1(n19012), .B2(n19000), .A(n18999), .ZN(P2_U2909) );
  AOI22_X1 U21979 ( .A1(n19005), .A2(n19001), .B1(P2_EAX_REG_9__SCAN_IN), .B2(
        n20780), .ZN(n19002) );
  OAI21_X1 U21980 ( .B1(n19012), .B2(n19003), .A(n19002), .ZN(P2_U2910) );
  AOI22_X1 U21981 ( .A1(n19005), .A2(n19004), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n20780), .ZN(n19010) );
  INV_X1 U21982 ( .A(n19006), .ZN(n19007) );
  NAND3_X1 U21983 ( .A1(n19008), .A2(n19007), .A3(n20791), .ZN(n19009) );
  OAI211_X1 U21984 ( .C1(n19012), .C2(n19011), .A(n19010), .B(n19009), .ZN(
        P2_U2914) );
  NOR2_X1 U21985 ( .A1(n19017), .A2(n19013), .ZN(P2_U2920) );
  INV_X1 U21986 ( .A(n19014), .ZN(n19015) );
  AOI22_X1 U21987 ( .A1(n19015), .A2(P2_EAX_REG_28__SCAN_IN), .B1(
        P2_UWORD_REG_12__SCAN_IN), .B2(n19045), .ZN(n19016) );
  OAI21_X1 U21988 ( .B1(n20929), .B2(n19017), .A(n19016), .ZN(P2_U2923) );
  AOI22_X1 U21989 ( .A1(n19045), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19018) );
  OAI21_X1 U21990 ( .B1(n19019), .B2(n19049), .A(n19018), .ZN(P2_U2936) );
  AOI22_X1 U21991 ( .A1(n19045), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19020) );
  OAI21_X1 U21992 ( .B1(n19021), .B2(n19049), .A(n19020), .ZN(P2_U2937) );
  AOI22_X1 U21993 ( .A1(n19045), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19022) );
  OAI21_X1 U21994 ( .B1(n19023), .B2(n19049), .A(n19022), .ZN(P2_U2938) );
  INV_X1 U21995 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19025) );
  AOI22_X1 U21996 ( .A1(n19045), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19024) );
  OAI21_X1 U21997 ( .B1(n19025), .B2(n19049), .A(n19024), .ZN(P2_U2939) );
  AOI22_X1 U21998 ( .A1(n19045), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19026) );
  OAI21_X1 U21999 ( .B1(n19027), .B2(n19049), .A(n19026), .ZN(P2_U2940) );
  AOI22_X1 U22000 ( .A1(n19045), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19028) );
  OAI21_X1 U22001 ( .B1(n19029), .B2(n19049), .A(n19028), .ZN(P2_U2941) );
  AOI22_X1 U22002 ( .A1(n19045), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19030) );
  OAI21_X1 U22003 ( .B1(n19031), .B2(n19049), .A(n19030), .ZN(P2_U2942) );
  AOI22_X1 U22004 ( .A1(n19045), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19032) );
  OAI21_X1 U22005 ( .B1(n19033), .B2(n19049), .A(n19032), .ZN(P2_U2943) );
  AOI22_X1 U22006 ( .A1(n19045), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19034) );
  OAI21_X1 U22007 ( .B1(n19035), .B2(n19049), .A(n19034), .ZN(P2_U2944) );
  AOI22_X1 U22008 ( .A1(n19045), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19036) );
  OAI21_X1 U22009 ( .B1(n19037), .B2(n19049), .A(n19036), .ZN(P2_U2945) );
  INV_X1 U22010 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19039) );
  AOI22_X1 U22011 ( .A1(n19045), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19038) );
  OAI21_X1 U22012 ( .B1(n19039), .B2(n19049), .A(n19038), .ZN(P2_U2946) );
  AOI22_X1 U22013 ( .A1(n19045), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19040) );
  OAI21_X1 U22014 ( .B1(n13417), .B2(n19049), .A(n19040), .ZN(P2_U2947) );
  INV_X1 U22015 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19042) );
  AOI22_X1 U22016 ( .A1(n19045), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19041) );
  OAI21_X1 U22017 ( .B1(n19042), .B2(n19049), .A(n19041), .ZN(P2_U2948) );
  INV_X1 U22018 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19044) );
  AOI22_X1 U22019 ( .A1(n19045), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19043) );
  OAI21_X1 U22020 ( .B1(n19044), .B2(n19049), .A(n19043), .ZN(P2_U2949) );
  AOI22_X1 U22021 ( .A1(n19045), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19046) );
  OAI21_X1 U22022 ( .B1(n12937), .B2(n19049), .A(n19046), .ZN(P2_U2950) );
  INV_X1 U22023 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19050) );
  AOI22_X1 U22024 ( .A1(n19045), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19047), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19048) );
  OAI21_X1 U22025 ( .B1(n19050), .B2(n19049), .A(n19048), .ZN(P2_U2951) );
  AOI22_X1 U22026 ( .A1(n19061), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n19084), .ZN(n19051) );
  OAI21_X1 U22027 ( .B1(n19109), .B2(n19086), .A(n19051), .ZN(P2_U2952) );
  AOI22_X1 U22028 ( .A1(n19061), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19084), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n19052) );
  OAI21_X1 U22029 ( .B1(n19121), .B2(n19086), .A(n19052), .ZN(P2_U2953) );
  INV_X1 U22030 ( .A(n19126), .ZN(n19069) );
  AOI22_X1 U22031 ( .A1(n19061), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n19084), .ZN(n19053) );
  OAI21_X1 U22032 ( .B1(n19069), .B2(n19086), .A(n19053), .ZN(P2_U2954) );
  AOI22_X1 U22033 ( .A1(n19061), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19084), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n19054) );
  OAI21_X1 U22034 ( .B1(n19133), .B2(n19086), .A(n19054), .ZN(P2_U2955) );
  AOI22_X1 U22035 ( .A1(n19061), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n19084), .ZN(n19055) );
  OAI21_X1 U22036 ( .B1(n19139), .B2(n19086), .A(n19055), .ZN(P2_U2956) );
  AOI22_X1 U22037 ( .A1(n19061), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19084), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n19056) );
  OAI21_X1 U22038 ( .B1(n19145), .B2(n19086), .A(n19056), .ZN(P2_U2957) );
  AOI22_X1 U22039 ( .A1(n19061), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n19084), .ZN(n19057) );
  OAI21_X1 U22040 ( .B1(n19152), .B2(n19086), .A(n19057), .ZN(P2_U2958) );
  AOI22_X1 U22041 ( .A1(n19061), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19084), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n19058) );
  OAI21_X1 U22042 ( .B1(n19161), .B2(n19086), .A(n19058), .ZN(P2_U2959) );
  AOI22_X1 U22043 ( .A1(n19081), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n19084), .ZN(n19059) );
  OAI21_X1 U22044 ( .B1(n19076), .B2(n19086), .A(n19059), .ZN(P2_U2960) );
  AOI22_X1 U22045 ( .A1(n19081), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n19084), .ZN(n19060) );
  OAI21_X1 U22046 ( .B1(n19078), .B2(n19086), .A(n19060), .ZN(P2_U2963) );
  AOI22_X1 U22047 ( .A1(n19061), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n19084), .ZN(n19064) );
  NAND2_X1 U22048 ( .A1(n19063), .A2(n19062), .ZN(n19079) );
  NAND2_X1 U22049 ( .A1(n19064), .A2(n19079), .ZN(P2_U2964) );
  AOI22_X1 U22050 ( .A1(n19061), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19084), .ZN(n19065) );
  OAI21_X1 U22051 ( .B1(n19083), .B2(n19086), .A(n19065), .ZN(P2_U2965) );
  AOI22_X1 U22052 ( .A1(n19081), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19084), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n19066) );
  OAI21_X1 U22053 ( .B1(n19109), .B2(n19086), .A(n19066), .ZN(P2_U2967) );
  AOI22_X1 U22054 ( .A1(n19081), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19084), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n19067) );
  OAI21_X1 U22055 ( .B1(n19121), .B2(n19086), .A(n19067), .ZN(P2_U2968) );
  AOI22_X1 U22056 ( .A1(n19081), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19084), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n19068) );
  OAI21_X1 U22057 ( .B1(n19069), .B2(n19086), .A(n19068), .ZN(P2_U2969) );
  AOI22_X1 U22058 ( .A1(n19081), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19084), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n19070) );
  OAI21_X1 U22059 ( .B1(n19133), .B2(n19086), .A(n19070), .ZN(P2_U2970) );
  AOI22_X1 U22060 ( .A1(n19081), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n19084), .ZN(n19071) );
  OAI21_X1 U22061 ( .B1(n19139), .B2(n19086), .A(n19071), .ZN(P2_U2971) );
  AOI22_X1 U22062 ( .A1(n19081), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19084), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n19072) );
  OAI21_X1 U22063 ( .B1(n19145), .B2(n19086), .A(n19072), .ZN(P2_U2972) );
  AOI22_X1 U22064 ( .A1(n19081), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19084), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n19073) );
  OAI21_X1 U22065 ( .B1(n19152), .B2(n19086), .A(n19073), .ZN(P2_U2973) );
  AOI22_X1 U22066 ( .A1(n19081), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19084), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n19074) );
  OAI21_X1 U22067 ( .B1(n19161), .B2(n19086), .A(n19074), .ZN(P2_U2974) );
  AOI22_X1 U22068 ( .A1(n19081), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19084), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n19075) );
  OAI21_X1 U22069 ( .B1(n19076), .B2(n19086), .A(n19075), .ZN(P2_U2975) );
  AOI22_X1 U22070 ( .A1(n19081), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19084), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n19077) );
  OAI21_X1 U22071 ( .B1(n19078), .B2(n19086), .A(n19077), .ZN(P2_U2978) );
  AOI22_X1 U22072 ( .A1(n19081), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n19084), .ZN(n19080) );
  NAND2_X1 U22073 ( .A1(n19080), .A2(n19079), .ZN(P2_U2979) );
  AOI22_X1 U22074 ( .A1(n19081), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n19084), .ZN(n19082) );
  OAI21_X1 U22075 ( .B1(n19083), .B2(n19086), .A(n19082), .ZN(P2_U2980) );
  AOI22_X1 U22076 ( .A1(n19081), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19084), 
        .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n19085) );
  OAI21_X1 U22077 ( .B1(n19087), .B2(n19086), .A(n19085), .ZN(P2_U2982) );
  AOI22_X1 U22078 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19090), .B1(n19089), 
        .B2(n19088), .ZN(n19098) );
  AOI222_X1 U22079 ( .A1(n19096), .A2(n19095), .B1(n19094), .B2(n19093), .C1(
        n19092), .C2(n19091), .ZN(n19097) );
  OAI211_X1 U22080 ( .C1(n19100), .C2(n19099), .A(n19098), .B(n19097), .ZN(
        P2_U3010) );
  AOI22_X2 U22081 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19156), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19155), .ZN(n19700) );
  OAI22_X2 U22082 ( .A1(n14325), .A2(n19150), .B1(n19104), .B2(n19148), .ZN(
        n19697) );
  OR2_X1 U22083 ( .A1(n19158), .A2(n11895), .ZN(n19626) );
  NOR2_X1 U22084 ( .A1(n19555), .A2(n19212), .ZN(n19110) );
  INV_X1 U22085 ( .A(n19110), .ZN(n19159) );
  OAI22_X1 U22086 ( .A1(n19737), .A2(n19627), .B1(n19626), .B2(n19159), .ZN(
        n19105) );
  INV_X1 U22087 ( .A(n19105), .ZN(n19116) );
  INV_X1 U22088 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19491) );
  NOR3_X1 U22089 ( .A1(n19111), .A2(n19110), .A3(n19491), .ZN(n19108) );
  NOR2_X1 U22090 ( .A1(n19744), .A2(n19206), .ZN(n19106) );
  OAI21_X1 U22091 ( .B1(n19106), .B2(n19630), .A(n19837), .ZN(n19114) );
  AOI221_X1 U22092 ( .B1(n19883), .B2(n19114), .C1(n19883), .C2(n19739), .A(
        n19110), .ZN(n19107) );
  OR2_X1 U22093 ( .A1(n19452), .A2(n19109), .ZN(n19168) );
  INV_X1 U22094 ( .A(n19168), .ZN(n19689) );
  NOR2_X1 U22095 ( .A1(n19739), .A2(n19110), .ZN(n19113) );
  OAI21_X1 U22096 ( .B1(n19111), .B2(n19110), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19112) );
  AOI22_X1 U22097 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19163), .B1(
        n19689), .B2(n19162), .ZN(n19115) );
  OAI211_X1 U22098 ( .C1(n19700), .C2(n19189), .A(n19116), .B(n19115), .ZN(
        P2_U3048) );
  AOI22_X1 U22099 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19156), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19155), .ZN(n19706) );
  OAI22_X1 U22100 ( .A1(n19118), .A2(n19150), .B1(n19117), .B2(n19148), .ZN(
        n19703) );
  OR2_X1 U22101 ( .A1(n19158), .A2(n19119), .ZN(n19645) );
  OAI22_X1 U22102 ( .A1(n19737), .A2(n19646), .B1(n19159), .B2(n19645), .ZN(
        n19120) );
  INV_X1 U22103 ( .A(n19120), .ZN(n19123) );
  OR2_X1 U22104 ( .A1(n19452), .A2(n19121), .ZN(n19177) );
  INV_X1 U22105 ( .A(n19177), .ZN(n19702) );
  AOI22_X1 U22106 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19163), .B1(
        n19702), .B2(n19162), .ZN(n19122) );
  OAI211_X1 U22107 ( .C1(n19706), .C2(n19189), .A(n19123), .B(n19122), .ZN(
        P2_U3049) );
  AOI22_X2 U22108 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19156), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19155), .ZN(n19712) );
  OAI22_X1 U22109 ( .A1(n19124), .A2(n19150), .B1(n14960), .B2(n19148), .ZN(
        n19709) );
  OR2_X1 U22110 ( .A1(n19158), .A2(n11916), .ZN(n19650) );
  OAI22_X1 U22111 ( .A1(n19737), .A2(n19654), .B1(n19159), .B2(n19650), .ZN(
        n19125) );
  INV_X1 U22112 ( .A(n19125), .ZN(n19128) );
  AOI22_X1 U22113 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19163), .B1(
        n19708), .B2(n19162), .ZN(n19127) );
  OAI211_X1 U22114 ( .C1(n19712), .C2(n19189), .A(n19128), .B(n19127), .ZN(
        P2_U3050) );
  OAI22_X1 U22115 ( .A1(n19130), .A2(n19150), .B1(n19129), .B2(n19148), .ZN(
        n19715) );
  AOI22_X1 U22116 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19156), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19155), .ZN(n19718) );
  OR2_X1 U22117 ( .A1(n19158), .A2(n19131), .ZN(n19655) );
  OAI22_X1 U22118 ( .A1(n19737), .A2(n19718), .B1(n19655), .B2(n19159), .ZN(
        n19132) );
  INV_X1 U22119 ( .A(n19132), .ZN(n19135) );
  OR2_X1 U22120 ( .A1(n19452), .A2(n19133), .ZN(n19185) );
  INV_X1 U22121 ( .A(n19185), .ZN(n19714) );
  AOI22_X1 U22122 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19163), .B1(
        n19714), .B2(n19162), .ZN(n19134) );
  OAI211_X1 U22123 ( .C1(n19656), .C2(n19189), .A(n19135), .B(n19134), .ZN(
        P2_U3051) );
  OAI22_X1 U22124 ( .A1(n19137), .A2(n19150), .B1(n19136), .B2(n19148), .ZN(
        n19609) );
  AOI22_X1 U22125 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19156), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19155), .ZN(n19664) );
  OR2_X1 U22126 ( .A1(n19158), .A2(n11423), .ZN(n19660) );
  OAI22_X1 U22127 ( .A1(n19737), .A2(n19664), .B1(n19660), .B2(n19159), .ZN(
        n19138) );
  INV_X1 U22128 ( .A(n19138), .ZN(n19141) );
  OR2_X1 U22129 ( .A1(n19452), .A2(n19139), .ZN(n19190) );
  INV_X1 U22130 ( .A(n19190), .ZN(n19720) );
  AOI22_X1 U22131 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19163), .B1(
        n19720), .B2(n19162), .ZN(n19140) );
  OAI211_X1 U22132 ( .C1(n19724), .C2(n19189), .A(n19141), .B(n19140), .ZN(
        P2_U3052) );
  OAI22_X1 U22133 ( .A1(n19143), .A2(n19150), .B1(n19142), .B2(n19148), .ZN(
        n19727) );
  INV_X1 U22134 ( .A(n19727), .ZN(n19669) );
  OR2_X1 U22135 ( .A1(n19158), .A2(n12321), .ZN(n19665) );
  OAI22_X1 U22136 ( .A1(n19737), .A2(n19730), .B1(n19665), .B2(n19159), .ZN(
        n19144) );
  INV_X1 U22137 ( .A(n19144), .ZN(n19147) );
  OR2_X1 U22138 ( .A1(n19452), .A2(n19145), .ZN(n19194) );
  INV_X1 U22139 ( .A(n19194), .ZN(n19726) );
  AOI22_X1 U22140 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19163), .B1(
        n19726), .B2(n19162), .ZN(n19146) );
  OAI211_X1 U22141 ( .C1(n19669), .C2(n19189), .A(n19147), .B(n19146), .ZN(
        P2_U3053) );
  AOI22_X2 U22142 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19156), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19155), .ZN(n19738) );
  OAI22_X1 U22143 ( .A1(n14072), .A2(n19150), .B1(n19149), .B2(n19148), .ZN(
        n19733) );
  INV_X1 U22144 ( .A(n19733), .ZN(n19674) );
  OR2_X1 U22145 ( .A1(n19158), .A2(n12798), .ZN(n19670) );
  OAI22_X1 U22146 ( .A1(n19737), .A2(n19674), .B1(n19670), .B2(n19159), .ZN(
        n19151) );
  INV_X1 U22147 ( .A(n19151), .ZN(n19154) );
  OR2_X1 U22148 ( .A1(n19452), .A2(n19152), .ZN(n19198) );
  INV_X1 U22149 ( .A(n19198), .ZN(n19732) );
  AOI22_X1 U22150 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19163), .B1(
        n19732), .B2(n19162), .ZN(n19153) );
  OAI211_X1 U22151 ( .C1(n19738), .C2(n19189), .A(n19154), .B(n19153), .ZN(
        P2_U3054) );
  AOI22_X2 U22152 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19156), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19155), .ZN(n19683) );
  AOI22_X1 U22153 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19156), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19155), .ZN(n19749) );
  OR2_X1 U22154 ( .A1(n19158), .A2(n19157), .ZN(n19676) );
  OAI22_X1 U22155 ( .A1(n19737), .A2(n19749), .B1(n19159), .B2(n19676), .ZN(
        n19160) );
  INV_X1 U22156 ( .A(n19160), .ZN(n19165) );
  OR2_X1 U22157 ( .A1(n19452), .A2(n19161), .ZN(n19203) );
  INV_X1 U22158 ( .A(n19203), .ZN(n19741) );
  AOI22_X1 U22159 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19163), .B1(
        n19741), .B2(n19162), .ZN(n19164) );
  OAI211_X1 U22160 ( .C1(n19683), .C2(n19189), .A(n19165), .B(n19164), .ZN(
        P2_U3055) );
  NAND2_X1 U22161 ( .A1(n19414), .A2(n19383), .ZN(n19210) );
  OR2_X1 U22162 ( .A1(n19212), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19170) );
  NOR2_X1 U22163 ( .A1(n19865), .A2(n19170), .ZN(n19174) );
  NOR2_X1 U22164 ( .A1(n19491), .A2(n19174), .ZN(n19166) );
  NAND2_X1 U22165 ( .A1(n11665), .A2(n19166), .ZN(n19171) );
  AOI21_X1 U22166 ( .B1(n19170), .B2(n19491), .A(n19593), .ZN(n19167) );
  NAND2_X1 U22167 ( .A1(n19171), .A2(n19167), .ZN(n19204) );
  INV_X1 U22168 ( .A(n19174), .ZN(n19202) );
  OAI22_X1 U22169 ( .A1(n19204), .A2(n19168), .B1(n19626), .B2(n19202), .ZN(
        n19169) );
  INV_X1 U22170 ( .A(n19169), .ZN(n19176) );
  INV_X1 U22171 ( .A(n19414), .ZN(n19462) );
  NAND2_X1 U22172 ( .A1(n19450), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19388) );
  OAI21_X1 U22173 ( .B1(n19462), .B2(n19388), .A(n19170), .ZN(n19172) );
  AND2_X1 U22174 ( .A1(n19172), .A2(n19171), .ZN(n19173) );
  OAI211_X1 U22175 ( .C1(n19174), .C2(n19883), .A(n19173), .B(n19695), .ZN(
        n19207) );
  AOI22_X1 U22176 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19207), .B1(
        n19206), .B2(n19697), .ZN(n19175) );
  OAI211_X1 U22177 ( .C1(n19700), .C2(n19210), .A(n19176), .B(n19175), .ZN(
        P2_U3056) );
  OAI22_X1 U22178 ( .A1(n19204), .A2(n19177), .B1(n19645), .B2(n19202), .ZN(
        n19178) );
  INV_X1 U22179 ( .A(n19178), .ZN(n19180) );
  INV_X1 U22180 ( .A(n19706), .ZN(n19601) );
  AOI22_X1 U22181 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19207), .B1(
        n19239), .B2(n19601), .ZN(n19179) );
  OAI211_X1 U22182 ( .C1(n19646), .C2(n19189), .A(n19180), .B(n19179), .ZN(
        P2_U3057) );
  INV_X1 U22183 ( .A(n19708), .ZN(n19181) );
  OAI22_X1 U22184 ( .A1(n19204), .A2(n19181), .B1(n19650), .B2(n19202), .ZN(
        n19182) );
  INV_X1 U22185 ( .A(n19182), .ZN(n19184) );
  INV_X1 U22186 ( .A(n19712), .ZN(n19535) );
  AOI22_X1 U22187 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19207), .B1(
        n19239), .B2(n19535), .ZN(n19183) );
  OAI211_X1 U22188 ( .C1(n19654), .C2(n19189), .A(n19184), .B(n19183), .ZN(
        P2_U3058) );
  OAI22_X1 U22189 ( .A1(n19204), .A2(n19185), .B1(n19655), .B2(n19202), .ZN(
        n19186) );
  INV_X1 U22190 ( .A(n19186), .ZN(n19188) );
  AOI22_X1 U22191 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19207), .B1(
        n19239), .B2(n19715), .ZN(n19187) );
  OAI211_X1 U22192 ( .C1(n19718), .C2(n19189), .A(n19188), .B(n19187), .ZN(
        P2_U3059) );
  OAI22_X1 U22193 ( .A1(n19204), .A2(n19190), .B1(n19660), .B2(n19202), .ZN(
        n19191) );
  INV_X1 U22194 ( .A(n19191), .ZN(n19193) );
  INV_X1 U22195 ( .A(n19664), .ZN(n19721) );
  AOI22_X1 U22196 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19207), .B1(
        n19206), .B2(n19721), .ZN(n19192) );
  OAI211_X1 U22197 ( .C1(n19724), .C2(n19210), .A(n19193), .B(n19192), .ZN(
        P2_U3060) );
  OAI22_X1 U22198 ( .A1(n19204), .A2(n19194), .B1(n19665), .B2(n19202), .ZN(
        n19195) );
  INV_X1 U22199 ( .A(n19195), .ZN(n19197) );
  INV_X1 U22200 ( .A(n19730), .ZN(n19577) );
  AOI22_X1 U22201 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19207), .B1(
        n19206), .B2(n19577), .ZN(n19196) );
  OAI211_X1 U22202 ( .C1(n19669), .C2(n19210), .A(n19197), .B(n19196), .ZN(
        P2_U3061) );
  OAI22_X1 U22203 ( .A1(n19204), .A2(n19198), .B1(n19670), .B2(n19202), .ZN(
        n19199) );
  INV_X1 U22204 ( .A(n19199), .ZN(n19201) );
  AOI22_X1 U22205 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19207), .B1(
        n19206), .B2(n19733), .ZN(n19200) );
  OAI211_X1 U22206 ( .C1(n19738), .C2(n19210), .A(n19201), .B(n19200), .ZN(
        P2_U3062) );
  OAI22_X1 U22207 ( .A1(n19204), .A2(n19203), .B1(n19676), .B2(n19202), .ZN(
        n19205) );
  INV_X1 U22208 ( .A(n19205), .ZN(n19209) );
  INV_X1 U22209 ( .A(n19749), .ZN(n19620) );
  AOI22_X1 U22210 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19207), .B1(
        n19206), .B2(n19620), .ZN(n19208) );
  OAI211_X1 U22211 ( .C1(n19683), .C2(n19210), .A(n19209), .B(n19208), .ZN(
        P2_U3063) );
  INV_X1 U22212 ( .A(n19211), .ZN(n19216) );
  NOR2_X1 U22213 ( .A1(n19857), .A2(n19212), .ZN(n19246) );
  NAND2_X1 U22214 ( .A1(n19246), .A2(n19865), .ZN(n19215) );
  AND2_X1 U22215 ( .A1(n19216), .A2(n19215), .ZN(n19214) );
  INV_X1 U22216 ( .A(n19489), .ZN(n19213) );
  INV_X1 U22217 ( .A(n19212), .ZN(n19243) );
  NAND2_X1 U22218 ( .A1(n19213), .A2(n19243), .ZN(n19218) );
  INV_X1 U22219 ( .A(n19626), .ZN(n19688) );
  INV_X1 U22220 ( .A(n19215), .ZN(n19237) );
  AOI22_X1 U22221 ( .A1(n19238), .A2(n19689), .B1(n19688), .B2(n19237), .ZN(
        n19224) );
  OAI21_X1 U22222 ( .B1(n19216), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19215), 
        .ZN(n19221) );
  INV_X1 U22223 ( .A(n19274), .ZN(n19217) );
  NOR2_X1 U22224 ( .A1(n19217), .A2(n19239), .ZN(n19219) );
  OAI21_X1 U22225 ( .B1(n19219), .B2(n19630), .A(n19218), .ZN(n19220) );
  MUX2_X1 U22226 ( .A(n19221), .B(n19220), .S(n19837), .Z(n19222) );
  NAND2_X1 U22227 ( .A1(n19222), .A2(n19695), .ZN(n19240) );
  AOI22_X1 U22228 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19240), .B1(
        n19239), .B2(n19697), .ZN(n19223) );
  OAI211_X1 U22229 ( .C1(n19700), .C2(n19274), .A(n19224), .B(n19223), .ZN(
        P2_U3064) );
  AOI22_X1 U22230 ( .A1(n19238), .A2(n19702), .B1(n19701), .B2(n19237), .ZN(
        n19226) );
  AOI22_X1 U22231 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19240), .B1(
        n19239), .B2(n19703), .ZN(n19225) );
  OAI211_X1 U22232 ( .C1(n19706), .C2(n19274), .A(n19226), .B(n19225), .ZN(
        P2_U3065) );
  INV_X1 U22233 ( .A(n19650), .ZN(n19707) );
  AOI22_X1 U22234 ( .A1(n19238), .A2(n19708), .B1(n19707), .B2(n19237), .ZN(
        n19228) );
  AOI22_X1 U22235 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19240), .B1(
        n19239), .B2(n19709), .ZN(n19227) );
  OAI211_X1 U22236 ( .C1(n19712), .C2(n19274), .A(n19228), .B(n19227), .ZN(
        P2_U3066) );
  INV_X1 U22237 ( .A(n19655), .ZN(n19713) );
  AOI22_X1 U22238 ( .A1(n19238), .A2(n19714), .B1(n19713), .B2(n19237), .ZN(
        n19230) );
  INV_X1 U22239 ( .A(n19718), .ZN(n19606) );
  AOI22_X1 U22240 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19240), .B1(
        n19239), .B2(n19606), .ZN(n19229) );
  OAI211_X1 U22241 ( .C1(n19656), .C2(n19274), .A(n19230), .B(n19229), .ZN(
        P2_U3067) );
  INV_X1 U22242 ( .A(n19660), .ZN(n19719) );
  AOI22_X1 U22243 ( .A1(n19238), .A2(n19720), .B1(n19719), .B2(n19237), .ZN(
        n19232) );
  AOI22_X1 U22244 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19240), .B1(
        n19239), .B2(n19721), .ZN(n19231) );
  OAI211_X1 U22245 ( .C1(n19724), .C2(n19274), .A(n19232), .B(n19231), .ZN(
        P2_U3068) );
  AOI22_X1 U22246 ( .A1(n19238), .A2(n19726), .B1(n19725), .B2(n19237), .ZN(
        n19234) );
  AOI22_X1 U22247 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19240), .B1(
        n19239), .B2(n19577), .ZN(n19233) );
  OAI211_X1 U22248 ( .C1(n19669), .C2(n19274), .A(n19234), .B(n19233), .ZN(
        P2_U3069) );
  INV_X1 U22249 ( .A(n19670), .ZN(n19731) );
  AOI22_X1 U22250 ( .A1(n19238), .A2(n19732), .B1(n19731), .B2(n19237), .ZN(
        n19236) );
  AOI22_X1 U22251 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19240), .B1(
        n19239), .B2(n19733), .ZN(n19235) );
  OAI211_X1 U22252 ( .C1(n19738), .C2(n19274), .A(n19236), .B(n19235), .ZN(
        P2_U3070) );
  AOI22_X1 U22253 ( .A1(n19238), .A2(n19741), .B1(n19740), .B2(n19237), .ZN(
        n19242) );
  AOI22_X1 U22254 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19240), .B1(
        n19239), .B2(n19620), .ZN(n19241) );
  OAI211_X1 U22255 ( .C1(n19683), .C2(n19274), .A(n19242), .B(n19241), .ZN(
        P2_U3071) );
  NAND2_X1 U22256 ( .A1(n19519), .A2(n19243), .ZN(n19273) );
  OAI22_X1 U22257 ( .A1(n19274), .A2(n19627), .B1(n19273), .B2(n19626), .ZN(
        n19244) );
  INV_X1 U22258 ( .A(n19244), .ZN(n19254) );
  OAI21_X1 U22259 ( .B1(n19517), .B2(n19388), .A(n19837), .ZN(n19252) );
  INV_X1 U22260 ( .A(n19837), .ZN(n19634) );
  OAI211_X1 U22261 ( .C1(n19247), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19273), 
        .B(n19634), .ZN(n19245) );
  OAI211_X1 U22262 ( .C1(n19252), .C2(n19246), .A(n19695), .B(n19245), .ZN(
        n19277) );
  INV_X1 U22263 ( .A(n19246), .ZN(n19251) );
  INV_X1 U22264 ( .A(n19247), .ZN(n19249) );
  INV_X1 U22265 ( .A(n19273), .ZN(n19248) );
  OAI21_X1 U22266 ( .B1(n19249), .B2(n19248), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19250) );
  AOI22_X1 U22267 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19277), .B1(
        n19689), .B2(n19276), .ZN(n19253) );
  OAI211_X1 U22268 ( .C1(n19700), .C2(n19317), .A(n19254), .B(n19253), .ZN(
        P2_U3072) );
  OAI22_X1 U22269 ( .A1(n19317), .A2(n19706), .B1(n19273), .B2(n19645), .ZN(
        n19255) );
  INV_X1 U22270 ( .A(n19255), .ZN(n19257) );
  AOI22_X1 U22271 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19277), .B1(
        n19702), .B2(n19276), .ZN(n19256) );
  OAI211_X1 U22272 ( .C1(n19646), .C2(n19274), .A(n19257), .B(n19256), .ZN(
        P2_U3073) );
  OAI22_X1 U22273 ( .A1(n19317), .A2(n19712), .B1(n19273), .B2(n19650), .ZN(
        n19258) );
  INV_X1 U22274 ( .A(n19258), .ZN(n19260) );
  AOI22_X1 U22275 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19277), .B1(
        n19708), .B2(n19276), .ZN(n19259) );
  OAI211_X1 U22276 ( .C1(n19654), .C2(n19274), .A(n19260), .B(n19259), .ZN(
        P2_U3074) );
  OAI22_X1 U22277 ( .A1(n19274), .A2(n19718), .B1(n19273), .B2(n19655), .ZN(
        n19261) );
  INV_X1 U22278 ( .A(n19261), .ZN(n19263) );
  AOI22_X1 U22279 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19277), .B1(
        n19714), .B2(n19276), .ZN(n19262) );
  OAI211_X1 U22280 ( .C1(n19656), .C2(n19317), .A(n19263), .B(n19262), .ZN(
        P2_U3075) );
  OAI22_X1 U22281 ( .A1(n19274), .A2(n19664), .B1(n19273), .B2(n19660), .ZN(
        n19264) );
  INV_X1 U22282 ( .A(n19264), .ZN(n19266) );
  AOI22_X1 U22283 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19277), .B1(
        n19720), .B2(n19276), .ZN(n19265) );
  OAI211_X1 U22284 ( .C1(n19724), .C2(n19317), .A(n19266), .B(n19265), .ZN(
        P2_U3076) );
  OAI22_X1 U22285 ( .A1(n19317), .A2(n19669), .B1(n19273), .B2(n19665), .ZN(
        n19267) );
  INV_X1 U22286 ( .A(n19267), .ZN(n19269) );
  AOI22_X1 U22287 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19277), .B1(
        n19726), .B2(n19276), .ZN(n19268) );
  OAI211_X1 U22288 ( .C1(n19730), .C2(n19274), .A(n19269), .B(n19268), .ZN(
        P2_U3077) );
  OAI22_X1 U22289 ( .A1(n19274), .A2(n19674), .B1(n19273), .B2(n19670), .ZN(
        n19270) );
  INV_X1 U22290 ( .A(n19270), .ZN(n19272) );
  AOI22_X1 U22291 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19277), .B1(
        n19732), .B2(n19276), .ZN(n19271) );
  OAI211_X1 U22292 ( .C1(n19738), .C2(n19317), .A(n19272), .B(n19271), .ZN(
        P2_U3078) );
  OAI22_X1 U22293 ( .A1(n19274), .A2(n19749), .B1(n19273), .B2(n19676), .ZN(
        n19275) );
  INV_X1 U22294 ( .A(n19275), .ZN(n19279) );
  AOI22_X1 U22295 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19277), .B1(
        n19741), .B2(n19276), .ZN(n19278) );
  OAI211_X1 U22296 ( .C1(n19683), .C2(n19317), .A(n19279), .B(n19278), .ZN(
        P2_U3079) );
  NOR2_X1 U22297 ( .A1(n19356), .A2(n19555), .ZN(n19291) );
  INV_X1 U22298 ( .A(n19291), .ZN(n19316) );
  OAI22_X1 U22299 ( .A1(n19317), .A2(n19627), .B1(n19626), .B2(n19316), .ZN(
        n19282) );
  INV_X1 U22300 ( .A(n19282), .ZN(n19297) );
  INV_X1 U22301 ( .A(n19353), .ZN(n19284) );
  INV_X1 U22302 ( .A(n19317), .ZN(n19283) );
  NOR2_X1 U22303 ( .A1(n19284), .A2(n19283), .ZN(n19285) );
  OAI21_X1 U22304 ( .B1(n19285), .B2(n19630), .A(n19837), .ZN(n19295) );
  INV_X1 U22305 ( .A(n19286), .ZN(n19632) );
  NAND2_X1 U22306 ( .A1(n19632), .A2(n19287), .ZN(n19561) );
  NOR2_X1 U22307 ( .A1(n19561), .A2(n19559), .ZN(n19290) );
  INV_X1 U22308 ( .A(n19292), .ZN(n19288) );
  OAI211_X1 U22309 ( .C1(n19288), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19316), 
        .B(n19634), .ZN(n19289) );
  OAI211_X1 U22310 ( .C1(n19295), .C2(n19290), .A(n19695), .B(n19289), .ZN(
        n19320) );
  INV_X1 U22311 ( .A(n19290), .ZN(n19294) );
  OAI21_X1 U22312 ( .B1(n19292), .B2(n19291), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19293) );
  AOI22_X1 U22313 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19320), .B1(
        n19689), .B2(n19319), .ZN(n19296) );
  OAI211_X1 U22314 ( .C1(n19700), .C2(n19353), .A(n19297), .B(n19296), .ZN(
        P2_U3080) );
  OAI22_X1 U22315 ( .A1(n19317), .A2(n19646), .B1(n19645), .B2(n19316), .ZN(
        n19298) );
  INV_X1 U22316 ( .A(n19298), .ZN(n19300) );
  AOI22_X1 U22317 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19320), .B1(
        n19702), .B2(n19319), .ZN(n19299) );
  OAI211_X1 U22318 ( .C1(n19706), .C2(n19353), .A(n19300), .B(n19299), .ZN(
        P2_U3081) );
  OAI22_X1 U22319 ( .A1(n19353), .A2(n19712), .B1(n19650), .B2(n19316), .ZN(
        n19301) );
  INV_X1 U22320 ( .A(n19301), .ZN(n19303) );
  AOI22_X1 U22321 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19320), .B1(
        n19708), .B2(n19319), .ZN(n19302) );
  OAI211_X1 U22322 ( .C1(n19654), .C2(n19317), .A(n19303), .B(n19302), .ZN(
        P2_U3082) );
  OAI22_X1 U22323 ( .A1(n19353), .A2(n19656), .B1(n19655), .B2(n19316), .ZN(
        n19304) );
  INV_X1 U22324 ( .A(n19304), .ZN(n19306) );
  AOI22_X1 U22325 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19320), .B1(
        n19714), .B2(n19319), .ZN(n19305) );
  OAI211_X1 U22326 ( .C1(n19718), .C2(n19317), .A(n19306), .B(n19305), .ZN(
        P2_U3083) );
  OAI22_X1 U22327 ( .A1(n19353), .A2(n19724), .B1(n19660), .B2(n19316), .ZN(
        n19307) );
  INV_X1 U22328 ( .A(n19307), .ZN(n19309) );
  AOI22_X1 U22329 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19320), .B1(
        n19720), .B2(n19319), .ZN(n19308) );
  OAI211_X1 U22330 ( .C1(n19664), .C2(n19317), .A(n19309), .B(n19308), .ZN(
        P2_U3084) );
  OAI22_X1 U22331 ( .A1(n19353), .A2(n19669), .B1(n19665), .B2(n19316), .ZN(
        n19310) );
  INV_X1 U22332 ( .A(n19310), .ZN(n19312) );
  AOI22_X1 U22333 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19320), .B1(
        n19726), .B2(n19319), .ZN(n19311) );
  OAI211_X1 U22334 ( .C1(n19730), .C2(n19317), .A(n19312), .B(n19311), .ZN(
        P2_U3085) );
  OAI22_X1 U22335 ( .A1(n19317), .A2(n19674), .B1(n19670), .B2(n19316), .ZN(
        n19313) );
  INV_X1 U22336 ( .A(n19313), .ZN(n19315) );
  AOI22_X1 U22337 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19320), .B1(
        n19732), .B2(n19319), .ZN(n19314) );
  OAI211_X1 U22338 ( .C1(n19738), .C2(n19353), .A(n19315), .B(n19314), .ZN(
        P2_U3086) );
  OAI22_X1 U22339 ( .A1(n19317), .A2(n19749), .B1(n19676), .B2(n19316), .ZN(
        n19318) );
  INV_X1 U22340 ( .A(n19318), .ZN(n19322) );
  AOI22_X1 U22341 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19320), .B1(
        n19741), .B2(n19319), .ZN(n19321) );
  OAI211_X1 U22342 ( .C1(n19683), .C2(n19353), .A(n19322), .B(n19321), .ZN(
        P2_U3087) );
  NOR2_X1 U22343 ( .A1(n19356), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19326) );
  INV_X1 U22344 ( .A(n19326), .ZN(n19330) );
  NOR2_X1 U22345 ( .A1(n19865), .A2(n19330), .ZN(n19348) );
  INV_X1 U22346 ( .A(n19348), .ZN(n19357) );
  OAI22_X1 U22347 ( .A1(n19353), .A2(n19627), .B1(n19626), .B2(n19357), .ZN(
        n19323) );
  INV_X1 U22348 ( .A(n19323), .ZN(n19333) );
  INV_X1 U22349 ( .A(n19594), .ZN(n19324) );
  OAI21_X1 U22350 ( .B1(n19388), .B2(n19324), .A(n19837), .ZN(n19331) );
  OAI211_X1 U22351 ( .C1(n19327), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19357), 
        .B(n19634), .ZN(n19325) );
  OAI211_X1 U22352 ( .C1(n19331), .C2(n19326), .A(n19695), .B(n19325), .ZN(
        n19350) );
  INV_X1 U22353 ( .A(n19327), .ZN(n19328) );
  OAI21_X1 U22354 ( .B1(n19328), .B2(n19348), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19329) );
  OAI21_X1 U22355 ( .B1(n19331), .B2(n19330), .A(n19329), .ZN(n19349) );
  AOI22_X1 U22356 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19350), .B1(
        n19689), .B2(n19349), .ZN(n19332) );
  OAI211_X1 U22357 ( .C1(n19700), .C2(n19358), .A(n19333), .B(n19332), .ZN(
        P2_U3088) );
  AOI22_X1 U22358 ( .A1(n19379), .A2(n19601), .B1(n19701), .B2(n19348), .ZN(
        n19335) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19350), .B1(
        n19702), .B2(n19349), .ZN(n19334) );
  OAI211_X1 U22360 ( .C1(n19646), .C2(n19353), .A(n19335), .B(n19334), .ZN(
        P2_U3089) );
  AOI22_X1 U22361 ( .A1(n19379), .A2(n19535), .B1(n19707), .B2(n19348), .ZN(
        n19337) );
  AOI22_X1 U22362 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19350), .B1(
        n19708), .B2(n19349), .ZN(n19336) );
  OAI211_X1 U22363 ( .C1(n19654), .C2(n19353), .A(n19337), .B(n19336), .ZN(
        P2_U3090) );
  OAI22_X1 U22364 ( .A1(n19353), .A2(n19718), .B1(n19655), .B2(n19357), .ZN(
        n19338) );
  INV_X1 U22365 ( .A(n19338), .ZN(n19340) );
  AOI22_X1 U22366 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19350), .B1(
        n19714), .B2(n19349), .ZN(n19339) );
  OAI211_X1 U22367 ( .C1(n19656), .C2(n19358), .A(n19340), .B(n19339), .ZN(
        P2_U3091) );
  AOI22_X1 U22368 ( .A1(n19379), .A2(n19609), .B1(n19719), .B2(n19348), .ZN(
        n19342) );
  AOI22_X1 U22369 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19350), .B1(
        n19720), .B2(n19349), .ZN(n19341) );
  OAI211_X1 U22370 ( .C1(n19664), .C2(n19353), .A(n19342), .B(n19341), .ZN(
        P2_U3092) );
  AOI22_X1 U22371 ( .A1(n19379), .A2(n19727), .B1(n19725), .B2(n19348), .ZN(
        n19344) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19350), .B1(
        n19726), .B2(n19349), .ZN(n19343) );
  OAI211_X1 U22373 ( .C1(n19730), .C2(n19353), .A(n19344), .B(n19343), .ZN(
        P2_U3093) );
  OAI22_X1 U22374 ( .A1(n19353), .A2(n19674), .B1(n19670), .B2(n19357), .ZN(
        n19345) );
  INV_X1 U22375 ( .A(n19345), .ZN(n19347) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19350), .B1(
        n19732), .B2(n19349), .ZN(n19346) );
  OAI211_X1 U22377 ( .C1(n19738), .C2(n19358), .A(n19347), .B(n19346), .ZN(
        P2_U3094) );
  INV_X1 U22378 ( .A(n19683), .ZN(n19743) );
  AOI22_X1 U22379 ( .A1(n19379), .A2(n19743), .B1(n19740), .B2(n19348), .ZN(
        n19352) );
  AOI22_X1 U22380 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19350), .B1(
        n19741), .B2(n19349), .ZN(n19351) );
  OAI211_X1 U22381 ( .C1(n19749), .C2(n19353), .A(n19352), .B(n19351), .ZN(
        P2_U3095) );
  NOR2_X1 U22382 ( .A1(n19857), .A2(n19356), .ZN(n19391) );
  INV_X1 U22383 ( .A(n19391), .ZN(n19386) );
  NOR2_X1 U22384 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19386), .ZN(
        n19377) );
  OAI21_X1 U22385 ( .B1(n19360), .B2(n19377), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19355) );
  AOI22_X1 U22386 ( .A1(n19378), .A2(n19689), .B1(n19688), .B2(n19377), .ZN(
        n19364) );
  OAI221_X1 U22387 ( .B1(n19630), .B2(n19358), .C1(n19630), .C2(n19406), .A(
        n19357), .ZN(n19359) );
  OAI211_X1 U22388 ( .C1(n19360), .C2(n19491), .A(n19359), .B(n19883), .ZN(
        n19361) );
  INV_X1 U22389 ( .A(n19361), .ZN(n19362) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19380), .B1(
        n19379), .B2(n19697), .ZN(n19363) );
  OAI211_X1 U22391 ( .C1(n19700), .C2(n19406), .A(n19364), .B(n19363), .ZN(
        P2_U3096) );
  AOI22_X1 U22392 ( .A1(n19378), .A2(n19702), .B1(n19701), .B2(n19377), .ZN(
        n19366) );
  AOI22_X1 U22393 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19380), .B1(
        n19379), .B2(n19703), .ZN(n19365) );
  OAI211_X1 U22394 ( .C1(n19706), .C2(n19406), .A(n19366), .B(n19365), .ZN(
        P2_U3097) );
  AOI22_X1 U22395 ( .A1(n19378), .A2(n19708), .B1(n19707), .B2(n19377), .ZN(
        n19368) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19380), .B1(
        n19379), .B2(n19709), .ZN(n19367) );
  OAI211_X1 U22397 ( .C1(n19712), .C2(n19406), .A(n19368), .B(n19367), .ZN(
        P2_U3098) );
  AOI22_X1 U22398 ( .A1(n19378), .A2(n19714), .B1(n19713), .B2(n19377), .ZN(
        n19370) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19380), .B1(
        n19379), .B2(n19606), .ZN(n19369) );
  OAI211_X1 U22400 ( .C1(n19656), .C2(n19406), .A(n19370), .B(n19369), .ZN(
        P2_U3099) );
  AOI22_X1 U22401 ( .A1(n19378), .A2(n19720), .B1(n19719), .B2(n19377), .ZN(
        n19372) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19380), .B1(
        n19379), .B2(n19721), .ZN(n19371) );
  OAI211_X1 U22403 ( .C1(n19724), .C2(n19406), .A(n19372), .B(n19371), .ZN(
        P2_U3100) );
  AOI22_X1 U22404 ( .A1(n19378), .A2(n19726), .B1(n19725), .B2(n19377), .ZN(
        n19374) );
  AOI22_X1 U22405 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19380), .B1(
        n19379), .B2(n19577), .ZN(n19373) );
  OAI211_X1 U22406 ( .C1(n19669), .C2(n19406), .A(n19374), .B(n19373), .ZN(
        P2_U3101) );
  AOI22_X1 U22407 ( .A1(n19378), .A2(n19732), .B1(n19731), .B2(n19377), .ZN(
        n19376) );
  AOI22_X1 U22408 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19380), .B1(
        n19379), .B2(n19733), .ZN(n19375) );
  OAI211_X1 U22409 ( .C1(n19738), .C2(n19406), .A(n19376), .B(n19375), .ZN(
        P2_U3102) );
  AOI22_X1 U22410 ( .A1(n19378), .A2(n19741), .B1(n19740), .B2(n19377), .ZN(
        n19382) );
  AOI22_X1 U22411 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19380), .B1(
        n19379), .B2(n19620), .ZN(n19381) );
  OAI211_X1 U22412 ( .C1(n19683), .C2(n19406), .A(n19382), .B(n19381), .ZN(
        P2_U3103) );
  INV_X1 U22413 ( .A(n19389), .ZN(n19384) );
  INV_X1 U22414 ( .A(n19423), .ZN(n19407) );
  OAI21_X1 U22415 ( .B1(n19384), .B2(n19407), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19385) );
  AOI22_X1 U22416 ( .A1(n19408), .A2(n19689), .B1(n19407), .B2(n19688), .ZN(
        n19393) );
  INV_X1 U22417 ( .A(n19690), .ZN(n19387) );
  NOR2_X1 U22418 ( .A1(n19388), .A2(n19387), .ZN(n19836) );
  OAI211_X1 U22419 ( .C1(n19389), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19423), 
        .B(n19634), .ZN(n19390) );
  OAI211_X1 U22420 ( .C1(n19836), .C2(n19391), .A(n19695), .B(n19390), .ZN(
        n19410) );
  INV_X1 U22421 ( .A(n19406), .ZN(n19409) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19410), .B1(
        n19409), .B2(n19697), .ZN(n19392) );
  OAI211_X1 U22423 ( .C1(n19700), .C2(n19441), .A(n19393), .B(n19392), .ZN(
        P2_U3104) );
  AOI22_X1 U22424 ( .A1(n19408), .A2(n19702), .B1(n19407), .B2(n19701), .ZN(
        n19395) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19410), .B1(
        n19445), .B2(n19601), .ZN(n19394) );
  OAI211_X1 U22426 ( .C1(n19646), .C2(n19406), .A(n19395), .B(n19394), .ZN(
        P2_U3105) );
  AOI22_X1 U22427 ( .A1(n19408), .A2(n19708), .B1(n19407), .B2(n19707), .ZN(
        n19397) );
  AOI22_X1 U22428 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19410), .B1(
        n19409), .B2(n19709), .ZN(n19396) );
  OAI211_X1 U22429 ( .C1(n19712), .C2(n19441), .A(n19397), .B(n19396), .ZN(
        P2_U3106) );
  AOI22_X1 U22430 ( .A1(n19408), .A2(n19714), .B1(n19407), .B2(n19713), .ZN(
        n19399) );
  AOI22_X1 U22431 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19410), .B1(
        n19409), .B2(n19606), .ZN(n19398) );
  OAI211_X1 U22432 ( .C1(n19656), .C2(n19441), .A(n19399), .B(n19398), .ZN(
        P2_U3107) );
  AOI22_X1 U22433 ( .A1(n19408), .A2(n19720), .B1(n19407), .B2(n19719), .ZN(
        n19401) );
  AOI22_X1 U22434 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19410), .B1(
        n19445), .B2(n19609), .ZN(n19400) );
  OAI211_X1 U22435 ( .C1(n19664), .C2(n19406), .A(n19401), .B(n19400), .ZN(
        P2_U3108) );
  AOI22_X1 U22436 ( .A1(n19408), .A2(n19726), .B1(n19407), .B2(n19725), .ZN(
        n19403) );
  AOI22_X1 U22437 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19410), .B1(
        n19445), .B2(n19727), .ZN(n19402) );
  OAI211_X1 U22438 ( .C1(n19730), .C2(n19406), .A(n19403), .B(n19402), .ZN(
        P2_U3109) );
  AOI22_X1 U22439 ( .A1(n19408), .A2(n19732), .B1(n19407), .B2(n19731), .ZN(
        n19405) );
  INV_X1 U22440 ( .A(n19738), .ZN(n19614) );
  AOI22_X1 U22441 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19410), .B1(
        n19445), .B2(n19614), .ZN(n19404) );
  OAI211_X1 U22442 ( .C1(n19674), .C2(n19406), .A(n19405), .B(n19404), .ZN(
        P2_U3110) );
  AOI22_X1 U22443 ( .A1(n19408), .A2(n19741), .B1(n19407), .B2(n19740), .ZN(
        n19412) );
  AOI22_X1 U22444 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19410), .B1(
        n19409), .B2(n19620), .ZN(n19411) );
  OAI211_X1 U22445 ( .C1(n19683), .C2(n19441), .A(n19412), .B(n19411), .ZN(
        P2_U3111) );
  NAND2_X1 U22446 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20880), .ZN(
        n19490) );
  NOR2_X1 U22447 ( .A1(n19555), .A2(n19490), .ZN(n19444) );
  AOI22_X1 U22448 ( .A1(n19445), .A2(n19697), .B1(n19444), .B2(n19688), .ZN(
        n19426) );
  NAND2_X1 U22449 ( .A1(n19441), .A2(n19486), .ZN(n19415) );
  AOI21_X1 U22450 ( .B1(n19415), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19634), 
        .ZN(n19421) );
  OAI21_X1 U22451 ( .B1(n19416), .B2(n19491), .A(n19883), .ZN(n19417) );
  AOI21_X1 U22452 ( .B1(n19421), .B2(n19423), .A(n19417), .ZN(n19418) );
  INV_X1 U22453 ( .A(n19421), .ZN(n19424) );
  NOR2_X1 U22454 ( .A1(n19419), .A2(n19491), .ZN(n19420) );
  OAI22_X1 U22455 ( .A1(n19421), .A2(P2_STATE2_REG_2__SCAN_IN), .B1(n19444), 
        .B2(n19420), .ZN(n19422) );
  AOI22_X1 U22456 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19447), .B1(
        n19689), .B2(n19446), .ZN(n19425) );
  OAI211_X1 U22457 ( .C1(n19700), .C2(n19486), .A(n19426), .B(n19425), .ZN(
        P2_U3112) );
  AOI22_X1 U22458 ( .A1(n19445), .A2(n19703), .B1(n19444), .B2(n19701), .ZN(
        n19428) );
  AOI22_X1 U22459 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19447), .B1(
        n19702), .B2(n19446), .ZN(n19427) );
  OAI211_X1 U22460 ( .C1(n19706), .C2(n19486), .A(n19428), .B(n19427), .ZN(
        P2_U3113) );
  AOI22_X1 U22461 ( .A1(n19445), .A2(n19709), .B1(n19444), .B2(n19707), .ZN(
        n19430) );
  AOI22_X1 U22462 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19447), .B1(
        n19708), .B2(n19446), .ZN(n19429) );
  OAI211_X1 U22463 ( .C1(n19712), .C2(n19486), .A(n19430), .B(n19429), .ZN(
        P2_U3114) );
  INV_X1 U22464 ( .A(n19444), .ZN(n19437) );
  OAI22_X1 U22465 ( .A1(n19486), .A2(n19656), .B1(n19437), .B2(n19655), .ZN(
        n19431) );
  INV_X1 U22466 ( .A(n19431), .ZN(n19433) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19447), .B1(
        n19714), .B2(n19446), .ZN(n19432) );
  OAI211_X1 U22468 ( .C1(n19718), .C2(n19441), .A(n19433), .B(n19432), .ZN(
        P2_U3115) );
  OAI22_X1 U22469 ( .A1(n19486), .A2(n19724), .B1(n19437), .B2(n19660), .ZN(
        n19434) );
  INV_X1 U22470 ( .A(n19434), .ZN(n19436) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19447), .B1(
        n19720), .B2(n19446), .ZN(n19435) );
  OAI211_X1 U22472 ( .C1(n19664), .C2(n19441), .A(n19436), .B(n19435), .ZN(
        P2_U3116) );
  OAI22_X1 U22473 ( .A1(n19486), .A2(n19669), .B1(n19437), .B2(n19665), .ZN(
        n19438) );
  INV_X1 U22474 ( .A(n19438), .ZN(n19440) );
  AOI22_X1 U22475 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19447), .B1(
        n19726), .B2(n19446), .ZN(n19439) );
  OAI211_X1 U22476 ( .C1(n19730), .C2(n19441), .A(n19440), .B(n19439), .ZN(
        P2_U3117) );
  AOI22_X1 U22477 ( .A1(n19445), .A2(n19733), .B1(n19444), .B2(n19731), .ZN(
        n19443) );
  AOI22_X1 U22478 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19447), .B1(
        n19732), .B2(n19446), .ZN(n19442) );
  OAI211_X1 U22479 ( .C1(n19738), .C2(n19486), .A(n19443), .B(n19442), .ZN(
        P2_U3118) );
  AOI22_X1 U22480 ( .A1(n19445), .A2(n19620), .B1(n19444), .B2(n19740), .ZN(
        n19449) );
  AOI22_X1 U22481 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19447), .B1(
        n19741), .B2(n19446), .ZN(n19448) );
  OAI211_X1 U22482 ( .C1(n19683), .C2(n19486), .A(n19449), .B(n19448), .ZN(
        P2_U3119) );
  OR2_X1 U22483 ( .A1(n19450), .A2(n19630), .ZN(n19526) );
  OAI21_X1 U22484 ( .B1(n19462), .B2(n19526), .A(n19837), .ZN(n19461) );
  INV_X1 U22485 ( .A(n19490), .ZN(n19522) );
  NAND2_X1 U22486 ( .A1(n19522), .A2(n19857), .ZN(n19460) );
  INV_X1 U22487 ( .A(n19460), .ZN(n19451) );
  OR2_X1 U22488 ( .A1(n19461), .A2(n19451), .ZN(n19456) );
  NAND2_X1 U22489 ( .A1(n19458), .A2(n19883), .ZN(n19454) );
  NOR3_X2 U22490 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19865), .A3(
        n19490), .ZN(n19493) );
  NOR2_X1 U22491 ( .A1(n19837), .A2(n19493), .ZN(n19453) );
  AOI21_X1 U22492 ( .B1(n19454), .B2(n19453), .A(n19452), .ZN(n19455) );
  INV_X1 U22493 ( .A(n19493), .ZN(n19477) );
  OAI22_X1 U22494 ( .A1(n19486), .A2(n19627), .B1(n19626), .B2(n19477), .ZN(
        n19457) );
  INV_X1 U22495 ( .A(n19457), .ZN(n19465) );
  OAI21_X1 U22496 ( .B1(n19458), .B2(n19493), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19459) );
  OAI21_X1 U22497 ( .B1(n19461), .B2(n19460), .A(n19459), .ZN(n19482) );
  INV_X1 U22498 ( .A(n19700), .ZN(n19463) );
  AOI22_X1 U22499 ( .A1(n19689), .A2(n19482), .B1(n19513), .B2(n19463), .ZN(
        n19464) );
  OAI211_X1 U22500 ( .C1(n19481), .C2(n19466), .A(n19465), .B(n19464), .ZN(
        P2_U3120) );
  AOI22_X1 U22501 ( .A1(n19513), .A2(n19601), .B1(n19493), .B2(n19701), .ZN(
        n19468) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19483), .B1(
        n19702), .B2(n19482), .ZN(n19467) );
  OAI211_X1 U22503 ( .C1(n19646), .C2(n19486), .A(n19468), .B(n19467), .ZN(
        P2_U3121) );
  AOI22_X1 U22504 ( .A1(n19513), .A2(n19535), .B1(n19493), .B2(n19707), .ZN(
        n19470) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19483), .B1(
        n19708), .B2(n19482), .ZN(n19469) );
  OAI211_X1 U22506 ( .C1(n19654), .C2(n19486), .A(n19470), .B(n19469), .ZN(
        P2_U3122) );
  AOI22_X1 U22507 ( .A1(n19513), .A2(n19715), .B1(n19713), .B2(n19493), .ZN(
        n19472) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19483), .B1(
        n19714), .B2(n19482), .ZN(n19471) );
  OAI211_X1 U22509 ( .C1(n19718), .C2(n19486), .A(n19472), .B(n19471), .ZN(
        P2_U3123) );
  AOI22_X1 U22510 ( .A1(n19513), .A2(n19609), .B1(n19719), .B2(n19493), .ZN(
        n19474) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19483), .B1(
        n19720), .B2(n19482), .ZN(n19473) );
  OAI211_X1 U22512 ( .C1(n19664), .C2(n19486), .A(n19474), .B(n19473), .ZN(
        P2_U3124) );
  AOI22_X1 U22513 ( .A1(n19513), .A2(n19727), .B1(n19725), .B2(n19493), .ZN(
        n19476) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19483), .B1(
        n19726), .B2(n19482), .ZN(n19475) );
  OAI211_X1 U22515 ( .C1(n19730), .C2(n19486), .A(n19476), .B(n19475), .ZN(
        P2_U3125) );
  OAI22_X1 U22516 ( .A1(n19486), .A2(n19674), .B1(n19477), .B2(n19670), .ZN(
        n19478) );
  INV_X1 U22517 ( .A(n19478), .ZN(n19480) );
  AOI22_X1 U22518 ( .A1(n19732), .A2(n19482), .B1(n19513), .B2(n19614), .ZN(
        n19479) );
  OAI211_X1 U22519 ( .C1(n19481), .C2(n20921), .A(n19480), .B(n19479), .ZN(
        P2_U3126) );
  AOI22_X1 U22520 ( .A1(n19513), .A2(n19743), .B1(n19493), .B2(n19740), .ZN(
        n19485) );
  AOI22_X1 U22521 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19483), .B1(
        n19741), .B2(n19482), .ZN(n19484) );
  OAI211_X1 U22522 ( .C1(n19749), .C2(n19486), .A(n19485), .B(n19484), .ZN(
        P2_U3127) );
  NOR3_X2 U22523 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19857), .A3(
        n19490), .ZN(n19511) );
  OAI21_X1 U22524 ( .B1(n19492), .B2(n19511), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19488) );
  AOI22_X1 U22525 ( .A1(n19512), .A2(n19689), .B1(n19688), .B2(n19511), .ZN(
        n19498) );
  NOR2_X1 U22526 ( .A1(n19492), .A2(n19491), .ZN(n19495) );
  AOI221_X1 U22527 ( .B1(n19549), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19513), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19493), .ZN(n19494) );
  NOR3_X1 U22528 ( .A1(n19495), .A2(n19494), .A3(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n19496) );
  AOI22_X1 U22529 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19697), .ZN(n19497) );
  OAI211_X1 U22530 ( .C1(n19700), .C2(n19544), .A(n19498), .B(n19497), .ZN(
        P2_U3128) );
  AOI22_X1 U22531 ( .A1(n19512), .A2(n19702), .B1(n19701), .B2(n19511), .ZN(
        n19500) );
  AOI22_X1 U22532 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19703), .ZN(n19499) );
  OAI211_X1 U22533 ( .C1(n19706), .C2(n19544), .A(n19500), .B(n19499), .ZN(
        P2_U3129) );
  AOI22_X1 U22534 ( .A1(n19512), .A2(n19708), .B1(n19707), .B2(n19511), .ZN(
        n19502) );
  AOI22_X1 U22535 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19709), .ZN(n19501) );
  OAI211_X1 U22536 ( .C1(n19712), .C2(n19544), .A(n19502), .B(n19501), .ZN(
        P2_U3130) );
  AOI22_X1 U22537 ( .A1(n19512), .A2(n19714), .B1(n19713), .B2(n19511), .ZN(
        n19504) );
  AOI22_X1 U22538 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19606), .ZN(n19503) );
  OAI211_X1 U22539 ( .C1(n19656), .C2(n19544), .A(n19504), .B(n19503), .ZN(
        P2_U3131) );
  AOI22_X1 U22540 ( .A1(n19512), .A2(n19720), .B1(n19719), .B2(n19511), .ZN(
        n19506) );
  AOI22_X1 U22541 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19721), .ZN(n19505) );
  OAI211_X1 U22542 ( .C1(n19724), .C2(n19544), .A(n19506), .B(n19505), .ZN(
        P2_U3132) );
  AOI22_X1 U22543 ( .A1(n19512), .A2(n19726), .B1(n19725), .B2(n19511), .ZN(
        n19508) );
  AOI22_X1 U22544 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19577), .ZN(n19507) );
  OAI211_X1 U22545 ( .C1(n19669), .C2(n19544), .A(n19508), .B(n19507), .ZN(
        P2_U3133) );
  AOI22_X1 U22546 ( .A1(n19512), .A2(n19732), .B1(n19731), .B2(n19511), .ZN(
        n19510) );
  AOI22_X1 U22547 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19733), .ZN(n19509) );
  OAI211_X1 U22548 ( .C1(n19738), .C2(n19544), .A(n19510), .B(n19509), .ZN(
        P2_U3134) );
  AOI22_X1 U22549 ( .A1(n19512), .A2(n19741), .B1(n19740), .B2(n19511), .ZN(
        n19516) );
  AOI22_X1 U22550 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19620), .ZN(n19515) );
  OAI211_X1 U22551 ( .C1(n19683), .C2(n19544), .A(n19516), .B(n19515), .ZN(
        P2_U3135) );
  INV_X1 U22552 ( .A(n19584), .ZN(n19553) );
  NAND2_X1 U22553 ( .A1(n19519), .A2(n19522), .ZN(n19524) );
  AND2_X1 U22554 ( .A1(n19524), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19520) );
  NAND2_X1 U22555 ( .A1(n19521), .A2(n19520), .ZN(n19527) );
  NAND2_X1 U22556 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19522), .ZN(
        n19525) );
  OAI21_X1 U22557 ( .B1(n19525), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19491), 
        .ZN(n19523) );
  AND2_X1 U22558 ( .A1(n19527), .A2(n19523), .ZN(n19548) );
  INV_X1 U22559 ( .A(n19524), .ZN(n19547) );
  AOI22_X1 U22560 ( .A1(n19548), .A2(n19689), .B1(n19688), .B2(n19547), .ZN(
        n19532) );
  INV_X1 U22561 ( .A(n19525), .ZN(n19530) );
  OAI211_X1 U22562 ( .C1(n19547), .C2(n19883), .A(n19527), .B(n19695), .ZN(
        n19528) );
  INV_X1 U22563 ( .A(n19528), .ZN(n19529) );
  OAI221_X1 U22564 ( .B1(n19530), .B2(n19832), .C1(n19530), .C2(n19691), .A(
        n19529), .ZN(n19550) );
  AOI22_X1 U22565 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19550), .B1(
        n19549), .B2(n19697), .ZN(n19531) );
  OAI211_X1 U22566 ( .C1(n19700), .C2(n19553), .A(n19532), .B(n19531), .ZN(
        P2_U3136) );
  AOI22_X1 U22567 ( .A1(n19548), .A2(n19702), .B1(n19701), .B2(n19547), .ZN(
        n19534) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19550), .B1(
        n19584), .B2(n19601), .ZN(n19533) );
  OAI211_X1 U22569 ( .C1(n19646), .C2(n19544), .A(n19534), .B(n19533), .ZN(
        P2_U3137) );
  AOI22_X1 U22570 ( .A1(n19548), .A2(n19708), .B1(n19707), .B2(n19547), .ZN(
        n19537) );
  AOI22_X1 U22571 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19550), .B1(
        n19584), .B2(n19535), .ZN(n19536) );
  OAI211_X1 U22572 ( .C1(n19654), .C2(n19544), .A(n19537), .B(n19536), .ZN(
        P2_U3138) );
  AOI22_X1 U22573 ( .A1(n19548), .A2(n19714), .B1(n19713), .B2(n19547), .ZN(
        n19539) );
  AOI22_X1 U22574 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19550), .B1(
        n19549), .B2(n19606), .ZN(n19538) );
  OAI211_X1 U22575 ( .C1(n19656), .C2(n19553), .A(n19539), .B(n19538), .ZN(
        P2_U3139) );
  AOI22_X1 U22576 ( .A1(n19548), .A2(n19720), .B1(n19719), .B2(n19547), .ZN(
        n19541) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19550), .B1(
        n19549), .B2(n19721), .ZN(n19540) );
  OAI211_X1 U22578 ( .C1(n19724), .C2(n19553), .A(n19541), .B(n19540), .ZN(
        P2_U3140) );
  AOI22_X1 U22579 ( .A1(n19548), .A2(n19726), .B1(n19725), .B2(n19547), .ZN(
        n19543) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19550), .B1(
        n19584), .B2(n19727), .ZN(n19542) );
  OAI211_X1 U22581 ( .C1(n19730), .C2(n19544), .A(n19543), .B(n19542), .ZN(
        P2_U3141) );
  AOI22_X1 U22582 ( .A1(n19548), .A2(n19732), .B1(n19731), .B2(n19547), .ZN(
        n19546) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19550), .B1(
        n19549), .B2(n19733), .ZN(n19545) );
  OAI211_X1 U22584 ( .C1(n19738), .C2(n19553), .A(n19546), .B(n19545), .ZN(
        P2_U3142) );
  AOI22_X1 U22585 ( .A1(n19548), .A2(n19741), .B1(n19740), .B2(n19547), .ZN(
        n19552) );
  AOI22_X1 U22586 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19550), .B1(
        n19549), .B2(n19620), .ZN(n19551) );
  OAI211_X1 U22587 ( .C1(n19683), .C2(n19553), .A(n19552), .B(n19551), .ZN(
        P2_U3143) );
  INV_X1 U22588 ( .A(n19554), .ZN(n19558) );
  INV_X1 U22589 ( .A(n19589), .ZN(n19633) );
  NOR2_X1 U22590 ( .A1(n19633), .A2(n19555), .ZN(n19582) );
  OAI21_X1 U22591 ( .B1(n19556), .B2(n19582), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19557) );
  AOI22_X1 U22592 ( .A1(n19583), .A2(n19689), .B1(n19688), .B2(n19582), .ZN(
        n19568) );
  INV_X1 U22593 ( .A(n19559), .ZN(n19562) );
  OAI21_X1 U22594 ( .B1(n19621), .B2(n19584), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19560) );
  OAI21_X1 U22595 ( .B1(n19562), .B2(n19561), .A(n19560), .ZN(n19566) );
  INV_X1 U22596 ( .A(n19582), .ZN(n19563) );
  OAI211_X1 U22597 ( .C1(n19564), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19563), 
        .B(n19634), .ZN(n19565) );
  NAND3_X1 U22598 ( .A1(n19566), .A2(n19695), .A3(n19565), .ZN(n19585) );
  AOI22_X1 U22599 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19585), .B1(
        n19584), .B2(n19697), .ZN(n19567) );
  OAI211_X1 U22600 ( .C1(n19700), .C2(n19617), .A(n19568), .B(n19567), .ZN(
        P2_U3144) );
  AOI22_X1 U22601 ( .A1(n19583), .A2(n19702), .B1(n19701), .B2(n19582), .ZN(
        n19570) );
  AOI22_X1 U22602 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19585), .B1(
        n19584), .B2(n19703), .ZN(n19569) );
  OAI211_X1 U22603 ( .C1(n19706), .C2(n19617), .A(n19570), .B(n19569), .ZN(
        P2_U3145) );
  AOI22_X1 U22604 ( .A1(n19583), .A2(n19708), .B1(n19707), .B2(n19582), .ZN(
        n19572) );
  AOI22_X1 U22605 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19585), .B1(
        n19584), .B2(n19709), .ZN(n19571) );
  OAI211_X1 U22606 ( .C1(n19712), .C2(n19617), .A(n19572), .B(n19571), .ZN(
        P2_U3146) );
  AOI22_X1 U22607 ( .A1(n19583), .A2(n19714), .B1(n19713), .B2(n19582), .ZN(
        n19574) );
  AOI22_X1 U22608 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19585), .B1(
        n19584), .B2(n19606), .ZN(n19573) );
  OAI211_X1 U22609 ( .C1(n19656), .C2(n19617), .A(n19574), .B(n19573), .ZN(
        P2_U3147) );
  AOI22_X1 U22610 ( .A1(n19583), .A2(n19720), .B1(n19719), .B2(n19582), .ZN(
        n19576) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19585), .B1(
        n19584), .B2(n19721), .ZN(n19575) );
  OAI211_X1 U22612 ( .C1(n19724), .C2(n19617), .A(n19576), .B(n19575), .ZN(
        P2_U3148) );
  AOI22_X1 U22613 ( .A1(n19583), .A2(n19726), .B1(n19725), .B2(n19582), .ZN(
        n19579) );
  AOI22_X1 U22614 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19585), .B1(
        n19584), .B2(n19577), .ZN(n19578) );
  OAI211_X1 U22615 ( .C1(n19669), .C2(n19617), .A(n19579), .B(n19578), .ZN(
        P2_U3149) );
  AOI22_X1 U22616 ( .A1(n19583), .A2(n19732), .B1(n19731), .B2(n19582), .ZN(
        n19581) );
  AOI22_X1 U22617 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19585), .B1(
        n19584), .B2(n19733), .ZN(n19580) );
  OAI211_X1 U22618 ( .C1(n19738), .C2(n19617), .A(n19581), .B(n19580), .ZN(
        P2_U3150) );
  AOI22_X1 U22619 ( .A1(n19583), .A2(n19741), .B1(n19740), .B2(n19582), .ZN(
        n19587) );
  AOI22_X1 U22620 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19585), .B1(
        n19584), .B2(n19620), .ZN(n19586) );
  OAI211_X1 U22621 ( .C1(n19683), .C2(n19617), .A(n19587), .B(n19586), .ZN(
        P2_U3151) );
  NAND2_X1 U22622 ( .A1(n19589), .A2(n19857), .ZN(n19596) );
  NOR2_X1 U22623 ( .A1(n19865), .A2(n19596), .ZN(n19618) );
  INV_X1 U22624 ( .A(n19618), .ZN(n19590) );
  NAND3_X1 U22625 ( .A1(n19591), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19590), 
        .ZN(n19597) );
  INV_X1 U22626 ( .A(n19597), .ZN(n19592) );
  AOI211_X2 U22627 ( .C1(n19491), .C2(n19596), .A(n19593), .B(n19592), .ZN(
        n19619) );
  AOI22_X1 U22628 ( .A1(n19619), .A2(n19689), .B1(n19688), .B2(n19618), .ZN(
        n19600) );
  NAND3_X1 U22629 ( .A1(n19594), .A2(n19691), .A3(n19883), .ZN(n19595) );
  OAI21_X1 U22630 ( .B1(n19862), .B2(n19596), .A(n19595), .ZN(n19598) );
  NAND3_X1 U22631 ( .A1(n19598), .A2(n19695), .A3(n19597), .ZN(n19622) );
  AOI22_X1 U22632 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19622), .B1(
        n19621), .B2(n19697), .ZN(n19599) );
  OAI211_X1 U22633 ( .C1(n19700), .C2(n19677), .A(n19600), .B(n19599), .ZN(
        P2_U3152) );
  AOI22_X1 U22634 ( .A1(n19619), .A2(n19702), .B1(n19701), .B2(n19618), .ZN(
        n19603) );
  AOI22_X1 U22635 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19622), .B1(
        n19629), .B2(n19601), .ZN(n19602) );
  OAI211_X1 U22636 ( .C1(n19646), .C2(n19617), .A(n19603), .B(n19602), .ZN(
        P2_U3153) );
  AOI22_X1 U22637 ( .A1(n19619), .A2(n19708), .B1(n19707), .B2(n19618), .ZN(
        n19605) );
  AOI22_X1 U22638 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19622), .B1(
        n19621), .B2(n19709), .ZN(n19604) );
  OAI211_X1 U22639 ( .C1(n19712), .C2(n19677), .A(n19605), .B(n19604), .ZN(
        P2_U3154) );
  AOI22_X1 U22640 ( .A1(n19619), .A2(n19714), .B1(n19713), .B2(n19618), .ZN(
        n19608) );
  AOI22_X1 U22641 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19622), .B1(
        n19621), .B2(n19606), .ZN(n19607) );
  OAI211_X1 U22642 ( .C1(n19656), .C2(n19677), .A(n19608), .B(n19607), .ZN(
        P2_U3155) );
  AOI22_X1 U22643 ( .A1(n19619), .A2(n19720), .B1(n19719), .B2(n19618), .ZN(
        n19611) );
  AOI22_X1 U22644 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19622), .B1(
        n19629), .B2(n19609), .ZN(n19610) );
  OAI211_X1 U22645 ( .C1(n19664), .C2(n19617), .A(n19611), .B(n19610), .ZN(
        P2_U3156) );
  AOI22_X1 U22646 ( .A1(n19619), .A2(n19726), .B1(n19725), .B2(n19618), .ZN(
        n19613) );
  AOI22_X1 U22647 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19622), .B1(
        n19629), .B2(n19727), .ZN(n19612) );
  OAI211_X1 U22648 ( .C1(n19730), .C2(n19617), .A(n19613), .B(n19612), .ZN(
        P2_U3157) );
  AOI22_X1 U22649 ( .A1(n19619), .A2(n19732), .B1(n19731), .B2(n19618), .ZN(
        n19616) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19622), .B1(
        n19629), .B2(n19614), .ZN(n19615) );
  OAI211_X1 U22651 ( .C1(n19674), .C2(n19617), .A(n19616), .B(n19615), .ZN(
        P2_U3158) );
  AOI22_X1 U22652 ( .A1(n19619), .A2(n19741), .B1(n19740), .B2(n19618), .ZN(
        n19624) );
  AOI22_X1 U22653 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19622), .B1(
        n19621), .B2(n19620), .ZN(n19623) );
  OAI211_X1 U22654 ( .C1(n19683), .C2(n19677), .A(n19624), .B(n19623), .ZN(
        P2_U3159) );
  NOR2_X1 U22655 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19693), .ZN(
        n19638) );
  INV_X1 U22656 ( .A(n19638), .ZN(n19675) );
  OAI22_X1 U22657 ( .A1(n19677), .A2(n19627), .B1(n19626), .B2(n19675), .ZN(
        n19628) );
  INV_X1 U22658 ( .A(n19628), .ZN(n19644) );
  NOR2_X1 U22659 ( .A1(n19734), .A2(n19629), .ZN(n19631) );
  OAI21_X1 U22660 ( .B1(n19631), .B2(n19630), .A(n19837), .ZN(n19642) );
  NOR2_X1 U22661 ( .A1(n19633), .A2(n19632), .ZN(n19637) );
  OAI211_X1 U22662 ( .C1(n19635), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19675), 
        .B(n19634), .ZN(n19636) );
  OAI211_X1 U22663 ( .C1(n19642), .C2(n19637), .A(n19695), .B(n19636), .ZN(
        n19680) );
  INV_X1 U22664 ( .A(n19637), .ZN(n19641) );
  OAI21_X1 U22665 ( .B1(n19639), .B2(n19638), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19640) );
  AOI22_X1 U22666 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19680), .B1(
        n19689), .B2(n19679), .ZN(n19643) );
  OAI211_X1 U22667 ( .C1(n19700), .C2(n19748), .A(n19644), .B(n19643), .ZN(
        P2_U3160) );
  OAI22_X1 U22668 ( .A1(n19677), .A2(n19646), .B1(n19645), .B2(n19675), .ZN(
        n19647) );
  INV_X1 U22669 ( .A(n19647), .ZN(n19649) );
  AOI22_X1 U22670 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19680), .B1(
        n19702), .B2(n19679), .ZN(n19648) );
  OAI211_X1 U22671 ( .C1(n19706), .C2(n19748), .A(n19649), .B(n19648), .ZN(
        P2_U3161) );
  OAI22_X1 U22672 ( .A1(n19748), .A2(n19712), .B1(n19650), .B2(n19675), .ZN(
        n19651) );
  INV_X1 U22673 ( .A(n19651), .ZN(n19653) );
  AOI22_X1 U22674 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19680), .B1(
        n19708), .B2(n19679), .ZN(n19652) );
  OAI211_X1 U22675 ( .C1(n19654), .C2(n19677), .A(n19653), .B(n19652), .ZN(
        P2_U3162) );
  OAI22_X1 U22676 ( .A1(n19748), .A2(n19656), .B1(n19655), .B2(n19675), .ZN(
        n19657) );
  INV_X1 U22677 ( .A(n19657), .ZN(n19659) );
  AOI22_X1 U22678 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19680), .B1(
        n19714), .B2(n19679), .ZN(n19658) );
  OAI211_X1 U22679 ( .C1(n19718), .C2(n19677), .A(n19659), .B(n19658), .ZN(
        P2_U3163) );
  OAI22_X1 U22680 ( .A1(n19748), .A2(n19724), .B1(n19660), .B2(n19675), .ZN(
        n19661) );
  INV_X1 U22681 ( .A(n19661), .ZN(n19663) );
  AOI22_X1 U22682 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19680), .B1(
        n19720), .B2(n19679), .ZN(n19662) );
  OAI211_X1 U22683 ( .C1(n19664), .C2(n19677), .A(n19663), .B(n19662), .ZN(
        P2_U3164) );
  OAI22_X1 U22684 ( .A1(n19677), .A2(n19730), .B1(n19665), .B2(n19675), .ZN(
        n19666) );
  INV_X1 U22685 ( .A(n19666), .ZN(n19668) );
  AOI22_X1 U22686 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19680), .B1(
        n19726), .B2(n19679), .ZN(n19667) );
  OAI211_X1 U22687 ( .C1(n19669), .C2(n19748), .A(n19668), .B(n19667), .ZN(
        P2_U3165) );
  OAI22_X1 U22688 ( .A1(n19748), .A2(n19738), .B1(n19670), .B2(n19675), .ZN(
        n19671) );
  INV_X1 U22689 ( .A(n19671), .ZN(n19673) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19680), .B1(
        n19732), .B2(n19679), .ZN(n19672) );
  OAI211_X1 U22691 ( .C1(n19674), .C2(n19677), .A(n19673), .B(n19672), .ZN(
        P2_U3166) );
  OAI22_X1 U22692 ( .A1(n19677), .A2(n19749), .B1(n19676), .B2(n19675), .ZN(
        n19678) );
  INV_X1 U22693 ( .A(n19678), .ZN(n19682) );
  AOI22_X1 U22694 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19680), .B1(
        n19741), .B2(n19679), .ZN(n19681) );
  OAI211_X1 U22695 ( .C1(n19683), .C2(n19748), .A(n19682), .B(n19681), .ZN(
        P2_U3167) );
  INV_X1 U22696 ( .A(n19684), .ZN(n19685) );
  NOR3_X1 U22697 ( .A1(n19685), .A2(n19739), .A3(n19491), .ZN(n19692) );
  INV_X1 U22698 ( .A(n19693), .ZN(n19686) );
  AOI21_X1 U22699 ( .B1(n19686), .B2(n19883), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19687) );
  AOI22_X1 U22700 ( .A1(n19742), .A2(n19689), .B1(n19688), .B2(n19739), .ZN(
        n19699) );
  NAND2_X1 U22701 ( .A1(n19691), .A2(n19690), .ZN(n19694) );
  AOI21_X1 U22702 ( .B1(n19694), .B2(n19693), .A(n19692), .ZN(n19696) );
  OAI211_X1 U22703 ( .C1(n19739), .C2(n19883), .A(n19696), .B(n19695), .ZN(
        n19745) );
  AOI22_X1 U22704 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19745), .B1(
        n19734), .B2(n19697), .ZN(n19698) );
  OAI211_X1 U22705 ( .C1(n19700), .C2(n19737), .A(n19699), .B(n19698), .ZN(
        P2_U3168) );
  AOI22_X1 U22706 ( .A1(n19742), .A2(n19702), .B1(n19701), .B2(n19739), .ZN(
        n19705) );
  AOI22_X1 U22707 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19745), .B1(
        n19734), .B2(n19703), .ZN(n19704) );
  OAI211_X1 U22708 ( .C1(n19706), .C2(n19737), .A(n19705), .B(n19704), .ZN(
        P2_U3169) );
  AOI22_X1 U22709 ( .A1(n19742), .A2(n19708), .B1(n19707), .B2(n19739), .ZN(
        n19711) );
  AOI22_X1 U22710 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19745), .B1(
        n19734), .B2(n19709), .ZN(n19710) );
  OAI211_X1 U22711 ( .C1(n19712), .C2(n19737), .A(n19711), .B(n19710), .ZN(
        P2_U3170) );
  AOI22_X1 U22712 ( .A1(n19742), .A2(n19714), .B1(n19713), .B2(n19739), .ZN(
        n19717) );
  AOI22_X1 U22713 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19745), .B1(
        n19744), .B2(n19715), .ZN(n19716) );
  OAI211_X1 U22714 ( .C1(n19718), .C2(n19748), .A(n19717), .B(n19716), .ZN(
        P2_U3171) );
  AOI22_X1 U22715 ( .A1(n19742), .A2(n19720), .B1(n19719), .B2(n19739), .ZN(
        n19723) );
  AOI22_X1 U22716 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19745), .B1(
        n19734), .B2(n19721), .ZN(n19722) );
  OAI211_X1 U22717 ( .C1(n19724), .C2(n19737), .A(n19723), .B(n19722), .ZN(
        P2_U3172) );
  AOI22_X1 U22718 ( .A1(n19742), .A2(n19726), .B1(n19725), .B2(n19739), .ZN(
        n19729) );
  AOI22_X1 U22719 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19745), .B1(
        n19744), .B2(n19727), .ZN(n19728) );
  OAI211_X1 U22720 ( .C1(n19730), .C2(n19748), .A(n19729), .B(n19728), .ZN(
        P2_U3173) );
  AOI22_X1 U22721 ( .A1(n19742), .A2(n19732), .B1(n19731), .B2(n19739), .ZN(
        n19736) );
  AOI22_X1 U22722 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19745), .B1(
        n19734), .B2(n19733), .ZN(n19735) );
  OAI211_X1 U22723 ( .C1(n19738), .C2(n19737), .A(n19736), .B(n19735), .ZN(
        P2_U3174) );
  AOI22_X1 U22724 ( .A1(n19742), .A2(n19741), .B1(n19740), .B2(n19739), .ZN(
        n19747) );
  AOI22_X1 U22725 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19745), .B1(
        n19744), .B2(n19743), .ZN(n19746) );
  OAI211_X1 U22726 ( .C1(n19749), .C2(n19748), .A(n19747), .B(n19746), .ZN(
        P2_U3175) );
  NAND2_X1 U22727 ( .A1(n19886), .A2(n19491), .ZN(n19750) );
  NAND4_X1 U22728 ( .A1(n19753), .A2(n19752), .A3(n19751), .A4(n19750), .ZN(
        n19754) );
  OAI221_X1 U22729 ( .B1(n19757), .B2(n19756), .C1(n19757), .C2(n19755), .A(
        n19754), .ZN(P2_U3177) );
  AND2_X1 U22730 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19758), .ZN(
        P2_U3179) );
  AND2_X1 U22731 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19758), .ZN(
        P2_U3180) );
  NOR2_X1 U22732 ( .A1(n20859), .A2(n19831), .ZN(P2_U3181) );
  AND2_X1 U22733 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19758), .ZN(
        P2_U3182) );
  AND2_X1 U22734 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19758), .ZN(
        P2_U3183) );
  NOR2_X1 U22735 ( .A1(n20845), .A2(n19831), .ZN(P2_U3184) );
  AND2_X1 U22736 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19758), .ZN(
        P2_U3185) );
  AND2_X1 U22737 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19758), .ZN(
        P2_U3186) );
  AND2_X1 U22738 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19758), .ZN(
        P2_U3187) );
  AND2_X1 U22739 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19758), .ZN(
        P2_U3188) );
  AND2_X1 U22740 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19758), .ZN(
        P2_U3189) );
  AND2_X1 U22741 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19758), .ZN(
        P2_U3190) );
  AND2_X1 U22742 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19758), .ZN(
        P2_U3191) );
  AND2_X1 U22743 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19758), .ZN(
        P2_U3192) );
  NOR2_X1 U22744 ( .A1(n20878), .A2(n19831), .ZN(P2_U3193) );
  AND2_X1 U22745 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19758), .ZN(
        P2_U3194) );
  AND2_X1 U22746 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19758), .ZN(
        P2_U3195) );
  AND2_X1 U22747 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19758), .ZN(
        P2_U3196) );
  INV_X1 U22748 ( .A(P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20864) );
  NOR2_X1 U22749 ( .A1(n20864), .A2(n19831), .ZN(P2_U3197) );
  NOR2_X1 U22750 ( .A1(n20836), .A2(n19831), .ZN(P2_U3198) );
  AND2_X1 U22751 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19758), .ZN(
        P2_U3199) );
  AND2_X1 U22752 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19758), .ZN(
        P2_U3200) );
  AND2_X1 U22753 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19758), .ZN(P2_U3201) );
  AND2_X1 U22754 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19758), .ZN(P2_U3202) );
  AND2_X1 U22755 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19758), .ZN(P2_U3203) );
  AND2_X1 U22756 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19758), .ZN(P2_U3204) );
  AND2_X1 U22757 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19758), .ZN(P2_U3205) );
  AND2_X1 U22758 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19758), .ZN(P2_U3206) );
  AND2_X1 U22759 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19758), .ZN(P2_U3207) );
  AND2_X1 U22760 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19758), .ZN(P2_U3208) );
  OAI21_X1 U22761 ( .B1(n20689), .B2(n19764), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19773) );
  INV_X1 U22762 ( .A(n19773), .ZN(n19761) );
  NAND2_X1 U22763 ( .A1(n19886), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19771) );
  INV_X1 U22764 ( .A(n19771), .ZN(n19762) );
  INV_X1 U22765 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19896) );
  NOR3_X1 U22766 ( .A1(n19762), .A2(n19896), .A3(n19763), .ZN(n19760) );
  OAI211_X1 U22767 ( .C1(HOLD), .C2(n19896), .A(n19897), .B(n19768), .ZN(
        n19759) );
  OAI21_X1 U22768 ( .B1(n19761), .B2(n19760), .A(n19759), .ZN(P2_U3209) );
  NOR2_X1 U22769 ( .A1(n19891), .A2(n19762), .ZN(n19766) );
  NOR2_X1 U22770 ( .A1(HOLD), .A2(n19763), .ZN(n19772) );
  OAI211_X1 U22771 ( .C1(n19772), .C2(n19774), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n19764), .ZN(n19765) );
  OAI211_X1 U22772 ( .C1(n19767), .C2(n20683), .A(n19766), .B(n19765), .ZN(
        P2_U3210) );
  OAI22_X1 U22773 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19768), .B1(NA), 
        .B2(n19771), .ZN(n19769) );
  OAI211_X1 U22774 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19769), .ZN(n19770) );
  OAI221_X1 U22775 ( .B1(n19773), .B2(n19772), .C1(n19773), .C2(n19771), .A(
        n19770), .ZN(P2_U3211) );
  NAND2_X1 U22776 ( .A1(n19813), .A2(n19774), .ZN(n19821) );
  CLKBUF_X1 U22777 ( .A(n19821), .Z(n19817) );
  OAI222_X1 U22778 ( .A1(n19818), .A2(n19776), .B1(n19775), .B2(n19813), .C1(
        n19777), .C2(n19817), .ZN(P2_U3212) );
  OAI222_X1 U22779 ( .A1(n19817), .A2(n13493), .B1(n19778), .B2(n19813), .C1(
        n19777), .C2(n19818), .ZN(P2_U3213) );
  OAI222_X1 U22780 ( .A1(n19821), .A2(n11948), .B1(n19779), .B2(n19813), .C1(
        n13493), .C2(n19818), .ZN(P2_U3214) );
  OAI222_X1 U22781 ( .A1(n19821), .A2(n13588), .B1(n19780), .B2(n19813), .C1(
        n11948), .C2(n19818), .ZN(P2_U3215) );
  OAI222_X1 U22782 ( .A1(n19821), .A2(n15526), .B1(n19781), .B2(n19813), .C1(
        n13588), .C2(n19818), .ZN(P2_U3216) );
  OAI222_X1 U22783 ( .A1(n19821), .A2(n15210), .B1(n19782), .B2(n19813), .C1(
        n15526), .C2(n19818), .ZN(P2_U3217) );
  OAI222_X1 U22784 ( .A1(n19821), .A2(n11961), .B1(n19783), .B2(n19813), .C1(
        n15210), .C2(n19818), .ZN(P2_U3218) );
  OAI222_X1 U22785 ( .A1(n19817), .A2(n11967), .B1(n19784), .B2(n19813), .C1(
        n11961), .C2(n19818), .ZN(P2_U3219) );
  OAI222_X1 U22786 ( .A1(n19817), .A2(n11970), .B1(n19785), .B2(n19813), .C1(
        n11967), .C2(n19818), .ZN(P2_U3220) );
  OAI222_X1 U22787 ( .A1(n19817), .A2(n11973), .B1(n19786), .B2(n19813), .C1(
        n11970), .C2(n19818), .ZN(P2_U3221) );
  OAI222_X1 U22788 ( .A1(n19817), .A2(n14817), .B1(n19787), .B2(n19813), .C1(
        n11973), .C2(n19818), .ZN(P2_U3222) );
  OAI222_X1 U22789 ( .A1(n19817), .A2(n15199), .B1(n19788), .B2(n19813), .C1(
        n14817), .C2(n19818), .ZN(P2_U3223) );
  OAI222_X1 U22790 ( .A1(n19817), .A2(n11980), .B1(n19789), .B2(n19813), .C1(
        n15199), .C2(n19818), .ZN(P2_U3224) );
  OAI222_X1 U22791 ( .A1(n19821), .A2(n15188), .B1(n19790), .B2(n19813), .C1(
        n11980), .C2(n19818), .ZN(P2_U3225) );
  OAI222_X1 U22792 ( .A1(n19821), .A2(n11986), .B1(n19791), .B2(n19813), .C1(
        n15188), .C2(n19818), .ZN(P2_U3226) );
  OAI222_X1 U22793 ( .A1(n19821), .A2(n20892), .B1(n19792), .B2(n19813), .C1(
        n11986), .C2(n19818), .ZN(P2_U3227) );
  OAI222_X1 U22794 ( .A1(n19821), .A2(n19794), .B1(n19793), .B2(n19813), .C1(
        n20892), .C2(n19818), .ZN(P2_U3228) );
  OAI222_X1 U22795 ( .A1(n19821), .A2(n19796), .B1(n19795), .B2(n19813), .C1(
        n19794), .C2(n19818), .ZN(P2_U3229) );
  OAI222_X1 U22796 ( .A1(n19821), .A2(n15128), .B1(n19797), .B2(n19813), .C1(
        n19796), .C2(n19818), .ZN(P2_U3230) );
  OAI222_X1 U22797 ( .A1(n19817), .A2(n19799), .B1(n19798), .B2(n19813), .C1(
        n15128), .C2(n19818), .ZN(P2_U3231) );
  OAI222_X1 U22798 ( .A1(n19817), .A2(n12007), .B1(n19800), .B2(n19813), .C1(
        n19799), .C2(n19818), .ZN(P2_U3232) );
  OAI222_X1 U22799 ( .A1(n19817), .A2(n19802), .B1(n19801), .B2(n19813), .C1(
        n12007), .C2(n19818), .ZN(P2_U3233) );
  OAI222_X1 U22800 ( .A1(n19817), .A2(n19804), .B1(n19803), .B2(n19813), .C1(
        n19802), .C2(n19818), .ZN(P2_U3234) );
  OAI222_X1 U22801 ( .A1(n19817), .A2(n19806), .B1(n19805), .B2(n19813), .C1(
        n19804), .C2(n19818), .ZN(P2_U3235) );
  OAI222_X1 U22802 ( .A1(n19817), .A2(n19808), .B1(n19807), .B2(n19813), .C1(
        n19806), .C2(n19818), .ZN(P2_U3236) );
  OAI222_X1 U22803 ( .A1(n19817), .A2(n19811), .B1(n19809), .B2(n19813), .C1(
        n19808), .C2(n19818), .ZN(P2_U3237) );
  OAI222_X1 U22804 ( .A1(n19818), .A2(n19811), .B1(n19810), .B2(n19813), .C1(
        n19812), .C2(n19817), .ZN(P2_U3238) );
  INV_X1 U22805 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19815) );
  OAI222_X1 U22806 ( .A1(n19817), .A2(n19815), .B1(n19814), .B2(n19813), .C1(
        n19812), .C2(n19818), .ZN(P2_U3239) );
  OAI222_X1 U22807 ( .A1(n19817), .A2(n12343), .B1(n19816), .B2(n19813), .C1(
        n19815), .C2(n19818), .ZN(P2_U3240) );
  OAI222_X1 U22808 ( .A1(n19821), .A2(n19820), .B1(n19819), .B2(n19813), .C1(
        n12343), .C2(n19818), .ZN(P2_U3241) );
  INV_X1 U22809 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19822) );
  AOI22_X1 U22810 ( .A1(n19813), .A2(n19823), .B1(n19822), .B2(n19897), .ZN(
        P2_U3585) );
  MUX2_X1 U22811 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19813), .Z(P2_U3586) );
  INV_X1 U22812 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19824) );
  AOI22_X1 U22813 ( .A1(n19813), .A2(n19825), .B1(n19824), .B2(n19897), .ZN(
        P2_U3587) );
  INV_X1 U22814 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19826) );
  AOI22_X1 U22815 ( .A1(n19813), .A2(n19827), .B1(n19826), .B2(n19897), .ZN(
        P2_U3588) );
  OAI21_X1 U22816 ( .B1(n19831), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19829), 
        .ZN(n19828) );
  INV_X1 U22817 ( .A(n19828), .ZN(P2_U3591) );
  OAI21_X1 U22818 ( .B1(n19831), .B2(n19830), .A(n19829), .ZN(P2_U3592) );
  INV_X1 U22819 ( .A(n19866), .ZN(n19858) );
  AND2_X1 U22820 ( .A1(n19837), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19853) );
  NAND2_X1 U22821 ( .A1(n19832), .A2(n19853), .ZN(n19843) );
  INV_X1 U22822 ( .A(n19833), .ZN(n19834) );
  NAND3_X1 U22823 ( .A1(n19851), .A2(n19834), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19835) );
  NAND2_X1 U22824 ( .A1(n19835), .A2(n19849), .ZN(n19844) );
  NAND2_X1 U22825 ( .A1(n19843), .A2(n19844), .ZN(n19840) );
  AOI222_X1 U22826 ( .A1(n19840), .A2(n19839), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19838), .C1(n19837), .C2(n19836), .ZN(n19841) );
  AOI22_X1 U22827 ( .A1(n19858), .A2(n19842), .B1(n19841), .B2(n19866), .ZN(
        P2_U3602) );
  OAI21_X1 U22828 ( .B1(n19845), .B2(n19844), .A(n19843), .ZN(n19846) );
  AOI21_X1 U22829 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19847), .A(n19846), 
        .ZN(n19848) );
  AOI22_X1 U22830 ( .A1(n19858), .A2(n20880), .B1(n19848), .B2(n19866), .ZN(
        P2_U3603) );
  INV_X1 U22831 ( .A(n19849), .ZN(n19860) );
  AND2_X1 U22832 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19850) );
  NOR2_X1 U22833 ( .A1(n19860), .A2(n19850), .ZN(n19852) );
  MUX2_X1 U22834 ( .A(n19853), .B(n19852), .S(n19851), .Z(n19854) );
  AOI21_X1 U22835 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19855), .A(n19854), 
        .ZN(n19856) );
  AOI22_X1 U22836 ( .A1(n19858), .A2(n19857), .B1(n19856), .B2(n19866), .ZN(
        P2_U3604) );
  OAI22_X1 U22837 ( .A1(n19861), .A2(n19860), .B1(n19491), .B2(n19859), .ZN(
        n19863) );
  OAI21_X1 U22838 ( .B1(n19863), .B2(n19862), .A(n19866), .ZN(n19864) );
  OAI21_X1 U22839 ( .B1(n19866), .B2(n19865), .A(n19864), .ZN(P2_U3605) );
  INV_X1 U22840 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19867) );
  AOI22_X1 U22841 ( .A1(n19813), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19867), 
        .B2(n19897), .ZN(P2_U3608) );
  INV_X1 U22842 ( .A(n19868), .ZN(n19874) );
  INV_X1 U22843 ( .A(n19869), .ZN(n19871) );
  AOI21_X1 U22844 ( .B1(n19872), .B2(n19871), .A(n19870), .ZN(n19873) );
  OAI21_X1 U22845 ( .B1(n19875), .B2(n19874), .A(n19873), .ZN(n19877) );
  MUX2_X1 U22846 ( .A(P2_MORE_REG_SCAN_IN), .B(n19877), .S(n19876), .Z(
        P2_U3609) );
  INV_X1 U22847 ( .A(n19878), .ZN(n19879) );
  OAI21_X1 U22848 ( .B1(n19886), .B2(n19880), .A(n19879), .ZN(n19881) );
  AOI21_X1 U22849 ( .B1(n19883), .B2(n19882), .A(n19881), .ZN(n19895) );
  NAND2_X1 U22850 ( .A1(n19884), .A2(n19890), .ZN(n19888) );
  OAI21_X1 U22851 ( .B1(n19886), .B2(n19491), .A(n19885), .ZN(n19887) );
  OAI21_X1 U22852 ( .B1(n19888), .B2(n19891), .A(n19887), .ZN(n19889) );
  INV_X1 U22853 ( .A(n19889), .ZN(n19894) );
  AOI211_X1 U22854 ( .C1(n19891), .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19890), 
        .B(n11422), .ZN(n19892) );
  NOR2_X1 U22855 ( .A1(n19895), .A2(n19892), .ZN(n19893) );
  AOI22_X1 U22856 ( .A1(n19896), .A2(n19895), .B1(n19894), .B2(n19893), .ZN(
        P2_U3610) );
  INV_X1 U22857 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19898) );
  AOI22_X1 U22858 ( .A1(n19813), .A2(n19899), .B1(n19898), .B2(n19897), .ZN(
        P2_U3611) );
  OAI21_X1 U22859 ( .B1(n20686), .B2(P1_STATE_REG_2__SCAN_IN), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n19906) );
  INV_X2 U22860 ( .A(n20765), .ZN(n20777) );
  OAI21_X1 U22861 ( .B1(n19906), .B2(P1_ADS_N_REG_SCAN_IN), .A(n20777), .ZN(
        n19900) );
  INV_X1 U22862 ( .A(n19900), .ZN(P1_U2802) );
  OAI21_X1 U22863 ( .B1(n19902), .B2(n19901), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19903) );
  OAI21_X1 U22864 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19904), .A(n19903), 
        .ZN(P1_U2803) );
  NOR2_X1 U22865 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19907) );
  OAI21_X1 U22866 ( .B1(n19907), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20777), .ZN(
        n19905) );
  OAI21_X1 U22867 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20777), .A(n19905), 
        .ZN(P1_U2804) );
  OAI21_X1 U22868 ( .B1(BS16), .B2(n19907), .A(n20757), .ZN(n20755) );
  OAI21_X1 U22869 ( .B1(n20757), .B2(n20254), .A(n20755), .ZN(P1_U2805) );
  OAI21_X1 U22870 ( .B1(n19910), .B2(n19909), .A(n19908), .ZN(P1_U2806) );
  NOR4_X1 U22871 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19914) );
  NOR4_X1 U22872 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19913) );
  NOR4_X1 U22873 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19912) );
  NOR4_X1 U22874 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19911) );
  NAND4_X1 U22875 ( .A1(n19914), .A2(n19913), .A3(n19912), .A4(n19911), .ZN(
        n19920) );
  NOR4_X1 U22876 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19918) );
  AOI211_X1 U22877 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19917) );
  NOR4_X1 U22878 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19916) );
  NOR4_X1 U22879 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19915) );
  NAND4_X1 U22880 ( .A1(n19918), .A2(n19917), .A3(n19916), .A4(n19915), .ZN(
        n19919) );
  NOR2_X1 U22881 ( .A1(n19920), .A2(n19919), .ZN(n20760) );
  INV_X1 U22882 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20750) );
  NOR3_X1 U22883 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19922) );
  OAI21_X1 U22884 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19922), .A(n20760), .ZN(
        n19921) );
  OAI21_X1 U22885 ( .B1(n20760), .B2(n20750), .A(n19921), .ZN(P1_U2807) );
  INV_X1 U22886 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20756) );
  AOI21_X1 U22887 ( .B1(n14227), .B2(n20756), .A(n19922), .ZN(n19923) );
  INV_X1 U22888 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20748) );
  INV_X1 U22889 ( .A(n20760), .ZN(n20762) );
  AOI22_X1 U22890 ( .A1(n20760), .A2(n19923), .B1(n20748), .B2(n20762), .ZN(
        P1_U2808) );
  NAND2_X1 U22891 ( .A1(n19925), .A2(n19924), .ZN(n19940) );
  INV_X1 U22892 ( .A(n19940), .ZN(n19961) );
  AOI21_X1 U22893 ( .B1(n19926), .B2(n19961), .A(P1_REIP_REG_9__SCAN_IN), .ZN(
        n19933) );
  OAI22_X1 U22894 ( .A1(n19928), .A2(n19927), .B1(n20002), .B2(n19936), .ZN(
        n19929) );
  AOI211_X1 U22895 ( .C1(n19983), .C2(n19998), .A(n19973), .B(n19929), .ZN(
        n19932) );
  AOI22_X1 U22896 ( .A1(n20000), .A2(n19955), .B1(n19993), .B2(n19930), .ZN(
        n19931) );
  OAI211_X1 U22897 ( .C1(n19934), .C2(n19933), .A(n19932), .B(n19931), .ZN(
        P1_U2831) );
  INV_X1 U22898 ( .A(n19935), .ZN(n19938) );
  OAI22_X1 U22899 ( .A1(n19938), .A2(n19971), .B1(n19937), .B2(n19936), .ZN(
        n19939) );
  AOI211_X1 U22900 ( .C1(n19986), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19973), .B(n19939), .ZN(n19946) );
  OAI21_X1 U22901 ( .B1(n19941), .B2(n19940), .A(n20704), .ZN(n19943) );
  AOI22_X1 U22902 ( .A1(n19944), .A2(n19955), .B1(n19943), .B2(n19942), .ZN(
        n19945) );
  OAI211_X1 U22903 ( .C1(n19947), .C2(n19981), .A(n19946), .B(n19945), .ZN(
        P1_U2833) );
  INV_X1 U22904 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20702) );
  AOI22_X1 U22905 ( .A1(n19983), .A2(n19948), .B1(n19982), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n19949) );
  OAI21_X1 U22906 ( .B1(n19950), .B2(n20702), .A(n19949), .ZN(n19951) );
  INV_X1 U22907 ( .A(n19951), .ZN(n19958) );
  NAND2_X1 U22908 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19961), .ZN(n19953) );
  AOI21_X1 U22909 ( .B1(n19986), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n19973), .ZN(n19952) );
  OAI21_X1 U22910 ( .B1(n19953), .B2(P1_REIP_REG_6__SCAN_IN), .A(n19952), .ZN(
        n19954) );
  AOI21_X1 U22911 ( .B1(n19956), .B2(n19955), .A(n19954), .ZN(n19957) );
  OAI211_X1 U22912 ( .C1(n19959), .C2(n19981), .A(n19958), .B(n19957), .ZN(
        P1_U2834) );
  INV_X1 U22913 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20700) );
  AOI22_X1 U22914 ( .A1(n19983), .A2(n19960), .B1(n19982), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n19968) );
  AOI22_X1 U22915 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19986), .B1(
        n19961), .B2(n20700), .ZN(n19963) );
  OAI211_X1 U22916 ( .C1(n19981), .C2(n19964), .A(n19963), .B(n19962), .ZN(
        n19965) );
  AOI21_X1 U22917 ( .B1(n19966), .B2(n19978), .A(n19965), .ZN(n19967) );
  OAI211_X1 U22918 ( .C1(n20700), .C2(n19975), .A(n19968), .B(n19967), .ZN(
        P1_U2835) );
  AOI22_X1 U22919 ( .A1(n19969), .A2(n19987), .B1(n19982), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n19970) );
  OAI21_X1 U22920 ( .B1(n19971), .B2(n20039), .A(n19970), .ZN(n19972) );
  AOI211_X1 U22921 ( .C1(n19986), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n19973), .B(n19972), .ZN(n19980) );
  INV_X1 U22922 ( .A(n19985), .ZN(n19974) );
  OAI21_X1 U22923 ( .B1(n19984), .B2(n19974), .A(n20697), .ZN(n19977) );
  INV_X1 U22924 ( .A(n19975), .ZN(n19976) );
  AOI22_X1 U22925 ( .A1(n20030), .A2(n19978), .B1(n19977), .B2(n19976), .ZN(
        n19979) );
  OAI211_X1 U22926 ( .C1(n20035), .C2(n19981), .A(n19980), .B(n19979), .ZN(
        P1_U2836) );
  AOI22_X1 U22927 ( .A1(n19983), .A2(n20047), .B1(n19982), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n19996) );
  OAI211_X1 U22928 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(P1_REIP_REG_2__SCAN_IN), 
        .A(n19985), .B(n19984), .ZN(n19989) );
  AOI22_X1 U22929 ( .A1(n9603), .A2(n19987), .B1(n19986), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19988) );
  OAI211_X1 U22930 ( .C1(n19991), .C2(n19990), .A(n19989), .B(n19988), .ZN(
        n19992) );
  AOI21_X1 U22931 ( .B1(n19994), .B2(n19993), .A(n19992), .ZN(n19995) );
  OAI211_X1 U22932 ( .C1(n19997), .C2(n13528), .A(n19996), .B(n19995), .ZN(
        P1_U2837) );
  AOI22_X1 U22933 ( .A1(n20000), .A2(n19999), .B1(n12418), .B2(n19998), .ZN(
        n20001) );
  OAI21_X1 U22934 ( .B1(n20003), .B2(n20002), .A(n20001), .ZN(P1_U2863) );
  INV_X1 U22935 ( .A(P1_UWORD_REG_13__SCAN_IN), .ZN(n20814) );
  AOI22_X1 U22936 ( .A1(n20009), .A2(P1_DATAO_REG_29__SCAN_IN), .B1(n20004), 
        .B2(P1_EAX_REG_29__SCAN_IN), .ZN(n20005) );
  OAI21_X1 U22937 ( .B1(n20814), .B2(n20011), .A(n20005), .ZN(P1_U2907) );
  AOI22_X1 U22938 ( .A1(n20008), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20769), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20006) );
  OAI21_X1 U22939 ( .B1(n20877), .B2(n20007), .A(n20006), .ZN(P1_U2923) );
  INV_X1 U22940 ( .A(P1_LWORD_REG_9__SCAN_IN), .ZN(n20848) );
  AOI22_X1 U22941 ( .A1(n20009), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(
        P1_EAX_REG_9__SCAN_IN), .B2(n20008), .ZN(n20010) );
  OAI21_X1 U22942 ( .B1(n20848), .B2(n20011), .A(n20010), .ZN(P1_U2927) );
  INV_X1 U22943 ( .A(n20012), .ZN(n20013) );
  NAND2_X1 U22944 ( .A1(n20014), .A2(n20013), .ZN(n20022) );
  INV_X1 U22945 ( .A(n20022), .ZN(n20015) );
  AOI21_X1 U22946 ( .B1(n20021), .B2(P1_EAX_REG_29__SCAN_IN), .A(n20015), .ZN(
        n20016) );
  OAI21_X1 U22947 ( .B1(n20019), .B2(n20814), .A(n20016), .ZN(P1_U2950) );
  AOI21_X1 U22948 ( .B1(n20021), .B2(P1_EAX_REG_9__SCAN_IN), .A(n20017), .ZN(
        n20018) );
  OAI21_X1 U22949 ( .B1(n20019), .B2(n20848), .A(n20018), .ZN(P1_U2961) );
  AOI22_X1 U22950 ( .A1(n20021), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20020), .ZN(n20023) );
  NAND2_X1 U22951 ( .A1(n20023), .A2(n20022), .ZN(P1_U2965) );
  AOI22_X1 U22952 ( .A1(n20025), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20024), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20034) );
  OAI21_X1 U22953 ( .B1(n20028), .B2(n20027), .A(n20026), .ZN(n20029) );
  INV_X1 U22954 ( .A(n20029), .ZN(n20043) );
  AOI22_X1 U22955 ( .A1(n20043), .A2(n20032), .B1(n20031), .B2(n20030), .ZN(
        n20033) );
  OAI211_X1 U22956 ( .C1(n20036), .C2(n20035), .A(n20034), .B(n20033), .ZN(
        P1_U2995) );
  NOR2_X1 U22957 ( .A1(n20057), .A2(n20037), .ZN(n20067) );
  AOI211_X1 U22958 ( .C1(n20061), .C2(n20038), .A(n20067), .B(n20059), .ZN(
        n20055) );
  OAI22_X1 U22959 ( .A1(n20079), .A2(n20039), .B1(n20697), .B2(n20065), .ZN(
        n20042) );
  AOI211_X1 U22960 ( .C1(n20045), .C2(n20054), .A(n20049), .B(n20040), .ZN(
        n20041) );
  AOI211_X1 U22961 ( .C1(n20043), .C2(n20062), .A(n20042), .B(n20041), .ZN(
        n20044) );
  OAI21_X1 U22962 ( .B1(n20055), .B2(n20045), .A(n20044), .ZN(P1_U3027) );
  AOI21_X1 U22963 ( .B1(n20048), .B2(n20047), .A(n20046), .ZN(n20053) );
  INV_X1 U22964 ( .A(n20049), .ZN(n20050) );
  AOI22_X1 U22965 ( .A1(n20051), .A2(n20062), .B1(n20050), .B2(n20054), .ZN(
        n20052) );
  OAI211_X1 U22966 ( .C1(n20055), .C2(n20054), .A(n20053), .B(n20052), .ZN(
        P1_U3028) );
  NAND2_X1 U22967 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20056), .ZN(
        n20072) );
  NOR3_X1 U22968 ( .A1(n20058), .A2(n20086), .A3(n20057), .ZN(n20060) );
  AOI211_X1 U22969 ( .C1(n20086), .C2(n20061), .A(n20060), .B(n20059), .ZN(
        n20070) );
  AND3_X1 U22970 ( .A1(n20063), .A2(n20062), .A3(n13469), .ZN(n20068) );
  OAI22_X1 U22971 ( .A1(n20079), .A2(n9864), .B1(n20695), .B2(n20065), .ZN(
        n20066) );
  NOR3_X1 U22972 ( .A1(n20068), .A2(n20067), .A3(n20066), .ZN(n20069) );
  OAI221_X1 U22973 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20072), .C1(
        n20071), .C2(n20070), .A(n20069), .ZN(P1_U3029) );
  NOR2_X1 U22974 ( .A1(n20074), .A2(n20073), .ZN(n20082) );
  NAND3_X1 U22975 ( .A1(n20086), .A2(n20076), .A3(n20075), .ZN(n20078) );
  OAI211_X1 U22976 ( .C1(n20080), .C2(n20079), .A(n20078), .B(n20077), .ZN(
        n20081) );
  AOI21_X1 U22977 ( .B1(n20082), .B2(n13152), .A(n20081), .ZN(n20083) );
  OAI221_X1 U22978 ( .B1(n20086), .B2(n20085), .C1(n20086), .C2(n20084), .A(
        n20083), .ZN(P1_U3030) );
  NOR2_X1 U22979 ( .A1(n20088), .A2(n20087), .ZN(P1_U3032) );
  AOI22_X2 U22980 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n9575), .B1(DATAI_16_), 
        .B2(n9574), .ZN(n20628) );
  INV_X1 U22981 ( .A(n20093), .ZN(n20094) );
  AOI22_X1 U22982 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n9575), .B1(DATAI_24_), 
        .B2(n9574), .ZN(n20577) );
  NAND2_X1 U22983 ( .A1(n20142), .A2(n10224), .ZN(n20426) );
  NAND3_X1 U22984 ( .A1(n20473), .A2(n20425), .A3(n20505), .ZN(n20151) );
  OR2_X1 U22985 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20151), .ZN(
        n20143) );
  OAI22_X1 U22986 ( .A1(n20674), .A2(n20577), .B1(n20426), .B2(n20143), .ZN(
        n20098) );
  INV_X1 U22987 ( .A(n20098), .ZN(n20112) );
  INV_X1 U22988 ( .A(n20099), .ZN(n20374) );
  INV_X1 U22989 ( .A(n20430), .ZN(n20100) );
  NOR2_X1 U22990 ( .A1(n20374), .A2(n20100), .ZN(n20108) );
  NAND2_X1 U22991 ( .A1(n20107), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20565) );
  INV_X1 U22992 ( .A(n20257), .ZN(n20101) );
  NAND3_X1 U22993 ( .A1(n20177), .A2(n20624), .A3(n20674), .ZN(n20102) );
  NAND2_X1 U22994 ( .A1(n20624), .A2(n20254), .ZN(n20507) );
  NAND2_X1 U22995 ( .A1(n20102), .A2(n20507), .ZN(n20106) );
  NOR2_X1 U22996 ( .A1(n9603), .A2(n20103), .ZN(n20216) );
  NAND2_X1 U22997 ( .A1(n20216), .A2(n13648), .ZN(n20109) );
  AOI22_X1 U22998 ( .A1(n20106), .A2(n20109), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20143), .ZN(n20104) );
  NOR2_X2 U22999 ( .A1(n20105), .A2(n20257), .ZN(n20616) );
  INV_X1 U23000 ( .A(n20106), .ZN(n20110) );
  NOR2_X1 U23001 ( .A1(n20107), .A2(n20613), .ZN(n20258) );
  INV_X1 U23002 ( .A(n20258), .ZN(n20436) );
  INV_X1 U23003 ( .A(n20108), .ZN(n20253) );
  AOI22_X1 U23004 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20147), .B1(
        n20616), .B2(n20146), .ZN(n20111) );
  OAI211_X1 U23005 ( .C1(n20628), .C2(n20177), .A(n20112), .B(n20111), .ZN(
        P1_U3033) );
  AOI22_X1 U23006 ( .A1(DATAI_17_), .A2(n9574), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n9575), .ZN(n20634) );
  NAND2_X1 U23007 ( .A1(n20142), .A2(n10222), .ZN(n20441) );
  OAI22_X1 U23008 ( .A1(n20674), .A2(n20581), .B1(n20441), .B2(n20143), .ZN(
        n20113) );
  INV_X1 U23009 ( .A(n20113), .ZN(n20116) );
  NOR2_X2 U23010 ( .A1(n20114), .A2(n20257), .ZN(n20630) );
  AOI22_X1 U23011 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20147), .B1(
        n20630), .B2(n20146), .ZN(n20115) );
  OAI211_X1 U23012 ( .C1(n20634), .C2(n20177), .A(n20116), .B(n20115), .ZN(
        P1_U3034) );
  AOI22_X2 U23013 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n9575), .B1(DATAI_18_), 
        .B2(n9574), .ZN(n20640) );
  AOI22_X1 U23014 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n9575), .B1(DATAI_26_), 
        .B2(n9574), .ZN(n20585) );
  NAND2_X1 U23015 ( .A1(n20142), .A2(n20117), .ZN(n20445) );
  OAI22_X1 U23016 ( .A1(n20674), .A2(n20585), .B1(n20445), .B2(n20143), .ZN(
        n20118) );
  INV_X1 U23017 ( .A(n20118), .ZN(n20121) );
  NOR2_X2 U23018 ( .A1(n20119), .A2(n20257), .ZN(n20636) );
  AOI22_X1 U23019 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20147), .B1(
        n20636), .B2(n20146), .ZN(n20120) );
  OAI211_X1 U23020 ( .C1(n20640), .C2(n20177), .A(n20121), .B(n20120), .ZN(
        P1_U3035) );
  AOI22_X1 U23021 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n9575), .B1(DATAI_27_), 
        .B2(n9574), .ZN(n20589) );
  NAND2_X1 U23022 ( .A1(n20142), .A2(n20122), .ZN(n20449) );
  OAI22_X1 U23023 ( .A1(n20674), .A2(n20589), .B1(n20449), .B2(n20143), .ZN(
        n20123) );
  INV_X1 U23024 ( .A(n20123), .ZN(n20126) );
  NOR2_X2 U23025 ( .A1(n20124), .A2(n20257), .ZN(n20642) );
  AOI22_X1 U23026 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20147), .B1(
        n20642), .B2(n20146), .ZN(n20125) );
  OAI211_X1 U23027 ( .C1(n20646), .C2(n20177), .A(n20126), .B(n20125), .ZN(
        P1_U3036) );
  AOI22_X1 U23028 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n9575), .B1(DATAI_28_), 
        .B2(n9574), .ZN(n20593) );
  NAND2_X1 U23029 ( .A1(n20142), .A2(n20127), .ZN(n20453) );
  OAI22_X1 U23030 ( .A1(n20674), .A2(n20593), .B1(n20453), .B2(n20143), .ZN(
        n20128) );
  INV_X1 U23031 ( .A(n20128), .ZN(n20131) );
  NOR2_X2 U23032 ( .A1(n20129), .A2(n20257), .ZN(n20648) );
  AOI22_X1 U23033 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20147), .B1(
        n20648), .B2(n20146), .ZN(n20130) );
  OAI211_X1 U23034 ( .C1(n20652), .C2(n20177), .A(n20131), .B(n20130), .ZN(
        P1_U3037) );
  AOI22_X1 U23035 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n9575), .B1(DATAI_29_), 
        .B2(n9574), .ZN(n20597) );
  NAND2_X1 U23036 ( .A1(n20142), .A2(n20132), .ZN(n20457) );
  OAI22_X1 U23037 ( .A1(n20674), .A2(n20597), .B1(n20457), .B2(n20143), .ZN(
        n20133) );
  INV_X1 U23038 ( .A(n20133), .ZN(n20136) );
  NOR2_X2 U23039 ( .A1(n20134), .A2(n20257), .ZN(n20654) );
  AOI22_X1 U23040 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20147), .B1(
        n20654), .B2(n20146), .ZN(n20135) );
  OAI211_X1 U23041 ( .C1(n20658), .C2(n20177), .A(n20136), .B(n20135), .ZN(
        P1_U3038) );
  AOI22_X1 U23042 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n9575), .B1(DATAI_30_), 
        .B2(n9574), .ZN(n20601) );
  NAND2_X1 U23043 ( .A1(n20142), .A2(n10209), .ZN(n20461) );
  OAI22_X1 U23044 ( .A1(n20674), .A2(n20601), .B1(n20461), .B2(n20143), .ZN(
        n20137) );
  INV_X1 U23045 ( .A(n20137), .ZN(n20140) );
  NOR2_X2 U23046 ( .A1(n20138), .A2(n20257), .ZN(n20660) );
  AOI22_X1 U23047 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20147), .B1(
        n20660), .B2(n20146), .ZN(n20139) );
  OAI211_X1 U23048 ( .C1(n20664), .C2(n20177), .A(n20140), .B(n20139), .ZN(
        P1_U3039) );
  AOI22_X1 U23049 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n9575), .B1(DATAI_23_), 
        .B2(n9574), .ZN(n20675) );
  NAND2_X1 U23050 ( .A1(n20142), .A2(n10229), .ZN(n20465) );
  OAI22_X1 U23051 ( .A1(n20674), .A2(n20609), .B1(n20465), .B2(n20143), .ZN(
        n20144) );
  INV_X1 U23052 ( .A(n20144), .ZN(n20149) );
  NOR2_X2 U23053 ( .A1(n20145), .A2(n20257), .ZN(n20668) );
  AOI22_X1 U23054 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20147), .B1(
        n20668), .B2(n20146), .ZN(n20148) );
  OAI211_X1 U23055 ( .C1(n20675), .C2(n20177), .A(n20149), .B(n20148), .ZN(
        P1_U3040) );
  INV_X1 U23056 ( .A(n20150), .ZN(n20537) );
  NOR2_X1 U23057 ( .A1(n20536), .A2(n20151), .ZN(n20171) );
  AOI21_X1 U23058 ( .B1(n20216), .B2(n20537), .A(n20171), .ZN(n20152) );
  OAI22_X1 U23059 ( .A1(n20152), .A2(n20622), .B1(n20151), .B2(n20613), .ZN(
        n20172) );
  AOI22_X1 U23060 ( .A1(n20616), .A2(n20172), .B1(n20615), .B2(n20171), .ZN(
        n20157) );
  INV_X1 U23061 ( .A(n20151), .ZN(n20155) );
  OAI21_X1 U23062 ( .B1(n20153), .B2(n20541), .A(n20152), .ZN(n20154) );
  OAI221_X1 U23063 ( .B1(n20624), .B2(n20155), .C1(n20622), .C2(n20154), .A(
        n20620), .ZN(n20174) );
  INV_X1 U23064 ( .A(n20177), .ZN(n20164) );
  INV_X1 U23065 ( .A(n20577), .ZN(n20625) );
  AOI22_X1 U23066 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20174), .B1(
        n20164), .B2(n20625), .ZN(n20156) );
  OAI211_X1 U23067 ( .C1(n20628), .C2(n20210), .A(n20157), .B(n20156), .ZN(
        P1_U3041) );
  AOI22_X1 U23068 ( .A1(n20630), .A2(n20172), .B1(n20629), .B2(n20171), .ZN(
        n20159) );
  INV_X1 U23069 ( .A(n20634), .ZN(n20578) );
  AOI22_X1 U23070 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20174), .B1(
        n20173), .B2(n20578), .ZN(n20158) );
  OAI211_X1 U23071 ( .C1(n20581), .C2(n20177), .A(n20159), .B(n20158), .ZN(
        P1_U3042) );
  AOI22_X1 U23072 ( .A1(n20636), .A2(n20172), .B1(n20635), .B2(n20171), .ZN(
        n20161) );
  INV_X1 U23073 ( .A(n20640), .ZN(n20582) );
  AOI22_X1 U23074 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20174), .B1(
        n20173), .B2(n20582), .ZN(n20160) );
  OAI211_X1 U23075 ( .C1(n20585), .C2(n20177), .A(n20161), .B(n20160), .ZN(
        P1_U3043) );
  AOI22_X1 U23076 ( .A1(n20642), .A2(n20172), .B1(n20641), .B2(n20171), .ZN(
        n20163) );
  INV_X1 U23077 ( .A(n20646), .ZN(n20586) );
  AOI22_X1 U23078 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20174), .B1(
        n20173), .B2(n20586), .ZN(n20162) );
  OAI211_X1 U23079 ( .C1(n20589), .C2(n20177), .A(n20163), .B(n20162), .ZN(
        P1_U3044) );
  AOI22_X1 U23080 ( .A1(n20648), .A2(n20172), .B1(n20647), .B2(n20171), .ZN(
        n20166) );
  INV_X1 U23081 ( .A(n20593), .ZN(n20649) );
  AOI22_X1 U23082 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20174), .B1(
        n20164), .B2(n20649), .ZN(n20165) );
  OAI211_X1 U23083 ( .C1(n20652), .C2(n20210), .A(n20166), .B(n20165), .ZN(
        P1_U3045) );
  AOI22_X1 U23084 ( .A1(n20654), .A2(n20172), .B1(n20653), .B2(n20171), .ZN(
        n20168) );
  INV_X1 U23085 ( .A(n20658), .ZN(n20594) );
  AOI22_X1 U23086 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20174), .B1(
        n20173), .B2(n20594), .ZN(n20167) );
  OAI211_X1 U23087 ( .C1(n20597), .C2(n20177), .A(n20168), .B(n20167), .ZN(
        P1_U3046) );
  AOI22_X1 U23088 ( .A1(n20660), .A2(n20172), .B1(n20659), .B2(n20171), .ZN(
        n20170) );
  INV_X1 U23089 ( .A(n20664), .ZN(n20598) );
  AOI22_X1 U23090 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20174), .B1(
        n20173), .B2(n20598), .ZN(n20169) );
  OAI211_X1 U23091 ( .C1(n20601), .C2(n20177), .A(n20170), .B(n20169), .ZN(
        P1_U3047) );
  AOI22_X1 U23092 ( .A1(n20668), .A2(n20172), .B1(n20665), .B2(n20171), .ZN(
        n20176) );
  INV_X1 U23093 ( .A(n20675), .ZN(n20604) );
  AOI22_X1 U23094 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20174), .B1(
        n20173), .B2(n20604), .ZN(n20175) );
  OAI211_X1 U23095 ( .C1(n20609), .C2(n20177), .A(n20176), .B(n20175), .ZN(
        P1_U3048) );
  NAND3_X1 U23096 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20473), .A3(
        n20425), .ZN(n20221) );
  OR2_X1 U23097 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20221), .ZN(
        n20204) );
  OAI22_X1 U23098 ( .A1(n20245), .A2(n20628), .B1(n20426), .B2(n20204), .ZN(
        n20178) );
  INV_X1 U23099 ( .A(n20178), .ZN(n20185) );
  NAND2_X1 U23100 ( .A1(n20245), .A2(n20210), .ZN(n20179) );
  AOI21_X1 U23101 ( .B1(n20179), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20622), 
        .ZN(n20181) );
  NAND2_X1 U23102 ( .A1(n20216), .A2(n20564), .ZN(n20182) );
  AOI22_X1 U23103 ( .A1(n20181), .A2(n20182), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20204), .ZN(n20180) );
  OR2_X1 U23104 ( .A1(n20430), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20312) );
  NAND2_X1 U23105 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20312), .ZN(n20309) );
  NAND3_X1 U23106 ( .A1(n20433), .A2(n20180), .A3(n20309), .ZN(n20207) );
  INV_X1 U23107 ( .A(n20181), .ZN(n20183) );
  AOI22_X1 U23108 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20207), .B1(
        n20616), .B2(n20206), .ZN(n20184) );
  OAI211_X1 U23109 ( .C1(n20577), .C2(n20210), .A(n20185), .B(n20184), .ZN(
        P1_U3049) );
  OAI22_X1 U23110 ( .A1(n20245), .A2(n20634), .B1(n20441), .B2(n20204), .ZN(
        n20186) );
  INV_X1 U23111 ( .A(n20186), .ZN(n20188) );
  AOI22_X1 U23112 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20207), .B1(
        n20630), .B2(n20206), .ZN(n20187) );
  OAI211_X1 U23113 ( .C1(n20581), .C2(n20210), .A(n20188), .B(n20187), .ZN(
        P1_U3050) );
  OAI22_X1 U23114 ( .A1(n20245), .A2(n20640), .B1(n20445), .B2(n20204), .ZN(
        n20189) );
  INV_X1 U23115 ( .A(n20189), .ZN(n20191) );
  AOI22_X1 U23116 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20207), .B1(
        n20636), .B2(n20206), .ZN(n20190) );
  OAI211_X1 U23117 ( .C1(n20585), .C2(n20210), .A(n20191), .B(n20190), .ZN(
        P1_U3051) );
  OAI22_X1 U23118 ( .A1(n20210), .A2(n20589), .B1(n20449), .B2(n20204), .ZN(
        n20192) );
  INV_X1 U23119 ( .A(n20192), .ZN(n20194) );
  AOI22_X1 U23120 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20207), .B1(
        n20642), .B2(n20206), .ZN(n20193) );
  OAI211_X1 U23121 ( .C1(n20646), .C2(n20245), .A(n20194), .B(n20193), .ZN(
        P1_U3052) );
  OAI22_X1 U23122 ( .A1(n20245), .A2(n20652), .B1(n20453), .B2(n20204), .ZN(
        n20195) );
  INV_X1 U23123 ( .A(n20195), .ZN(n20197) );
  AOI22_X1 U23124 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20207), .B1(
        n20648), .B2(n20206), .ZN(n20196) );
  OAI211_X1 U23125 ( .C1(n20593), .C2(n20210), .A(n20197), .B(n20196), .ZN(
        P1_U3053) );
  OAI22_X1 U23126 ( .A1(n20245), .A2(n20658), .B1(n20457), .B2(n20204), .ZN(
        n20198) );
  INV_X1 U23127 ( .A(n20198), .ZN(n20200) );
  AOI22_X1 U23128 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20207), .B1(
        n20654), .B2(n20206), .ZN(n20199) );
  OAI211_X1 U23129 ( .C1(n20597), .C2(n20210), .A(n20200), .B(n20199), .ZN(
        P1_U3054) );
  OAI22_X1 U23130 ( .A1(n20210), .A2(n20601), .B1(n20461), .B2(n20204), .ZN(
        n20201) );
  INV_X1 U23131 ( .A(n20201), .ZN(n20203) );
  AOI22_X1 U23132 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20207), .B1(
        n20660), .B2(n20206), .ZN(n20202) );
  OAI211_X1 U23133 ( .C1(n20664), .C2(n20245), .A(n20203), .B(n20202), .ZN(
        P1_U3055) );
  OAI22_X1 U23134 ( .A1(n20245), .A2(n20675), .B1(n20465), .B2(n20204), .ZN(
        n20205) );
  INV_X1 U23135 ( .A(n20205), .ZN(n20209) );
  AOI22_X1 U23136 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20207), .B1(
        n20668), .B2(n20206), .ZN(n20208) );
  OAI211_X1 U23137 ( .C1(n20609), .C2(n20210), .A(n20209), .B(n20208), .ZN(
        P1_U3056) );
  INV_X1 U23138 ( .A(n20474), .ZN(n20211) );
  NAND2_X1 U23139 ( .A1(n20211), .A2(n20473), .ZN(n20244) );
  OAI22_X1 U23140 ( .A1(n20245), .A2(n20577), .B1(n20426), .B2(n20244), .ZN(
        n20212) );
  INV_X1 U23141 ( .A(n20212), .ZN(n20225) );
  NOR2_X1 U23142 ( .A1(n20214), .A2(n9591), .ZN(n20611) );
  INV_X1 U23143 ( .A(n20244), .ZN(n20215) );
  AOI21_X1 U23144 ( .B1(n20216), .B2(n20611), .A(n20215), .ZN(n20223) );
  AOI21_X1 U23145 ( .B1(n20218), .B2(n20217), .A(n20622), .ZN(n20220) );
  AOI22_X1 U23146 ( .A1(n20223), .A2(n20220), .B1(n20622), .B2(n20221), .ZN(
        n20219) );
  NAND2_X1 U23147 ( .A1(n20620), .A2(n20219), .ZN(n20248) );
  INV_X1 U23148 ( .A(n20220), .ZN(n20222) );
  OAI22_X1 U23149 ( .A1(n20223), .A2(n20222), .B1(n20613), .B2(n20221), .ZN(
        n20247) );
  AOI22_X1 U23150 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20248), .B1(
        n20616), .B2(n20247), .ZN(n20224) );
  OAI211_X1 U23151 ( .C1(n20628), .C2(n20260), .A(n20225), .B(n20224), .ZN(
        P1_U3057) );
  OAI22_X1 U23152 ( .A1(n20245), .A2(n20581), .B1(n20441), .B2(n20244), .ZN(
        n20226) );
  INV_X1 U23153 ( .A(n20226), .ZN(n20228) );
  AOI22_X1 U23154 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20248), .B1(
        n20630), .B2(n20247), .ZN(n20227) );
  OAI211_X1 U23155 ( .C1(n20634), .C2(n20260), .A(n20228), .B(n20227), .ZN(
        P1_U3058) );
  OAI22_X1 U23156 ( .A1(n20245), .A2(n20585), .B1(n20445), .B2(n20244), .ZN(
        n20229) );
  INV_X1 U23157 ( .A(n20229), .ZN(n20231) );
  AOI22_X1 U23158 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20248), .B1(
        n20636), .B2(n20247), .ZN(n20230) );
  OAI211_X1 U23159 ( .C1(n20640), .C2(n20260), .A(n20231), .B(n20230), .ZN(
        P1_U3059) );
  OAI22_X1 U23160 ( .A1(n20260), .A2(n20646), .B1(n20449), .B2(n20244), .ZN(
        n20232) );
  INV_X1 U23161 ( .A(n20232), .ZN(n20234) );
  AOI22_X1 U23162 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20248), .B1(
        n20642), .B2(n20247), .ZN(n20233) );
  OAI211_X1 U23163 ( .C1(n20589), .C2(n20245), .A(n20234), .B(n20233), .ZN(
        P1_U3060) );
  OAI22_X1 U23164 ( .A1(n20245), .A2(n20593), .B1(n20453), .B2(n20244), .ZN(
        n20235) );
  INV_X1 U23165 ( .A(n20235), .ZN(n20237) );
  AOI22_X1 U23166 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20248), .B1(
        n20648), .B2(n20247), .ZN(n20236) );
  OAI211_X1 U23167 ( .C1(n20652), .C2(n20260), .A(n20237), .B(n20236), .ZN(
        P1_U3061) );
  OAI22_X1 U23168 ( .A1(n20245), .A2(n20597), .B1(n20457), .B2(n20244), .ZN(
        n20238) );
  INV_X1 U23169 ( .A(n20238), .ZN(n20240) );
  AOI22_X1 U23170 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20248), .B1(
        n20654), .B2(n20247), .ZN(n20239) );
  OAI211_X1 U23171 ( .C1(n20658), .C2(n20260), .A(n20240), .B(n20239), .ZN(
        P1_U3062) );
  OAI22_X1 U23172 ( .A1(n20260), .A2(n20664), .B1(n20461), .B2(n20244), .ZN(
        n20241) );
  INV_X1 U23173 ( .A(n20241), .ZN(n20243) );
  AOI22_X1 U23174 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20248), .B1(
        n20660), .B2(n20247), .ZN(n20242) );
  OAI211_X1 U23175 ( .C1(n20601), .C2(n20245), .A(n20243), .B(n20242), .ZN(
        P1_U3063) );
  OAI22_X1 U23176 ( .A1(n20245), .A2(n20609), .B1(n20465), .B2(n20244), .ZN(
        n20246) );
  INV_X1 U23177 ( .A(n20246), .ZN(n20250) );
  AOI22_X1 U23178 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20248), .B1(
        n20668), .B2(n20247), .ZN(n20249) );
  OAI211_X1 U23179 ( .C1(n20675), .C2(n20260), .A(n20250), .B(n20249), .ZN(
        P1_U3064) );
  NOR2_X1 U23180 ( .A1(n12965), .A2(n20251), .ZN(n20345) );
  NAND3_X1 U23181 ( .A1(n20345), .A2(n20624), .A3(n13648), .ZN(n20252) );
  OAI21_X1 U23182 ( .B1(n20565), .B2(n20253), .A(n20252), .ZN(n20276) );
  NAND3_X1 U23183 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20473), .A3(
        n20505), .ZN(n20281) );
  NOR2_X1 U23184 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20281), .ZN(
        n20275) );
  AOI22_X1 U23185 ( .A1(n20616), .A2(n20276), .B1(n20615), .B2(n20275), .ZN(
        n20262) );
  AOI21_X1 U23186 ( .B1(n20260), .B2(n20300), .A(n20254), .ZN(n20255) );
  AOI21_X1 U23187 ( .B1(n20345), .B2(n13648), .A(n20255), .ZN(n20256) );
  NOR2_X1 U23188 ( .A1(n20256), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20259) );
  AOI22_X1 U23189 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20625), .ZN(n20261) );
  OAI211_X1 U23190 ( .C1(n20628), .C2(n20300), .A(n20262), .B(n20261), .ZN(
        P1_U3065) );
  AOI22_X1 U23191 ( .A1(n20630), .A2(n20276), .B1(n20629), .B2(n20275), .ZN(
        n20264) );
  INV_X1 U23192 ( .A(n20581), .ZN(n20631) );
  AOI22_X1 U23193 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20631), .ZN(n20263) );
  OAI211_X1 U23194 ( .C1(n20634), .C2(n20300), .A(n20264), .B(n20263), .ZN(
        P1_U3066) );
  AOI22_X1 U23195 ( .A1(n20636), .A2(n20276), .B1(n20635), .B2(n20275), .ZN(
        n20266) );
  INV_X1 U23196 ( .A(n20585), .ZN(n20637) );
  AOI22_X1 U23197 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20637), .ZN(n20265) );
  OAI211_X1 U23198 ( .C1(n20640), .C2(n20300), .A(n20266), .B(n20265), .ZN(
        P1_U3067) );
  AOI22_X1 U23199 ( .A1(n20642), .A2(n20276), .B1(n20641), .B2(n20275), .ZN(
        n20268) );
  INV_X1 U23200 ( .A(n20589), .ZN(n20643) );
  AOI22_X1 U23201 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20643), .ZN(n20267) );
  OAI211_X1 U23202 ( .C1(n20646), .C2(n20300), .A(n20268), .B(n20267), .ZN(
        P1_U3068) );
  AOI22_X1 U23203 ( .A1(n20648), .A2(n20276), .B1(n20647), .B2(n20275), .ZN(
        n20270) );
  AOI22_X1 U23204 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20649), .ZN(n20269) );
  OAI211_X1 U23205 ( .C1(n20652), .C2(n20300), .A(n20270), .B(n20269), .ZN(
        P1_U3069) );
  AOI22_X1 U23206 ( .A1(n20654), .A2(n20276), .B1(n20653), .B2(n20275), .ZN(
        n20272) );
  INV_X1 U23207 ( .A(n20597), .ZN(n20655) );
  AOI22_X1 U23208 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20655), .ZN(n20271) );
  OAI211_X1 U23209 ( .C1(n20658), .C2(n20300), .A(n20272), .B(n20271), .ZN(
        P1_U3070) );
  AOI22_X1 U23210 ( .A1(n20660), .A2(n20276), .B1(n20659), .B2(n20275), .ZN(
        n20274) );
  INV_X1 U23211 ( .A(n20601), .ZN(n20661) );
  AOI22_X1 U23212 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20661), .ZN(n20273) );
  OAI211_X1 U23213 ( .C1(n20664), .C2(n20300), .A(n20274), .B(n20273), .ZN(
        P1_U3071) );
  AOI22_X1 U23214 ( .A1(n20668), .A2(n20276), .B1(n20665), .B2(n20275), .ZN(
        n20280) );
  INV_X1 U23215 ( .A(n20609), .ZN(n20669) );
  AOI22_X1 U23216 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20278), .B1(
        n20277), .B2(n20669), .ZN(n20279) );
  OAI211_X1 U23217 ( .C1(n20675), .C2(n20300), .A(n20280), .B(n20279), .ZN(
        P1_U3072) );
  NOR2_X1 U23218 ( .A1(n20536), .A2(n20281), .ZN(n20301) );
  AOI21_X1 U23219 ( .B1(n20345), .B2(n20537), .A(n20301), .ZN(n20282) );
  OAI22_X1 U23220 ( .A1(n20282), .A2(n20622), .B1(n20281), .B2(n20613), .ZN(
        n20302) );
  AOI22_X1 U23221 ( .A1(n20616), .A2(n20302), .B1(n20615), .B2(n20301), .ZN(
        n20286) );
  INV_X1 U23222 ( .A(n20281), .ZN(n20284) );
  INV_X1 U23223 ( .A(n20343), .ZN(n20348) );
  OAI21_X1 U23224 ( .B1(n20348), .B2(n20541), .A(n20282), .ZN(n20283) );
  OAI221_X1 U23225 ( .B1(n20624), .B2(n20284), .C1(n20622), .C2(n20283), .A(
        n20620), .ZN(n20304) );
  INV_X1 U23226 ( .A(n20300), .ZN(n20303) );
  AOI22_X1 U23227 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20304), .B1(
        n20303), .B2(n20625), .ZN(n20285) );
  OAI211_X1 U23228 ( .C1(n20628), .C2(n20341), .A(n20286), .B(n20285), .ZN(
        P1_U3073) );
  AOI22_X1 U23229 ( .A1(n20630), .A2(n20302), .B1(n20629), .B2(n20301), .ZN(
        n20288) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20304), .B1(
        n20303), .B2(n20631), .ZN(n20287) );
  OAI211_X1 U23231 ( .C1(n20634), .C2(n20341), .A(n20288), .B(n20287), .ZN(
        P1_U3074) );
  AOI22_X1 U23232 ( .A1(n20636), .A2(n20302), .B1(n20635), .B2(n20301), .ZN(
        n20290) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20304), .B1(
        n20303), .B2(n20637), .ZN(n20289) );
  OAI211_X1 U23234 ( .C1(n20640), .C2(n20341), .A(n20290), .B(n20289), .ZN(
        P1_U3075) );
  AOI22_X1 U23235 ( .A1(n20642), .A2(n20302), .B1(n20641), .B2(n20301), .ZN(
        n20292) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20304), .B1(
        n20303), .B2(n20643), .ZN(n20291) );
  OAI211_X1 U23237 ( .C1(n20646), .C2(n20341), .A(n20292), .B(n20291), .ZN(
        P1_U3076) );
  AOI22_X1 U23238 ( .A1(n20648), .A2(n20302), .B1(n20647), .B2(n20301), .ZN(
        n20294) );
  INV_X1 U23239 ( .A(n20341), .ZN(n20297) );
  INV_X1 U23240 ( .A(n20652), .ZN(n20590) );
  AOI22_X1 U23241 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20304), .B1(
        n20297), .B2(n20590), .ZN(n20293) );
  OAI211_X1 U23242 ( .C1(n20593), .C2(n20300), .A(n20294), .B(n20293), .ZN(
        P1_U3077) );
  AOI22_X1 U23243 ( .A1(n20654), .A2(n20302), .B1(n20653), .B2(n20301), .ZN(
        n20296) );
  AOI22_X1 U23244 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20304), .B1(
        n20297), .B2(n20594), .ZN(n20295) );
  OAI211_X1 U23245 ( .C1(n20597), .C2(n20300), .A(n20296), .B(n20295), .ZN(
        P1_U3078) );
  AOI22_X1 U23246 ( .A1(n20660), .A2(n20302), .B1(n20659), .B2(n20301), .ZN(
        n20299) );
  AOI22_X1 U23247 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20304), .B1(
        n20297), .B2(n20598), .ZN(n20298) );
  OAI211_X1 U23248 ( .C1(n20601), .C2(n20300), .A(n20299), .B(n20298), .ZN(
        P1_U3079) );
  AOI22_X1 U23249 ( .A1(n20668), .A2(n20302), .B1(n20665), .B2(n20301), .ZN(
        n20306) );
  AOI22_X1 U23250 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20304), .B1(
        n20303), .B2(n20669), .ZN(n20305) );
  OAI211_X1 U23251 ( .C1(n20675), .C2(n20341), .A(n20306), .B(n20305), .ZN(
        P1_U3080) );
  INV_X1 U23252 ( .A(n20349), .ZN(n20346) );
  OR2_X1 U23253 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20346), .ZN(
        n20335) );
  OAI22_X1 U23254 ( .A1(n20372), .A2(n20628), .B1(n20426), .B2(n20335), .ZN(
        n20307) );
  INV_X1 U23255 ( .A(n20307), .ZN(n20316) );
  NAND3_X1 U23256 ( .A1(n20372), .A2(n20341), .A3(n20624), .ZN(n20308) );
  NAND2_X1 U23257 ( .A1(n20308), .A2(n20507), .ZN(n20311) );
  NAND2_X1 U23258 ( .A1(n20345), .A2(n20564), .ZN(n20313) );
  AOI22_X1 U23259 ( .A1(n20311), .A2(n20313), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20335), .ZN(n20310) );
  NAND3_X1 U23260 ( .A1(n20572), .A2(n20310), .A3(n20309), .ZN(n20338) );
  INV_X1 U23261 ( .A(n20311), .ZN(n20314) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20338), .B1(
        n20616), .B2(n20337), .ZN(n20315) );
  OAI211_X1 U23263 ( .C1(n20577), .C2(n20341), .A(n20316), .B(n20315), .ZN(
        P1_U3081) );
  OAI22_X1 U23264 ( .A1(n20341), .A2(n20581), .B1(n20441), .B2(n20335), .ZN(
        n20317) );
  INV_X1 U23265 ( .A(n20317), .ZN(n20319) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20338), .B1(
        n20630), .B2(n20337), .ZN(n20318) );
  OAI211_X1 U23267 ( .C1(n20634), .C2(n20372), .A(n20319), .B(n20318), .ZN(
        P1_U3082) );
  OAI22_X1 U23268 ( .A1(n20372), .A2(n20640), .B1(n20335), .B2(n20445), .ZN(
        n20320) );
  INV_X1 U23269 ( .A(n20320), .ZN(n20322) );
  AOI22_X1 U23270 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20338), .B1(
        n20636), .B2(n20337), .ZN(n20321) );
  OAI211_X1 U23271 ( .C1(n20585), .C2(n20341), .A(n20322), .B(n20321), .ZN(
        P1_U3083) );
  OAI22_X1 U23272 ( .A1(n20372), .A2(n20646), .B1(n20335), .B2(n20449), .ZN(
        n20323) );
  INV_X1 U23273 ( .A(n20323), .ZN(n20325) );
  AOI22_X1 U23274 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20338), .B1(
        n20642), .B2(n20337), .ZN(n20324) );
  OAI211_X1 U23275 ( .C1(n20589), .C2(n20341), .A(n20325), .B(n20324), .ZN(
        P1_U3084) );
  OAI22_X1 U23276 ( .A1(n20372), .A2(n20652), .B1(n20335), .B2(n20453), .ZN(
        n20326) );
  INV_X1 U23277 ( .A(n20326), .ZN(n20328) );
  AOI22_X1 U23278 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20338), .B1(
        n20648), .B2(n20337), .ZN(n20327) );
  OAI211_X1 U23279 ( .C1(n20593), .C2(n20341), .A(n20328), .B(n20327), .ZN(
        P1_U3085) );
  OAI22_X1 U23280 ( .A1(n20341), .A2(n20597), .B1(n20457), .B2(n20335), .ZN(
        n20329) );
  INV_X1 U23281 ( .A(n20329), .ZN(n20331) );
  AOI22_X1 U23282 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20338), .B1(
        n20654), .B2(n20337), .ZN(n20330) );
  OAI211_X1 U23283 ( .C1(n20658), .C2(n20372), .A(n20331), .B(n20330), .ZN(
        P1_U3086) );
  OAI22_X1 U23284 ( .A1(n20372), .A2(n20664), .B1(n20335), .B2(n20461), .ZN(
        n20332) );
  INV_X1 U23285 ( .A(n20332), .ZN(n20334) );
  AOI22_X1 U23286 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20338), .B1(
        n20660), .B2(n20337), .ZN(n20333) );
  OAI211_X1 U23287 ( .C1(n20601), .C2(n20341), .A(n20334), .B(n20333), .ZN(
        P1_U3087) );
  OAI22_X1 U23288 ( .A1(n20372), .A2(n20675), .B1(n20465), .B2(n20335), .ZN(
        n20336) );
  INV_X1 U23289 ( .A(n20336), .ZN(n20340) );
  AOI22_X1 U23290 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20338), .B1(
        n20668), .B2(n20337), .ZN(n20339) );
  OAI211_X1 U23291 ( .C1(n20609), .C2(n20341), .A(n20340), .B(n20339), .ZN(
        P1_U3088) );
  INV_X1 U23292 ( .A(n20344), .ZN(n20367) );
  AOI21_X1 U23293 ( .B1(n20345), .B2(n20611), .A(n20367), .ZN(n20347) );
  OAI22_X1 U23294 ( .A1(n20347), .A2(n20622), .B1(n20346), .B2(n20613), .ZN(
        n20368) );
  AOI22_X1 U23295 ( .A1(n20616), .A2(n20368), .B1(n20367), .B2(n20615), .ZN(
        n20352) );
  NOR3_X1 U23296 ( .A1(n20348), .A2(n20622), .A3(n20618), .ZN(n20350) );
  OAI21_X1 U23297 ( .B1(n20350), .B2(n20349), .A(n20620), .ZN(n20369) );
  INV_X1 U23298 ( .A(n20372), .ZN(n20363) );
  AOI22_X1 U23299 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20369), .B1(
        n20363), .B2(n20625), .ZN(n20351) );
  OAI211_X1 U23300 ( .C1(n20628), .C2(n20366), .A(n20352), .B(n20351), .ZN(
        P1_U3089) );
  AOI22_X1 U23301 ( .A1(n20630), .A2(n20368), .B1(n20367), .B2(n20629), .ZN(
        n20354) );
  AOI22_X1 U23302 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20369), .B1(
        n20395), .B2(n20578), .ZN(n20353) );
  OAI211_X1 U23303 ( .C1(n20581), .C2(n20372), .A(n20354), .B(n20353), .ZN(
        P1_U3090) );
  AOI22_X1 U23304 ( .A1(n20636), .A2(n20368), .B1(n20367), .B2(n20635), .ZN(
        n20356) );
  AOI22_X1 U23305 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20369), .B1(
        n20363), .B2(n20637), .ZN(n20355) );
  OAI211_X1 U23306 ( .C1(n20640), .C2(n20366), .A(n20356), .B(n20355), .ZN(
        P1_U3091) );
  AOI22_X1 U23307 ( .A1(n20642), .A2(n20368), .B1(n20367), .B2(n20641), .ZN(
        n20358) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20369), .B1(
        n20395), .B2(n20586), .ZN(n20357) );
  OAI211_X1 U23309 ( .C1(n20589), .C2(n20372), .A(n20358), .B(n20357), .ZN(
        P1_U3092) );
  AOI22_X1 U23310 ( .A1(n20648), .A2(n20368), .B1(n20367), .B2(n20647), .ZN(
        n20360) );
  AOI22_X1 U23311 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20369), .B1(
        n20363), .B2(n20649), .ZN(n20359) );
  OAI211_X1 U23312 ( .C1(n20652), .C2(n20366), .A(n20360), .B(n20359), .ZN(
        P1_U3093) );
  AOI22_X1 U23313 ( .A1(n20654), .A2(n20368), .B1(n20367), .B2(n20653), .ZN(
        n20362) );
  AOI22_X1 U23314 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20369), .B1(
        n20363), .B2(n20655), .ZN(n20361) );
  OAI211_X1 U23315 ( .C1(n20658), .C2(n20366), .A(n20362), .B(n20361), .ZN(
        P1_U3094) );
  AOI22_X1 U23316 ( .A1(n20660), .A2(n20368), .B1(n20367), .B2(n20659), .ZN(
        n20365) );
  AOI22_X1 U23317 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20369), .B1(
        n20363), .B2(n20661), .ZN(n20364) );
  OAI211_X1 U23318 ( .C1(n20664), .C2(n20366), .A(n20365), .B(n20364), .ZN(
        P1_U3095) );
  AOI22_X1 U23319 ( .A1(n20668), .A2(n20368), .B1(n20367), .B2(n20665), .ZN(
        n20371) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20369), .B1(
        n20395), .B2(n20604), .ZN(n20370) );
  OAI211_X1 U23321 ( .C1(n20609), .C2(n20372), .A(n20371), .B(n20370), .ZN(
        P1_U3096) );
  INV_X1 U23322 ( .A(n20481), .ZN(n20373) );
  AND2_X1 U23323 ( .A1(n9603), .A2(n12965), .ZN(n20475) );
  NAND3_X1 U23324 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20425), .A3(
        n20505), .ZN(n20399) );
  NOR2_X1 U23325 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20399), .ZN(
        n20393) );
  AOI21_X1 U23326 ( .B1(n20475), .B2(n13648), .A(n20393), .ZN(n20376) );
  NAND2_X1 U23327 ( .A1(n20374), .A2(n20430), .ZN(n20512) );
  OAI22_X1 U23328 ( .A1(n20376), .A2(n20622), .B1(n20436), .B2(n20512), .ZN(
        n20394) );
  AOI22_X1 U23329 ( .A1(n20616), .A2(n20394), .B1(n20615), .B2(n20393), .ZN(
        n20380) );
  INV_X1 U23330 ( .A(n20423), .ZN(n20375) );
  OAI21_X1 U23331 ( .B1(n20375), .B2(n20395), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20377) );
  NAND2_X1 U23332 ( .A1(n20377), .A2(n20376), .ZN(n20378) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20625), .ZN(n20379) );
  OAI211_X1 U23334 ( .C1(n20628), .C2(n20423), .A(n20380), .B(n20379), .ZN(
        P1_U3097) );
  AOI22_X1 U23335 ( .A1(n20630), .A2(n20394), .B1(n20629), .B2(n20393), .ZN(
        n20382) );
  AOI22_X1 U23336 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20631), .ZN(n20381) );
  OAI211_X1 U23337 ( .C1(n20634), .C2(n20423), .A(n20382), .B(n20381), .ZN(
        P1_U3098) );
  AOI22_X1 U23338 ( .A1(n20636), .A2(n20394), .B1(n20635), .B2(n20393), .ZN(
        n20384) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20637), .ZN(n20383) );
  OAI211_X1 U23340 ( .C1(n20640), .C2(n20423), .A(n20384), .B(n20383), .ZN(
        P1_U3099) );
  AOI22_X1 U23341 ( .A1(n20642), .A2(n20394), .B1(n20641), .B2(n20393), .ZN(
        n20386) );
  AOI22_X1 U23342 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20643), .ZN(n20385) );
  OAI211_X1 U23343 ( .C1(n20646), .C2(n20423), .A(n20386), .B(n20385), .ZN(
        P1_U3100) );
  AOI22_X1 U23344 ( .A1(n20648), .A2(n20394), .B1(n20647), .B2(n20393), .ZN(
        n20388) );
  AOI22_X1 U23345 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20649), .ZN(n20387) );
  OAI211_X1 U23346 ( .C1(n20652), .C2(n20423), .A(n20388), .B(n20387), .ZN(
        P1_U3101) );
  AOI22_X1 U23347 ( .A1(n20654), .A2(n20394), .B1(n20653), .B2(n20393), .ZN(
        n20390) );
  AOI22_X1 U23348 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20655), .ZN(n20389) );
  OAI211_X1 U23349 ( .C1(n20658), .C2(n20423), .A(n20390), .B(n20389), .ZN(
        P1_U3102) );
  AOI22_X1 U23350 ( .A1(n20660), .A2(n20394), .B1(n20659), .B2(n20393), .ZN(
        n20392) );
  AOI22_X1 U23351 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20661), .ZN(n20391) );
  OAI211_X1 U23352 ( .C1(n20664), .C2(n20423), .A(n20392), .B(n20391), .ZN(
        P1_U3103) );
  AOI22_X1 U23353 ( .A1(n20668), .A2(n20394), .B1(n20665), .B2(n20393), .ZN(
        n20398) );
  AOI22_X1 U23354 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20669), .ZN(n20397) );
  OAI211_X1 U23355 ( .C1(n20675), .C2(n20423), .A(n20398), .B(n20397), .ZN(
        P1_U3104) );
  NOR2_X1 U23356 ( .A1(n20536), .A2(n20399), .ZN(n20418) );
  AOI21_X1 U23357 ( .B1(n20475), .B2(n20537), .A(n20418), .ZN(n20400) );
  OAI22_X1 U23358 ( .A1(n20400), .A2(n20622), .B1(n20399), .B2(n20613), .ZN(
        n20419) );
  AOI22_X1 U23359 ( .A1(n20616), .A2(n20419), .B1(n20615), .B2(n20418), .ZN(
        n20405) );
  INV_X1 U23360 ( .A(n20399), .ZN(n20402) );
  OAI21_X1 U23361 ( .B1(n20481), .B2(n20541), .A(n20400), .ZN(n20401) );
  OAI221_X1 U23362 ( .B1(n20624), .B2(n20402), .C1(n20622), .C2(n20401), .A(
        n20620), .ZN(n20420) );
  INV_X1 U23363 ( .A(n20535), .ZN(n20403) );
  INV_X1 U23364 ( .A(n20628), .ZN(n20574) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20420), .B1(
        n20428), .B2(n20574), .ZN(n20404) );
  OAI211_X1 U23366 ( .C1(n20577), .C2(n20423), .A(n20405), .B(n20404), .ZN(
        P1_U3105) );
  AOI22_X1 U23367 ( .A1(n20630), .A2(n20419), .B1(n20629), .B2(n20418), .ZN(
        n20407) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20420), .B1(
        n20428), .B2(n20578), .ZN(n20406) );
  OAI211_X1 U23369 ( .C1(n20581), .C2(n20423), .A(n20407), .B(n20406), .ZN(
        P1_U3106) );
  AOI22_X1 U23370 ( .A1(n20636), .A2(n20419), .B1(n20635), .B2(n20418), .ZN(
        n20409) );
  AOI22_X1 U23371 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20420), .B1(
        n20428), .B2(n20582), .ZN(n20408) );
  OAI211_X1 U23372 ( .C1(n20585), .C2(n20423), .A(n20409), .B(n20408), .ZN(
        P1_U3107) );
  AOI22_X1 U23373 ( .A1(n20642), .A2(n20419), .B1(n20641), .B2(n20418), .ZN(
        n20411) );
  AOI22_X1 U23374 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20420), .B1(
        n20428), .B2(n20586), .ZN(n20410) );
  OAI211_X1 U23375 ( .C1(n20589), .C2(n20423), .A(n20411), .B(n20410), .ZN(
        P1_U3108) );
  AOI22_X1 U23376 ( .A1(n20648), .A2(n20419), .B1(n20647), .B2(n20418), .ZN(
        n20413) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20420), .B1(
        n20428), .B2(n20590), .ZN(n20412) );
  OAI211_X1 U23378 ( .C1(n20593), .C2(n20423), .A(n20413), .B(n20412), .ZN(
        P1_U3109) );
  AOI22_X1 U23379 ( .A1(n20654), .A2(n20419), .B1(n20653), .B2(n20418), .ZN(
        n20415) );
  AOI22_X1 U23380 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20420), .B1(
        n20428), .B2(n20594), .ZN(n20414) );
  OAI211_X1 U23381 ( .C1(n20597), .C2(n20423), .A(n20415), .B(n20414), .ZN(
        P1_U3110) );
  AOI22_X1 U23382 ( .A1(n20660), .A2(n20419), .B1(n20659), .B2(n20418), .ZN(
        n20417) );
  AOI22_X1 U23383 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20420), .B1(
        n20428), .B2(n20598), .ZN(n20416) );
  OAI211_X1 U23384 ( .C1(n20601), .C2(n20423), .A(n20417), .B(n20416), .ZN(
        P1_U3111) );
  AOI22_X1 U23385 ( .A1(n20668), .A2(n20419), .B1(n20665), .B2(n20418), .ZN(
        n20422) );
  AOI22_X1 U23386 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20420), .B1(
        n20428), .B2(n20604), .ZN(n20421) );
  OAI211_X1 U23387 ( .C1(n20609), .C2(n20423), .A(n20422), .B(n20421), .ZN(
        P1_U3112) );
  NAND3_X1 U23388 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20425), .ZN(n20476) );
  NOR2_X1 U23389 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20476), .ZN(
        n20431) );
  INV_X1 U23390 ( .A(n20431), .ZN(n20466) );
  OAI22_X1 U23391 ( .A1(n20467), .A2(n20577), .B1(n20466), .B2(n20426), .ZN(
        n20427) );
  INV_X1 U23392 ( .A(n20427), .ZN(n20440) );
  OAI21_X1 U23393 ( .B1(n20494), .B2(n20428), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20429) );
  NAND2_X1 U23394 ( .A1(n20429), .A2(n20624), .ZN(n20438) );
  AND2_X1 U23395 ( .A1(n20475), .A2(n20564), .ZN(n20435) );
  OR2_X1 U23396 ( .A1(n20430), .A2(n20473), .ZN(n20566) );
  NAND2_X1 U23397 ( .A1(n20566), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20571) );
  OAI21_X1 U23398 ( .B1(n20510), .B2(n20431), .A(n20571), .ZN(n20432) );
  INV_X1 U23399 ( .A(n20432), .ZN(n20434) );
  INV_X1 U23400 ( .A(n20435), .ZN(n20437) );
  AOI22_X1 U23401 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20470), .B1(
        n20616), .B2(n20469), .ZN(n20439) );
  OAI211_X1 U23402 ( .C1(n20628), .C2(n20503), .A(n20440), .B(n20439), .ZN(
        P1_U3113) );
  OAI22_X1 U23403 ( .A1(n20503), .A2(n20634), .B1(n20441), .B2(n20466), .ZN(
        n20442) );
  INV_X1 U23404 ( .A(n20442), .ZN(n20444) );
  AOI22_X1 U23405 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20470), .B1(
        n20630), .B2(n20469), .ZN(n20443) );
  OAI211_X1 U23406 ( .C1(n20581), .C2(n20467), .A(n20444), .B(n20443), .ZN(
        P1_U3114) );
  OAI22_X1 U23407 ( .A1(n20503), .A2(n20640), .B1(n20466), .B2(n20445), .ZN(
        n20446) );
  INV_X1 U23408 ( .A(n20446), .ZN(n20448) );
  AOI22_X1 U23409 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20470), .B1(
        n20636), .B2(n20469), .ZN(n20447) );
  OAI211_X1 U23410 ( .C1(n20585), .C2(n20467), .A(n20448), .B(n20447), .ZN(
        P1_U3115) );
  OAI22_X1 U23411 ( .A1(n20503), .A2(n20646), .B1(n20466), .B2(n20449), .ZN(
        n20450) );
  INV_X1 U23412 ( .A(n20450), .ZN(n20452) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20470), .B1(
        n20642), .B2(n20469), .ZN(n20451) );
  OAI211_X1 U23414 ( .C1(n20589), .C2(n20467), .A(n20452), .B(n20451), .ZN(
        P1_U3116) );
  OAI22_X1 U23415 ( .A1(n20503), .A2(n20652), .B1(n20466), .B2(n20453), .ZN(
        n20454) );
  INV_X1 U23416 ( .A(n20454), .ZN(n20456) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20470), .B1(
        n20648), .B2(n20469), .ZN(n20455) );
  OAI211_X1 U23418 ( .C1(n20593), .C2(n20467), .A(n20456), .B(n20455), .ZN(
        P1_U3117) );
  OAI22_X1 U23419 ( .A1(n20503), .A2(n20658), .B1(n20466), .B2(n20457), .ZN(
        n20458) );
  INV_X1 U23420 ( .A(n20458), .ZN(n20460) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20470), .B1(
        n20654), .B2(n20469), .ZN(n20459) );
  OAI211_X1 U23422 ( .C1(n20597), .C2(n20467), .A(n20460), .B(n20459), .ZN(
        P1_U3118) );
  OAI22_X1 U23423 ( .A1(n20503), .A2(n20664), .B1(n20466), .B2(n20461), .ZN(
        n20462) );
  INV_X1 U23424 ( .A(n20462), .ZN(n20464) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20470), .B1(
        n20660), .B2(n20469), .ZN(n20463) );
  OAI211_X1 U23426 ( .C1(n20601), .C2(n20467), .A(n20464), .B(n20463), .ZN(
        P1_U3119) );
  OAI22_X1 U23427 ( .A1(n20467), .A2(n20609), .B1(n20466), .B2(n20465), .ZN(
        n20468) );
  INV_X1 U23428 ( .A(n20468), .ZN(n20472) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20470), .B1(
        n20668), .B2(n20469), .ZN(n20471) );
  OAI211_X1 U23430 ( .C1(n20675), .C2(n20503), .A(n20472), .B(n20471), .ZN(
        P1_U3120) );
  NOR2_X1 U23431 ( .A1(n20474), .A2(n20473), .ZN(n20497) );
  AOI21_X1 U23432 ( .B1(n20475), .B2(n20611), .A(n20497), .ZN(n20477) );
  OAI22_X1 U23433 ( .A1(n20477), .A2(n20622), .B1(n20476), .B2(n20613), .ZN(
        n20498) );
  AOI22_X1 U23434 ( .A1(n20616), .A2(n20498), .B1(n20615), .B2(n20497), .ZN(
        n20483) );
  INV_X1 U23435 ( .A(n20476), .ZN(n20479) );
  OAI21_X1 U23436 ( .B1(n20481), .B2(n20618), .A(n20477), .ZN(n20478) );
  OAI221_X1 U23437 ( .B1(n20624), .B2(n20479), .C1(n20622), .C2(n20478), .A(
        n20620), .ZN(n20500) );
  INV_X1 U23438 ( .A(n20534), .ZN(n20499) );
  AOI22_X1 U23439 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20500), .B1(
        n20499), .B2(n20574), .ZN(n20482) );
  OAI211_X1 U23440 ( .C1(n20577), .C2(n20503), .A(n20483), .B(n20482), .ZN(
        P1_U3121) );
  AOI22_X1 U23441 ( .A1(n20630), .A2(n20498), .B1(n20629), .B2(n20497), .ZN(
        n20485) );
  AOI22_X1 U23442 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20500), .B1(
        n20499), .B2(n20578), .ZN(n20484) );
  OAI211_X1 U23443 ( .C1(n20581), .C2(n20503), .A(n20485), .B(n20484), .ZN(
        P1_U3122) );
  AOI22_X1 U23444 ( .A1(n20636), .A2(n20498), .B1(n20635), .B2(n20497), .ZN(
        n20487) );
  AOI22_X1 U23445 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20500), .B1(
        n20494), .B2(n20637), .ZN(n20486) );
  OAI211_X1 U23446 ( .C1(n20640), .C2(n20534), .A(n20487), .B(n20486), .ZN(
        P1_U3123) );
  AOI22_X1 U23447 ( .A1(n20642), .A2(n20498), .B1(n20641), .B2(n20497), .ZN(
        n20489) );
  AOI22_X1 U23448 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20500), .B1(
        n20494), .B2(n20643), .ZN(n20488) );
  OAI211_X1 U23449 ( .C1(n20646), .C2(n20534), .A(n20489), .B(n20488), .ZN(
        P1_U3124) );
  AOI22_X1 U23450 ( .A1(n20648), .A2(n20498), .B1(n20647), .B2(n20497), .ZN(
        n20491) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20500), .B1(
        n20499), .B2(n20590), .ZN(n20490) );
  OAI211_X1 U23452 ( .C1(n20593), .C2(n20503), .A(n20491), .B(n20490), .ZN(
        P1_U3125) );
  AOI22_X1 U23453 ( .A1(n20654), .A2(n20498), .B1(n20653), .B2(n20497), .ZN(
        n20493) );
  AOI22_X1 U23454 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20500), .B1(
        n20494), .B2(n20655), .ZN(n20492) );
  OAI211_X1 U23455 ( .C1(n20658), .C2(n20534), .A(n20493), .B(n20492), .ZN(
        P1_U3126) );
  AOI22_X1 U23456 ( .A1(n20660), .A2(n20498), .B1(n20659), .B2(n20497), .ZN(
        n20496) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20500), .B1(
        n20494), .B2(n20661), .ZN(n20495) );
  OAI211_X1 U23458 ( .C1(n20664), .C2(n20534), .A(n20496), .B(n20495), .ZN(
        P1_U3127) );
  AOI22_X1 U23459 ( .A1(n20668), .A2(n20498), .B1(n20665), .B2(n20497), .ZN(
        n20502) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20500), .B1(
        n20499), .B2(n20604), .ZN(n20501) );
  OAI211_X1 U23461 ( .C1(n20609), .C2(n20503), .A(n20502), .B(n20501), .ZN(
        P1_U3128) );
  NAND3_X1 U23462 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20505), .ZN(n20538) );
  NOR2_X1 U23463 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20538), .ZN(
        n20529) );
  AOI22_X1 U23464 ( .A1(n20560), .A2(n20574), .B1(n20615), .B2(n20529), .ZN(
        n20516) );
  INV_X1 U23465 ( .A(n20560), .ZN(n20506) );
  NAND3_X1 U23466 ( .A1(n20506), .A2(n20624), .A3(n20534), .ZN(n20508) );
  NAND2_X1 U23467 ( .A1(n20508), .A2(n20507), .ZN(n20511) );
  NOR2_X1 U23468 ( .A1(n12965), .A2(n9846), .ZN(n20612) );
  NAND2_X1 U23469 ( .A1(n20612), .A2(n13648), .ZN(n20513) );
  AOI22_X1 U23470 ( .A1(n20511), .A2(n20513), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20512), .ZN(n20509) );
  OAI211_X1 U23471 ( .C1(n20529), .C2(n20510), .A(n20572), .B(n20509), .ZN(
        n20531) );
  INV_X1 U23472 ( .A(n20511), .ZN(n20514) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20531), .B1(
        n20616), .B2(n20530), .ZN(n20515) );
  OAI211_X1 U23474 ( .C1(n20577), .C2(n20534), .A(n20516), .B(n20515), .ZN(
        P1_U3129) );
  AOI22_X1 U23475 ( .A1(n20560), .A2(n20578), .B1(n20629), .B2(n20529), .ZN(
        n20518) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20531), .B1(
        n20630), .B2(n20530), .ZN(n20517) );
  OAI211_X1 U23477 ( .C1(n20581), .C2(n20534), .A(n20518), .B(n20517), .ZN(
        P1_U3130) );
  AOI22_X1 U23478 ( .A1(n20560), .A2(n20582), .B1(n20635), .B2(n20529), .ZN(
        n20520) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20531), .B1(
        n20636), .B2(n20530), .ZN(n20519) );
  OAI211_X1 U23480 ( .C1(n20585), .C2(n20534), .A(n20520), .B(n20519), .ZN(
        P1_U3131) );
  AOI22_X1 U23481 ( .A1(n20560), .A2(n20586), .B1(n20641), .B2(n20529), .ZN(
        n20522) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20531), .B1(
        n20642), .B2(n20530), .ZN(n20521) );
  OAI211_X1 U23483 ( .C1(n20589), .C2(n20534), .A(n20522), .B(n20521), .ZN(
        P1_U3132) );
  AOI22_X1 U23484 ( .A1(n20560), .A2(n20590), .B1(n20647), .B2(n20529), .ZN(
        n20524) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20531), .B1(
        n20648), .B2(n20530), .ZN(n20523) );
  OAI211_X1 U23486 ( .C1(n20593), .C2(n20534), .A(n20524), .B(n20523), .ZN(
        P1_U3133) );
  AOI22_X1 U23487 ( .A1(n20560), .A2(n20594), .B1(n20653), .B2(n20529), .ZN(
        n20526) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20531), .B1(
        n20654), .B2(n20530), .ZN(n20525) );
  OAI211_X1 U23489 ( .C1(n20597), .C2(n20534), .A(n20526), .B(n20525), .ZN(
        P1_U3134) );
  AOI22_X1 U23490 ( .A1(n20560), .A2(n20598), .B1(n20659), .B2(n20529), .ZN(
        n20528) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20531), .B1(
        n20660), .B2(n20530), .ZN(n20527) );
  OAI211_X1 U23492 ( .C1(n20601), .C2(n20534), .A(n20528), .B(n20527), .ZN(
        P1_U3135) );
  AOI22_X1 U23493 ( .A1(n20560), .A2(n20604), .B1(n20665), .B2(n20529), .ZN(
        n20533) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20531), .B1(
        n20668), .B2(n20530), .ZN(n20532) );
  OAI211_X1 U23495 ( .C1(n20609), .C2(n20534), .A(n20533), .B(n20532), .ZN(
        P1_U3136) );
  NOR2_X1 U23496 ( .A1(n20536), .A2(n20538), .ZN(n20558) );
  AOI21_X1 U23497 ( .B1(n20612), .B2(n20537), .A(n20558), .ZN(n20540) );
  OAI22_X1 U23498 ( .A1(n20540), .A2(n20622), .B1(n20538), .B2(n20613), .ZN(
        n20559) );
  AOI22_X1 U23499 ( .A1(n20616), .A2(n20559), .B1(n20615), .B2(n20558), .ZN(
        n20545) );
  INV_X1 U23500 ( .A(n20538), .ZN(n20543) );
  INV_X1 U23501 ( .A(n20539), .ZN(n20619) );
  OAI21_X1 U23502 ( .B1(n20619), .B2(n20541), .A(n20540), .ZN(n20542) );
  OAI221_X1 U23503 ( .B1(n20624), .B2(n20543), .C1(n20622), .C2(n20542), .A(
        n20620), .ZN(n20561) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20561), .B1(
        n20560), .B2(n20625), .ZN(n20544) );
  OAI211_X1 U23505 ( .C1(n20628), .C2(n20608), .A(n20545), .B(n20544), .ZN(
        P1_U3137) );
  AOI22_X1 U23506 ( .A1(n20630), .A2(n20559), .B1(n20629), .B2(n20558), .ZN(
        n20547) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20561), .B1(
        n20560), .B2(n20631), .ZN(n20546) );
  OAI211_X1 U23508 ( .C1(n20634), .C2(n20608), .A(n20547), .B(n20546), .ZN(
        P1_U3138) );
  AOI22_X1 U23509 ( .A1(n20636), .A2(n20559), .B1(n20635), .B2(n20558), .ZN(
        n20549) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20561), .B1(
        n20560), .B2(n20637), .ZN(n20548) );
  OAI211_X1 U23511 ( .C1(n20640), .C2(n20608), .A(n20549), .B(n20548), .ZN(
        P1_U3139) );
  AOI22_X1 U23512 ( .A1(n20642), .A2(n20559), .B1(n20641), .B2(n20558), .ZN(
        n20551) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20561), .B1(
        n20560), .B2(n20643), .ZN(n20550) );
  OAI211_X1 U23514 ( .C1(n20646), .C2(n20608), .A(n20551), .B(n20550), .ZN(
        P1_U3140) );
  AOI22_X1 U23515 ( .A1(n20648), .A2(n20559), .B1(n20647), .B2(n20558), .ZN(
        n20553) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20561), .B1(
        n20560), .B2(n20649), .ZN(n20552) );
  OAI211_X1 U23517 ( .C1(n20652), .C2(n20608), .A(n20553), .B(n20552), .ZN(
        P1_U3141) );
  AOI22_X1 U23518 ( .A1(n20654), .A2(n20559), .B1(n20653), .B2(n20558), .ZN(
        n20555) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20561), .B1(
        n20560), .B2(n20655), .ZN(n20554) );
  OAI211_X1 U23520 ( .C1(n20658), .C2(n20608), .A(n20555), .B(n20554), .ZN(
        P1_U3142) );
  AOI22_X1 U23521 ( .A1(n20660), .A2(n20559), .B1(n20659), .B2(n20558), .ZN(
        n20557) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20561), .B1(
        n20560), .B2(n20661), .ZN(n20556) );
  OAI211_X1 U23523 ( .C1(n20664), .C2(n20608), .A(n20557), .B(n20556), .ZN(
        P1_U3143) );
  AOI22_X1 U23524 ( .A1(n20668), .A2(n20559), .B1(n20665), .B2(n20558), .ZN(
        n20563) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20561), .B1(
        n20560), .B2(n20669), .ZN(n20562) );
  OAI211_X1 U23526 ( .C1(n20675), .C2(n20608), .A(n20563), .B(n20562), .ZN(
        P1_U3144) );
  NAND2_X1 U23527 ( .A1(n20612), .A2(n20564), .ZN(n20569) );
  OAI22_X1 U23528 ( .A1(n20569), .A2(n20622), .B1(n20566), .B2(n20565), .ZN(
        n20603) );
  NOR2_X1 U23529 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20614), .ZN(
        n20602) );
  AOI22_X1 U23530 ( .A1(n20616), .A2(n20603), .B1(n20615), .B2(n20602), .ZN(
        n20576) );
  INV_X1 U23531 ( .A(n20608), .ZN(n20568) );
  OAI21_X1 U23532 ( .B1(n20670), .B2(n20568), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20570) );
  AOI21_X1 U23533 ( .B1(n20570), .B2(n20569), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20573) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20605), .B1(
        n20670), .B2(n20574), .ZN(n20575) );
  OAI211_X1 U23535 ( .C1(n20577), .C2(n20608), .A(n20576), .B(n20575), .ZN(
        P1_U3145) );
  AOI22_X1 U23536 ( .A1(n20630), .A2(n20603), .B1(n20629), .B2(n20602), .ZN(
        n20580) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20605), .B1(
        n20670), .B2(n20578), .ZN(n20579) );
  OAI211_X1 U23538 ( .C1(n20581), .C2(n20608), .A(n20580), .B(n20579), .ZN(
        P1_U3146) );
  AOI22_X1 U23539 ( .A1(n20636), .A2(n20603), .B1(n20635), .B2(n20602), .ZN(
        n20584) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20605), .B1(
        n20670), .B2(n20582), .ZN(n20583) );
  OAI211_X1 U23541 ( .C1(n20585), .C2(n20608), .A(n20584), .B(n20583), .ZN(
        P1_U3147) );
  AOI22_X1 U23542 ( .A1(n20642), .A2(n20603), .B1(n20641), .B2(n20602), .ZN(
        n20588) );
  AOI22_X1 U23543 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20605), .B1(
        n20670), .B2(n20586), .ZN(n20587) );
  OAI211_X1 U23544 ( .C1(n20589), .C2(n20608), .A(n20588), .B(n20587), .ZN(
        P1_U3148) );
  AOI22_X1 U23545 ( .A1(n20648), .A2(n20603), .B1(n20647), .B2(n20602), .ZN(
        n20592) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20605), .B1(
        n20670), .B2(n20590), .ZN(n20591) );
  OAI211_X1 U23547 ( .C1(n20593), .C2(n20608), .A(n20592), .B(n20591), .ZN(
        P1_U3149) );
  AOI22_X1 U23548 ( .A1(n20654), .A2(n20603), .B1(n20653), .B2(n20602), .ZN(
        n20596) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20605), .B1(
        n20670), .B2(n20594), .ZN(n20595) );
  OAI211_X1 U23550 ( .C1(n20597), .C2(n20608), .A(n20596), .B(n20595), .ZN(
        P1_U3150) );
  AOI22_X1 U23551 ( .A1(n20660), .A2(n20603), .B1(n20659), .B2(n20602), .ZN(
        n20600) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20605), .B1(
        n20670), .B2(n20598), .ZN(n20599) );
  OAI211_X1 U23553 ( .C1(n20601), .C2(n20608), .A(n20600), .B(n20599), .ZN(
        P1_U3151) );
  AOI22_X1 U23554 ( .A1(n20668), .A2(n20603), .B1(n20665), .B2(n20602), .ZN(
        n20607) );
  AOI22_X1 U23555 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20605), .B1(
        n20670), .B2(n20604), .ZN(n20606) );
  OAI211_X1 U23556 ( .C1(n20609), .C2(n20608), .A(n20607), .B(n20606), .ZN(
        P1_U3152) );
  INV_X1 U23557 ( .A(n20610), .ZN(n20666) );
  AOI21_X1 U23558 ( .B1(n20612), .B2(n20611), .A(n20666), .ZN(n20617) );
  OAI22_X1 U23559 ( .A1(n20617), .A2(n20622), .B1(n20614), .B2(n20613), .ZN(
        n20667) );
  AOI22_X1 U23560 ( .A1(n20616), .A2(n20667), .B1(n20666), .B2(n20615), .ZN(
        n20627) );
  OAI21_X1 U23561 ( .B1(n20619), .B2(n20618), .A(n20617), .ZN(n20621) );
  OAI221_X1 U23562 ( .B1(n20624), .B2(n20623), .C1(n20622), .C2(n20621), .A(
        n20620), .ZN(n20671) );
  AOI22_X1 U23563 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20625), .ZN(n20626) );
  OAI211_X1 U23564 ( .C1(n20628), .C2(n20674), .A(n20627), .B(n20626), .ZN(
        P1_U3153) );
  AOI22_X1 U23565 ( .A1(n20630), .A2(n20667), .B1(n20666), .B2(n20629), .ZN(
        n20633) );
  AOI22_X1 U23566 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20631), .ZN(n20632) );
  OAI211_X1 U23567 ( .C1(n20634), .C2(n20674), .A(n20633), .B(n20632), .ZN(
        P1_U3154) );
  AOI22_X1 U23568 ( .A1(n20636), .A2(n20667), .B1(n20666), .B2(n20635), .ZN(
        n20639) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20637), .ZN(n20638) );
  OAI211_X1 U23570 ( .C1(n20640), .C2(n20674), .A(n20639), .B(n20638), .ZN(
        P1_U3155) );
  AOI22_X1 U23571 ( .A1(n20642), .A2(n20667), .B1(n20666), .B2(n20641), .ZN(
        n20645) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20643), .ZN(n20644) );
  OAI211_X1 U23573 ( .C1(n20646), .C2(n20674), .A(n20645), .B(n20644), .ZN(
        P1_U3156) );
  AOI22_X1 U23574 ( .A1(n20648), .A2(n20667), .B1(n20666), .B2(n20647), .ZN(
        n20651) );
  AOI22_X1 U23575 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20649), .ZN(n20650) );
  OAI211_X1 U23576 ( .C1(n20652), .C2(n20674), .A(n20651), .B(n20650), .ZN(
        P1_U3157) );
  AOI22_X1 U23577 ( .A1(n20654), .A2(n20667), .B1(n20666), .B2(n20653), .ZN(
        n20657) );
  AOI22_X1 U23578 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20655), .ZN(n20656) );
  OAI211_X1 U23579 ( .C1(n20658), .C2(n20674), .A(n20657), .B(n20656), .ZN(
        P1_U3158) );
  AOI22_X1 U23580 ( .A1(n20660), .A2(n20667), .B1(n20666), .B2(n20659), .ZN(
        n20663) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20661), .ZN(n20662) );
  OAI211_X1 U23582 ( .C1(n20664), .C2(n20674), .A(n20663), .B(n20662), .ZN(
        P1_U3159) );
  AOI22_X1 U23583 ( .A1(n20668), .A2(n20667), .B1(n20666), .B2(n20665), .ZN(
        n20673) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20671), .B1(
        n20670), .B2(n20669), .ZN(n20672) );
  OAI211_X1 U23585 ( .C1(n20675), .C2(n20674), .A(n20673), .B(n20672), .ZN(
        P1_U3160) );
  OR2_X1 U23586 ( .A1(n20677), .A2(n20676), .ZN(P1_U3163) );
  INV_X1 U23587 ( .A(n20757), .ZN(n20753) );
  AND2_X1 U23588 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20753), .ZN(
        P1_U3164) );
  AND2_X1 U23589 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20753), .ZN(
        P1_U3165) );
  AND2_X1 U23590 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20753), .ZN(
        P1_U3166) );
  AND2_X1 U23591 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20753), .ZN(
        P1_U3167) );
  AND2_X1 U23592 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20753), .ZN(
        P1_U3168) );
  AND2_X1 U23593 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20753), .ZN(
        P1_U3169) );
  AND2_X1 U23594 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20753), .ZN(
        P1_U3170) );
  AND2_X1 U23595 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20753), .ZN(
        P1_U3171) );
  AND2_X1 U23596 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20753), .ZN(
        P1_U3172) );
  AND2_X1 U23597 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20753), .ZN(
        P1_U3173) );
  AND2_X1 U23598 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20753), .ZN(
        P1_U3174) );
  AND2_X1 U23599 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20753), .ZN(
        P1_U3175) );
  AND2_X1 U23600 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20753), .ZN(
        P1_U3176) );
  AND2_X1 U23601 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20753), .ZN(
        P1_U3177) );
  AND2_X1 U23602 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20753), .ZN(
        P1_U3178) );
  AND2_X1 U23603 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20753), .ZN(
        P1_U3179) );
  AND2_X1 U23604 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20753), .ZN(
        P1_U3180) );
  AND2_X1 U23605 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20753), .ZN(
        P1_U3181) );
  AND2_X1 U23606 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20753), .ZN(
        P1_U3182) );
  AND2_X1 U23607 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20753), .ZN(
        P1_U3183) );
  AND2_X1 U23608 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20753), .ZN(
        P1_U3184) );
  AND2_X1 U23609 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20753), .ZN(
        P1_U3185) );
  AND2_X1 U23610 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20753), .ZN(P1_U3186) );
  AND2_X1 U23611 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20753), .ZN(P1_U3187) );
  AND2_X1 U23612 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20753), .ZN(P1_U3188) );
  AND2_X1 U23613 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20753), .ZN(P1_U3189) );
  AND2_X1 U23614 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20753), .ZN(P1_U3190) );
  AND2_X1 U23615 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20753), .ZN(P1_U3191) );
  AND2_X1 U23616 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20753), .ZN(P1_U3192) );
  AND2_X1 U23617 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20753), .ZN(P1_U3193) );
  NAND2_X1 U23618 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20678), .ZN(n20688) );
  INV_X1 U23619 ( .A(n20688), .ZN(n20682) );
  OAI21_X1 U23620 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20689), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20679) );
  AOI211_X1 U23621 ( .C1(HOLD), .C2(P1_STATE_REG_1__SCAN_IN), .A(n20680), .B(
        n20679), .ZN(n20681) );
  OAI22_X1 U23622 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20682), .B1(n20765), 
        .B2(n20681), .ZN(P1_U3194) );
  AOI21_X1 U23623 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20693), .A(n20683), .ZN(n20685) );
  OAI221_X1 U23624 ( .B1(n20685), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .C1(
        n20685), .C2(n20684), .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20692) );
  AOI211_X1 U23625 ( .C1(n20687), .C2(n20689), .A(P1_STATE_REG_2__SCAN_IN), 
        .B(n20686), .ZN(n20691) );
  OAI211_X1 U23626 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20689), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20688), .ZN(n20690) );
  OAI21_X1 U23627 ( .B1(n20692), .B2(n20691), .A(n20690), .ZN(P1_U3196) );
  NAND2_X1 U23628 ( .A1(n20765), .A2(n20693), .ZN(n20746) );
  INV_X1 U23629 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20817) );
  NAND2_X1 U23630 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20765), .ZN(n20742) );
  OAI222_X1 U23631 ( .A1(n20746), .A2(n20695), .B1(n20817), .B2(n20779), .C1(
        n14227), .C2(n20742), .ZN(P1_U3197) );
  INV_X1 U23632 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20694) );
  OAI222_X1 U23633 ( .A1(n20742), .A2(n20695), .B1(n20694), .B2(n20765), .C1(
        n13528), .C2(n20746), .ZN(P1_U3198) );
  INV_X1 U23634 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20696) );
  OAI222_X1 U23635 ( .A1(n20742), .A2(n13528), .B1(n20696), .B2(n20765), .C1(
        n20697), .C2(n20746), .ZN(P1_U3199) );
  OAI222_X1 U23636 ( .A1(n20746), .A2(n20700), .B1(n20698), .B2(n20765), .C1(
        n20697), .C2(n20742), .ZN(P1_U3200) );
  INV_X1 U23637 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20699) );
  OAI222_X1 U23638 ( .A1(n20742), .A2(n20700), .B1(n20699), .B2(n20779), .C1(
        n20702), .C2(n20746), .ZN(P1_U3201) );
  INV_X1 U23639 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20701) );
  OAI222_X1 U23640 ( .A1(n20742), .A2(n20702), .B1(n20701), .B2(n20779), .C1(
        n20704), .C2(n20746), .ZN(P1_U3202) );
  INV_X1 U23641 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20703) );
  OAI222_X1 U23642 ( .A1(n20742), .A2(n20704), .B1(n20703), .B2(n20765), .C1(
        n20706), .C2(n20746), .ZN(P1_U3203) );
  INV_X1 U23643 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20705) );
  OAI222_X1 U23644 ( .A1(n20742), .A2(n20706), .B1(n20705), .B2(n20765), .C1(
        n20708), .C2(n20746), .ZN(P1_U3204) );
  AOI22_X1 U23645 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n20777), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n20740), .ZN(n20707) );
  OAI21_X1 U23646 ( .B1(n20708), .B2(n20742), .A(n20707), .ZN(P1_U3205) );
  INV_X1 U23647 ( .A(n20742), .ZN(n20744) );
  AOI22_X1 U23648 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n20777), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n20744), .ZN(n20709) );
  OAI21_X1 U23649 ( .B1(n20710), .B2(n20746), .A(n20709), .ZN(P1_U3206) );
  AOI222_X1 U23650 ( .A1(n20744), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20777), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20740), .ZN(n20711) );
  INV_X1 U23651 ( .A(n20711), .ZN(P1_U3207) );
  AOI222_X1 U23652 ( .A1(n20740), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20777), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20744), .ZN(n20712) );
  INV_X1 U23653 ( .A(n20712), .ZN(P1_U3208) );
  INV_X1 U23654 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20713) );
  OAI222_X1 U23655 ( .A1(n20742), .A2(n20714), .B1(n20713), .B2(n20765), .C1(
        n20716), .C2(n20746), .ZN(P1_U3209) );
  AOI22_X1 U23656 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20777), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n20740), .ZN(n20715) );
  OAI21_X1 U23657 ( .B1(n20716), .B2(n20742), .A(n20715), .ZN(P1_U3210) );
  INV_X1 U23658 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20718) );
  AOI22_X1 U23659 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n20777), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20740), .ZN(n20717) );
  OAI21_X1 U23660 ( .B1(n20718), .B2(n20742), .A(n20717), .ZN(P1_U3211) );
  AOI22_X1 U23661 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20777), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20744), .ZN(n20719) );
  OAI21_X1 U23662 ( .B1(n20721), .B2(n20746), .A(n20719), .ZN(P1_U3212) );
  AOI22_X1 U23663 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20777), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n20740), .ZN(n20720) );
  OAI21_X1 U23664 ( .B1(n20721), .B2(n20742), .A(n20720), .ZN(P1_U3213) );
  AOI22_X1 U23665 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20777), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n20744), .ZN(n20722) );
  OAI21_X1 U23666 ( .B1(n20724), .B2(n20746), .A(n20722), .ZN(P1_U3214) );
  AOI22_X1 U23667 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20777), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20740), .ZN(n20723) );
  OAI21_X1 U23668 ( .B1(n20724), .B2(n20742), .A(n20723), .ZN(P1_U3215) );
  AOI22_X1 U23669 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20777), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20744), .ZN(n20725) );
  OAI21_X1 U23670 ( .B1(n20727), .B2(n20746), .A(n20725), .ZN(P1_U3216) );
  INV_X1 U23671 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20726) );
  OAI222_X1 U23672 ( .A1(n20742), .A2(n20727), .B1(n20726), .B2(n20765), .C1(
        n20729), .C2(n20746), .ZN(P1_U3217) );
  INV_X1 U23673 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20728) );
  OAI222_X1 U23674 ( .A1(n20742), .A2(n20729), .B1(n20728), .B2(n20779), .C1(
        n20731), .C2(n20746), .ZN(P1_U3218) );
  INV_X1 U23675 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20730) );
  OAI222_X1 U23676 ( .A1(n20742), .A2(n20731), .B1(n20730), .B2(n20779), .C1(
        n20734), .C2(n20746), .ZN(P1_U3219) );
  INV_X1 U23677 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20733) );
  OAI222_X1 U23678 ( .A1(n20742), .A2(n20734), .B1(n20733), .B2(n20779), .C1(
        n20732), .C2(n20746), .ZN(P1_U3220) );
  AOI222_X1 U23679 ( .A1(n20744), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20777), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20740), .ZN(n20735) );
  INV_X1 U23680 ( .A(n20735), .ZN(P1_U3221) );
  AOI222_X1 U23681 ( .A1(n20744), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20777), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20740), .ZN(n20736) );
  INV_X1 U23682 ( .A(n20736), .ZN(P1_U3222) );
  AOI22_X1 U23683 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20740), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20777), .ZN(n20737) );
  OAI21_X1 U23684 ( .B1(n20738), .B2(n20742), .A(n20737), .ZN(P1_U3223) );
  INV_X1 U23685 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20739) );
  INV_X1 U23686 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20846) );
  OAI222_X1 U23687 ( .A1(n20742), .A2(n20739), .B1(n20846), .B2(n20779), .C1(
        n20743), .C2(n20746), .ZN(P1_U3224) );
  AOI22_X1 U23688 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20740), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20777), .ZN(n20741) );
  OAI21_X1 U23689 ( .B1(n20743), .B2(n20742), .A(n20741), .ZN(P1_U3225) );
  AOI22_X1 U23690 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20744), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20777), .ZN(n20745) );
  OAI21_X1 U23691 ( .B1(n20747), .B2(n20746), .A(n20745), .ZN(P1_U3226) );
  INV_X1 U23692 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20823) );
  AOI22_X1 U23693 ( .A1(n20779), .A2(n20748), .B1(n20823), .B2(n20777), .ZN(
        P1_U3458) );
  INV_X1 U23694 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20901) );
  INV_X1 U23695 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20749) );
  AOI22_X1 U23696 ( .A1(n20779), .A2(n20901), .B1(n20749), .B2(n20777), .ZN(
        P1_U3459) );
  INV_X1 U23697 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20851) );
  AOI22_X1 U23698 ( .A1(n20765), .A2(n20750), .B1(n20851), .B2(n20777), .ZN(
        P1_U3460) );
  INV_X1 U23699 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20763) );
  INV_X1 U23700 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20751) );
  AOI22_X1 U23701 ( .A1(n20765), .A2(n20763), .B1(n20751), .B2(n20777), .ZN(
        P1_U3461) );
  INV_X1 U23702 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20754) );
  INV_X1 U23703 ( .A(n20755), .ZN(n20752) );
  AOI21_X1 U23704 ( .B1(n20754), .B2(n20753), .A(n20752), .ZN(P1_U3464) );
  OAI21_X1 U23705 ( .B1(n20757), .B2(n20756), .A(n20755), .ZN(P1_U3465) );
  AOI21_X1 U23706 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20758) );
  AOI22_X1 U23707 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20758), .B2(n14227), .ZN(n20759) );
  AOI22_X1 U23708 ( .A1(n20760), .A2(n20759), .B1(n20901), .B2(n20762), .ZN(
        P1_U3481) );
  NOR2_X1 U23709 ( .A1(n20762), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20761) );
  AOI22_X1 U23710 ( .A1(n20763), .A2(n20762), .B1(n13023), .B2(n20761), .ZN(
        P1_U3482) );
  AOI22_X1 U23711 ( .A1(n20765), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20764), 
        .B2(n20777), .ZN(P1_U3483) );
  AOI211_X1 U23712 ( .C1(n20769), .C2(n20768), .A(n20767), .B(n20766), .ZN(
        n20776) );
  OAI211_X1 U23713 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20771), .A(n20770), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20773) );
  AOI21_X1 U23714 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20773), .A(n20772), 
        .ZN(n20775) );
  NAND2_X1 U23715 ( .A1(n20776), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20774) );
  OAI21_X1 U23716 ( .B1(n20776), .B2(n20775), .A(n20774), .ZN(P1_U3485) );
  AOI22_X1 U23717 ( .A1(n20779), .A2(n20832), .B1(n20778), .B2(n20777), .ZN(
        P1_U3486) );
  AOI22_X1 U23718 ( .A1(n20782), .A2(n20781), .B1(n20780), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n20786) );
  AOI22_X1 U23719 ( .A1(n20784), .A2(BUF2_REG_19__SCAN_IN), .B1(n20783), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n20785) );
  OAI211_X1 U23720 ( .C1(n20788), .C2(n20787), .A(n20786), .B(n20785), .ZN(
        n20789) );
  AOI21_X1 U23721 ( .B1(n20791), .B2(n20790), .A(n20789), .ZN(n20944) );
  NOR4_X1 U23722 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_BE_N_REG_1__SCAN_IN), .A4(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20795) );
  NOR4_X1 U23723 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(
        P1_DATAO_REG_13__SCAN_IN), .A3(P1_BYTEENABLE_REG_2__SCAN_IN), .A4(
        DATAI_0_), .ZN(n20794) );
  NOR4_X1 U23724 ( .A1(BUF1_REG_13__SCAN_IN), .A2(P1_EAX_REG_3__SCAN_IN), .A3(
        P1_UWORD_REG_13__SCAN_IN), .A4(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(
        n20793) );
  NOR4_X1 U23725 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_10__6__SCAN_IN), .A3(P3_REIP_REG_2__SCAN_IN), .A4(
        P3_DATAO_REG_26__SCAN_IN), .ZN(n20792) );
  NAND4_X1 U23726 ( .A1(n20795), .A2(n20794), .A3(n20793), .A4(n20792), .ZN(
        n20812) );
  INV_X1 U23727 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n20913) );
  NAND4_X1 U23728 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(
        P3_MEMORYFETCH_REG_SCAN_IN), .A3(P1_BE_N_REG_3__SCAN_IN), .A4(n20913), 
        .ZN(n20811) );
  NOR4_X1 U23729 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_15__SCAN_IN), .A4(P3_EBX_REG_29__SCAN_IN), .ZN(n20798)
         );
  NOR4_X1 U23730 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(
        BUF2_REG_26__SCAN_IN), .A3(BUF2_REG_22__SCAN_IN), .A4(
        P2_DATAO_REG_28__SCAN_IN), .ZN(n20797) );
  NOR4_X1 U23731 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(DATAI_29_), .A3(
        DATAI_22_), .A4(P1_READREQUEST_REG_SCAN_IN), .ZN(n20796) );
  NAND3_X1 U23732 ( .A1(n20798), .A2(n20797), .A3(n20796), .ZN(n20810) );
  NOR4_X1 U23733 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_7__1__SCAN_IN), .A3(P2_REIP_REG_17__SCAN_IN), .A4(
        n14003), .ZN(n20808) );
  NOR4_X1 U23734 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11704), .A3(
        n20921), .A4(n15174), .ZN(n20807) );
  INV_X1 U23735 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n20850) );
  INV_X1 U23736 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n20886) );
  NAND4_X1 U23737 ( .A1(n20861), .A2(n20886), .A3(n11515), .A4(n20815), .ZN(
        n20799) );
  NOR4_X1 U23738 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20850), .A3(
        n20800), .A4(n20799), .ZN(n20806) );
  NAND4_X1 U23739 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A3(P1_DATAO_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(n20804) );
  NAND4_X1 U23740 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_3__5__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), 
        .A4(P3_DATAO_REG_15__SCAN_IN), .ZN(n20803) );
  NAND4_X1 U23741 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(DATAI_21_), 
        .A3(P3_EAX_REG_21__SCAN_IN), .A4(BUF2_REG_18__SCAN_IN), .ZN(n20802) );
  NAND4_X1 U23742 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_9__4__SCAN_IN), .A3(P1_EBX_REG_17__SCAN_IN), .A4(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20801) );
  NOR4_X1 U23743 ( .A1(n20804), .A2(n20803), .A3(n20802), .A4(n20801), .ZN(
        n20805) );
  NAND4_X1 U23744 ( .A1(n20808), .A2(n20807), .A3(n20806), .A4(n20805), .ZN(
        n20809) );
  NOR4_X1 U23745 ( .A1(n20812), .A2(n20811), .A3(n20810), .A4(n20809), .ZN(
        n20942) );
  AOI22_X1 U23746 ( .A1(n20815), .A2(keyinput38), .B1(keyinput53), .B2(n20814), 
        .ZN(n20813) );
  OAI221_X1 U23747 ( .B1(n20815), .B2(keyinput38), .C1(n20814), .C2(keyinput53), .A(n20813), .ZN(n20827) );
  AOI22_X1 U23748 ( .A1(n20817), .A2(keyinput49), .B1(n14960), .B2(keyinput24), 
        .ZN(n20816) );
  OAI221_X1 U23749 ( .B1(n20817), .B2(keyinput49), .C1(n14960), .C2(keyinput24), .A(n20816), .ZN(n20826) );
  AOI22_X1 U23750 ( .A1(n20820), .A2(keyinput51), .B1(keyinput20), .B2(n20819), 
        .ZN(n20818) );
  OAI221_X1 U23751 ( .B1(n20820), .B2(keyinput51), .C1(n20819), .C2(keyinput20), .A(n20818), .ZN(n20825) );
  AOI22_X1 U23752 ( .A1(n20823), .A2(keyinput35), .B1(keyinput37), .B2(n20822), 
        .ZN(n20821) );
  OAI221_X1 U23753 ( .B1(n20823), .B2(keyinput35), .C1(n20822), .C2(keyinput37), .A(n20821), .ZN(n20824) );
  NOR4_X1 U23754 ( .A1(n20827), .A2(n20826), .A3(n20825), .A4(n20824), .ZN(
        n20875) );
  INV_X1 U23755 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n20829) );
  AOI22_X1 U23756 ( .A1(n20830), .A2(keyinput39), .B1(keyinput6), .B2(n20829), 
        .ZN(n20828) );
  OAI221_X1 U23757 ( .B1(n20830), .B2(keyinput39), .C1(n20829), .C2(keyinput6), 
        .A(n20828), .ZN(n20843) );
  INV_X1 U23758 ( .A(DATAI_29_), .ZN(n20833) );
  AOI22_X1 U23759 ( .A1(n20833), .A2(keyinput9), .B1(keyinput27), .B2(n20832), 
        .ZN(n20831) );
  OAI221_X1 U23760 ( .B1(n20833), .B2(keyinput9), .C1(n20832), .C2(keyinput27), 
        .A(n20831), .ZN(n20842) );
  AOI22_X1 U23761 ( .A1(n20836), .A2(keyinput28), .B1(keyinput46), .B2(n20835), 
        .ZN(n20834) );
  OAI221_X1 U23762 ( .B1(n20836), .B2(keyinput28), .C1(n20835), .C2(keyinput46), .A(n20834), .ZN(n20841) );
  AOI22_X1 U23763 ( .A1(n20839), .A2(keyinput1), .B1(n20838), .B2(keyinput15), 
        .ZN(n20837) );
  OAI221_X1 U23764 ( .B1(n20839), .B2(keyinput1), .C1(n20838), .C2(keyinput15), 
        .A(n20837), .ZN(n20840) );
  NOR4_X1 U23765 ( .A1(n20843), .A2(n20842), .A3(n20841), .A4(n20840), .ZN(
        n20874) );
  AOI22_X1 U23766 ( .A1(n20846), .A2(keyinput4), .B1(keyinput59), .B2(n20845), 
        .ZN(n20844) );
  OAI221_X1 U23767 ( .B1(n20846), .B2(keyinput4), .C1(n20845), .C2(keyinput59), 
        .A(n20844), .ZN(n20857) );
  AOI22_X1 U23768 ( .A1(n20848), .A2(keyinput0), .B1(n10089), .B2(keyinput32), 
        .ZN(n20847) );
  OAI221_X1 U23769 ( .B1(n20848), .B2(keyinput0), .C1(n10089), .C2(keyinput32), 
        .A(n20847), .ZN(n20856) );
  AOI22_X1 U23770 ( .A1(n20851), .A2(keyinput10), .B1(n20850), .B2(keyinput44), 
        .ZN(n20849) );
  OAI221_X1 U23771 ( .B1(n20851), .B2(keyinput10), .C1(n20850), .C2(keyinput44), .A(n20849), .ZN(n20855) );
  XOR2_X1 U23772 ( .A(n11704), .B(keyinput61), .Z(n20853) );
  XNOR2_X1 U23773 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B(keyinput54), .ZN(
        n20852) );
  NAND2_X1 U23774 ( .A1(n20853), .A2(n20852), .ZN(n20854) );
  NOR4_X1 U23775 ( .A1(n20857), .A2(n20856), .A3(n20855), .A4(n20854), .ZN(
        n20873) );
  AOI22_X1 U23776 ( .A1(n20859), .A2(keyinput12), .B1(n14299), .B2(keyinput56), 
        .ZN(n20858) );
  OAI221_X1 U23777 ( .B1(n20859), .B2(keyinput12), .C1(n14299), .C2(keyinput56), .A(n20858), .ZN(n20871) );
  AOI22_X1 U23778 ( .A1(n20862), .A2(keyinput13), .B1(n20861), .B2(keyinput47), 
        .ZN(n20860) );
  OAI221_X1 U23779 ( .B1(n20862), .B2(keyinput13), .C1(n20861), .C2(keyinput47), .A(n20860), .ZN(n20870) );
  AOI22_X1 U23780 ( .A1(n20865), .A2(keyinput58), .B1(keyinput36), .B2(n20864), 
        .ZN(n20863) );
  OAI221_X1 U23781 ( .B1(n20865), .B2(keyinput58), .C1(n20864), .C2(keyinput36), .A(n20863), .ZN(n20869) );
  AOI22_X1 U23782 ( .A1(n20867), .A2(keyinput2), .B1(n13889), .B2(keyinput22), 
        .ZN(n20866) );
  OAI221_X1 U23783 ( .B1(n20867), .B2(keyinput2), .C1(n13889), .C2(keyinput22), 
        .A(n20866), .ZN(n20868) );
  NOR4_X1 U23784 ( .A1(n20871), .A2(n20870), .A3(n20869), .A4(n20868), .ZN(
        n20872) );
  NAND4_X1 U23785 ( .A1(n20875), .A2(n20874), .A3(n20873), .A4(n20872), .ZN(
        n20940) );
  AOI22_X1 U23786 ( .A1(n20878), .A2(keyinput21), .B1(n20877), .B2(keyinput11), 
        .ZN(n20876) );
  OAI221_X1 U23787 ( .B1(n20878), .B2(keyinput21), .C1(n20877), .C2(keyinput11), .A(n20876), .ZN(n20890) );
  AOI22_X1 U23788 ( .A1(n20881), .A2(keyinput41), .B1(n20880), .B2(keyinput40), 
        .ZN(n20879) );
  OAI221_X1 U23789 ( .B1(n20881), .B2(keyinput41), .C1(n20880), .C2(keyinput40), .A(n20879), .ZN(n20889) );
  INV_X1 U23790 ( .A(DATAI_21_), .ZN(n20883) );
  AOI22_X1 U23791 ( .A1(n20883), .A2(keyinput45), .B1(n14003), .B2(keyinput34), 
        .ZN(n20882) );
  OAI221_X1 U23792 ( .B1(n20883), .B2(keyinput45), .C1(n14003), .C2(keyinput34), .A(n20882), .ZN(n20888) );
  AOI22_X1 U23793 ( .A1(n20886), .A2(keyinput3), .B1(keyinput63), .B2(n20885), 
        .ZN(n20884) );
  OAI221_X1 U23794 ( .B1(n20886), .B2(keyinput3), .C1(n20885), .C2(keyinput63), 
        .A(n20884), .ZN(n20887) );
  NOR4_X1 U23795 ( .A1(n20890), .A2(n20889), .A3(n20888), .A4(n20887), .ZN(
        n20938) );
  AOI22_X1 U23796 ( .A1(n20893), .A2(keyinput57), .B1(n20892), .B2(keyinput50), 
        .ZN(n20891) );
  OAI221_X1 U23797 ( .B1(n20893), .B2(keyinput57), .C1(n20892), .C2(keyinput50), .A(n20891), .ZN(n20897) );
  XNOR2_X1 U23798 ( .A(n20894), .B(keyinput33), .ZN(n20896) );
  XOR2_X1 U23799 ( .A(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B(keyinput7), .Z(
        n20895) );
  OR3_X1 U23800 ( .A1(n20897), .A2(n20896), .A3(n20895), .ZN(n20905) );
  INV_X1 U23801 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n20899) );
  AOI22_X1 U23802 ( .A1(n20899), .A2(keyinput23), .B1(n11515), .B2(keyinput62), 
        .ZN(n20898) );
  OAI221_X1 U23803 ( .B1(n20899), .B2(keyinput23), .C1(n11515), .C2(keyinput62), .A(n20898), .ZN(n20904) );
  AOI22_X1 U23804 ( .A1(n20902), .A2(keyinput19), .B1(n20901), .B2(keyinput5), 
        .ZN(n20900) );
  OAI221_X1 U23805 ( .B1(n20902), .B2(keyinput19), .C1(n20901), .C2(keyinput5), 
        .A(n20900), .ZN(n20903) );
  NOR3_X1 U23806 ( .A1(n20905), .A2(n20904), .A3(n20903), .ZN(n20937) );
  AOI22_X1 U23807 ( .A1(n20907), .A2(keyinput42), .B1(n14014), .B2(keyinput14), 
        .ZN(n20906) );
  OAI221_X1 U23808 ( .B1(n20907), .B2(keyinput42), .C1(n14014), .C2(keyinput14), .A(n20906), .ZN(n20919) );
  INV_X1 U23809 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n20909) );
  AOI22_X1 U23810 ( .A1(n20910), .A2(keyinput43), .B1(n20909), .B2(keyinput26), 
        .ZN(n20908) );
  OAI221_X1 U23811 ( .B1(n20910), .B2(keyinput43), .C1(n20909), .C2(keyinput26), .A(n20908), .ZN(n20918) );
  INV_X1 U23812 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n20912) );
  AOI22_X1 U23813 ( .A1(n20913), .A2(keyinput16), .B1(keyinput31), .B2(n20912), 
        .ZN(n20911) );
  OAI221_X1 U23814 ( .B1(n20913), .B2(keyinput16), .C1(n20912), .C2(keyinput31), .A(n20911), .ZN(n20917) );
  AOI22_X1 U23815 ( .A1(n15174), .A2(keyinput25), .B1(keyinput30), .B2(n20915), 
        .ZN(n20914) );
  OAI221_X1 U23816 ( .B1(n15174), .B2(keyinput25), .C1(n20915), .C2(keyinput30), .A(n20914), .ZN(n20916) );
  NOR4_X1 U23817 ( .A1(n20919), .A2(n20918), .A3(n20917), .A4(n20916), .ZN(
        n20936) );
  AOI22_X1 U23818 ( .A1(n9892), .A2(keyinput52), .B1(n20921), .B2(keyinput8), 
        .ZN(n20920) );
  OAI221_X1 U23819 ( .B1(n9892), .B2(keyinput52), .C1(n20921), .C2(keyinput8), 
        .A(n20920), .ZN(n20934) );
  AOI22_X1 U23820 ( .A1(n20924), .A2(keyinput18), .B1(keyinput17), .B2(n20923), 
        .ZN(n20922) );
  OAI221_X1 U23821 ( .B1(n20924), .B2(keyinput18), .C1(n20923), .C2(keyinput17), .A(n20922), .ZN(n20933) );
  INV_X1 U23822 ( .A(DATAI_0_), .ZN(n20926) );
  AOI22_X1 U23823 ( .A1(n20927), .A2(keyinput55), .B1(keyinput48), .B2(n20926), 
        .ZN(n20925) );
  OAI221_X1 U23824 ( .B1(n20927), .B2(keyinput55), .C1(n20926), .C2(keyinput48), .A(n20925), .ZN(n20932) );
  INV_X1 U23825 ( .A(DATAI_22_), .ZN(n20930) );
  AOI22_X1 U23826 ( .A1(n20930), .A2(keyinput60), .B1(keyinput29), .B2(n20929), 
        .ZN(n20928) );
  OAI221_X1 U23827 ( .B1(n20930), .B2(keyinput60), .C1(n20929), .C2(keyinput29), .A(n20928), .ZN(n20931) );
  NOR4_X1 U23828 ( .A1(n20934), .A2(n20933), .A3(n20932), .A4(n20931), .ZN(
        n20935) );
  NAND4_X1 U23829 ( .A1(n20938), .A2(n20937), .A3(n20936), .A4(n20935), .ZN(
        n20939) );
  NOR2_X1 U23830 ( .A1(n20940), .A2(n20939), .ZN(n20941) );
  XOR2_X1 U23831 ( .A(n20942), .B(n20941), .Z(n20943) );
  XNOR2_X1 U23832 ( .A(n20944), .B(n20943), .ZN(P2_U2900) );
  INV_X1 U15504 ( .A(n10015), .ZN(n17063) );
  CLKBUF_X3 U12798 ( .A(n12515), .Z(n17054) );
  BUF_X2 U11099 ( .A(n15856), .Z(n9582) );
  XNOR2_X1 U11123 ( .A(n13964), .B(n13961), .ZN(n14882) );
  INV_X1 U11054 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18690) );
  CLKBUF_X1 U11042 ( .A(n9604), .Z(n9619) );
  OR2_X1 U11067 ( .A1(n12426), .A2(n18517), .ZN(n12438) );
  CLKBUF_X1 U11093 ( .A(n11737), .Z(n12077) );
  NAND2_X1 U11096 ( .A1(n11336), .A2(n11335), .ZN(n11423) );
  CLKBUF_X1 U11102 ( .A(n12470), .Z(n16813) );
  AND2_X1 U11130 ( .A1(n9662), .A2(n17853), .ZN(n9904) );
  INV_X1 U11133 ( .A(n17246), .ZN(n12509) );
  CLKBUF_X1 U11171 ( .A(n14474), .Z(n15893) );
  CLKBUF_X1 U11421 ( .A(n11521), .Z(n19890) );
  NAND2_X1 U11438 ( .A1(n11429), .A2(n11428), .ZN(n11883) );
  CLKBUF_X1 U12103 ( .A(n14388), .Z(n14389) );
  CLKBUF_X1 U12184 ( .A(n13478), .Z(n20093) );
  CLKBUF_X1 U12278 ( .A(n18495), .Z(n9580) );
  CLKBUF_X1 U12590 ( .A(n16376), .Z(n16381) );
endmodule

