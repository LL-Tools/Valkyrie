

module b21_C_gen_AntiSAT_k_256_5 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67, 
        keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72, 
        keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77, 
        keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82, 
        keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87, 
        keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92, 
        keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97, 
        keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499;

  AND3_X1 U4985 ( .A1(n5899), .A2(n5898), .A3(n5897), .ZN(n10304) );
  CLKBUF_X2 U4986 ( .A(n5591), .Z(n4487) );
  CLKBUF_X2 U4987 ( .A(n5591), .Z(n4486) );
  NAND2_X1 U4988 ( .A1(n9615), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U4989 ( .A1(n5164), .A2(n4509), .ZN(n8552) );
  NAND2_X1 U4990 ( .A1(n7668), .A2(n5322), .ZN(n7736) );
  INV_X2 U4991 ( .A(n5210), .ZN(n5453) );
  NAND2_X2 U4992 ( .A1(n5673), .A2(n8552), .ZN(n5210) );
  OAI21_X1 U4993 ( .B1(n7802), .B2(n7922), .A(n7885), .ZN(n7916) );
  INV_X1 U4994 ( .A(n5739), .ZN(n5737) );
  BUF_X1 U4995 ( .A(n7547), .Z(n4482) );
  AOI21_X1 U4996 ( .B1(n5682), .B2(n10357), .A(n5681), .ZN(n7957) );
  NAND4_X1 U4997 ( .A1(n5743), .A2(n5742), .A3(n5741), .A4(n5740), .ZN(n9168)
         );
  XNOR2_X1 U4998 ( .A(n5284), .B(n5283), .ZN(n6685) );
  NAND2_X2 U4999 ( .A1(n7832), .A2(n8111), .ZN(n10111) );
  OAI211_X1 U5000 ( .C1(n8357), .C2(n6667), .A(n5238), .B(n5237), .ZN(n7351)
         );
  INV_X2 U5001 ( .A(n8576), .ZN(n6399) );
  NAND3_X2 U5002 ( .A1(n5219), .A2(n5218), .A3(n5217), .ZN(n8576) );
  NAND2_X2 U5003 ( .A1(n5088), .A2(n5087), .ZN(n5284) );
  XNOR2_X2 U5004 ( .A(n5642), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8407) );
  NAND3_X2 U5005 ( .A1(n5208), .A2(n5207), .A3(n5206), .ZN(n8579) );
  NAND2_X1 U5006 ( .A1(n4827), .A2(n4826), .ZN(n4480) );
  NAND2_X1 U5007 ( .A1(n4827), .A2(n4826), .ZN(n4481) );
  NAND2_X1 U5008 ( .A1(n4827), .A2(n4826), .ZN(n5222) );
  AOI21_X2 U5009 ( .B1(n8793), .B2(n5465), .A(n5464), .ZN(n8778) );
  NAND2_X2 U5010 ( .A1(n8820), .A2(n5448), .ZN(n8793) );
  XNOR2_X2 U5011 ( .A(n5736), .B(n5735), .ZN(n5739) );
  OR2_X2 U5012 ( .A1(n5173), .A2(n9022), .ZN(n5171) );
  XNOR2_X2 U5013 ( .A(n7062), .B(n7274), .ZN(n8105) );
  NAND4_X4 U5014 ( .A1(n5813), .A2(n5812), .A3(n5811), .A4(n5810), .ZN(n7062)
         );
  OR2_X1 U5015 ( .A1(n6547), .A2(n8348), .ZN(n4821) );
  AND3_X1 U5016 ( .A1(n6506), .A2(n6505), .A3(n4915), .ZN(n6547) );
  AND2_X1 U5017 ( .A1(n5016), .A2(n4548), .ZN(n8709) );
  AND2_X1 U5018 ( .A1(n5613), .A2(n5590), .ZN(n8669) );
  OR2_X1 U5019 ( .A1(n5589), .A2(n9779), .ZN(n5613) );
  NAND2_X1 U5020 ( .A1(n7110), .A2(n7112), .ZN(n7111) );
  NAND2_X1 U5021 ( .A1(n8160), .A2(n7457), .ZN(n7444) );
  INV_X2 U5022 ( .A(n9508), .ZN(n4483) );
  INV_X2 U5023 ( .A(n7231), .ZN(n7233) );
  INV_X2 U5024 ( .A(n5852), .ZN(n6332) );
  INV_X1 U5025 ( .A(n5803), .ZN(n6306) );
  INV_X2 U5027 ( .A(n5615), .ZN(n5195) );
  NAND2_X1 U5028 ( .A1(n5210), .A2(n6660), .ZN(n8357) );
  AND2_X1 U5029 ( .A1(n9027), .A2(n5175), .ZN(n5591) );
  MUX2_X1 U5030 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5160), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5161) );
  AND2_X1 U5031 ( .A1(n5874), .A2(n5729), .ZN(n5895) );
  INV_X2 U5032 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U5033 ( .A1(n4727), .A2(n4723), .ZN(n8558) );
  OR2_X1 U5034 ( .A1(n6586), .A2(n6358), .ZN(n6389) );
  NOR2_X1 U5035 ( .A1(n4725), .A2(n4926), .ZN(n4724) );
  OAI21_X1 U5036 ( .B1(n6586), .B2(n4759), .A(n10101), .ZN(n6593) );
  CLKBUF_X1 U5037 ( .A(n9060), .Z(n9137) );
  OR2_X1 U5038 ( .A1(n5007), .A2(n9034), .ZN(n5005) );
  AND2_X1 U5039 ( .A1(n4744), .A2(n4550), .ZN(n9098) );
  NAND2_X1 U5040 ( .A1(n6503), .A2(n6502), .ZN(n6506) );
  NAND2_X1 U5041 ( .A1(n8657), .A2(n5671), .ZN(n8661) );
  NAND2_X1 U5042 ( .A1(n4584), .A2(n9109), .ZN(n9053) );
  NAND2_X1 U5043 ( .A1(n4585), .A2(n4998), .ZN(n6147) );
  NAND2_X1 U5044 ( .A1(n7877), .A2(n8464), .ZN(n7876) );
  OR2_X1 U5045 ( .A1(n5055), .A2(n5663), .ZN(n4947) );
  AND2_X1 U5046 ( .A1(n7795), .A2(n8461), .ZN(n7877) );
  NAND2_X1 U5047 ( .A1(n4583), .A2(n5008), .ZN(n10100) );
  AND2_X1 U5048 ( .A1(n7782), .A2(n4689), .ZN(n4688) );
  NAND2_X1 U5049 ( .A1(n7798), .A2(n5037), .ZN(n5035) );
  NAND2_X1 U5050 ( .A1(n7648), .A2(n4683), .ZN(n7779) );
  AND2_X1 U5051 ( .A1(n7621), .A2(n5308), .ZN(n7670) );
  NAND2_X1 U5052 ( .A1(n5169), .A2(n5168), .ZN(n8946) );
  NAND2_X1 U5053 ( .A1(n7550), .A2(n7549), .ZN(n7548) );
  NAND2_X1 U5054 ( .A1(n7377), .A2(n5273), .ZN(n7550) );
  AOI21_X1 U5055 ( .B1(n4943), .B2(n7549), .A(n4942), .ZN(n4941) );
  NAND2_X1 U5056 ( .A1(n5361), .A2(n5360), .ZN(n7805) );
  NAND2_X1 U5057 ( .A1(n5989), .A2(n5988), .ZN(n10163) );
  INV_X1 U5058 ( .A(n7173), .ZN(n7174) );
  AND2_X1 U5059 ( .A1(n4818), .A2(n6422), .ZN(n5057) );
  AOI21_X1 U5060 ( .B1(n8430), .B2(n4945), .A(n4944), .ZN(n4943) );
  NAND2_X1 U5061 ( .A1(n5971), .A2(n5970), .ZN(n7831) );
  NAND2_X1 U5062 ( .A1(n5948), .A2(n5947), .ZN(n10277) );
  AND2_X1 U5063 ( .A1(n7592), .A2(n10316), .ZN(n10280) );
  NAND2_X2 U5064 ( .A1(n7473), .A2(n9505), .ZN(n9508) );
  INV_X1 U5065 ( .A(n7351), .ZN(n10419) );
  NAND2_X1 U5066 ( .A1(n5084), .A2(n5083), .ZN(n4814) );
  NAND2_X1 U5067 ( .A1(n5080), .A2(n5079), .ZN(n5257) );
  NAND4_X1 U5068 ( .A1(n5833), .A2(n5832), .A3(n5831), .A4(n5830), .ZN(n9167)
         );
  NAND3_X1 U5069 ( .A1(n5197), .A2(n4511), .A3(n5196), .ZN(n8577) );
  AND4_X1 U5070 ( .A1(n5267), .A2(n5266), .A3(n5265), .A4(n5264), .ZN(n7423)
         );
  AND2_X1 U5071 ( .A1(n4681), .A2(n4680), .ZN(n6835) );
  OR2_X1 U5072 ( .A1(n6848), .A2(n4682), .ZN(n4681) );
  CLKBUF_X2 U5073 ( .A(n5888), .Z(n4484) );
  INV_X2 U5074 ( .A(n8357), .ZN(n8352) );
  CLKBUF_X1 U5075 ( .A(n5214), .Z(n5637) );
  NAND2_X2 U5076 ( .A1(n9031), .A2(n9027), .ZN(n5615) );
  INV_X2 U5077 ( .A(n5798), .ZN(n6629) );
  XNOR2_X1 U5078 ( .A(n5768), .B(n5767), .ZN(n5786) );
  NAND2_X2 U5079 ( .A1(n4917), .A2(n5175), .ZN(n5229) );
  INV_X1 U5080 ( .A(n9027), .ZN(n4917) );
  XNOR2_X1 U5081 ( .A(n5761), .B(P1_IR_REG_25__SCAN_IN), .ZN(n7825) );
  NAND2_X1 U5082 ( .A1(n5754), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5761) );
  AOI21_X1 U5083 ( .B1(n4612), .B2(n4524), .A(n4611), .ZN(n4581) );
  MUX2_X1 U5084 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5163), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5164) );
  MUX2_X1 U5085 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5172), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5174) );
  OR2_X1 U5086 ( .A1(n5771), .A2(n5755), .ZN(n4588) );
  AND2_X1 U5087 ( .A1(n5773), .A2(n4497), .ZN(n5771) );
  OR2_X2 U5088 ( .A1(n7982), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6706) );
  INV_X1 U5089 ( .A(n4889), .ZN(n5773) );
  AND2_X1 U5090 ( .A1(n5748), .A2(n4764), .ZN(n5756) );
  INV_X1 U5091 ( .A(n5747), .ZN(n5748) );
  AND2_X1 U5092 ( .A1(n4766), .A2(n4765), .ZN(n4764) );
  NAND2_X1 U5093 ( .A1(n5796), .A2(n4972), .ZN(n5065) );
  AND2_X1 U5094 ( .A1(n5015), .A2(n5733), .ZN(n5014) );
  NOR2_X1 U5095 ( .A1(n4490), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n4766) );
  AND2_X1 U5096 ( .A1(n4885), .A2(n5753), .ZN(n5015) );
  AND2_X1 U5097 ( .A1(n5155), .A2(n5259), .ZN(n4961) );
  AND2_X1 U5098 ( .A1(n5029), .A2(n5166), .ZN(n4962) );
  AND3_X1 U5099 ( .A1(n4587), .A2(n5731), .A3(n5732), .ZN(n5733) );
  NAND2_X1 U5100 ( .A1(n10014), .A2(n4973), .ZN(n4643) );
  AND4_X1 U5101 ( .A1(n5153), .A2(n5355), .A3(n5373), .A4(n5389), .ZN(n5155)
         );
  AND2_X1 U5102 ( .A1(n4887), .A2(n4886), .ZN(n4885) );
  AND4_X1 U5103 ( .A1(n4825), .A2(n4824), .A3(n4823), .A4(n4822), .ZN(n5156)
         );
  AND2_X1 U5104 ( .A1(n5031), .A2(n5030), .ZN(n5029) );
  AND2_X1 U5105 ( .A1(n5730), .A2(n5967), .ZN(n4587) );
  AND3_X1 U5106 ( .A1(n4758), .A2(n4757), .A3(n4756), .ZN(n5874) );
  AND2_X1 U5107 ( .A1(n5223), .A2(n5154), .ZN(n5259) );
  NOR2_X1 U5108 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4771) );
  NOR2_X1 U5109 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5154) );
  NOR2_X1 U5110 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4769) );
  NOR2_X1 U5111 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4772) );
  NOR2_X1 U5112 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5223) );
  CLKBUF_X1 U5113 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n10355) );
  NOR2_X1 U5114 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4757) );
  NOR2_X1 U5115 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4758) );
  AND2_X1 U5116 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n10014) );
  INV_X2 U5117 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U5118 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5355) );
  INV_X1 U5119 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9992) );
  NOR2_X1 U5120 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n4611) );
  INV_X1 U5121 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5967) );
  NOR2_X1 U5122 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4824) );
  INV_X1 U5123 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5389) );
  INV_X1 U5124 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5757) );
  NOR2_X1 U5125 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5153) );
  INV_X1 U5126 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5373) );
  INV_X1 U5127 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5749) );
  NOR2_X1 U5128 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4825) );
  NOR2_X1 U5129 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n4822) );
  INV_X1 U5130 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5031) );
  NOR2_X1 U5131 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4823) );
  NOR2_X2 U5132 ( .A1(n9504), .A2(n9483), .ZN(n9482) );
  NAND2_X1 U5133 ( .A1(n6399), .A2(n7231), .ZN(n8421) );
  XNOR2_X1 U5134 ( .A(n5235), .B(n5234), .ZN(n6667) );
  XNOR2_X1 U5135 ( .A(n5074), .B(n5073), .ZN(n5235) );
  OAI21_X2 U5136 ( .B1(n7736), .B2(n5351), .A(n5350), .ZN(n7798) );
  NAND2_X1 U5138 ( .A1(n5737), .A2(n5738), .ZN(n5888) );
  OAI222_X1 U5139 ( .A1(n9622), .A2(n6668), .B1(n9624), .B2(n6667), .C1(
        P1_U3084), .C2(n6666), .ZN(P1_U3350) );
  XNOR2_X2 U5140 ( .A(n5200), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10023) );
  AOI211_X2 U5141 ( .C1(n10164), .C2(n10146), .A(n10145), .B(n10144), .ZN(
        n10173) );
  INV_X1 U5142 ( .A(n5416), .ZN(n4977) );
  OR2_X1 U5143 ( .A1(n7954), .A2(n8649), .ZN(n8532) );
  NOR2_X1 U5144 ( .A1(n8377), .A2(n5021), .ZN(n5020) );
  INV_X1 U5145 ( .A(n5023), .ZN(n5021) );
  NAND2_X1 U5146 ( .A1(n8750), .A2(n8737), .ZN(n5027) );
  NAND2_X1 U5147 ( .A1(n9304), .A2(n9239), .ZN(n4876) );
  OR2_X1 U5148 ( .A1(n9531), .A2(n9239), .ZN(n9264) );
  OAI21_X1 U5149 ( .B1(n5518), .B2(n5517), .A(n5516), .ZN(n5527) );
  NOR2_X1 U5150 ( .A1(n5131), .A2(n4983), .ZN(n4982) );
  INV_X1 U5151 ( .A(n5126), .ZN(n4983) );
  INV_X1 U5152 ( .A(n5385), .ZN(n5131) );
  NAND2_X1 U5153 ( .A1(n5372), .A2(n5371), .ZN(n5127) );
  XNOR2_X1 U5154 ( .A(n8388), .B(n8650), .ZN(n8379) );
  NAND2_X1 U5155 ( .A1(n5210), .A2(n4831), .ZN(n4832) );
  NAND2_X1 U5156 ( .A1(n4743), .A2(n4566), .ZN(n4744) );
  INV_X1 U5157 ( .A(n8520), .ZN(n4722) );
  OR2_X1 U5158 ( .A1(n5599), .A2(n5598), .ZN(n5601) );
  NOR2_X1 U5159 ( .A1(n8542), .A2(n8387), .ZN(n8538) );
  OR2_X1 U5160 ( .A1(n8722), .A2(n8738), .ZN(n8500) );
  AND2_X1 U5161 ( .A1(n8713), .A2(n8499), .ZN(n8377) );
  OR2_X1 U5162 ( .A1(n7805), .A2(n7878), .ZN(n8461) );
  AND2_X1 U5163 ( .A1(n5156), .A2(n4959), .ZN(n4958) );
  INV_X1 U5164 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4959) );
  INV_X1 U5165 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U5166 ( .A1(n4755), .A2(n4753), .ZN(n4752) );
  INV_X1 U5167 ( .A(n5926), .ZN(n4753) );
  NOR2_X1 U5168 ( .A1(n7860), .A2(n4763), .ZN(n4762) );
  INV_X1 U5169 ( .A(n7725), .ZN(n4763) );
  NAND2_X1 U5170 ( .A1(n7254), .A2(n5864), .ZN(n5886) );
  OR2_X1 U5171 ( .A1(n6043), .A2(n5011), .ZN(n5010) );
  INV_X1 U5172 ( .A(n6023), .ZN(n5011) );
  AND2_X1 U5173 ( .A1(n8067), .A2(n8066), .ZN(n8081) );
  OR2_X1 U5174 ( .A1(n9523), .A2(n8092), .ZN(n8127) );
  NAND2_X1 U5175 ( .A1(n9547), .A2(n9234), .ZN(n9258) );
  INV_X1 U5176 ( .A(n8076), .ZN(n6372) );
  NAND2_X1 U5177 ( .A1(n7689), .A2(n7688), .ZN(n4864) );
  NAND2_X1 U5178 ( .A1(n6336), .A2(n9322), .ZN(n7058) );
  NAND2_X1 U5179 ( .A1(n5629), .A2(n5628), .ZN(n7974) );
  NAND2_X1 U5180 ( .A1(n4987), .A2(n4985), .ZN(n5629) );
  NAND2_X1 U5181 ( .A1(n5527), .A2(n5526), .ZN(n5538) );
  NAND2_X1 U5182 ( .A1(n4669), .A2(n4667), .ZN(n5503) );
  AOI21_X1 U5183 ( .B1(n4671), .B2(n4673), .A(n4668), .ZN(n4667) );
  INV_X1 U5184 ( .A(n5487), .ZN(n4668) );
  AND2_X1 U5185 ( .A1(n5487), .A2(n5472), .ZN(n5485) );
  AND2_X1 U5186 ( .A1(n5142), .A2(n5141), .ZN(n5416) );
  NAND2_X1 U5187 ( .A1(n5136), .A2(n5135), .ZN(n5402) );
  XNOR2_X1 U5188 ( .A(n5129), .B(n5128), .ZN(n5385) );
  OAI21_X1 U5189 ( .B1(n4966), .B2(n4489), .A(n4963), .ZN(n5372) );
  INV_X1 U5190 ( .A(n4964), .ZN(n4963) );
  OAI21_X1 U5191 ( .B1(n4489), .B2(n4969), .A(n5121), .ZN(n4964) );
  AND2_X1 U5192 ( .A1(n5126), .A2(n5125), .ZN(n5371) );
  XNOR2_X1 U5193 ( .A(n5113), .B(SI_11_), .ZN(n5335) );
  NAND2_X1 U5194 ( .A1(n5098), .A2(n5097), .ZN(n5298) );
  NAND2_X1 U5195 ( .A1(n8577), .A2(n10436), .ZN(n6395) );
  OR2_X1 U5196 ( .A1(n5559), .A2(n5558), .ZN(n5589) );
  NOR2_X1 U5197 ( .A1(n4906), .A2(n4905), .ZN(n4904) );
  AOI21_X1 U5198 ( .B1(n4899), .B2(n4901), .A(n4536), .ZN(n4897) );
  NAND2_X1 U5199 ( .A1(n8337), .A2(n8338), .ZN(n6461) );
  OAI21_X1 U5200 ( .B1(n4928), .B2(n8359), .A(n4923), .ZN(n4725) );
  NAND2_X1 U5201 ( .A1(n4531), .A2(n8551), .ZN(n4928) );
  INV_X1 U5202 ( .A(n4487), .ZN(n5476) );
  INV_X1 U5203 ( .A(n5229), .ZN(n5634) );
  INV_X1 U5204 ( .A(n5214), .ZN(n5674) );
  AND2_X1 U5205 ( .A1(n6853), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4682) );
  NAND2_X1 U5206 ( .A1(n7652), .A2(n5394), .ZN(n4683) );
  NAND2_X1 U5207 ( .A1(n8661), .A2(n8515), .ZN(n6559) );
  AND2_X1 U5208 ( .A1(n5042), .A2(n6555), .ZN(n5041) );
  NAND2_X1 U5209 ( .A1(n8677), .A2(n5043), .ZN(n5042) );
  INV_X1 U5210 ( .A(n5548), .ZN(n5043) );
  AND2_X1 U5211 ( .A1(n5669), .A2(n8505), .ZN(n4920) );
  NAND2_X1 U5212 ( .A1(n4545), .A2(n5027), .ZN(n5023) );
  OAI21_X1 U5213 ( .B1(n8782), .B2(n8321), .A(n5466), .ZN(n8758) );
  NAND2_X1 U5214 ( .A1(n5034), .A2(n4521), .ZN(n8820) );
  AND2_X1 U5215 ( .A1(n8878), .A2(n8458), .ZN(n4957) );
  NAND2_X1 U5216 ( .A1(n4922), .A2(n4921), .ZN(n7795) );
  AND2_X1 U5217 ( .A1(n7797), .A2(n8456), .ZN(n4921) );
  NOR2_X1 U5218 ( .A1(n5051), .A2(n5061), .ZN(n5350) );
  NAND2_X1 U5219 ( .A1(n7548), .A2(n4527), .ZN(n7621) );
  NAND2_X1 U5220 ( .A1(n7243), .A2(n5248), .ZN(n7409) );
  NAND2_X1 U5221 ( .A1(n4829), .A2(n5161), .ZN(n4826) );
  NAND2_X1 U5222 ( .A1(n4828), .A2(n7982), .ZN(n4827) );
  NOR2_X1 U5223 ( .A1(n4830), .A2(n6660), .ZN(n4829) );
  NAND2_X1 U5224 ( .A1(n9053), .A2(n9054), .ZN(n6225) );
  OAI21_X1 U5225 ( .B1(n9034), .B2(n5003), .A(n5004), .ZN(n9060) );
  NAND2_X1 U5226 ( .A1(n5006), .A2(n6264), .ZN(n5004) );
  OR2_X1 U5227 ( .A1(n9098), .A2(n4557), .ZN(n5003) );
  NAND2_X1 U5228 ( .A1(n6268), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6285) );
  OR2_X1 U5229 ( .A1(n6285), .A2(n9140), .ZN(n6319) );
  NOR2_X1 U5230 ( .A1(n7128), .A2(n7129), .ZN(n9169) );
  NAND2_X1 U5231 ( .A1(n4544), .A2(n4876), .ZN(n4873) );
  AOI21_X1 U5232 ( .B1(n4873), .B2(n4871), .A(n9265), .ZN(n4870) );
  INV_X1 U5233 ( .A(n4874), .ZN(n4871) );
  INV_X1 U5234 ( .A(n4873), .ZN(n4872) );
  OR2_X1 U5235 ( .A1(n9540), .A2(n9316), .ZN(n9237) );
  AND2_X1 U5236 ( .A1(n5798), .A2(n7982), .ZN(n5834) );
  NAND2_X2 U5237 ( .A1(n6365), .A2(n6955), .ZN(n5798) );
  NAND2_X1 U5238 ( .A1(n4614), .A2(n4514), .ZN(n4613) );
  OAI21_X1 U5239 ( .B1(n7998), .B2(n8000), .A(n4616), .ZN(n4615) );
  AOI21_X1 U5240 ( .B1(n8220), .B2(n8160), .A(n8061), .ZN(n4616) );
  OAI21_X1 U5241 ( .B1(n4594), .B2(n4593), .A(n8061), .ZN(n4592) );
  NAND2_X1 U5242 ( .A1(n8020), .A2(n8015), .ZN(n4593) );
  AOI21_X1 U5243 ( .B1(n4595), .B2(n4520), .A(n8169), .ZN(n4594) );
  NAND2_X1 U5244 ( .A1(n4597), .A2(n8039), .ZN(n4596) );
  OAI21_X1 U5245 ( .B1(n4599), .B2(n8148), .A(n4598), .ZN(n4597) );
  AND2_X1 U5246 ( .A1(n8017), .A2(n8147), .ZN(n4598) );
  AOI21_X1 U5247 ( .B1(n8013), .B2(n8146), .A(n8011), .ZN(n4599) );
  OR2_X1 U5248 ( .A1(n8176), .A2(n8170), .ZN(n4601) );
  NAND2_X1 U5249 ( .A1(n8145), .A2(n8151), .ZN(n8023) );
  NAND2_X1 U5250 ( .A1(n4714), .A2(n4713), .ZN(n4712) );
  AND2_X1 U5251 ( .A1(n8473), .A2(n8472), .ZN(n4713) );
  NAND2_X1 U5252 ( .A1(n4609), .A2(n8033), .ZN(n4608) );
  NAND2_X1 U5253 ( .A1(n4707), .A2(n4700), .ZN(n8504) );
  OAI21_X1 U5254 ( .B1(n4708), .B2(n4705), .A(n8523), .ZN(n4707) );
  NOR2_X1 U5255 ( .A1(n4703), .A2(n4701), .ZN(n4700) );
  AOI21_X1 U5256 ( .B1(n8497), .B2(n4709), .A(n4542), .ZN(n4708) );
  AND2_X1 U5257 ( .A1(n4718), .A2(n5595), .ZN(n4717) );
  OR2_X1 U5258 ( .A1(n4722), .A2(n4719), .ZN(n4718) );
  AND2_X1 U5259 ( .A1(n8509), .A2(n8508), .ZN(n4719) );
  NAND2_X1 U5260 ( .A1(n4622), .A2(n8048), .ZN(n8058) );
  NAND2_X1 U5261 ( .A1(n8047), .A2(n4623), .ZN(n4622) );
  AOI21_X1 U5262 ( .B1(n8040), .B2(n8039), .A(n8142), .ZN(n4623) );
  NOR2_X1 U5263 ( .A1(n8668), .A2(n8685), .ZN(n4841) );
  NAND2_X1 U5264 ( .A1(n4819), .A2(n7419), .ZN(n4818) );
  INV_X1 U5265 ( .A(n7420), .ZN(n4819) );
  NAND2_X1 U5266 ( .A1(n8326), .A2(n6492), .ZN(n6496) );
  INV_X1 U5267 ( .A(n8393), .ZN(n4956) );
  OR2_X1 U5268 ( .A1(n8905), .A2(n8524), .ZN(n8521) );
  AND2_X1 U5269 ( .A1(n4841), .A2(n4840), .ZN(n4839) );
  AND2_X1 U5270 ( .A1(n5597), .A2(n5596), .ZN(n5602) );
  OR2_X1 U5271 ( .A1(n8668), .A2(n8284), .ZN(n8516) );
  OR2_X1 U5272 ( .A1(n8940), .A2(n8275), .ZN(n8493) );
  NOR2_X1 U5273 ( .A1(n8886), .A2(n8967), .ZN(n4835) );
  OR2_X1 U5274 ( .A1(n8967), .A2(n8891), .ZN(n8475) );
  OR2_X1 U5275 ( .A1(n8886), .A2(n8860), .ZN(n8470) );
  NAND2_X1 U5276 ( .A1(n6910), .A2(n6391), .ZN(n5649) );
  NAND2_X1 U5277 ( .A1(n8696), .A2(n4841), .ZN(n8666) );
  OR2_X1 U5278 ( .A1(n7801), .A2(n7805), .ZN(n7885) );
  NAND2_X1 U5279 ( .A1(n7661), .A2(n8355), .ZN(n8385) );
  AND2_X1 U5280 ( .A1(n5157), .A2(n5158), .ZN(n5046) );
  INV_X1 U5281 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5158) );
  AND2_X1 U5282 ( .A1(n6257), .A2(n6256), .ZN(n6259) );
  AND2_X1 U5283 ( .A1(n10065), .A2(n6005), .ZN(n5012) );
  INV_X1 U5284 ( .A(n5010), .ZN(n4761) );
  NAND2_X1 U5285 ( .A1(n4621), .A2(n4620), .ZN(n4619) );
  AOI21_X1 U5286 ( .B1(n8069), .B2(n9276), .A(n4493), .ZN(n4621) );
  NAND2_X1 U5287 ( .A1(n8068), .A2(n9523), .ZN(n4620) );
  OR2_X1 U5288 ( .A1(n9284), .A2(n9269), .ZN(n8126) );
  OAI21_X1 U5289 ( .B1(n9261), .B2(n4798), .A(n4510), .ZN(n4797) );
  INV_X1 U5290 ( .A(n9263), .ZN(n4798) );
  NAND2_X1 U5291 ( .A1(n4510), .A2(n4800), .ZN(n4799) );
  INV_X1 U5292 ( .A(n4799), .ZN(n4794) );
  NOR2_X1 U5293 ( .A1(n9536), .A2(n9540), .ZN(n4894) );
  NOR2_X1 U5294 ( .A1(n9259), .A2(n4801), .ZN(n4800) );
  INV_X1 U5295 ( .A(n9262), .ZN(n4801) );
  OR2_X1 U5296 ( .A1(n9536), .A2(n8093), .ZN(n9263) );
  OR2_X1 U5297 ( .A1(n7831), .A2(n10130), .ZN(n8147) );
  OR2_X1 U5298 ( .A1(n9165), .A2(n9081), .ZN(n8160) );
  OR2_X1 U5299 ( .A1(n9166), .A2(n7940), .ZN(n8157) );
  OR2_X1 U5300 ( .A1(n9168), .A2(n7333), .ZN(n8213) );
  AOI21_X1 U5301 ( .B1(n4862), .B2(n4861), .A(n4534), .ZN(n4860) );
  INV_X1 U5302 ( .A(n7688), .ZN(n4861) );
  OAI21_X1 U5303 ( .B1(n7974), .B2(n7973), .A(n7976), .ZN(n7979) );
  XNOR2_X1 U5304 ( .A(n7979), .B(n4994), .ZN(n7977) );
  INV_X1 U5305 ( .A(n7978), .ZN(n4994) );
  NOR2_X1 U5306 ( .A1(n4768), .A2(n4770), .ZN(n4586) );
  AOI21_X1 U5307 ( .B1(n4651), .B2(n4650), .A(n4648), .ZN(n4647) );
  INV_X1 U5308 ( .A(n4650), .ZN(n4649) );
  INV_X1 U5309 ( .A(n5566), .ZN(n4648) );
  NAND2_X1 U5310 ( .A1(n5549), .A2(n5537), .ZN(n4651) );
  OAI21_X1 U5311 ( .B1(n5503), .B2(n5502), .A(n5501), .ZN(n5518) );
  AOI21_X1 U5312 ( .B1(n4976), .B2(n4979), .A(n4655), .ZN(n4654) );
  INV_X1 U5313 ( .A(n5142), .ZN(n4655) );
  INV_X1 U5314 ( .A(n5130), .ZN(n4980) );
  INV_X1 U5315 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4887) );
  NAND2_X1 U5316 ( .A1(n5121), .A2(n5120), .ZN(n5352) );
  AOI21_X1 U5317 ( .B1(n4971), .B2(n4969), .A(n4541), .ZN(n4967) );
  INV_X1 U5318 ( .A(n5323), .ZN(n4971) );
  NAND2_X1 U5319 ( .A1(n5108), .A2(n5107), .ZN(n5111) );
  NAND2_X1 U5320 ( .A1(n4659), .A2(n4662), .ZN(n5105) );
  INV_X1 U5321 ( .A(n4663), .ZN(n4662) );
  NOR2_X1 U5322 ( .A1(n5298), .A2(n4666), .ZN(n4665) );
  INV_X1 U5323 ( .A(n5093), .ZN(n4666) );
  AND2_X1 U5324 ( .A1(n5104), .A2(n5103), .ZN(n5318) );
  INV_X1 U5325 ( .A(n6572), .ZN(n4916) );
  NAND2_X1 U5326 ( .A1(n4817), .A2(n4815), .ZN(n4907) );
  NAND2_X1 U5327 ( .A1(n4516), .A2(n4816), .ZN(n4815) );
  INV_X1 U5328 ( .A(n5057), .ZN(n4817) );
  AND2_X1 U5329 ( .A1(n7485), .A2(n6422), .ZN(n4816) );
  NAND2_X1 U5330 ( .A1(n5183), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5442) );
  INV_X1 U5331 ( .A(n5429), .ZN(n5183) );
  OR2_X1 U5332 ( .A1(n5532), .A2(n5531), .ZN(n5542) );
  AND2_X1 U5333 ( .A1(n6408), .A2(n6405), .ZN(n4911) );
  INV_X1 U5334 ( .A(n7175), .ZN(n6408) );
  NAND2_X1 U5335 ( .A1(n5179), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5310) );
  INV_X1 U5336 ( .A(n5291), .ZN(n5179) );
  NAND2_X1 U5337 ( .A1(n5509), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5532) );
  INV_X1 U5338 ( .A(n5511), .ZN(n5509) );
  OR2_X1 U5339 ( .A1(n5493), .A2(n9955), .ZN(n5511) );
  NAND2_X1 U5340 ( .A1(n4537), .A2(n6438), .ZN(n4809) );
  OR2_X1 U5341 ( .A1(n5442), .A2(n5441), .ZN(n5456) );
  INV_X1 U5342 ( .A(n6467), .ZN(n4808) );
  INV_X1 U5343 ( .A(n8294), .ZN(n4806) );
  NAND2_X1 U5344 ( .A1(n7846), .A2(n4526), .ZN(n8337) );
  INV_X1 U5345 ( .A(n8366), .ZN(n8546) );
  XNOR2_X1 U5346 ( .A(n4992), .B(n8622), .ZN(n8383) );
  NOR2_X1 U5347 ( .A1(n8382), .A2(n8381), .ZN(n4993) );
  NOR2_X1 U5348 ( .A1(n4929), .A2(n4927), .ZN(n4926) );
  OAI21_X1 U5349 ( .B1(n4932), .B2(n8390), .A(n4930), .ZN(n4929) );
  NAND2_X1 U5350 ( .A1(n4932), .A2(n4931), .ZN(n4930) );
  NAND2_X1 U5351 ( .A1(n4935), .A2(n8622), .ZN(n4931) );
  NAND2_X1 U5352 ( .A1(n4487), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4734) );
  OR2_X1 U5353 ( .A1(n5214), .A2(n6800), .ZN(n5193) );
  OR2_X1 U5354 ( .A1(n10038), .A2(n10039), .ZN(n4692) );
  INV_X1 U5355 ( .A(n7783), .ZN(n4689) );
  OR2_X1 U5356 ( .A1(n8920), .A2(n8257), .ZN(n8676) );
  AND2_X1 U5357 ( .A1(n5565), .A2(n5564), .ZN(n8702) );
  NOR2_X1 U5358 ( .A1(n8720), .A2(n8920), .ZN(n8696) );
  NAND2_X1 U5359 ( .A1(n8676), .A2(n8506), .ZN(n8701) );
  AOI21_X1 U5360 ( .B1(n5020), .B2(n5018), .A(n4570), .ZN(n5017) );
  INV_X1 U5361 ( .A(n5024), .ZN(n5018) );
  INV_X1 U5362 ( .A(n5020), .ZN(n5019) );
  INV_X1 U5363 ( .A(n8772), .ZN(n8737) );
  AND2_X1 U5364 ( .A1(n5027), .A2(n8771), .ZN(n5024) );
  NOR2_X1 U5365 ( .A1(n8950), .A2(n8814), .ZN(n5464) );
  OR2_X1 U5366 ( .A1(n8825), .A2(n8842), .ZN(n8800) );
  OR2_X1 U5367 ( .A1(n8823), .A2(n8950), .ZN(n8794) );
  NOR2_X1 U5368 ( .A1(n8834), .A2(n5033), .ZN(n5032) );
  INV_X1 U5369 ( .A(n5415), .ZN(n5033) );
  NAND2_X1 U5370 ( .A1(n5182), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5429) );
  INV_X1 U5371 ( .A(n5409), .ZN(n5182) );
  NOR2_X1 U5372 ( .A1(n7885), .A2(n10079), .ZN(n8881) );
  AOI21_X1 U5373 ( .B1(n5037), .B2(n7797), .A(n4530), .ZN(n5036) );
  OR2_X1 U5374 ( .A1(n8566), .A2(n7805), .ZN(n5370) );
  NOR2_X1 U5375 ( .A1(n8464), .A2(n5038), .ZN(n5037) );
  INV_X1 U5376 ( .A(n5370), .ZN(n5038) );
  OR2_X1 U5377 ( .A1(n7798), .A2(n7797), .ZN(n5039) );
  NAND2_X1 U5378 ( .A1(n7759), .A2(n5349), .ZN(n4922) );
  AND2_X1 U5379 ( .A1(n8461), .A2(n8463), .ZN(n7797) );
  OR2_X1 U5380 ( .A1(n5310), .A2(n5309), .ZN(n5329) );
  NAND2_X1 U5381 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5249) );
  INV_X1 U5382 ( .A(n8890), .ZN(n8815) );
  INV_X1 U5383 ( .A(n8574), .ZN(n7407) );
  AND4_X1 U5384 ( .A1(n5233), .A2(n5232), .A3(n5231), .A4(n5230), .ZN(n7198)
         );
  INV_X1 U5385 ( .A(n10357), .ZN(n8889) );
  NAND2_X1 U5386 ( .A1(n8418), .A2(n10408), .ZN(n8363) );
  OAI22_X1 U5387 ( .A1(n8357), .A2(n9619), .B1(n6719), .B2(n8356), .ZN(n8628)
         );
  OAI211_X1 U5388 ( .C1(n8357), .C2(n6680), .A(n5247), .B(n5246), .ZN(n7362)
         );
  INV_X1 U5389 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4729) );
  INV_X1 U5390 ( .A(n4732), .ZN(n4730) );
  AOI21_X1 U5391 ( .B1(n4744), .B2(n4746), .A(n6243), .ZN(n9036) );
  OR2_X1 U5392 ( .A1(n7274), .A2(n6306), .ZN(n5820) );
  INV_X1 U5393 ( .A(n5001), .ZN(n5000) );
  OAI21_X1 U5394 ( .B1(n6104), .B2(n5002), .A(n9091), .ZN(n5001) );
  INV_X1 U5395 ( .A(n9068), .ZN(n6105) );
  NAND2_X1 U5396 ( .A1(n6105), .A2(n6104), .ZN(n9069) );
  XNOR2_X1 U5397 ( .A(n4579), .B(n7437), .ZN(n5863) );
  NAND2_X1 U5398 ( .A1(n5859), .A2(n5860), .ZN(n4579) );
  AOI21_X1 U5399 ( .B1(n5927), .B2(n5926), .A(n4517), .ZN(n4755) );
  NAND2_X1 U5400 ( .A1(n7381), .A2(n7382), .ZN(n4580) );
  OR2_X1 U5401 ( .A1(n5882), .A2(n7070), .ZN(n5801) );
  NAND2_X1 U5402 ( .A1(n4742), .A2(n4741), .ZN(n4740) );
  INV_X1 U5403 ( .A(n5829), .ZN(n4742) );
  INV_X1 U5404 ( .A(n5828), .ZN(n4741) );
  AND2_X1 U5405 ( .A1(n5829), .A2(n5828), .ZN(n4739) );
  AND2_X1 U5406 ( .A1(n6305), .A2(n6304), .ZN(n9239) );
  OR2_X1 U5407 ( .A1(n4485), .A2(n5788), .ZN(n5792) );
  INV_X1 U5408 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U5409 ( .A1(n6892), .A2(n6893), .ZN(n6964) );
  OR2_X1 U5410 ( .A1(n9169), .A2(n4574), .ZN(n4635) );
  AND2_X1 U5411 ( .A1(n4635), .A2(n4634), .ZN(n10182) );
  INV_X1 U5412 ( .A(n10183), .ZN(n4634) );
  OAI21_X1 U5413 ( .B1(n10209), .B2(n4627), .A(n4626), .ZN(n10219) );
  NAND2_X1 U5414 ( .A1(n4630), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4627) );
  NAND2_X1 U5415 ( .A1(n9174), .A2(n4630), .ZN(n4626) );
  INV_X1 U5416 ( .A(n10220), .ZN(n4630) );
  OR2_X1 U5417 ( .A1(n10209), .A2(n9507), .ZN(n4629) );
  XNOR2_X1 U5418 ( .A(n9178), .B(n9431), .ZN(n9196) );
  AND2_X1 U5419 ( .A1(n4876), .A2(n5059), .ZN(n4874) );
  INV_X1 U5420 ( .A(n4800), .ZN(n4796) );
  AND2_X1 U5421 ( .A1(n4510), .A2(n9263), .ZN(n9314) );
  NAND2_X1 U5422 ( .A1(n9260), .A2(n9262), .ZN(n9337) );
  OAI21_X1 U5423 ( .B1(n9364), .B2(n9365), .A(n9257), .ZN(n9346) );
  INV_X1 U5424 ( .A(n6211), .ZN(n6209) );
  AND3_X1 U5425 ( .A1(n6199), .A2(n6198), .A3(n6197), .ZN(n9377) );
  OAI21_X1 U5426 ( .B1(n9246), .B2(n4776), .A(n4773), .ZN(n9434) );
  INV_X1 U5427 ( .A(n9248), .ZN(n4776) );
  AOI21_X1 U5428 ( .B1(n9248), .B2(n4775), .A(n4774), .ZN(n4773) );
  INV_X1 U5429 ( .A(n9249), .ZN(n4774) );
  NOR2_X1 U5430 ( .A1(n9247), .A2(n4778), .ZN(n4777) );
  AOI21_X1 U5431 ( .B1(n4882), .B2(n4884), .A(n4535), .ZN(n4880) );
  AND2_X1 U5432 ( .A1(n8030), .A2(n9450), .ZN(n9465) );
  OR2_X1 U5433 ( .A1(n9510), .A2(n9220), .ZN(n9221) );
  AND2_X1 U5434 ( .A1(n8178), .A2(n9245), .ZN(n9479) );
  NAND2_X1 U5435 ( .A1(n6086), .A2(n6085), .ZN(n9483) );
  AND4_X1 U5436 ( .A1(n6094), .A2(n6093), .A3(n6092), .A4(n6091), .ZN(n9496)
         );
  OR2_X1 U5437 ( .A1(n9163), .A2(n10312), .ZN(n8006) );
  NAND2_X1 U5438 ( .A1(n7507), .A2(n7468), .ZN(n7469) );
  AND2_X1 U5439 ( .A1(n7444), .A2(n7439), .ZN(n4854) );
  NAND2_X1 U5440 ( .A1(n7305), .A2(n8104), .ZN(n7440) );
  AND2_X1 U5441 ( .A1(n7069), .A2(n8195), .ZN(n10263) );
  AND2_X1 U5442 ( .A1(n7069), .A2(n6958), .ZN(n10264) );
  NAND2_X1 U5443 ( .A1(n7064), .A2(n8105), .ZN(n7261) );
  NOR2_X1 U5444 ( .A1(n7063), .A2(n7273), .ZN(n7065) );
  INV_X1 U5445 ( .A(n10263), .ZN(n10129) );
  INV_X1 U5446 ( .A(n10264), .ZN(n10128) );
  AND2_X1 U5447 ( .A1(n9523), .A2(n10164), .ZN(n4785) );
  INV_X1 U5448 ( .A(n9356), .ZN(n9547) );
  NAND2_X1 U5449 ( .A1(n6110), .A2(n6109), .ZN(n9581) );
  XNOR2_X1 U5450 ( .A(n8071), .B(SI_30_), .ZN(n9026) );
  INV_X1 U5451 ( .A(n7977), .ZN(n8071) );
  NAND2_X1 U5452 ( .A1(n5586), .A2(n5585), .ZN(n5573) );
  XNOR2_X1 U5453 ( .A(n5552), .B(n5549), .ZN(n7789) );
  NAND2_X1 U5454 ( .A1(n5538), .A2(n5537), .ZN(n5552) );
  INV_X1 U5455 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5764) );
  OAI21_X1 U5456 ( .B1(n4503), .B2(n5013), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5765) );
  NAND2_X1 U5457 ( .A1(n5749), .A2(n5769), .ZN(n5013) );
  OAI21_X1 U5458 ( .B1(n4503), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U5459 ( .A1(n4670), .A2(n5469), .ZN(n5486) );
  NAND2_X1 U5460 ( .A1(n4981), .A2(n5130), .ZN(n5403) );
  NAND2_X1 U5461 ( .A1(n5127), .A2(n4982), .ZN(n4981) );
  NAND2_X1 U5462 ( .A1(n5127), .A2(n5126), .ZN(n5386) );
  NAND2_X1 U5463 ( .A1(n4660), .A2(n5093), .ZN(n5299) );
  XNOR2_X1 U5464 ( .A(n5091), .B(SI_7_), .ZN(n5283) );
  XNOR2_X1 U5465 ( .A(n5086), .B(n5085), .ZN(n5268) );
  NAND2_X1 U5466 ( .A1(n5530), .A2(n5529), .ZN(n8722) );
  INV_X1 U5467 ( .A(n8579), .ZN(n8418) );
  INV_X1 U5468 ( .A(n6395), .ZN(n6392) );
  NAND2_X1 U5469 ( .A1(n5490), .A2(n5489), .ZN(n8935) );
  AND4_X1 U5470 ( .A1(n5348), .A2(n5347), .A3(n5346), .A4(n5345), .ZN(n7793)
         );
  AND4_X1 U5471 ( .A1(n5383), .A2(n5382), .A3(n5381), .A4(n5380), .ZN(n8893)
         );
  NAND2_X1 U5472 ( .A1(n7148), .A2(n7147), .ZN(n4912) );
  NAND2_X1 U5473 ( .A1(n5341), .A2(n5340), .ZN(n7766) );
  AND4_X1 U5474 ( .A1(n5282), .A2(n5281), .A3(n5280), .A4(n5279), .ZN(n7625)
         );
  AND4_X1 U5475 ( .A1(n5255), .A2(n5254), .A3(n5253), .A4(n5252), .ZN(n7489)
         );
  INV_X1 U5476 ( .A(n6836), .ZN(n4680) );
  NOR2_X1 U5477 ( .A1(n7094), .A2(n4690), .ZN(n7095) );
  AND2_X1 U5478 ( .A1(n7098), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4690) );
  NAND2_X1 U5479 ( .A1(n7095), .A2(n7096), .ZN(n7166) );
  NAND2_X1 U5480 ( .A1(n8619), .A2(n8618), .ZN(n4699) );
  OAI22_X1 U5481 ( .A1(n8621), .A2(n10347), .B1(n8620), .B2(n10344), .ZN(n4697) );
  NAND2_X1 U5482 ( .A1(n5633), .A2(n5632), .ZN(n7954) );
  AOI21_X1 U5483 ( .B1(n7947), .B2(n10440), .A(n5684), .ZN(n6546) );
  NAND2_X1 U5484 ( .A1(n7927), .A2(n8352), .ZN(n5581) );
  AOI21_X1 U5485 ( .B1(n9139), .B2(n6585), .A(n6584), .ZN(n4759) );
  AND2_X1 U5486 ( .A1(n6253), .A2(n6252), .ZN(n9234) );
  NAND2_X1 U5487 ( .A1(n6153), .A2(n6152), .ZN(n9573) );
  NAND2_X1 U5488 ( .A1(n9107), .A2(n9108), .ZN(n4584) );
  AND4_X1 U5489 ( .A1(n6142), .A2(n6141), .A3(n6140), .A4(n6139), .ZN(n9437)
         );
  AND2_X1 U5490 ( .A1(n6276), .A2(n6275), .ZN(n9350) );
  NAND2_X1 U5491 ( .A1(n4679), .A2(n4676), .ZN(n8205) );
  NOR2_X1 U5492 ( .A1(n8088), .A2(n4677), .ZN(n4676) );
  NAND2_X1 U5493 ( .A1(n4617), .A2(n8190), .ZN(n4679) );
  INV_X1 U5494 ( .A(n9239), .ZN(n9317) );
  NAND2_X1 U5495 ( .A1(n6292), .A2(n6291), .ZN(n9339) );
  INV_X1 U5496 ( .A(n6676), .ZN(n7007) );
  NOR2_X1 U5497 ( .A1(n5780), .A2(n5779), .ZN(n7020) );
  NOR2_X1 U5498 ( .A1(n6762), .A2(n6763), .ZN(n6761) );
  NAND2_X1 U5499 ( .A1(n5748), .A2(n4886), .ZN(n6025) );
  OAI21_X1 U5500 ( .B1(n9196), .B2(n10245), .A(n4641), .ZN(n4640) );
  OR2_X1 U5501 ( .A1(n9197), .A2(n10257), .ZN(n4641) );
  NAND2_X1 U5502 ( .A1(n7988), .A2(n7987), .ZN(n9516) );
  OR2_X1 U5503 ( .A1(n9619), .A2(n6024), .ZN(n7988) );
  AOI21_X1 U5504 ( .B1(n4870), .B2(n4872), .A(n4569), .ZN(n4868) );
  NAND2_X1 U5505 ( .A1(n4789), .A2(n4787), .ZN(n9521) );
  INV_X1 U5506 ( .A(n4788), .ZN(n4787) );
  NAND2_X1 U5507 ( .A1(n4790), .A2(n10266), .ZN(n4789) );
  OAI22_X1 U5508 ( .A1(n9269), .A2(n10129), .B1(n9271), .B2(n9270), .ZN(n4788)
         );
  INV_X1 U5509 ( .A(n7074), .ZN(n8244) );
  NAND2_X1 U5510 ( .A1(n8013), .A2(n8167), .ZN(n4595) );
  NAND2_X1 U5511 ( .A1(n8469), .A2(n8543), .ZN(n4716) );
  NAND2_X1 U5512 ( .A1(n8468), .A2(n8523), .ZN(n4715) );
  OAI21_X1 U5513 ( .B1(n8023), .B2(n8018), .A(n8039), .ZN(n4590) );
  NAND2_X1 U5514 ( .A1(n4601), .A2(n8061), .ZN(n4600) );
  NAND2_X1 U5515 ( .A1(n4711), .A2(n8478), .ZN(n8480) );
  NAND2_X1 U5516 ( .A1(n4712), .A2(n4528), .ZN(n4711) );
  NAND2_X1 U5517 ( .A1(n4608), .A2(n8134), .ZN(n4604) );
  NOR2_X1 U5518 ( .A1(n8037), .A2(n8039), .ZN(n4603) );
  NAND2_X1 U5519 ( .A1(n4608), .A2(n8035), .ZN(n4607) );
  NOR2_X1 U5520 ( .A1(n4710), .A2(n5660), .ZN(n4709) );
  INV_X1 U5521 ( .A(n8495), .ZN(n4710) );
  AOI211_X1 U5522 ( .C1(n8487), .C2(n4706), .A(n4705), .B(n4704), .ZN(n4703)
         );
  NAND2_X1 U5523 ( .A1(n8495), .A2(n8543), .ZN(n4704) );
  AND2_X1 U5524 ( .A1(n8498), .A2(n8493), .ZN(n4706) );
  NAND2_X1 U5525 ( .A1(n8711), .A2(n4702), .ZN(n4701) );
  NAND2_X1 U5526 ( .A1(n5666), .A2(n8543), .ZN(n4702) );
  NAND2_X1 U5527 ( .A1(n4605), .A2(n4602), .ZN(n8042) );
  NAND2_X1 U5528 ( .A1(n4607), .A2(n4606), .ZN(n4605) );
  NAND2_X1 U5529 ( .A1(n4604), .A2(n4603), .ZN(n4602) );
  NOR2_X1 U5530 ( .A1(n8034), .A2(n8061), .ZN(n4606) );
  NAND2_X1 U5531 ( .A1(n7992), .A2(n7991), .ZN(n7995) );
  AND2_X1 U5532 ( .A1(n9260), .A2(n8061), .ZN(n7991) );
  OAI21_X1 U5533 ( .B1(n8511), .B2(n4720), .A(n4717), .ZN(n4721) );
  OR2_X1 U5534 ( .A1(n4722), .A2(n8510), .ZN(n4720) );
  INV_X1 U5535 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5730) );
  NOR2_X1 U5536 ( .A1(n8060), .A2(n8059), .ZN(n8063) );
  NAND2_X1 U5537 ( .A1(n9241), .A2(n8019), .ZN(n8176) );
  AOI21_X1 U5538 ( .B1(n4988), .B2(n4991), .A(n4986), .ZN(n4985) );
  INV_X1 U5539 ( .A(n5623), .ZN(n4986) );
  NOR2_X1 U5540 ( .A1(n5567), .A2(n4564), .ZN(n4650) );
  INV_X1 U5541 ( .A(n4672), .ZN(n4671) );
  OAI21_X1 U5542 ( .B1(n4674), .B2(n4673), .A(n5485), .ZN(n4672) );
  INV_X1 U5543 ( .A(n5469), .ZN(n4673) );
  INV_X1 U5544 ( .A(n5352), .ZN(n4965) );
  NAND2_X1 U5545 ( .A1(n5118), .A2(n5117), .ZN(n5121) );
  OAI21_X1 U5546 ( .B1(n4665), .B2(n4664), .A(n5318), .ZN(n4663) );
  INV_X1 U5547 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4974) );
  INV_X1 U5548 ( .A(n7499), .ZN(n4905) );
  INV_X1 U5549 ( .A(n4900), .ZN(n4899) );
  OAI21_X1 U5550 ( .B1(n6621), .B2(n4901), .A(n6600), .ZN(n4900) );
  INV_X1 U5551 ( .A(n6442), .ZN(n4901) );
  INV_X1 U5552 ( .A(n6433), .ZN(n4811) );
  AND2_X1 U5553 ( .A1(n4934), .A2(n4925), .ZN(n4924) );
  NOR2_X1 U5554 ( .A1(n4927), .A2(n8622), .ZN(n4925) );
  NAND2_X1 U5555 ( .A1(n10436), .A2(n8361), .ZN(n8551) );
  INV_X1 U5556 ( .A(n8551), .ZN(n4927) );
  NAND2_X1 U5557 ( .A1(n8627), .A2(n4939), .ZN(n4936) );
  AOI21_X1 U5558 ( .B1(n4934), .B2(n4937), .A(n4933), .ZN(n4932) );
  INV_X1 U5559 ( .A(n8545), .ZN(n4933) );
  AND2_X1 U5560 ( .A1(n8541), .A2(n4938), .ZN(n4937) );
  INV_X1 U5561 ( .A(n4939), .ZN(n4938) );
  NAND2_X1 U5562 ( .A1(n8628), .A2(n8360), .ZN(n8545) );
  AND2_X1 U5563 ( .A1(n4694), .A2(n4693), .ZN(n10020) );
  NOR2_X1 U5564 ( .A1(n10353), .A2(n10360), .ZN(n4693) );
  INV_X1 U5565 ( .A(n10019), .ZN(n4694) );
  AOI21_X1 U5566 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n8594), .A(n8593), .ZN(
        n8609) );
  NOR2_X1 U5567 ( .A1(n8905), .A2(n4838), .ZN(n4837) );
  INV_X1 U5568 ( .A(n4839), .ZN(n4838) );
  NOR2_X1 U5569 ( .A1(n5055), .A2(n4950), .ZN(n4948) );
  NAND2_X1 U5570 ( .A1(n4850), .A2(n8750), .ZN(n4849) );
  NOR2_X1 U5571 ( .A1(n8940), .A2(n8946), .ZN(n4850) );
  OR2_X1 U5572 ( .A1(n7766), .A2(n7793), .ZN(n8460) );
  INV_X1 U5573 ( .A(n8433), .ZN(n4944) );
  INV_X1 U5574 ( .A(n8432), .ZN(n4945) );
  NOR2_X1 U5575 ( .A1(n6391), .A2(n10408), .ZN(n7200) );
  NAND2_X1 U5576 ( .A1(n5649), .A2(n8363), .ZN(n8410) );
  NOR2_X1 U5577 ( .A1(n6677), .A2(n7982), .ZN(n4831) );
  INV_X1 U5578 ( .A(n5170), .ZN(n4830) );
  NAND2_X1 U5579 ( .A1(n8696), .A2(n8999), .ZN(n8682) );
  NOR2_X1 U5580 ( .A1(n4732), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4731) );
  NAND2_X1 U5581 ( .A1(n4509), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5160) );
  NAND2_X1 U5582 ( .A1(n5159), .A2(n4733), .ZN(n4732) );
  INV_X1 U5583 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4733) );
  INV_X1 U5584 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5159) );
  OR2_X1 U5585 ( .A1(n5000), .A2(n4999), .ZN(n4998) );
  NAND2_X1 U5586 ( .A1(n9068), .A2(n4525), .ZN(n4585) );
  INV_X1 U5587 ( .A(n6127), .ZN(n4999) );
  NOR2_X1 U5588 ( .A1(n10182), .A2(n4632), .ZN(n9171) );
  NOR2_X1 U5589 ( .A1(n4633), .A2(n6031), .ZN(n4632) );
  NAND2_X1 U5590 ( .A1(n9531), .A2(n9239), .ZN(n8128) );
  AND2_X1 U5591 ( .A1(n9304), .A2(n4894), .ZN(n4893) );
  OR2_X1 U5592 ( .A1(n9547), .A2(n9234), .ZN(n8094) );
  INV_X1 U5593 ( .A(n9256), .ZN(n4782) );
  NOR2_X1 U5594 ( .A1(n9252), .A2(n8185), .ZN(n4783) );
  INV_X1 U5595 ( .A(n4777), .ZN(n4775) );
  OR2_X1 U5596 ( .A1(n9164), .A2(n10304), .ZN(n8161) );
  NOR2_X1 U5597 ( .A1(n7562), .A2(n7307), .ZN(n7449) );
  NAND2_X1 U5598 ( .A1(n7267), .A2(n7266), .ZN(n4767) );
  NAND2_X1 U5599 ( .A1(n9413), .A2(n9409), .ZN(n9403) );
  AOI21_X1 U5600 ( .B1(n5578), .B2(n4990), .A(n4989), .ZN(n4988) );
  INV_X1 U5601 ( .A(n5607), .ZN(n4989) );
  INV_X1 U5602 ( .A(n5578), .ZN(n4991) );
  AND2_X1 U5603 ( .A1(n5572), .A2(n5571), .ZN(n5585) );
  NOR2_X1 U5604 ( .A1(n5468), .A2(n4675), .ZN(n4674) );
  INV_X1 U5605 ( .A(n5148), .ZN(n4675) );
  NAND2_X1 U5606 ( .A1(n5123), .A2(n5122), .ZN(n5126) );
  INV_X1 U5607 ( .A(n5111), .ZN(n4970) );
  OR2_X1 U5608 ( .A1(n5945), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5966) );
  INV_X1 U5609 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U5610 ( .A1(n5178), .A2(n5177), .ZN(n5291) );
  AND2_X1 U5611 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5177) );
  INV_X1 U5612 ( .A(n5277), .ZN(n5178) );
  OR2_X1 U5613 ( .A1(n7625), .A2(n8951), .ZN(n6424) );
  INV_X1 U5614 ( .A(n7848), .ZN(n4803) );
  OR2_X1 U5615 ( .A1(n8312), .A2(n8311), .ZN(n6494) );
  NAND2_X1 U5616 ( .A1(n6461), .A2(n8336), .ZN(n8293) );
  NAND2_X1 U5617 ( .A1(n8293), .A2(n8294), .ZN(n8292) );
  INV_X1 U5618 ( .A(n5542), .ZN(n5541) );
  INV_X1 U5619 ( .A(n5478), .ZN(n5477) );
  NAND2_X1 U5620 ( .A1(n5184), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5458) );
  AND2_X1 U5621 ( .A1(n4909), .A2(n4516), .ZN(n7484) );
  NAND2_X1 U5622 ( .A1(n4910), .A2(n6414), .ZN(n4909) );
  AND2_X1 U5623 ( .A1(n5621), .A2(n5620), .ZN(n8524) );
  AND3_X1 U5624 ( .A1(n5515), .A2(n5514), .A3(n5513), .ZN(n8274) );
  AND4_X1 U5625 ( .A1(n5297), .A2(n5296), .A3(n5295), .A4(n5294), .ZN(n7613)
         );
  AOI21_X1 U5626 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7040), .A(n7039), .ZN(
        n8582) );
  AND2_X1 U5627 ( .A1(n7295), .A2(n7294), .ZN(n7296) );
  NAND2_X1 U5628 ( .A1(n7296), .A2(n7297), .ZN(n7394) );
  NAND2_X1 U5629 ( .A1(n7394), .A2(n4684), .ZN(n7396) );
  OR2_X1 U5630 ( .A1(n7395), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4684) );
  NAND2_X1 U5631 ( .A1(n7396), .A2(n7397), .ZN(n7648) );
  OR2_X1 U5632 ( .A1(n5683), .A2(n7954), .ZN(n8634) );
  NAND2_X1 U5633 ( .A1(n4953), .A2(n4951), .ZN(n8648) );
  NAND2_X1 U5634 ( .A1(n4952), .A2(n4956), .ZN(n4951) );
  INV_X1 U5635 ( .A(n4954), .ZN(n4952) );
  NAND2_X1 U5636 ( .A1(n8521), .A2(n8522), .ZN(n8647) );
  INV_X1 U5637 ( .A(n8647), .ZN(n8639) );
  OR2_X1 U5638 ( .A1(n5604), .A2(n5603), .ZN(n5605) );
  NOR2_X1 U5639 ( .A1(n8379), .A2(n4955), .ZN(n4954) );
  INV_X1 U5640 ( .A(n8515), .ZN(n4955) );
  OR2_X1 U5641 ( .A1(n8730), .A2(n8722), .ZN(n8720) );
  NOR2_X1 U5642 ( .A1(n8709), .A2(n5062), .ZN(n8694) );
  NOR2_X1 U5643 ( .A1(n8794), .A2(n4848), .ZN(n8759) );
  INV_X1 U5644 ( .A(n4850), .ZN(n4848) );
  AND2_X1 U5645 ( .A1(n8492), .A2(n8490), .ZN(n8787) );
  NOR2_X1 U5646 ( .A1(n8794), .A2(n8946), .ZN(n8779) );
  OR2_X1 U5647 ( .A1(n8825), .A2(n8803), .ZN(n5448) );
  NAND2_X1 U5648 ( .A1(n8881), .A2(n4532), .ZN(n8823) );
  NAND2_X1 U5649 ( .A1(n8862), .A2(n8475), .ZN(n8839) );
  NAND2_X1 U5650 ( .A1(n8862), .A2(n4949), .ZN(n8841) );
  NAND2_X1 U5651 ( .A1(n8881), .A2(n4835), .ZN(n8867) );
  AND4_X1 U5652 ( .A1(n5435), .A2(n5434), .A3(n5433), .A4(n5432), .ZN(n8859)
         );
  NAND2_X1 U5653 ( .A1(n8881), .A2(n9020), .ZN(n8880) );
  OR2_X1 U5654 ( .A1(n7746), .A2(n7766), .ZN(n7801) );
  NAND2_X1 U5655 ( .A1(n5180), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5343) );
  AND2_X1 U5656 ( .A1(n8449), .A2(n8448), .ZN(n8444) );
  AND2_X1 U5657 ( .A1(n5328), .A2(n5327), .ZN(n7748) );
  AND2_X1 U5658 ( .A1(n4843), .A2(n7411), .ZN(n7745) );
  NOR2_X1 U5659 ( .A1(n4845), .A2(n7675), .ZN(n4843) );
  AND2_X1 U5660 ( .A1(n8440), .A2(n8450), .ZN(n8443) );
  NAND2_X1 U5661 ( .A1(n7370), .A2(n8432), .ZN(n7539) );
  NAND2_X1 U5662 ( .A1(n7539), .A2(n8430), .ZN(n7622) );
  NAND2_X1 U5663 ( .A1(n7411), .A2(n4508), .ZN(n7628) );
  AND2_X1 U5664 ( .A1(n7410), .A2(n7573), .ZN(n7411) );
  NAND2_X1 U5665 ( .A1(n7411), .A2(n7606), .ZN(n7543) );
  NAND2_X1 U5666 ( .A1(n7344), .A2(n4918), .ZN(n7404) );
  NOR2_X1 U5667 ( .A1(n5652), .A2(n4919), .ZN(n4918) );
  INV_X1 U5668 ( .A(n8402), .ZN(n4919) );
  NOR2_X1 U5669 ( .A1(n7353), .A2(n7362), .ZN(n7410) );
  NAND2_X1 U5670 ( .A1(n7200), .A2(n7233), .ZN(n7352) );
  OR2_X1 U5671 ( .A1(n7352), .A2(n7351), .ZN(n7353) );
  NAND2_X1 U5672 ( .A1(n5588), .A2(n5587), .ZN(n8668) );
  NAND2_X1 U5673 ( .A1(n5508), .A2(n5507), .ZN(n8930) );
  NAND2_X1 U5674 ( .A1(n8864), .A2(n5415), .ZN(n8835) );
  INV_X1 U5675 ( .A(n10434), .ZN(n8982) );
  INV_X1 U5676 ( .A(n5046), .ZN(n5045) );
  AND2_X1 U5677 ( .A1(n4962), .A2(n5156), .ZN(n4960) );
  INV_X1 U5678 ( .A(n5696), .ZN(n5705) );
  AND2_X1 U5679 ( .A1(n4960), .A2(n4961), .ZN(n5643) );
  INV_X1 U5680 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5907) );
  AND2_X1 U5681 ( .A1(n4748), .A2(n4747), .ZN(n4746) );
  OR2_X1 U5682 ( .A1(n6224), .A2(n6221), .ZN(n4747) );
  OR2_X1 U5683 ( .A1(n6222), .A2(n4749), .ZN(n4748) );
  INV_X1 U5684 ( .A(n9119), .ZN(n4749) );
  AND2_X1 U5685 ( .A1(n6314), .A2(n6313), .ZN(n6582) );
  NOR2_X1 U5686 ( .A1(n5908), .A2(n5907), .ZN(n5928) );
  INV_X1 U5687 ( .A(n6089), .ZN(n6087) );
  OR2_X1 U5688 ( .A1(n9098), .A2(n9097), .ZN(n5007) );
  NAND2_X1 U5689 ( .A1(n4512), .A2(n4995), .ZN(n7254) );
  INV_X1 U5690 ( .A(n7256), .ZN(n5861) );
  OR2_X1 U5691 ( .A1(n5950), .A2(n5949), .ZN(n5972) );
  INV_X1 U5692 ( .A(n4755), .ZN(n4754) );
  AND2_X1 U5693 ( .A1(n4558), .A2(n4752), .ZN(n4751) );
  NAND2_X1 U5694 ( .A1(n5983), .A2(n4762), .ZN(n7857) );
  NAND2_X1 U5695 ( .A1(n5889), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5908) );
  AND3_X1 U5696 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5889) );
  NAND2_X1 U5697 ( .A1(n6047), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6070) );
  OR2_X1 U5698 ( .A1(n6070), .A2(n6069), .ZN(n6089) );
  INV_X1 U5699 ( .A(n5009), .ZN(n5008) );
  OAI21_X1 U5700 ( .B1(n5010), .B2(n5012), .A(n6042), .ZN(n5009) );
  NAND2_X1 U5701 ( .A1(n4618), .A2(n8083), .ZN(n4617) );
  NAND2_X1 U5702 ( .A1(n4619), .A2(n8193), .ZN(n4618) );
  AND2_X1 U5703 ( .A1(n8085), .A2(n4678), .ZN(n4677) );
  INV_X1 U5704 ( .A(n8190), .ZN(n4678) );
  INV_X1 U5705 ( .A(n4484), .ZN(n6299) );
  NOR2_X1 U5706 ( .A1(n7017), .A2(n7016), .ZN(n7015) );
  OR2_X1 U5707 ( .A1(n6761), .A2(n4631), .ZN(n6729) );
  NOR2_X1 U5708 ( .A1(n6768), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4631) );
  OR2_X1 U5709 ( .A1(n6890), .A2(n4638), .ZN(n6892) );
  OAI22_X1 U5710 ( .A1(n6890), .A2(n4637), .B1(n6893), .B2(n4636), .ZN(n6966)
         );
  NAND2_X1 U5711 ( .A1(n6891), .A2(n6963), .ZN(n4637) );
  INV_X1 U5712 ( .A(n6963), .ZN(n4636) );
  XNOR2_X1 U5713 ( .A(n9171), .B(n9184), .ZN(n10196) );
  NAND2_X1 U5714 ( .A1(n5014), .A2(n5895), .ZN(n6107) );
  AOI21_X1 U5715 ( .B1(n10236), .B2(P1_REG2_REG_17__SCAN_IN), .A(n10231), .ZN(
        n10248) );
  OR2_X1 U5716 ( .A1(n6598), .A2(n6627), .ZN(n6655) );
  XNOR2_X1 U5717 ( .A(n9268), .B(n9267), .ZN(n4790) );
  AND2_X1 U5718 ( .A1(n9351), .A2(n4891), .ZN(n9283) );
  NOR2_X1 U5719 ( .A1(n9284), .A2(n4892), .ZN(n4891) );
  INV_X1 U5720 ( .A(n4893), .ZN(n4892) );
  NAND2_X1 U5721 ( .A1(n4793), .A2(n4791), .ZN(n9306) );
  INV_X1 U5722 ( .A(n4792), .ZN(n4791) );
  OAI21_X1 U5723 ( .B1(n4799), .B2(n4802), .A(n4797), .ZN(n4792) );
  NAND2_X1 U5724 ( .A1(n9264), .A2(n8128), .ZN(n9305) );
  NAND2_X1 U5725 ( .A1(n9351), .A2(n4894), .ZN(n9319) );
  NAND2_X1 U5726 ( .A1(n9351), .A2(n9336), .ZN(n9330) );
  OR2_X1 U5727 ( .A1(n6246), .A2(n9102), .ZN(n6269) );
  AND2_X1 U5728 ( .A1(n4780), .A2(n4779), .ZN(n9364) );
  INV_X1 U5729 ( .A(n4781), .ZN(n4780) );
  NAND2_X1 U5730 ( .A1(n9251), .A2(n4522), .ZN(n4779) );
  OAI21_X1 U5731 ( .B1(n9254), .B2(n4782), .A(n8139), .ZN(n4781) );
  OR2_X1 U5732 ( .A1(n9403), .A2(n9390), .ZN(n9385) );
  OR2_X1 U5733 ( .A1(n9255), .A2(n8097), .ZN(n9380) );
  AND2_X1 U5734 ( .A1(n6208), .A2(n6207), .ZN(n9230) );
  OR2_X1 U5735 ( .A1(n6176), .A2(n9111), .ZN(n6193) );
  OR2_X1 U5736 ( .A1(n6193), .A2(n6192), .ZN(n6211) );
  AND2_X1 U5737 ( .A1(n6218), .A2(n6217), .ZN(n9402) );
  NAND2_X1 U5738 ( .A1(n9251), .A2(n4783), .ZN(n9396) );
  NAND2_X1 U5739 ( .A1(n9396), .A2(n9254), .ZN(n9397) );
  AND2_X1 U5740 ( .A1(n9428), .A2(n9418), .ZN(n9413) );
  NAND2_X1 U5741 ( .A1(n6154), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6176) );
  INV_X1 U5742 ( .A(n6156), .ZN(n6154) );
  OR2_X1 U5743 ( .A1(n6113), .A2(n6112), .ZN(n6137) );
  NAND2_X1 U5744 ( .A1(n6135), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6156) );
  INV_X1 U5745 ( .A(n6137), .ZN(n6135) );
  NAND2_X1 U5746 ( .A1(n9482), .A2(n9464), .ZN(n9458) );
  AND2_X1 U5747 ( .A1(n9473), .A2(n9243), .ZN(n9497) );
  NAND2_X1 U5748 ( .A1(n4890), .A2(n9592), .ZN(n9504) );
  INV_X1 U5749 ( .A(n4890), .ZN(n9502) );
  NAND2_X1 U5750 ( .A1(n10108), .A2(n10113), .ZN(n10107) );
  NAND2_X1 U5751 ( .A1(n4855), .A2(n4856), .ZN(n7832) );
  AOI21_X1 U5752 ( .B1(n4488), .B2(n4863), .A(n4495), .ZN(n4856) );
  NAND2_X1 U5753 ( .A1(n6008), .A2(n6007), .ZN(n7893) );
  AND2_X1 U5754 ( .A1(n10138), .A2(n10066), .ZN(n10119) );
  NOR2_X1 U5755 ( .A1(n5991), .A2(n5990), .ZN(n6010) );
  OR2_X1 U5756 ( .A1(n5972), .A2(n6894), .ZN(n5991) );
  NAND2_X1 U5757 ( .A1(n7834), .A2(n8147), .ZN(n10126) );
  AND4_X1 U5758 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .ZN(n10130)
         );
  OR2_X1 U5759 ( .A1(n10279), .A2(n7831), .ZN(n10139) );
  AND2_X1 U5760 ( .A1(n8014), .A2(n8012), .ZN(n10268) );
  NAND2_X1 U5761 ( .A1(n4888), .A2(n10304), .ZN(n7518) );
  NOR2_X1 U5762 ( .A1(n7518), .A2(n7476), .ZN(n7592) );
  OAI21_X1 U5763 ( .B1(n4854), .B2(n4853), .A(n4852), .ZN(n7508) );
  INV_X1 U5764 ( .A(n7466), .ZN(n4853) );
  AND2_X1 U5765 ( .A1(n8104), .A2(n7466), .ZN(n4851) );
  AND3_X1 U5766 ( .A1(n5878), .A2(n5877), .A3(n5876), .ZN(n9081) );
  NAND2_X1 U5767 ( .A1(n7311), .A2(n8215), .ZN(n8000) );
  INV_X1 U5768 ( .A(n4767), .ZN(n8214) );
  AND3_X2 U5769 ( .A1(n5819), .A2(n5818), .A3(n5817), .ZN(n7274) );
  AND2_X1 U5770 ( .A1(n7061), .A2(n7060), .ZN(n10272) );
  OR2_X1 U5771 ( .A1(n7326), .A2(n7325), .ZN(n7473) );
  NAND2_X1 U5772 ( .A1(n6284), .A2(n6283), .ZN(n9536) );
  NAND2_X1 U5773 ( .A1(n7912), .A2(n8072), .ZN(n6284) );
  NAND2_X1 U5774 ( .A1(n6228), .A2(n6227), .ZN(n9550) );
  NAND2_X1 U5775 ( .A1(n4858), .A2(n4860), .ZN(n10132) );
  NAND2_X1 U5776 ( .A1(n4859), .A2(n4862), .ZN(n4858) );
  INV_X1 U5777 ( .A(n10261), .ZN(n4859) );
  INV_X1 U5778 ( .A(n10323), .ZN(n10164) );
  INV_X1 U5779 ( .A(n7823), .ZN(n6341) );
  OR2_X1 U5780 ( .A1(n6340), .A2(n6339), .ZN(n10287) );
  XNOR2_X1 U5781 ( .A(n7974), .B(n5631), .ZN(n9029) );
  CLKBUF_X1 U5782 ( .A(n6365), .Z(n6958) );
  XNOR2_X1 U5783 ( .A(n5624), .B(n5623), .ZN(n7931) );
  NAND2_X1 U5784 ( .A1(n4984), .A2(n4988), .ZN(n5624) );
  OR2_X1 U5785 ( .A1(n5573), .A2(n4991), .ZN(n4984) );
  NAND2_X1 U5786 ( .A1(n4889), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5774) );
  XNOR2_X1 U5787 ( .A(n5586), .B(n5585), .ZN(n7912) );
  INV_X1 U5788 ( .A(n4645), .ZN(n5568) );
  AOI21_X1 U5789 ( .B1(n5538), .B2(n4646), .A(n4564), .ZN(n4645) );
  INV_X1 U5790 ( .A(n4651), .ZN(n4646) );
  OAI21_X1 U5791 ( .B1(n5127), .B2(n4656), .A(n4654), .ZN(n5437) );
  NAND2_X1 U5792 ( .A1(n4975), .A2(n4978), .ZN(n5417) );
  OR2_X1 U5793 ( .A1(n5127), .A2(n4504), .ZN(n4975) );
  NOR2_X1 U5794 ( .A1(n5747), .A2(n4589), .ZN(n6044) );
  INV_X1 U5795 ( .A(n4885), .ZN(n4589) );
  OAI21_X1 U5796 ( .B1(n4966), .B2(n4971), .A(n5111), .ZN(n5336) );
  INV_X1 U5797 ( .A(n4661), .ZN(n5319) );
  AOI21_X1 U5798 ( .B1(n4660), .B2(n4665), .A(n4664), .ZN(n4661) );
  OR2_X1 U5799 ( .A1(n5935), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U5800 ( .A1(n5076), .A2(n5075), .ZN(n5244) );
  NOR2_X1 U5801 ( .A1(n6547), .A2(n6510), .ZN(n6571) );
  INV_X1 U5802 ( .A(n7846), .ZN(n6456) );
  NAND2_X1 U5803 ( .A1(n6450), .A2(n6449), .ZN(n7847) );
  CLKBUF_X1 U5804 ( .A(n8255), .Z(n8256) );
  AND4_X1 U5805 ( .A1(n5316), .A2(n5315), .A3(n5314), .A4(n5313), .ZN(n7742)
         );
  INV_X1 U5806 ( .A(n7748), .ZN(n8981) );
  NAND2_X1 U5807 ( .A1(n7610), .A2(n6433), .ZN(n6614) );
  AND4_X1 U5808 ( .A1(n5484), .A2(n5483), .A3(n5482), .A4(n5481), .ZN(n8275)
         );
  NAND2_X1 U5809 ( .A1(n4916), .A2(n6510), .ZN(n4914) );
  NAND2_X1 U5810 ( .A1(n4910), .A2(n4908), .ZN(n4902) );
  NAND2_X1 U5811 ( .A1(n6620), .A2(n6621), .ZN(n4898) );
  AND4_X1 U5812 ( .A1(n5414), .A2(n5413), .A3(n5412), .A4(n5411), .ZN(n8891)
         );
  NAND2_X1 U5813 ( .A1(n8292), .A2(n6467), .ZN(n8303) );
  NAND2_X1 U5814 ( .A1(n5540), .A2(n5539), .ZN(n8920) );
  NAND2_X1 U5815 ( .A1(n7789), .A2(n8352), .ZN(n5540) );
  AND4_X1 U5816 ( .A1(n5400), .A2(n5399), .A3(n5398), .A4(n5397), .ZN(n8860)
         );
  AND4_X1 U5817 ( .A1(n5369), .A2(n5368), .A3(n5367), .A4(n5366), .ZN(n7878)
         );
  NAND2_X1 U5818 ( .A1(n4804), .A2(n4805), .ZN(n7968) );
  AOI21_X1 U5819 ( .B1(n4806), .B2(n4807), .A(n4523), .ZN(n4805) );
  OR2_X1 U5820 ( .A1(n6919), .A2(n8890), .ZN(n8342) );
  OR2_X1 U5821 ( .A1(n6919), .A2(n8892), .ZN(n8343) );
  NOR2_X2 U5822 ( .A1(n6532), .A2(n6519), .ZN(n8329) );
  NAND2_X1 U5823 ( .A1(n6526), .A2(n10358), .ZN(n8346) );
  NAND2_X1 U5824 ( .A1(n5407), .A2(n5406), .ZN(n8967) );
  OAI21_X1 U5825 ( .B1(n8549), .B2(n4726), .A(n4724), .ZN(n4723) );
  INV_X1 U5826 ( .A(n8550), .ZN(n4726) );
  NOR2_X1 U5827 ( .A1(n4728), .A2(n4578), .ZN(n4727) );
  INV_X1 U5828 ( .A(n8549), .ZN(n4728) );
  OR2_X1 U5829 ( .A1(n5497), .A2(n5496), .ZN(n8772) );
  INV_X1 U5830 ( .A(n7613), .ZN(n8570) );
  NAND2_X1 U5831 ( .A1(n5674), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4735) );
  OR2_X1 U5832 ( .A1(n5615), .A2(n5212), .ZN(n5219) );
  OR2_X1 U5833 ( .A1(n5229), .A2(n5213), .ZN(n5218) );
  NAND2_X1 U5834 ( .A1(n5195), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5196) );
  OR2_X1 U5835 ( .A1(n5229), .A2(n5202), .ZN(n5208) );
  OR2_X1 U5836 ( .A1(n5615), .A2(n10359), .ZN(n5207) );
  AND2_X1 U5837 ( .A1(n4692), .A2(n4691), .ZN(n6850) );
  INV_X1 U5838 ( .A(n4681), .ZN(n6837) );
  NOR2_X1 U5839 ( .A1(n6835), .A2(n4565), .ZN(n6877) );
  AOI21_X1 U5840 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n6880), .A(n4515), .ZN(
        n6825) );
  AOI21_X1 U5841 ( .B1(n6983), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6979), .ZN(
        n6981) );
  NOR2_X1 U5842 ( .A1(n7045), .A2(n7044), .ZN(n7094) );
  AND2_X1 U5843 ( .A1(n7166), .A2(n7167), .ZN(n7168) );
  NAND2_X1 U5844 ( .A1(n7650), .A2(n8871), .ZN(n7781) );
  OR2_X1 U5845 ( .A1(n7777), .A2(n7776), .ZN(n7813) );
  OR2_X1 U5846 ( .A1(n4688), .A2(n4502), .ZN(n4686) );
  NOR2_X1 U5847 ( .A1(n4502), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4687) );
  OR2_X1 U5848 ( .A1(n5680), .A2(n5679), .ZN(n5681) );
  XNOR2_X1 U5849 ( .A(n8656), .B(n8659), .ZN(n8912) );
  NAND2_X1 U5850 ( .A1(n5668), .A2(n8505), .ZN(n8700) );
  NAND2_X1 U5851 ( .A1(n5016), .A2(n5017), .ZN(n8710) );
  NAND2_X1 U5852 ( .A1(n5022), .A2(n5023), .ZN(n8729) );
  NAND2_X1 U5853 ( .A1(n8758), .A2(n5024), .ZN(n5022) );
  INV_X1 U5854 ( .A(n8935), .ZN(n8750) );
  AND2_X1 U5855 ( .A1(n5025), .A2(n5028), .ZN(n8744) );
  NAND2_X1 U5856 ( .A1(n8758), .A2(n8771), .ZN(n5025) );
  AND2_X1 U5857 ( .A1(n5034), .A2(n4499), .ZN(n8822) );
  NAND2_X1 U5858 ( .A1(n5035), .A2(n5036), .ZN(n8879) );
  NAND2_X1 U5859 ( .A1(n5376), .A2(n5375), .ZN(n10079) );
  NAND2_X1 U5860 ( .A1(n5039), .A2(n5037), .ZN(n7875) );
  NAND2_X1 U5861 ( .A1(n5039), .A2(n5370), .ZN(n7873) );
  NAND2_X1 U5862 ( .A1(n4922), .A2(n8456), .ZN(n7792) );
  NAND2_X1 U5863 ( .A1(n7548), .A2(n5290), .ZN(n7619) );
  NAND2_X1 U5864 ( .A1(n7344), .A2(n8402), .ZN(n7237) );
  OR2_X1 U5865 ( .A1(n10368), .A2(n6527), .ZN(n10358) );
  INV_X1 U5866 ( .A(n8809), .ZN(n10366) );
  OAI211_X1 U5867 ( .C1(n8357), .C2(n6682), .A(n5272), .B(n5271), .ZN(n7603)
         );
  NAND2_X1 U5868 ( .A1(n6565), .A2(n6564), .ZN(n6566) );
  INV_X1 U5869 ( .A(n7959), .ZN(n6564) );
  INV_X1 U5870 ( .A(n7964), .ZN(n6565) );
  INV_X1 U5871 ( .A(n7603), .ZN(n7606) );
  INV_X1 U5872 ( .A(n5175), .ZN(n9031) );
  XNOR2_X1 U5873 ( .A(n5703), .B(n5702), .ZN(n7791) );
  INV_X1 U5874 ( .A(n8554), .ZN(n7661) );
  INV_X1 U5875 ( .A(n8407), .ZN(n8355) );
  INV_X1 U5876 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6687) );
  AND3_X2 U5877 ( .A1(n5919), .A2(n5918), .A3(n5917), .ZN(n10312) );
  AND4_X1 U5878 ( .A1(n6075), .A2(n6074), .A3(n6073), .A4(n6072), .ZN(n10093)
         );
  NAND2_X1 U5879 ( .A1(n6046), .A2(n6045), .ZN(n10096) );
  NAND2_X1 U5880 ( .A1(n5835), .A2(n5834), .ZN(n5839) );
  AND2_X1 U5881 ( .A1(n5938), .A2(n5937), .ZN(n10316) );
  NAND2_X1 U5882 ( .A1(n6191), .A2(n6190), .ZN(n9563) );
  OR2_X1 U5883 ( .A1(n6380), .A2(n8195), .ZN(n10092) );
  OAI21_X1 U5884 ( .B1(n6105), .B2(n5002), .A(n5000), .ZN(n9089) );
  NAND2_X1 U5885 ( .A1(n9069), .A2(n6106), .ZN(n9090) );
  INV_X1 U5886 ( .A(n5005), .ZN(n9101) );
  NAND2_X1 U5887 ( .A1(n4997), .A2(n5944), .ZN(n7706) );
  NAND2_X1 U5888 ( .A1(n4750), .A2(n4755), .ZN(n4997) );
  NAND2_X1 U5889 ( .A1(n7527), .A2(n5926), .ZN(n4750) );
  NAND2_X1 U5890 ( .A1(n6173), .A2(n6172), .ZN(n9566) );
  NAND2_X1 U5891 ( .A1(n6225), .A2(n6222), .ZN(n9118) );
  NAND2_X1 U5892 ( .A1(n6225), .A2(n6224), .ZN(n4745) );
  AND2_X1 U5893 ( .A1(n6362), .A2(n6370), .ZN(n10067) );
  NAND2_X1 U5894 ( .A1(n5983), .A2(n7725), .ZN(n7859) );
  INV_X1 U5895 ( .A(n4739), .ZN(n4738) );
  NAND2_X1 U5896 ( .A1(n6133), .A2(n6132), .ZN(n9578) );
  OR2_X1 U5897 ( .A1(n6380), .A2(n6958), .ZN(n10061) );
  OR2_X1 U5898 ( .A1(n9135), .A2(n9136), .ZN(n4760) );
  AND2_X1 U5899 ( .A1(n6357), .A2(n6364), .ZN(n10101) );
  AND2_X1 U5900 ( .A1(n6319), .A2(n6286), .ZN(n9321) );
  INV_X1 U5901 ( .A(n9402), .ZN(n9366) );
  OR2_X1 U5902 ( .A1(n6376), .A2(n6639), .ZN(n5740) );
  OR2_X1 U5903 ( .A1(n6376), .A2(n5808), .ZN(n5813) );
  OR2_X1 U5904 ( .A1(n8076), .A2(n5789), .ZN(n5791) );
  NAND2_X1 U5905 ( .A1(n4996), .A2(n5776), .ZN(n5854) );
  AND2_X1 U5906 ( .A1(n5727), .A2(n5728), .ZN(n4996) );
  AOI21_X1 U5907 ( .B1(n6633), .B2(n6679), .A(n6948), .ZN(n6752) );
  NAND2_X1 U5908 ( .A1(n6927), .A2(n4567), .ZN(n6762) );
  NOR2_X1 U5909 ( .A1(n6638), .A2(n6637), .ZN(n6890) );
  INV_X1 U5910 ( .A(n4635), .ZN(n10184) );
  INV_X1 U5911 ( .A(n4629), .ZN(n10208) );
  INV_X1 U5912 ( .A(n9174), .ZN(n4628) );
  NAND2_X1 U5913 ( .A1(n8074), .A2(n8073), .ZN(n10146) );
  NAND2_X1 U5914 ( .A1(n4869), .A2(n4873), .ZN(n9282) );
  OAI21_X1 U5915 ( .B1(n9238), .B2(n4872), .A(n4870), .ZN(n9281) );
  INV_X1 U5916 ( .A(n4795), .ZN(n9315) );
  OAI21_X1 U5917 ( .B1(n9345), .B2(n4796), .A(n9260), .ZN(n4795) );
  NOR2_X1 U5918 ( .A1(n9345), .A2(n9259), .ZN(n9338) );
  AND2_X1 U5919 ( .A1(n6245), .A2(n6244), .ZN(n9356) );
  INV_X1 U5920 ( .A(n9230), .ZN(n9390) );
  INV_X1 U5921 ( .A(n9563), .ZN(n9409) );
  NAND2_X1 U5922 ( .A1(n9251), .A2(n9250), .ZN(n9420) );
  NAND2_X1 U5923 ( .A1(n9246), .A2(n4777), .ZN(n9451) );
  OAI21_X1 U5924 ( .B1(n9480), .B2(n4881), .A(n4880), .ZN(n9442) );
  NAND2_X1 U5925 ( .A1(n9246), .A2(n9245), .ZN(n9466) );
  INV_X1 U5926 ( .A(n9581), .ZN(n9464) );
  NOR2_X1 U5927 ( .A1(n9587), .A2(n4884), .ZN(n9457) );
  NOR2_X1 U5928 ( .A1(n9480), .A2(n9479), .ZN(n9587) );
  NAND2_X1 U5929 ( .A1(n6028), .A2(n6027), .ZN(n10122) );
  NAND2_X1 U5930 ( .A1(n4854), .A2(n7440), .ZN(n7467) );
  AND2_X1 U5931 ( .A1(n7440), .A2(n7439), .ZN(n7441) );
  OR2_X1 U5932 ( .A1(n4483), .A2(n7330), .ZN(n9512) );
  NAND2_X1 U5933 ( .A1(n5834), .A2(n5775), .ZN(n5783) );
  OR2_X1 U5934 ( .A1(n4483), .A2(n7331), .ZN(n9484) );
  OR2_X1 U5935 ( .A1(n10325), .A2(n7327), .ZN(n9505) );
  INV_X1 U5936 ( .A(n9521), .ZN(n4786) );
  NOR2_X1 U5937 ( .A1(n9522), .A2(n4785), .ZN(n4784) );
  INV_X2 U5938 ( .A(n10331), .ZN(n10333) );
  XNOR2_X1 U5939 ( .A(n7986), .B(n7985), .ZN(n9619) );
  INV_X1 U5940 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4865) );
  NAND2_X1 U5941 ( .A1(n5608), .A2(n5579), .ZN(n7927) );
  NAND2_X1 U5942 ( .A1(n5573), .A2(n4658), .ZN(n5579) );
  NOR2_X1 U5943 ( .A1(n5578), .A2(n4990), .ZN(n4658) );
  XNOR2_X1 U5944 ( .A(n5758), .B(n5757), .ZN(n7823) );
  OR2_X1 U5945 ( .A1(n5756), .A2(n5755), .ZN(n5758) );
  NAND2_X1 U5946 ( .A1(n5766), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5768) );
  INV_X1 U5947 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9792) );
  INV_X1 U5948 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6726) );
  INV_X1 U5949 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9805) );
  INV_X1 U5950 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6703) );
  INV_X1 U5951 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U5952 ( .A1(n5816), .A2(n4624), .ZN(n6676) );
  AOI22_X1 U5953 ( .A1(n4543), .A2(P1_IR_REG_0__SCAN_IN), .B1(n4625), .B2(
        n5755), .ZN(n4624) );
  NOR2_X1 U5954 ( .A1(n9651), .A2(n10481), .ZN(n10480) );
  AOI21_X1 U5955 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10478), .ZN(n10477) );
  NOR2_X1 U5956 ( .A1(n10477), .A2(n10476), .ZN(n10475) );
  NOR2_X2 U5957 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n10015) );
  INV_X1 U5958 ( .A(n8626), .ZN(n4695) );
  NAND2_X1 U5959 ( .A1(n4697), .A2(n8622), .ZN(n4696) );
  NAND2_X1 U5960 ( .A1(n4699), .A2(n8390), .ZN(n4698) );
  NOR2_X1 U5961 ( .A1(n6544), .A2(n5048), .ZN(n6545) );
  OAI21_X1 U5962 ( .B1(n5724), .B2(n9019), .A(n5723), .ZN(n5725) );
  AOI21_X1 U5963 ( .B1(n8252), .B2(n4610), .A(n8251), .ZN(P1_U3240) );
  AOI211_X1 U5964 ( .C1(n8205), .C2(n4491), .A(n8201), .B(n4576), .ZN(n4610)
         );
  NAND2_X1 U5965 ( .A1(n4642), .A2(n4639), .ZN(P1_U3260) );
  AOI21_X1 U5966 ( .B1(n4640), .B2(n9322), .A(n9204), .ZN(n4639) );
  NAND2_X1 U5967 ( .A1(n9201), .A2(n9200), .ZN(n4642) );
  NOR2_X1 U5968 ( .A1(n9346), .A2(n9347), .ZN(n9345) );
  AND2_X1 U5969 ( .A1(n4860), .A2(n4857), .ZN(n4488) );
  INV_X2 U5970 ( .A(n5814), .ZN(n5852) );
  NAND2_X1 U5971 ( .A1(n4967), .A2(n4965), .ZN(n4489) );
  NAND2_X1 U5972 ( .A1(n8110), .A2(n4864), .ZN(n4863) );
  OR2_X1 U5973 ( .A1(n9540), .A2(n9350), .ZN(n9260) );
  INV_X1 U5974 ( .A(n5882), .ZN(n6308) );
  INV_X1 U5975 ( .A(n6660), .ZN(n5165) );
  AND2_X1 U5976 ( .A1(n7334), .A2(n6598), .ZN(n5814) );
  AND2_X1 U5977 ( .A1(n5696), .A2(n4555), .ZN(n5173) );
  XNOR2_X1 U5978 ( .A(n8685), .B(n8702), .ZN(n8677) );
  INV_X1 U5979 ( .A(n8677), .ZN(n8508) );
  OAI211_X1 U5980 ( .C1(n8356), .C2(n6687), .A(n5307), .B(n5306), .ZN(n7631)
         );
  INV_X1 U5981 ( .A(n8388), .ZN(n4840) );
  NAND4_X1 U5982 ( .A1(n5056), .A2(n5753), .A3(n5752), .A4(n5751), .ZN(n4490)
         );
  AOI21_X1 U5983 ( .B1(n4978), .B2(n4504), .A(n4977), .ZN(n4976) );
  XNOR2_X1 U5984 ( .A(n5144), .B(n5143), .ZN(n5436) );
  INV_X1 U5985 ( .A(n9441), .ZN(n4879) );
  AND2_X1 U5986 ( .A1(n8091), .A2(n8089), .ZN(n4491) );
  NOR2_X1 U5987 ( .A1(n10122), .A2(n10089), .ZN(n4492) );
  AND2_X1 U5988 ( .A1(n8070), .A2(n8039), .ZN(n4493) );
  AND2_X1 U5989 ( .A1(n5005), .A2(n6263), .ZN(n4494) );
  INV_X1 U5990 ( .A(n4884), .ZN(n4883) );
  AND2_X1 U5991 ( .A1(n9483), .A2(n9467), .ZN(n4884) );
  AND2_X1 U5992 ( .A1(n10163), .A2(n9161), .ZN(n4495) );
  NAND2_X1 U5993 ( .A1(n5105), .A2(n5104), .ZN(n5324) );
  INV_X1 U5994 ( .A(n5324), .ZN(n4966) );
  OR2_X1 U5995 ( .A1(n8930), .A2(n8274), .ZN(n8713) );
  AND2_X1 U5996 ( .A1(n4882), .A2(n9441), .ZN(n4496) );
  AND2_X1 U5997 ( .A1(n5734), .A2(n4866), .ZN(n4497) );
  INV_X1 U5998 ( .A(n8878), .ZN(n5040) );
  AND2_X1 U5999 ( .A1(n4835), .A2(n4834), .ZN(n4498) );
  NAND2_X1 U6000 ( .A1(n8850), .A2(n8817), .ZN(n4499) );
  AND2_X1 U6001 ( .A1(n4653), .A2(n5145), .ZN(n4500) );
  AND2_X1 U6002 ( .A1(n4803), .A2(n6449), .ZN(n4501) );
  NAND2_X1 U6003 ( .A1(n7857), .A2(n5012), .ZN(n10064) );
  INV_X1 U6004 ( .A(n10131), .ZN(n4857) );
  INV_X1 U6005 ( .A(n4863), .ZN(n4862) );
  AND2_X1 U6006 ( .A1(n7811), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4502) );
  OR2_X1 U6007 ( .A1(n6107), .A2(n5745), .ZN(n4503) );
  AND2_X1 U6008 ( .A1(n5798), .A2(n6660), .ZN(n5873) );
  CLKBUF_X3 U6009 ( .A(n5873), .Z(n6265) );
  NAND2_X1 U6010 ( .A1(n4917), .A2(n9031), .ZN(n5214) );
  INV_X1 U6011 ( .A(n5222), .ZN(n8356) );
  OR2_X1 U6012 ( .A1(n5402), .A2(n4980), .ZN(n4504) );
  NAND2_X1 U6013 ( .A1(n5776), .A2(n5727), .ZN(n5778) );
  OAI211_X1 U6014 ( .C1(n8357), .C2(n6685), .A(n5289), .B(n5288), .ZN(n7547)
         );
  NAND2_X1 U6015 ( .A1(n5643), .A2(n5157), .ZN(n4505) );
  OR2_X1 U6016 ( .A1(n8320), .A2(n8319), .ZN(n4506) );
  OR3_X1 U6017 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n4507) );
  AND2_X1 U6018 ( .A1(n7606), .A2(n10426), .ZN(n4508) );
  NAND2_X1 U6019 ( .A1(n5696), .A2(n4730), .ZN(n4509) );
  NAND2_X1 U6020 ( .A1(n9536), .A2(n8093), .ZN(n4510) );
  AND2_X1 U6021 ( .A1(n5194), .A2(n5193), .ZN(n4511) );
  AND2_X1 U6022 ( .A1(n5861), .A2(n5846), .ZN(n4512) );
  AND2_X1 U6023 ( .A1(n4833), .A2(n4832), .ZN(n4513) );
  NAND2_X1 U6024 ( .A1(n5174), .A2(n9023), .ZN(n5175) );
  NAND2_X1 U6025 ( .A1(n5557), .A2(n5556), .ZN(n8685) );
  AND2_X1 U6026 ( .A1(n8001), .A2(n8061), .ZN(n4514) );
  NOR2_X1 U6027 ( .A1(n6877), .A2(n6876), .ZN(n4515) );
  NAND2_X1 U6028 ( .A1(n6413), .A2(n6412), .ZN(n4516) );
  INV_X1 U6029 ( .A(n8530), .ZN(n8382) );
  AND2_X1 U6030 ( .A1(n8532), .A2(n8533), .ZN(n8530) );
  NAND4_X1 U6031 ( .A1(n5793), .A2(n5792), .A3(n5791), .A4(n5790), .ZN(n7063)
         );
  AND2_X1 U6032 ( .A1(n8127), .A2(n8131), .ZN(n9267) );
  NOR2_X1 U6033 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5776) );
  AND2_X1 U6034 ( .A1(n7638), .A2(n7637), .ZN(n4517) );
  NAND2_X1 U6035 ( .A1(n5393), .A2(n5392), .ZN(n8886) );
  OR3_X1 U6036 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        n10355), .ZN(n4518) );
  NAND2_X1 U6037 ( .A1(n4745), .A2(n6226), .ZN(n9117) );
  AND2_X1 U6038 ( .A1(n6337), .A2(n8244), .ZN(n7334) );
  AND2_X1 U6039 ( .A1(n8935), .A2(n8772), .ZN(n4519) );
  INV_X1 U6040 ( .A(n9061), .ZN(n5006) );
  AND2_X1 U6041 ( .A1(n8012), .A2(n8146), .ZN(n4520) );
  AND2_X1 U6042 ( .A1(n8821), .A2(n4499), .ZN(n4521) );
  AND2_X1 U6043 ( .A1(n9256), .A2(n4783), .ZN(n4522) );
  AND2_X1 U6044 ( .A1(n6469), .A2(n6468), .ZN(n4523) );
  NAND2_X1 U6045 ( .A1(n5643), .A2(n5046), .ZN(n5641) );
  INV_X1 U6046 ( .A(n7208), .ZN(n6414) );
  INV_X1 U6047 ( .A(n4979), .ZN(n4978) );
  OAI21_X1 U6048 ( .B1(n4982), .B2(n4504), .A(n5136), .ZN(n4979) );
  INV_X1 U6049 ( .A(n6106), .ZN(n5002) );
  NAND2_X1 U6050 ( .A1(n5610), .A2(n5609), .ZN(n8905) );
  NAND2_X1 U6051 ( .A1(n6267), .A2(n6266), .ZN(n9540) );
  NAND2_X1 U6052 ( .A1(n5474), .A2(n5473), .ZN(n8940) );
  AND2_X1 U6053 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n4524) );
  NAND2_X1 U6054 ( .A1(n6316), .A2(n6315), .ZN(n9284) );
  AND2_X1 U6055 ( .A1(n6127), .A2(n6106), .ZN(n4525) );
  AND2_X1 U6056 ( .A1(n8500), .A2(n8505), .ZN(n8711) );
  NAND2_X1 U6057 ( .A1(n9351), .A2(n4893), .ZN(n4895) );
  INV_X1 U6058 ( .A(n9592), .ZN(n9510) );
  AND2_X1 U6059 ( .A1(n6067), .A2(n6066), .ZN(n9592) );
  AND2_X1 U6060 ( .A1(n8466), .A2(n8458), .ZN(n8464) );
  NAND2_X1 U6061 ( .A1(n8696), .A2(n4839), .ZN(n4842) );
  NAND2_X1 U6062 ( .A1(n5440), .A2(n5439), .ZN(n8825) );
  AND2_X1 U6063 ( .A1(n6458), .A2(n6457), .ZN(n4526) );
  AND2_X1 U6064 ( .A1(n4942), .A2(n5290), .ZN(n4527) );
  AND2_X1 U6065 ( .A1(n8476), .A2(n8834), .ZN(n4528) );
  AND2_X1 U6066 ( .A1(n4688), .A2(n7781), .ZN(n4529) );
  INV_X1 U6067 ( .A(n5098), .ZN(n4664) );
  NAND2_X1 U6068 ( .A1(n5095), .A2(n5094), .ZN(n5098) );
  AND2_X1 U6069 ( .A1(n10079), .A2(n8565), .ZN(n4530) );
  AND2_X1 U6070 ( .A1(n4932), .A2(n8622), .ZN(n4531) );
  AND2_X1 U6071 ( .A1(n4498), .A2(n9013), .ZN(n4532) );
  AND2_X1 U6072 ( .A1(n10023), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4533) );
  INV_X1 U6073 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5769) );
  INV_X1 U6074 ( .A(n4969), .ZN(n4968) );
  NOR2_X1 U6075 ( .A1(n5115), .A2(n4970), .ZN(n4969) );
  NOR2_X1 U6076 ( .A1(n7831), .A2(n10265), .ZN(n4534) );
  NOR2_X1 U6077 ( .A1(n9464), .A2(n9478), .ZN(n4535) );
  NAND2_X1 U6078 ( .A1(n8126), .A2(n9266), .ZN(n9289) );
  INV_X1 U6079 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4737) );
  INV_X1 U6080 ( .A(n4845), .ZN(n4844) );
  NAND2_X1 U6081 ( .A1(n4508), .A2(n7715), .ZN(n4845) );
  AND2_X1 U6082 ( .A1(n6445), .A2(n6444), .ZN(n4536) );
  AND2_X1 U6083 ( .A1(n9206), .A2(n8086), .ZN(n8191) );
  OR2_X1 U6084 ( .A1(n6613), .A2(n4811), .ZN(n4537) );
  OR2_X1 U6085 ( .A1(n5324), .A2(n4968), .ZN(n4538) );
  NAND4_X1 U6086 ( .A1(n5156), .A2(n5259), .A3(n5155), .A4(n5029), .ZN(n4539)
         );
  INV_X1 U6087 ( .A(n4882), .ZN(n4881) );
  AOI21_X1 U6088 ( .B1(n9479), .B2(n4883), .A(n9224), .ZN(n4882) );
  INV_X1 U6089 ( .A(n4950), .ZN(n4949) );
  NAND2_X1 U6090 ( .A1(n8834), .A2(n8475), .ZN(n4950) );
  NAND2_X1 U6091 ( .A1(n9578), .A2(n9468), .ZN(n4540) );
  AND2_X1 U6092 ( .A1(n5114), .A2(SI_11_), .ZN(n4541) );
  NAND2_X1 U6093 ( .A1(n8713), .A2(n8498), .ZN(n4542) );
  AND2_X1 U6094 ( .A1(n8354), .A2(n8353), .ZN(n10073) );
  INV_X1 U6095 ( .A(n9347), .ZN(n4802) );
  AND2_X1 U6096 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4543) );
  AND2_X1 U6097 ( .A1(n8477), .A2(n8810), .ZN(n8834) );
  NAND2_X1 U6098 ( .A1(n9305), .A2(n4875), .ZN(n4544) );
  INV_X1 U6099 ( .A(n4935), .ZN(n4934) );
  NAND2_X1 U6100 ( .A1(n8538), .A2(n4936), .ZN(n4935) );
  OR2_X1 U6101 ( .A1(n4519), .A2(n5026), .ZN(n4545) );
  NAND2_X1 U6102 ( .A1(n6298), .A2(n6297), .ZN(n9531) );
  INV_X1 U6103 ( .A(n9531), .ZN(n9304) );
  AND2_X1 U6104 ( .A1(n5671), .A2(n4956), .ZN(n4546) );
  OR2_X1 U6105 ( .A1(n6427), .A2(n6426), .ZN(n4547) );
  AND2_X1 U6106 ( .A1(n5017), .A2(n8714), .ZN(n4548) );
  NOR2_X1 U6107 ( .A1(n6583), .A2(n6582), .ZN(n4549) );
  AND2_X1 U6108 ( .A1(n4746), .A2(n6243), .ZN(n4550) );
  AND2_X1 U6109 ( .A1(n5036), .A2(n5040), .ZN(n4551) );
  AND2_X1 U6110 ( .A1(n5283), .A2(n5098), .ZN(n4552) );
  AND2_X1 U6111 ( .A1(n8661), .A2(n4954), .ZN(n4553) );
  AND2_X1 U6112 ( .A1(n4762), .A2(n4761), .ZN(n4554) );
  AND2_X1 U6113 ( .A1(n4731), .A2(n4729), .ZN(n4555) );
  AND2_X1 U6114 ( .A1(n7611), .A2(n6438), .ZN(n4556) );
  OR2_X1 U6115 ( .A1(n9061), .A2(n9097), .ZN(n4557) );
  AND2_X1 U6116 ( .A1(n5964), .A2(n5944), .ZN(n4558) );
  NOR2_X1 U6117 ( .A1(n8302), .A2(n4808), .ZN(n4807) );
  AND2_X1 U6118 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4559) );
  AND2_X1 U6119 ( .A1(n8470), .A2(n8471), .ZN(n8878) );
  AND2_X1 U6120 ( .A1(n8362), .A2(n8545), .ZN(n4560) );
  OAI21_X1 U6121 ( .B1(n4880), .B2(n4879), .A(n4540), .ZN(n4878) );
  AND2_X1 U6122 ( .A1(n4497), .A2(n4865), .ZN(n4561) );
  AND2_X1 U6123 ( .A1(n4916), .A2(n4915), .ZN(n4562) );
  INV_X1 U6124 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U6125 ( .A1(n4654), .A2(n5436), .ZN(n4563) );
  INV_X1 U6126 ( .A(n6195), .ZN(n6134) );
  INV_X1 U6127 ( .A(n5834), .ZN(n6024) );
  NAND2_X1 U6128 ( .A1(n5581), .A2(n5580), .ZN(n8388) );
  AND2_X1 U6129 ( .A1(n5551), .A2(SI_24_), .ZN(n4564) );
  AND2_X1 U6130 ( .A1(n6840), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4565) );
  INV_X1 U6131 ( .A(n6548), .ZN(n4915) );
  NAND2_X1 U6132 ( .A1(n4582), .A2(n6061), .ZN(n9147) );
  NAND2_X1 U6133 ( .A1(n10064), .A2(n6023), .ZN(n7864) );
  NAND2_X1 U6134 ( .A1(n4898), .A2(n6442), .ZN(n6599) );
  INV_X1 U6135 ( .A(n9245), .ZN(n4778) );
  OR2_X1 U6136 ( .A1(n9119), .A2(n6226), .ZN(n4566) );
  INV_X1 U6137 ( .A(n8499), .ZN(n4705) );
  NAND2_X1 U6138 ( .A1(n6083), .A2(n6082), .ZN(n9068) );
  NAND2_X1 U6139 ( .A1(n7990), .A2(n7989), .ZN(n9523) );
  NAND2_X1 U6140 ( .A1(n7876), .A2(n8458), .ZN(n8888) );
  AND4_X1 U6141 ( .A1(n4961), .A2(n4962), .A3(n5044), .A4(n4958), .ZN(n5696)
         );
  NAND2_X1 U6142 ( .A1(n5455), .A2(n5454), .ZN(n8950) );
  NOR3_X1 U6143 ( .A1(n8794), .A2(n8930), .A3(n4849), .ZN(n4846) );
  NAND2_X1 U6144 ( .A1(n8881), .A2(n4498), .ZN(n4836) );
  OR2_X1 U6145 ( .A1(n6924), .A2(n7515), .ZN(n4567) );
  AND2_X1 U6146 ( .A1(n4629), .A2(n4628), .ZN(n4568) );
  INV_X1 U6147 ( .A(n4847), .ZN(n8745) );
  NOR2_X1 U6148 ( .A1(n8794), .A2(n4849), .ZN(n4847) );
  AND2_X1 U6149 ( .A1(n9284), .A2(n9307), .ZN(n4569) );
  NOR2_X1 U6150 ( .A1(n8930), .A2(n8753), .ZN(n4570) );
  INV_X1 U6151 ( .A(n6891), .ZN(n4638) );
  NAND2_X1 U6152 ( .A1(n6151), .A2(n9126), .ZN(n9044) );
  AND2_X1 U6153 ( .A1(n6220), .A2(n6219), .ZN(n6226) );
  AND2_X1 U6154 ( .A1(n6554), .A2(n6553), .ZN(n4571) );
  NAND2_X1 U6155 ( .A1(n6450), .A2(n4501), .ZN(n7846) );
  AND2_X1 U6156 ( .A1(n7857), .A2(n6005), .ZN(n4572) );
  INV_X1 U6157 ( .A(n5028), .ZN(n5026) );
  NAND2_X1 U6158 ( .A1(n8940), .A2(n8788), .ZN(n5028) );
  INV_X1 U6159 ( .A(n5058), .ZN(n4875) );
  AND2_X1 U6160 ( .A1(n9536), .A2(n9339), .ZN(n5058) );
  INV_X1 U6161 ( .A(n7209), .ZN(n4910) );
  INV_X1 U6162 ( .A(n10187), .ZN(n4633) );
  NAND2_X1 U6163 ( .A1(n5426), .A2(n5425), .ZN(n8850) );
  INV_X1 U6164 ( .A(n8850), .ZN(n4834) );
  AND2_X1 U6165 ( .A1(n7411), .A2(n4844), .ZN(n4573) );
  NAND2_X1 U6166 ( .A1(n4580), .A2(n5906), .ZN(n7527) );
  AND2_X1 U6167 ( .A1(n4810), .A2(n4809), .ZN(n6620) );
  NAND2_X1 U6168 ( .A1(n7704), .A2(n5965), .ZN(n7724) );
  NAND2_X1 U6169 ( .A1(n4902), .A2(n4907), .ZN(n7498) );
  INV_X1 U6170 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5030) );
  INV_X1 U6171 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4765) );
  AND2_X1 U6172 ( .A1(n9179), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4574) );
  INV_X1 U6173 ( .A(n5786), .ZN(n6336) );
  NAND2_X1 U6174 ( .A1(n4995), .A2(n5846), .ZN(n7253) );
  INV_X1 U6175 ( .A(n5572), .ZN(n4990) );
  NAND2_X1 U6176 ( .A1(n4912), .A2(n6405), .ZN(n7172) );
  AND2_X1 U6177 ( .A1(n8438), .A2(n8439), .ZN(n8436) );
  INV_X1 U6178 ( .A(n8436), .ZN(n4942) );
  AND2_X1 U6179 ( .A1(n4813), .A2(n4812), .ZN(n4575) );
  NAND2_X1 U6180 ( .A1(n5748), .A2(n4766), .ZN(n6354) );
  NAND2_X1 U6181 ( .A1(n5161), .A2(n5170), .ZN(n5673) );
  AND2_X2 U6182 ( .A1(n6542), .A2(n6541), .ZN(n10452) );
  NAND2_X1 U6183 ( .A1(n7068), .A2(n7067), .ZN(n10266) );
  NAND2_X1 U6184 ( .A1(n7221), .A2(n5211), .ZN(n7191) );
  AOI21_X1 U6185 ( .B1(n6992), .B2(n4740), .A(n4739), .ZN(n7081) );
  INV_X1 U6186 ( .A(n7262), .ZN(n8100) );
  NAND2_X1 U6187 ( .A1(n8213), .A2(n8217), .ZN(n7262) );
  NAND2_X1 U6188 ( .A1(n8410), .A2(n5650), .ZN(n7194) );
  NAND2_X1 U6189 ( .A1(n7449), .A2(n9081), .ZN(n7516) );
  INV_X1 U6190 ( .A(n7516), .ZN(n4888) );
  OR2_X1 U6191 ( .A1(n8249), .A2(n8244), .ZN(n4576) );
  AND2_X1 U6192 ( .A1(n4738), .A2(n4740), .ZN(n4577) );
  AND2_X1 U6193 ( .A1(n6396), .A2(n6398), .ZN(n7110) );
  INV_X1 U6194 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4625) );
  INV_X1 U6195 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4866) );
  INV_X1 U6196 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6128) );
  INV_X1 U6197 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5727) );
  INV_X1 U6198 ( .A(n9322), .ZN(n9200) );
  OR2_X1 U6199 ( .A1(n8386), .A2(n10407), .ZN(n4578) );
  INV_X1 U6200 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4756) );
  XNOR2_X1 U6201 ( .A(n5863), .B(n5862), .ZN(n7256) );
  OAI21_X2 U6202 ( .B1(n7527), .B2(n4754), .A(n4751), .ZN(n7704) );
  NAND2_X1 U6203 ( .A1(n5772), .A2(n4581), .ZN(n6365) );
  NAND2_X1 U6204 ( .A1(n10100), .A2(n6058), .ZN(n4582) );
  NAND2_X1 U6205 ( .A1(n5983), .A2(n4554), .ZN(n4583) );
  NAND2_X1 U6206 ( .A1(n4736), .A2(n9045), .ZN(n9107) );
  XNOR2_X1 U6207 ( .A(n5886), .B(n5884), .ZN(n9079) );
  NAND2_X1 U6208 ( .A1(n6147), .A2(n6148), .ZN(n9127) );
  NOR2_X2 U6209 ( .A1(n9036), .A2(n9035), .ZN(n9034) );
  NAND3_X1 U6210 ( .A1(n5895), .A2(n5014), .A3(n4586), .ZN(n4889) );
  NAND2_X2 U6211 ( .A1(n5738), .A2(n5739), .ZN(n6376) );
  XNOR2_X2 U6212 ( .A(n4588), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5738) );
  NAND3_X1 U6213 ( .A1(n4600), .A2(n4591), .A3(n4590), .ZN(n8027) );
  NAND3_X1 U6214 ( .A1(n4596), .A2(n4592), .A3(n10131), .ZN(n4591) );
  NAND3_X1 U6215 ( .A1(n8032), .A2(n8031), .A3(n9465), .ZN(n4609) );
  NAND2_X1 U6216 ( .A1(n5773), .A2(n5734), .ZN(n4612) );
  NAND3_X1 U6217 ( .A1(n8107), .A2(n4615), .A3(n4613), .ZN(n8010) );
  NAND3_X1 U6218 ( .A1(n8000), .A2(n7999), .A3(n8101), .ZN(n4614) );
  XNOR2_X1 U6219 ( .A(n9173), .B(n9186), .ZN(n10209) );
  NAND2_X2 U6220 ( .A1(n4644), .A2(n4643), .ZN(n5072) );
  NAND2_X1 U6221 ( .A1(n10015), .A2(n4974), .ZN(n4644) );
  NAND3_X1 U6222 ( .A1(n4644), .A2(n4643), .A3(n4559), .ZN(n4972) );
  OAI21_X1 U6223 ( .B1(n5538), .B2(n4649), .A(n4647), .ZN(n5586) );
  INV_X1 U6224 ( .A(n5127), .ZN(n4652) );
  OAI21_X1 U6225 ( .B1(n4652), .B2(n4563), .A(n4500), .ZN(n5450) );
  NAND3_X1 U6226 ( .A1(n4654), .A2(n4656), .A3(n5436), .ZN(n4653) );
  INV_X1 U6227 ( .A(n4976), .ZN(n4656) );
  INV_X1 U6228 ( .A(n5573), .ZN(n4657) );
  OAI21_X1 U6229 ( .B1(n4657), .B2(n4990), .A(n5578), .ZN(n5608) );
  NAND2_X1 U6230 ( .A1(n5284), .A2(n4552), .ZN(n4659) );
  NAND2_X1 U6231 ( .A1(n5284), .A2(n5283), .ZN(n4660) );
  NAND2_X1 U6232 ( .A1(n5149), .A2(n4671), .ZN(n4669) );
  NAND2_X1 U6233 ( .A1(n5149), .A2(n4674), .ZN(n4670) );
  NAND2_X1 U6234 ( .A1(n5149), .A2(n5148), .ZN(n5467) );
  NAND2_X1 U6235 ( .A1(n4686), .A2(n4685), .ZN(n7810) );
  NAND2_X1 U6236 ( .A1(n7650), .A2(n4687), .ZN(n4685) );
  NAND2_X1 U6237 ( .A1(n7781), .A2(n7782), .ZN(n7784) );
  INV_X1 U6238 ( .A(n4692), .ZN(n10037) );
  NAND2_X1 U6239 ( .A1(n10041), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4691) );
  NOR2_X1 U6240 ( .A1(n10020), .A2(n4533), .ZN(n10039) );
  NAND3_X1 U6241 ( .A1(n4698), .A2(n4696), .A3(n4695), .ZN(P2_U3264) );
  NAND3_X1 U6242 ( .A1(n4716), .A2(n4715), .A3(n8878), .ZN(n4714) );
  NAND2_X1 U6243 ( .A1(n4721), .A2(n8521), .ZN(n8528) );
  NAND2_X1 U6244 ( .A1(n5696), .A2(n4731), .ZN(n5170) );
  NAND2_X1 U6245 ( .A1(n5696), .A2(n5159), .ZN(n5162) );
  NAND4_X1 U6246 ( .A1(n5242), .A2(n5241), .A3(n4735), .A4(n4734), .ZN(n8574)
         );
  NAND2_X1 U6247 ( .A1(n9044), .A2(n9046), .ZN(n4736) );
  INV_X1 U6248 ( .A(n6353), .ZN(n6339) );
  AND2_X2 U6249 ( .A1(n6598), .A2(n5763), .ZN(n5803) );
  NAND3_X2 U6250 ( .A1(n6353), .A2(n7825), .A3(n6341), .ZN(n6598) );
  XNOR2_X2 U6251 ( .A(n5762), .B(n4737), .ZN(n6353) );
  XNOR2_X1 U6252 ( .A(n6992), .B(n4577), .ZN(n6997) );
  INV_X1 U6253 ( .A(n6225), .ZN(n4743) );
  OAI21_X1 U6254 ( .B1(n7527), .B2(n5927), .A(n5926), .ZN(n7636) );
  AND2_X2 U6255 ( .A1(n9139), .A2(n4549), .ZN(n6586) );
  OR2_X2 U6256 ( .A1(n9060), .A2(n4760), .ZN(n9139) );
  NAND2_X1 U6257 ( .A1(n4767), .A2(n8100), .ZN(n7309) );
  XNOR2_X1 U6258 ( .A(n8214), .B(n7262), .ZN(n7270) );
  NAND4_X1 U6259 ( .A1(n4769), .A2(n5769), .A3(n5757), .A4(n6128), .ZN(n4768)
         );
  NAND4_X1 U6260 ( .A1(n4772), .A2(n4771), .A3(n4737), .A4(n9992), .ZN(n4770)
         );
  NAND3_X1 U6261 ( .A1(n9524), .A2(n4786), .A3(n4784), .ZN(n9600) );
  NAND2_X1 U6262 ( .A1(n9346), .A2(n4794), .ZN(n4793) );
  NAND2_X1 U6263 ( .A1(n7846), .A2(n6457), .ZN(n6460) );
  NAND3_X1 U6264 ( .A1(n6461), .A2(n4807), .A3(n8336), .ZN(n4804) );
  NAND3_X1 U6265 ( .A1(n4813), .A2(n4812), .A3(n7611), .ZN(n7610) );
  NAND3_X1 U6266 ( .A1(n4813), .A2(n4812), .A3(n4556), .ZN(n4810) );
  NAND2_X1 U6267 ( .A1(n4904), .A2(n4910), .ZN(n4812) );
  INV_X1 U6268 ( .A(n4903), .ZN(n4813) );
  NAND2_X1 U6269 ( .A1(n4814), .A2(n5268), .ZN(n5088) );
  XNOR2_X1 U6270 ( .A(n4814), .B(n5268), .ZN(n6682) );
  OAI21_X1 U6271 ( .B1(n4821), .B2(n4820), .A(n4571), .ZN(P2_U3242) );
  AOI21_X1 U6272 ( .B1(n6506), .B2(n6505), .A(n4915), .ZN(n4820) );
  AOI21_X1 U6273 ( .B1(n4506), .B2(n6487), .A(n5052), .ZN(n6491) );
  AOI21_X1 U6274 ( .B1(n7968), .B2(n7967), .A(n6473), .ZN(n8265) );
  NAND2_X1 U6275 ( .A1(n5067), .A2(n5066), .ZN(n5221) );
  INV_X1 U6276 ( .A(n8105), .ZN(n7066) );
  NAND2_X1 U6277 ( .A1(n7462), .A2(n7463), .ZN(n7587) );
  OAI21_X1 U6278 ( .B1(n4907), .B2(n4905), .A(n4547), .ZN(n4903) );
  INV_X1 U6279 ( .A(n4908), .ZN(n4906) );
  AOI21_X1 U6280 ( .B1(n8309), .B2(n6494), .A(n5053), .ZN(n6500) );
  NAND2_X1 U6281 ( .A1(n5071), .A2(n5070), .ZN(n5234) );
  XNOR2_X1 U6282 ( .A(n5065), .B(n5064), .ZN(n5199) );
  NAND2_X1 U6283 ( .A1(n4480), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4833) );
  INV_X1 U6284 ( .A(n8552), .ZN(n4828) );
  INV_X1 U6285 ( .A(n4836), .ZN(n8846) );
  NAND2_X1 U6286 ( .A1(n8696), .A2(n4837), .ZN(n5683) );
  INV_X1 U6287 ( .A(n4842), .ZN(n8640) );
  INV_X1 U6288 ( .A(n4846), .ZN(n8730) );
  NAND2_X1 U6289 ( .A1(n7305), .A2(n4851), .ZN(n4852) );
  NAND2_X1 U6290 ( .A1(n4488), .A2(n10261), .ZN(n4855) );
  OAI21_X1 U6291 ( .B1(n10261), .B2(n7689), .A(n7688), .ZN(n7830) );
  NAND2_X1 U6292 ( .A1(n5773), .A2(n4561), .ZN(n9615) );
  NAND2_X1 U6293 ( .A1(n9238), .A2(n4870), .ZN(n4867) );
  AOI21_X1 U6294 ( .B1(n9238), .B2(n5059), .A(n5058), .ZN(n9300) );
  NAND2_X1 U6295 ( .A1(n4867), .A2(n4868), .ZN(n9240) );
  NAND2_X1 U6296 ( .A1(n9238), .A2(n4874), .ZN(n4869) );
  INV_X1 U6297 ( .A(n9480), .ZN(n4877) );
  AOI21_X1 U6298 ( .B1(n4877), .B2(n4496), .A(n4878), .ZN(n9427) );
  INV_X2 U6299 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4886) );
  NAND2_X1 U6300 ( .A1(n5853), .A2(n5834), .ZN(n5858) );
  NAND2_X1 U6301 ( .A1(n5872), .A2(n8072), .ZN(n5878) );
  NAND2_X1 U6302 ( .A1(n5894), .A2(n8072), .ZN(n5899) );
  NAND2_X1 U6303 ( .A1(n6686), .A2(n8072), .ZN(n5938) );
  NAND2_X1 U6304 ( .A1(n6693), .A2(n8072), .ZN(n5948) );
  NAND2_X1 U6305 ( .A1(n6704), .A2(n8072), .ZN(n5971) );
  NAND2_X1 U6306 ( .A1(n6707), .A2(n8072), .ZN(n5989) );
  NAND2_X1 U6307 ( .A1(n6720), .A2(n8072), .ZN(n6008) );
  NOR2_X2 U6308 ( .A1(n9385), .A2(n9550), .ZN(n9360) );
  NOR2_X2 U6309 ( .A1(n7905), .A2(n10096), .ZN(n4890) );
  INV_X1 U6310 ( .A(n4895), .ZN(n9301) );
  NAND2_X1 U6311 ( .A1(n6620), .A2(n4899), .ZN(n4896) );
  NAND2_X1 U6312 ( .A1(n4896), .A2(n4897), .ZN(n6606) );
  NOR2_X1 U6313 ( .A1(n5057), .A2(n7208), .ZN(n4908) );
  NAND2_X1 U6314 ( .A1(n4912), .A2(n4911), .ZN(n7173) );
  NAND2_X1 U6315 ( .A1(n4913), .A2(n4914), .ZN(n6521) );
  NAND3_X1 U6316 ( .A1(n6506), .A2(n4562), .A3(n6505), .ZN(n4913) );
  INV_X2 U6317 ( .A(n10436), .ZN(n8951) );
  NAND2_X1 U6318 ( .A1(n7345), .A2(n8413), .ZN(n7344) );
  NAND2_X1 U6319 ( .A1(n7404), .A2(n8398), .ZN(n7371) );
  NAND2_X1 U6320 ( .A1(n5668), .A2(n4920), .ZN(n8704) );
  NAND2_X1 U6321 ( .A1(n8704), .A2(n8676), .ZN(n5670) );
  NAND2_X1 U6322 ( .A1(n8359), .A2(n4924), .ZN(n4923) );
  NOR2_X1 U6323 ( .A1(n8631), .A2(n8355), .ZN(n4939) );
  NAND2_X1 U6324 ( .A1(n7370), .A2(n4943), .ZN(n4940) );
  NAND2_X1 U6325 ( .A1(n4940), .A2(n4941), .ZN(n7624) );
  NAND2_X1 U6326 ( .A1(n8862), .A2(n4948), .ZN(n4946) );
  NAND2_X1 U6327 ( .A1(n4946), .A2(n4947), .ZN(n5664) );
  NAND2_X1 U6328 ( .A1(n8657), .A2(n4546), .ZN(n4953) );
  NAND2_X1 U6329 ( .A1(n7876), .A2(n4957), .ZN(n8895) );
  NAND3_X1 U6330 ( .A1(n4960), .A2(n4961), .A3(n5044), .ZN(n5694) );
  NAND2_X1 U6331 ( .A1(n4538), .A2(n4967), .ZN(n5353) );
  NAND2_X1 U6332 ( .A1(n5072), .A2(n5063), .ZN(n5796) );
  INV_X1 U6333 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4973) );
  NAND2_X1 U6334 ( .A1(n5573), .A2(n4988), .ZN(n4987) );
  NAND3_X1 U6335 ( .A1(n8538), .A2(n4560), .A3(n4993), .ZN(n4992) );
  NAND2_X1 U6336 ( .A1(n7081), .A2(n7082), .ZN(n4995) );
  NAND2_X2 U6337 ( .A1(n5803), .A2(n7059), .ZN(n5882) );
  XNOR2_X1 U6338 ( .A(n5765), .B(n5764), .ZN(n6335) );
  NAND2_X1 U6339 ( .A1(n5895), .A2(n5733), .ZN(n5747) );
  OAI21_X2 U6340 ( .B1(n7191), .B2(n7193), .A(n5227), .ZN(n7343) );
  OR2_X2 U6341 ( .A1(n8758), .A2(n5019), .ZN(n5016) );
  NAND4_X1 U6342 ( .A1(n5156), .A2(n5259), .A3(n5031), .A4(n5155), .ZN(n5451)
         );
  NAND3_X1 U6343 ( .A1(n5156), .A2(n5155), .A3(n5259), .ZN(n5418) );
  NAND2_X1 U6344 ( .A1(n8864), .A2(n5032), .ZN(n5034) );
  INV_X1 U6345 ( .A(n5034), .ZN(n8837) );
  NAND2_X1 U6346 ( .A1(n5035), .A2(n4551), .ZN(n5047) );
  NAND2_X1 U6347 ( .A1(n8693), .A2(n5548), .ZN(n8675) );
  OAI21_X2 U6348 ( .B1(n8693), .B2(n8508), .A(n5041), .ZN(n8656) );
  NOR2_X2 U6349 ( .A1(n5045), .A2(n4507), .ZN(n5044) );
  AOI21_X1 U6350 ( .B1(n8638), .B2(n8647), .A(n5622), .ZN(n5640) );
  XNOR2_X1 U6351 ( .A(n8638), .B(n8639), .ZN(n8909) );
  AOI21_X2 U6352 ( .B1(n9344), .B2(n9236), .A(n9235), .ZN(n9328) );
  AOI21_X2 U6353 ( .B1(n9359), .B2(n9233), .A(n9232), .ZN(n9344) );
  AOI22_X2 U6354 ( .A1(n9381), .A2(n9231), .B1(n9366), .B2(n9390), .ZN(n9359)
         );
  INV_X1 U6355 ( .A(n8685), .ZN(n8999) );
  INV_X1 U6356 ( .A(n8280), .ZN(n6504) );
  INV_X1 U6357 ( .A(n8367), .ZN(n8413) );
  AOI21_X1 U6358 ( .B1(n8351), .B2(n8532), .A(n8350), .ZN(n8359) );
  AND2_X4 U6359 ( .A1(n5739), .A2(n9625), .ZN(n6195) );
  INV_X1 U6360 ( .A(n8577), .ZN(n6910) );
  OR2_X1 U6361 ( .A1(n6491), .A2(n6490), .ZN(n6492) );
  CLKBUF_X1 U6362 ( .A(n6335), .Z(n8253) );
  NAND2_X1 U6363 ( .A1(n5827), .A2(n7050), .ZN(n6992) );
  OAI22_X2 U6364 ( .A1(n9427), .A2(n9225), .B1(n9454), .B2(n9429), .ZN(n9412)
         );
  OAI22_X1 U6365 ( .A1(n7137), .A2(n7138), .B1(n6401), .B2(n6400), .ZN(n7148)
         );
  NOR2_X2 U6366 ( .A1(n8646), .A2(n5672), .ZN(n8351) );
  AND2_X1 U6367 ( .A1(n10452), .A2(n8982), .ZN(n7604) );
  AND2_X2 U6368 ( .A1(n6542), .A2(n7182), .ZN(n10444) );
  INV_X1 U6369 ( .A(n8464), .ZN(n5384) );
  AND2_X1 U6370 ( .A1(n7954), .A2(n7604), .ZN(n5048) );
  AND2_X1 U6371 ( .A1(n6538), .A2(n6537), .ZN(n5049) );
  AND2_X1 U6372 ( .A1(n6522), .A2(n8329), .ZN(n5050) );
  NOR2_X1 U6373 ( .A1(n5349), .A2(n7755), .ZN(n5051) );
  NOR2_X1 U6374 ( .A1(n6486), .A2(n8272), .ZN(n5052) );
  AND2_X1 U6375 ( .A1(n8312), .A2(n8311), .ZN(n5053) );
  AND2_X1 U6376 ( .A1(n6520), .A2(n5050), .ZN(n5054) );
  NAND2_X1 U6377 ( .A1(n5662), .A2(n5661), .ZN(n5055) );
  AND4_X1 U6378 ( .A1(n9992), .A2(n5750), .A3(n5764), .A4(n5749), .ZN(n5056)
         );
  INV_X1 U6379 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6380 ( .A1(n8421), .A2(n8423), .ZN(n7192) );
  INV_X1 U6381 ( .A(n9566), .ZN(n9418) );
  OR2_X1 U6382 ( .A1(n9536), .A2(n9339), .ZN(n5059) );
  INV_X1 U6383 ( .A(n8257), .ZN(n8562) );
  AND3_X1 U6384 ( .A1(n5546), .A2(n5545), .A3(n5544), .ZN(n8257) );
  INV_X1 U6385 ( .A(n7797), .ZN(n8372) );
  INV_X1 U6386 ( .A(n8377), .ZN(n8735) );
  AND2_X1 U6387 ( .A1(n7766), .A2(n8567), .ZN(n5061) );
  INV_X1 U6388 ( .A(n8920), .ZN(n5547) );
  XNOR2_X1 U6389 ( .A(n8920), .B(n6513), .ZN(n8312) );
  AND2_X1 U6390 ( .A1(n8722), .A2(n6933), .ZN(n5062) );
  INV_X1 U6391 ( .A(n8061), .ZN(n8039) );
  NAND2_X1 U6392 ( .A1(n8046), .A2(n8061), .ZN(n8047) );
  OAI21_X1 U6393 ( .B1(n8312), .B2(n8562), .A(n8310), .ZN(n6497) );
  INV_X1 U6394 ( .A(n6497), .ZN(n6498) );
  NAND2_X1 U6395 ( .A1(n6392), .A2(n6393), .ZN(n6396) );
  INV_X1 U6396 ( .A(n6306), .ZN(n6317) );
  INV_X1 U6397 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5734) );
  NOR2_X1 U6398 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5753) );
  INV_X1 U6399 ( .A(n5456), .ZN(n5184) );
  NAND2_X1 U6400 ( .A1(n5547), .A2(n8257), .ZN(n5548) );
  INV_X1 U6401 ( .A(n5249), .ZN(n5176) );
  INV_X1 U6402 ( .A(n6598), .ZN(n5799) );
  INV_X1 U6403 ( .A(n6269), .ZN(n6268) );
  NAND2_X1 U6404 ( .A1(n8125), .A2(n8039), .ZN(n8087) );
  INV_X1 U6405 ( .A(n6231), .ZN(n6229) );
  INV_X1 U6406 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6894) );
  INV_X1 U6407 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5949) );
  OR2_X1 U6408 ( .A1(n5395), .A2(n9755), .ZN(n5409) );
  INV_X1 U6409 ( .A(n5329), .ZN(n5180) );
  INV_X1 U6410 ( .A(n5363), .ZN(n5181) );
  NAND2_X1 U6411 ( .A1(n5541), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U6412 ( .A1(n5477), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5493) );
  OR2_X1 U6413 ( .A1(n5458), .A2(n5185), .ZN(n5478) );
  INV_X1 U6414 ( .A(n10073), .ZN(n8627) );
  NAND2_X1 U6415 ( .A1(n5176), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5277) );
  OR2_X1 U6416 ( .A1(n5304), .A2(n5303), .ZN(n5317) );
  INV_X1 U6417 ( .A(n7707), .ZN(n5964) );
  NAND2_X1 U6418 ( .A1(n8087), .A2(n8091), .ZN(n8088) );
  NAND2_X1 U6419 ( .A1(n6229), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U6420 ( .A1(n6209), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U6421 ( .A1(n6087), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6113) );
  INV_X1 U6422 ( .A(n7444), .ZN(n8101) );
  INV_X2 U6423 ( .A(n6024), .ZN(n8072) );
  OR2_X1 U6424 ( .A1(n8204), .A2(n8242), .ZN(n6367) );
  NAND2_X1 U6425 ( .A1(n5133), .A2(n5132), .ZN(n5136) );
  INV_X1 U6426 ( .A(n5335), .ZN(n5115) );
  AND2_X1 U6427 ( .A1(n6479), .A2(n6478), .ZN(n8264) );
  OAI21_X1 U6428 ( .B1(n6512), .B2(n6511), .A(n6522), .ZN(n6572) );
  NAND2_X1 U6429 ( .A1(n5181), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5378) );
  OR2_X1 U6430 ( .A1(n5378), .A2(n7282), .ZN(n5395) );
  OR2_X1 U6431 ( .A1(n5343), .A2(n5342), .ZN(n5363) );
  OR2_X1 U6432 ( .A1(n6528), .A2(n10368), .ZN(n6532) );
  AND3_X1 U6433 ( .A1(n5536), .A2(n5535), .A3(n5534), .ZN(n8738) );
  AND2_X1 U6434 ( .A1(n8559), .A2(n8630), .ZN(n5679) );
  OR2_X1 U6435 ( .A1(n7736), .A2(n8444), .ZN(n7756) );
  OR2_X1 U6436 ( .A1(n10436), .A2(n8622), .ZN(n6527) );
  INV_X1 U6437 ( .A(n7576), .ZN(n7573) );
  OR2_X1 U6438 ( .A1(n8385), .A2(n6533), .ZN(n10434) );
  INV_X1 U6439 ( .A(n7192), .ZN(n7193) );
  AND2_X1 U6440 ( .A1(n6029), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6047) );
  INV_X1 U6441 ( .A(n5852), .ZN(n6309) );
  AND2_X1 U6442 ( .A1(n8244), .A2(n9322), .ZN(n8242) );
  OR2_X1 U6443 ( .A1(n6888), .A2(n6887), .ZN(n6974) );
  OR2_X1 U6444 ( .A1(n6650), .A2(n7924), .ZN(n6654) );
  NOR2_X1 U6445 ( .A1(n9566), .A2(n9226), .ZN(n9227) );
  AND2_X1 U6446 ( .A1(n8019), .A2(n8151), .ZN(n10113) );
  INV_X1 U6447 ( .A(n6958), .ZN(n8195) );
  INV_X1 U6448 ( .A(n9223), .ZN(n9478) );
  INV_X1 U6449 ( .A(n10266), .ZN(n9477) );
  OR2_X1 U6450 ( .A1(n7329), .A2(n8242), .ZN(n10323) );
  AND2_X1 U6451 ( .A1(n5111), .A2(n5110), .ZN(n5323) );
  INV_X2 U6452 ( .A(n5072), .ZN(n6660) );
  OAI21_X1 U6453 ( .B1(n4840), .B2(n8335), .A(n6578), .ZN(n6579) );
  NAND2_X1 U6454 ( .A1(n6530), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8341) );
  INV_X1 U6455 ( .A(n6552), .ZN(n6553) );
  INV_X1 U6456 ( .A(n8816), .ZN(n8892) );
  AND4_X1 U6457 ( .A1(n5447), .A2(n5446), .A3(n5445), .A4(n5444), .ZN(n8842)
         );
  AND2_X1 U6458 ( .A1(n7756), .A2(n7737), .ZN(n8980) );
  INV_X1 U6459 ( .A(n10362), .ZN(n8885) );
  AND2_X1 U6460 ( .A1(n5719), .A2(n6516), .ZN(n6542) );
  NOR2_X1 U6461 ( .A1(n5708), .A2(n7914), .ZN(n10369) );
  INV_X1 U6462 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5166) );
  AND2_X1 U6463 ( .A1(n6010), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6029) );
  INV_X1 U6464 ( .A(n10061), .ZN(n10090) );
  INV_X1 U6465 ( .A(n10092), .ZN(n9152) );
  INV_X1 U6466 ( .A(n9146), .ZN(n10095) );
  AND2_X1 U6467 ( .A1(n6328), .A2(n6327), .ZN(n9269) );
  AND4_X1 U6468 ( .A1(n6015), .A2(n6014), .A3(n6013), .A4(n6012), .ZN(n10127)
         );
  AND2_X1 U6469 ( .A1(n6652), .A2(n6651), .ZN(n10238) );
  INV_X1 U6470 ( .A(n9516), .ZN(n9206) );
  INV_X1 U6471 ( .A(n9305), .ZN(n9299) );
  AND2_X1 U6472 ( .A1(n8135), .A2(n9250), .ZN(n9435) );
  INV_X1 U6473 ( .A(n7845), .ZN(n10283) );
  INV_X1 U6474 ( .A(n9484), .ZN(n10276) );
  AND2_X1 U6475 ( .A1(n10272), .A2(n10170), .ZN(n10298) );
  OR2_X1 U6476 ( .A1(n6902), .A2(n7326), .ZN(n7079) );
  AND2_X1 U6477 ( .A1(n5969), .A2(n5984), .ZN(n6962) );
  INV_X4 U6478 ( .A(n6660), .ZN(n7982) );
  INV_X1 U6479 ( .A(n10026), .ZN(n10350) );
  INV_X1 U6480 ( .A(n7675), .ZN(n10429) );
  INV_X1 U6481 ( .A(n8346), .ZN(n8335) );
  INV_X1 U6482 ( .A(n8329), .ZN(n8348) );
  AOI21_X1 U6483 ( .B1(n8669), .B2(n5195), .A(n5594), .ZN(n8284) );
  OR2_X1 U6484 ( .A1(n8877), .A2(n7199), .ZN(n10362) );
  AND2_X1 U6485 ( .A1(n7202), .A2(n10358), .ZN(n8877) );
  OR2_X1 U6486 ( .A1(n8877), .A2(n7190), .ZN(n8809) );
  INV_X1 U6487 ( .A(n7604), .ZN(n8979) );
  INV_X1 U6488 ( .A(n10452), .ZN(n10450) );
  INV_X1 U6489 ( .A(n5725), .ZN(n5726) );
  INV_X1 U6490 ( .A(n10444), .ZN(n10442) );
  CLKBUF_X1 U6491 ( .A(n10383), .Z(n10405) );
  INV_X1 U6492 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6786) );
  AND2_X1 U6493 ( .A1(n6371), .A2(n6370), .ZN(n10106) );
  INV_X1 U6494 ( .A(n10101), .ZN(n9156) );
  INV_X1 U6495 ( .A(n9269), .ZN(n9307) );
  INV_X1 U6496 ( .A(n9350), .ZN(n9316) );
  INV_X1 U6497 ( .A(n10130), .ZN(n10265) );
  INV_X1 U6498 ( .A(n9195), .ZN(n10245) );
  INV_X1 U6499 ( .A(n10238), .ZN(n10257) );
  OR2_X1 U6500 ( .A1(P1_U3083), .A2(n6656), .ZN(n10260) );
  OR2_X1 U6501 ( .A1(n4483), .A2(n7438), .ZN(n9481) );
  OR2_X1 U6502 ( .A1(n7079), .A2(n7078), .ZN(n10339) );
  INV_X2 U6503 ( .A(n10339), .ZN(n10341) );
  OR4_X1 U6504 ( .A1(n9591), .A2(n9590), .A3(n9589), .A4(n9588), .ZN(n9613) );
  OR2_X1 U6505 ( .A1(n7079), .A2(n7324), .ZN(n10331) );
  AND2_X1 U6506 ( .A1(n6598), .A2(n6356), .ZN(n10288) );
  INV_X1 U6507 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9804) );
  INV_X1 U6508 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6709) );
  NOR2_X1 U6509 ( .A1(n10483), .A2(n10482), .ZN(n10481) );
  NOR2_X1 U6510 ( .A1(n10480), .A2(n10479), .ZN(n10478) );
  OAI21_X1 U6511 ( .B1(n6546), .B2(n10450), .A(n6545), .ZN(P2_U3549) );
  OAI21_X1 U6512 ( .B1(n6546), .B2(n10442), .A(n5726), .ZN(P2_U3517) );
  INV_X1 U6513 ( .A(n9159), .ZN(P1_U4006) );
  AND2_X1 U6514 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5063) );
  INV_X1 U6515 ( .A(SI_1_), .ZN(n5064) );
  MUX2_X1 U6516 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5072), .Z(n5198) );
  NAND2_X1 U6517 ( .A1(n5199), .A2(n5198), .ZN(n5067) );
  NAND2_X1 U6518 ( .A1(n5065), .A2(SI_1_), .ZN(n5066) );
  MUX2_X1 U6519 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5072), .Z(n5069) );
  INV_X1 U6520 ( .A(SI_2_), .ZN(n5068) );
  XNOR2_X1 U6521 ( .A(n5069), .B(n5068), .ZN(n5220) );
  NAND2_X1 U6522 ( .A1(n5221), .A2(n5220), .ZN(n5071) );
  NAND2_X1 U6523 ( .A1(n5069), .A2(SI_2_), .ZN(n5070) );
  MUX2_X1 U6524 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5165), .Z(n5074) );
  INV_X1 U6525 ( .A(SI_3_), .ZN(n5073) );
  NAND2_X1 U6526 ( .A1(n5234), .A2(n5235), .ZN(n5076) );
  NAND2_X1 U6527 ( .A1(n5074), .A2(SI_3_), .ZN(n5075) );
  MUX2_X1 U6528 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5165), .Z(n5078) );
  INV_X1 U6529 ( .A(SI_4_), .ZN(n5077) );
  XNOR2_X1 U6530 ( .A(n5078), .B(n5077), .ZN(n5243) );
  NAND2_X1 U6531 ( .A1(n5244), .A2(n5243), .ZN(n5080) );
  NAND2_X1 U6532 ( .A1(n5078), .A2(SI_4_), .ZN(n5079) );
  MUX2_X1 U6533 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7982), .Z(n5082) );
  INV_X1 U6534 ( .A(SI_5_), .ZN(n5081) );
  XNOR2_X1 U6535 ( .A(n5082), .B(n5081), .ZN(n5256) );
  NAND2_X1 U6536 ( .A1(n5257), .A2(n5256), .ZN(n5084) );
  NAND2_X1 U6537 ( .A1(n5082), .A2(SI_5_), .ZN(n5083) );
  MUX2_X1 U6538 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7982), .Z(n5086) );
  INV_X1 U6539 ( .A(SI_6_), .ZN(n5085) );
  NAND2_X1 U6540 ( .A1(n5086), .A2(SI_6_), .ZN(n5087) );
  INV_X1 U6541 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n5090) );
  INV_X1 U6542 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5089) );
  MUX2_X1 U6543 ( .A(n5090), .B(n5089), .S(n7982), .Z(n5091) );
  INV_X1 U6544 ( .A(n5091), .ZN(n5092) );
  NAND2_X1 U6545 ( .A1(n5092), .A2(SI_7_), .ZN(n5093) );
  MUX2_X1 U6546 ( .A(n6687), .B(n9987), .S(n7982), .Z(n5095) );
  INV_X1 U6547 ( .A(SI_8_), .ZN(n5094) );
  INV_X1 U6548 ( .A(n5095), .ZN(n5096) );
  NAND2_X1 U6549 ( .A1(n5096), .A2(SI_8_), .ZN(n5097) );
  INV_X1 U6550 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5099) );
  MUX2_X1 U6551 ( .A(n5099), .B(n6703), .S(n7982), .Z(n5101) );
  INV_X1 U6552 ( .A(SI_9_), .ZN(n5100) );
  NAND2_X1 U6553 ( .A1(n5101), .A2(n5100), .ZN(n5104) );
  INV_X1 U6554 ( .A(n5101), .ZN(n5102) );
  NAND2_X1 U6555 ( .A1(n5102), .A2(SI_9_), .ZN(n5103) );
  INV_X1 U6556 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5106) );
  MUX2_X1 U6557 ( .A(n5106), .B(n6709), .S(n7982), .Z(n5108) );
  INV_X1 U6558 ( .A(SI_10_), .ZN(n5107) );
  INV_X1 U6559 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U6560 ( .A1(n5109), .A2(SI_10_), .ZN(n5110) );
  INV_X1 U6561 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5112) );
  MUX2_X1 U6562 ( .A(n5112), .B(n9805), .S(n7982), .Z(n5113) );
  INV_X1 U6563 ( .A(n5113), .ZN(n5114) );
  INV_X1 U6564 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5116) );
  MUX2_X1 U6565 ( .A(n5116), .B(n6726), .S(n7982), .Z(n5118) );
  INV_X1 U6566 ( .A(SI_12_), .ZN(n5117) );
  INV_X1 U6567 ( .A(n5118), .ZN(n5119) );
  NAND2_X1 U6568 ( .A1(n5119), .A2(SI_12_), .ZN(n5120) );
  MUX2_X1 U6569 ( .A(n6786), .B(n9792), .S(n7982), .Z(n5123) );
  INV_X1 U6570 ( .A(SI_13_), .ZN(n5122) );
  INV_X1 U6571 ( .A(n5123), .ZN(n5124) );
  NAND2_X1 U6572 ( .A1(n5124), .A2(SI_13_), .ZN(n5125) );
  MUX2_X1 U6573 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7982), .Z(n5129) );
  INV_X1 U6574 ( .A(SI_14_), .ZN(n5128) );
  NAND2_X1 U6575 ( .A1(n5129), .A2(SI_14_), .ZN(n5130) );
  INV_X1 U6576 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7027) );
  INV_X1 U6577 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7025) );
  MUX2_X1 U6578 ( .A(n7027), .B(n7025), .S(n7982), .Z(n5133) );
  INV_X1 U6579 ( .A(SI_15_), .ZN(n5132) );
  INV_X1 U6580 ( .A(n5133), .ZN(n5134) );
  NAND2_X1 U6581 ( .A1(n5134), .A2(SI_15_), .ZN(n5135) );
  INV_X1 U6582 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5137) );
  MUX2_X1 U6583 ( .A(n5137), .B(n9804), .S(n7982), .Z(n5139) );
  INV_X1 U6584 ( .A(SI_16_), .ZN(n5138) );
  NAND2_X1 U6585 ( .A1(n5139), .A2(n5138), .ZN(n5142) );
  INV_X1 U6586 ( .A(n5139), .ZN(n5140) );
  NAND2_X1 U6587 ( .A1(n5140), .A2(SI_16_), .ZN(n5141) );
  MUX2_X1 U6588 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n7982), .Z(n5144) );
  INV_X1 U6589 ( .A(SI_17_), .ZN(n5143) );
  NAND2_X1 U6590 ( .A1(n5144), .A2(SI_17_), .ZN(n5145) );
  MUX2_X1 U6591 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7982), .Z(n5147) );
  XNOR2_X1 U6592 ( .A(n5147), .B(SI_18_), .ZN(n5449) );
  INV_X1 U6593 ( .A(n5449), .ZN(n5146) );
  NAND2_X1 U6594 ( .A1(n5450), .A2(n5146), .ZN(n5149) );
  NAND2_X1 U6595 ( .A1(n5147), .A2(SI_18_), .ZN(n5148) );
  INV_X1 U6596 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7321) );
  INV_X1 U6597 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9950) );
  MUX2_X1 U6598 ( .A(n7321), .B(n9950), .S(n7982), .Z(n5150) );
  INV_X1 U6599 ( .A(SI_19_), .ZN(n9742) );
  NAND2_X1 U6600 ( .A1(n5150), .A2(n9742), .ZN(n5469) );
  INV_X1 U6601 ( .A(n5150), .ZN(n5151) );
  NAND2_X1 U6602 ( .A1(n5151), .A2(SI_19_), .ZN(n5152) );
  NAND2_X1 U6603 ( .A1(n5469), .A2(n5152), .ZN(n5468) );
  XNOR2_X1 U6604 ( .A(n5467), .B(n5468), .ZN(n7320) );
  NAND2_X1 U6605 ( .A1(n5162), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5163) );
  NAND2_X1 U6606 ( .A1(n7320), .A2(n8352), .ZN(n5169) );
  NAND2_X1 U6607 ( .A1(n4539), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5167) );
  XNOR2_X1 U6608 ( .A(n5167), .B(n5166), .ZN(n8622) );
  INV_X1 U6609 ( .A(n8622), .ZN(n8390) );
  AOI22_X1 U6610 ( .A1(n5222), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5453), .B2(
        n8390), .ZN(n5168) );
  INV_X1 U6611 ( .A(n8946), .ZN(n8782) );
  XNOR2_X2 U6612 ( .A(n5171), .B(P2_IR_REG_30__SCAN_IN), .ZN(n9027) );
  NAND2_X1 U6613 ( .A1(n5170), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5172) );
  INV_X1 U6614 ( .A(n5173), .ZN(n9023) );
  NAND2_X1 U6615 ( .A1(n5634), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5191) );
  INV_X1 U6616 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5342) );
  INV_X1 U6617 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7282) );
  INV_X1 U6618 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9755) );
  INV_X1 U6619 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5441) );
  INV_X1 U6620 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6621 ( .A1(n5458), .A2(n5185), .ZN(n5186) );
  NAND2_X1 U6622 ( .A1(n5478), .A2(n5186), .ZN(n8267) );
  OR2_X1 U6623 ( .A1(n5615), .A2(n8267), .ZN(n5190) );
  INV_X1 U6624 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5187) );
  OR2_X1 U6625 ( .A1(n5637), .A2(n5187), .ZN(n5189) );
  INV_X1 U6626 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8612) );
  OR2_X1 U6627 ( .A1(n5476), .A2(n8612), .ZN(n5188) );
  NAND4_X1 U6628 ( .A1(n5191), .A2(n5190), .A3(n5189), .A4(n5188), .ZN(n8804)
         );
  INV_X1 U6629 ( .A(n8804), .ZN(n8321) );
  INV_X1 U6630 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5192) );
  OR2_X1 U6631 ( .A1(n5229), .A2(n5192), .ZN(n5197) );
  NAND2_X1 U6632 ( .A1(n5591), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5194) );
  INV_X1 U6633 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6800) );
  XNOR2_X1 U6634 ( .A(n5199), .B(n5198), .ZN(n6677) );
  NAND2_X1 U6635 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n10355), .ZN(n5200) );
  NAND2_X1 U6636 ( .A1(n5453), .A2(n10023), .ZN(n5201) );
  NAND2_X2 U6637 ( .A1(n4513), .A2(n5201), .ZN(n6391) );
  INV_X1 U6638 ( .A(n6391), .ZN(n10413) );
  NAND2_X1 U6639 ( .A1(n10413), .A2(n8577), .ZN(n5650) );
  NAND2_X1 U6640 ( .A1(n5649), .A2(n5650), .ZN(n7215) );
  INV_X1 U6641 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5202) );
  INV_X1 U6642 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10359) );
  INV_X1 U6643 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5203) );
  OR2_X1 U6644 ( .A1(n5214), .A2(n5203), .ZN(n5205) );
  NAND2_X1 U6645 ( .A1(n4486), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5204) );
  AND2_X1 U6646 ( .A1(n5205), .A2(n5204), .ZN(n5206) );
  NAND2_X1 U6647 ( .A1(n6660), .A2(SI_0_), .ZN(n5209) );
  XNOR2_X1 U6648 ( .A(n5209), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9033) );
  MUX2_X1 U6649 ( .A(n10355), .B(n9033), .S(n5210), .Z(n10408) );
  AND2_X1 U6650 ( .A1(n8579), .A2(n10408), .ZN(n7219) );
  NAND2_X1 U6651 ( .A1(n7215), .A2(n7219), .ZN(n7221) );
  NAND2_X1 U6652 ( .A1(n8577), .A2(n6391), .ZN(n5211) );
  INV_X1 U6653 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5212) );
  INV_X1 U6654 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5213) );
  INV_X1 U6655 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6799) );
  OR2_X1 U6656 ( .A1(n5214), .A2(n6799), .ZN(n5216) );
  NAND2_X1 U6657 ( .A1(n4487), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5215) );
  AND2_X1 U6658 ( .A1(n5216), .A2(n5215), .ZN(n5217) );
  XNOR2_X1 U6659 ( .A(n5221), .B(n5220), .ZN(n6664) );
  NAND2_X1 U6660 ( .A1(n4481), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5226) );
  OR2_X1 U6661 ( .A1(n5223), .A2(n9022), .ZN(n5224) );
  XNOR2_X1 U6662 ( .A(n5224), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10041) );
  NAND2_X1 U6663 ( .A1(n5453), .A2(n10041), .ZN(n5225) );
  OAI211_X2 U6664 ( .C1(n8357), .C2(n6664), .A(n5226), .B(n5225), .ZN(n7231)
         );
  NAND2_X1 U6665 ( .A1(n8576), .A2(n7233), .ZN(n8423) );
  NAND2_X1 U6666 ( .A1(n6399), .A2(n7233), .ZN(n5227) );
  NAND2_X1 U6667 ( .A1(n4487), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5233) );
  INV_X1 U6668 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6798) );
  OR2_X1 U6669 ( .A1(n5214), .A2(n6798), .ZN(n5232) );
  OR2_X1 U6670 ( .A1(n5615), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5231) );
  INV_X1 U6671 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5228) );
  OR2_X1 U6672 ( .A1(n5229), .A2(n5228), .ZN(n5230) );
  NAND2_X1 U6673 ( .A1(n5222), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6674 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4518), .ZN(n5236) );
  XNOR2_X1 U6675 ( .A(n5236), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6853) );
  NAND2_X1 U6676 ( .A1(n5453), .A2(n6853), .ZN(n5237) );
  NAND2_X1 U6677 ( .A1(n7198), .A2(n7351), .ZN(n8402) );
  INV_X1 U6678 ( .A(n7198), .ZN(n8575) );
  NAND2_X1 U6679 ( .A1(n8575), .A2(n10419), .ZN(n8397) );
  NAND2_X1 U6680 ( .A1(n8402), .A2(n8397), .ZN(n8367) );
  NAND2_X1 U6681 ( .A1(n7343), .A2(n8367), .ZN(n7342) );
  NAND2_X1 U6682 ( .A1(n7198), .A2(n10419), .ZN(n5239) );
  NAND2_X1 U6683 ( .A1(n7342), .A2(n5239), .ZN(n7244) );
  INV_X1 U6684 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6815) );
  OAI21_X1 U6685 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5249), .ZN(n7240) );
  OR2_X1 U6686 ( .A1(n5615), .A2(n7240), .ZN(n5242) );
  INV_X1 U6687 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5240) );
  OR2_X1 U6688 ( .A1(n5229), .A2(n5240), .ZN(n5241) );
  XNOR2_X1 U6689 ( .A(n5244), .B(n5243), .ZN(n6680) );
  NAND2_X1 U6690 ( .A1(n5222), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5247) );
  OR2_X1 U6691 ( .A1(n5259), .A2(n9022), .ZN(n5245) );
  XNOR2_X1 U6692 ( .A(n5245), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6840) );
  NAND2_X1 U6693 ( .A1(n5453), .A2(n6840), .ZN(n5246) );
  NAND2_X1 U6694 ( .A1(n7407), .A2(n7362), .ZN(n8403) );
  INV_X1 U6695 ( .A(n7362), .ZN(n7239) );
  NAND2_X1 U6696 ( .A1(n8574), .A2(n7239), .ZN(n7403) );
  NAND2_X1 U6697 ( .A1(n8403), .A2(n7403), .ZN(n8364) );
  NAND2_X1 U6698 ( .A1(n7244), .A2(n8364), .ZN(n7243) );
  NAND2_X1 U6699 ( .A1(n7407), .A2(n7239), .ZN(n5248) );
  NAND2_X1 U6700 ( .A1(n4487), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5255) );
  INV_X1 U6701 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6806) );
  OR2_X1 U6702 ( .A1(n5637), .A2(n6806), .ZN(n5254) );
  INV_X1 U6703 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9924) );
  NAND2_X1 U6704 ( .A1(n5249), .A2(n9924), .ZN(n5250) );
  NAND2_X1 U6705 ( .A1(n5277), .A2(n5250), .ZN(n7210) );
  OR2_X1 U6706 ( .A1(n5615), .A2(n7210), .ZN(n5253) );
  INV_X1 U6707 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5251) );
  OR2_X1 U6708 ( .A1(n5229), .A2(n5251), .ZN(n5252) );
  XNOR2_X1 U6709 ( .A(n5257), .B(n5256), .ZN(n6673) );
  NAND2_X1 U6710 ( .A1(n5222), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5261) );
  INV_X1 U6711 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5258) );
  NAND2_X1 U6712 ( .A1(n5259), .A2(n5258), .ZN(n5304) );
  NAND2_X1 U6713 ( .A1(n5304), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5269) );
  XNOR2_X1 U6714 ( .A(n5269), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6880) );
  NAND2_X1 U6715 ( .A1(n5453), .A2(n6880), .ZN(n5260) );
  OAI211_X1 U6716 ( .C1(n8357), .C2(n6673), .A(n5261), .B(n5260), .ZN(n7576)
         );
  NAND2_X1 U6717 ( .A1(n7489), .A2(n7576), .ZN(n8404) );
  INV_X1 U6718 ( .A(n7489), .ZN(n8573) );
  NAND2_X1 U6719 ( .A1(n8573), .A2(n7573), .ZN(n8395) );
  NAND2_X1 U6720 ( .A1(n8404), .A2(n8395), .ZN(n8365) );
  NAND2_X1 U6721 ( .A1(n7409), .A2(n8365), .ZN(n7408) );
  NAND2_X1 U6722 ( .A1(n7489), .A2(n7573), .ZN(n5262) );
  NAND2_X1 U6723 ( .A1(n7408), .A2(n5262), .ZN(n7378) );
  NAND2_X1 U6724 ( .A1(n4486), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5267) );
  INV_X1 U6725 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6809) );
  OR2_X1 U6726 ( .A1(n5637), .A2(n6809), .ZN(n5266) );
  INV_X1 U6727 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5276) );
  XNOR2_X1 U6728 ( .A(n5277), .B(n5276), .ZN(n7488) );
  OR2_X1 U6729 ( .A1(n5615), .A2(n7488), .ZN(n5265) );
  INV_X1 U6730 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5263) );
  OR2_X1 U6731 ( .A1(n5229), .A2(n5263), .ZN(n5264) );
  NAND2_X1 U6732 ( .A1(n5222), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5272) );
  INV_X1 U6733 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5301) );
  NAND2_X1 U6734 ( .A1(n5269), .A2(n5301), .ZN(n5270) );
  NAND2_X1 U6735 ( .A1(n5270), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5285) );
  XNOR2_X1 U6736 ( .A(n5285), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6864) );
  NAND2_X1 U6737 ( .A1(n5453), .A2(n6864), .ZN(n5271) );
  NAND2_X1 U6738 ( .A1(n7423), .A2(n7603), .ZN(n8432) );
  INV_X1 U6739 ( .A(n7423), .ZN(n8572) );
  NAND2_X1 U6740 ( .A1(n8572), .A2(n7606), .ZN(n8426) );
  NAND2_X1 U6741 ( .A1(n8432), .A2(n8426), .ZN(n8368) );
  NAND2_X1 U6742 ( .A1(n7378), .A2(n8368), .ZN(n7377) );
  NAND2_X1 U6743 ( .A1(n7423), .A2(n7606), .ZN(n5273) );
  NAND2_X1 U6744 ( .A1(n4486), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5282) );
  INV_X1 U6745 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5274) );
  OR2_X1 U6746 ( .A1(n5229), .A2(n5274), .ZN(n5281) );
  INV_X1 U6747 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5275) );
  OAI21_X1 U6748 ( .B1(n5277), .B2(n5276), .A(n5275), .ZN(n5278) );
  NAND2_X1 U6749 ( .A1(n5278), .A2(n5291), .ZN(n7541) );
  OR2_X1 U6750 ( .A1(n5615), .A2(n7541), .ZN(n5280) );
  INV_X1 U6751 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6857) );
  OR2_X1 U6752 ( .A1(n5214), .A2(n6857), .ZN(n5279) );
  NAND2_X1 U6753 ( .A1(n5222), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5289) );
  INV_X1 U6754 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5302) );
  NAND2_X1 U6755 ( .A1(n5285), .A2(n5302), .ZN(n5286) );
  NAND2_X1 U6756 ( .A1(n5286), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5287) );
  XNOR2_X1 U6757 ( .A(n5287), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6983) );
  NAND2_X1 U6758 ( .A1(n5453), .A2(n6983), .ZN(n5288) );
  NAND2_X1 U6759 ( .A1(n7625), .A2(n4482), .ZN(n8433) );
  INV_X1 U6760 ( .A(n7625), .ZN(n8571) );
  INV_X1 U6761 ( .A(n4482), .ZN(n10426) );
  NAND2_X1 U6762 ( .A1(n8571), .A2(n10426), .ZN(n8434) );
  NAND2_X1 U6763 ( .A1(n8433), .A2(n8434), .ZN(n7549) );
  NAND2_X1 U6764 ( .A1(n7625), .A2(n10426), .ZN(n5290) );
  NAND2_X1 U6765 ( .A1(n4486), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5297) );
  INV_X1 U6766 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7032) );
  OR2_X1 U6767 ( .A1(n5637), .A2(n7032), .ZN(n5296) );
  INV_X1 U6768 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7502) );
  NAND2_X1 U6769 ( .A1(n5291), .A2(n7502), .ZN(n5292) );
  NAND2_X1 U6770 ( .A1(n5310), .A2(n5292), .ZN(n7500) );
  OR2_X1 U6771 ( .A1(n5615), .A2(n7500), .ZN(n5295) );
  INV_X1 U6772 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5293) );
  OR2_X1 U6773 ( .A1(n5229), .A2(n5293), .ZN(n5294) );
  XNOR2_X1 U6774 ( .A(n5299), .B(n5298), .ZN(n6686) );
  NAND2_X1 U6775 ( .A1(n8352), .A2(n6686), .ZN(n5307) );
  INV_X1 U6776 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5300) );
  NAND3_X1 U6777 ( .A1(n5302), .A2(n5301), .A3(n5300), .ZN(n5303) );
  NAND2_X1 U6778 ( .A1(n5317), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5305) );
  XNOR2_X1 U6779 ( .A(n5305), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7040) );
  NAND2_X1 U6780 ( .A1(n5453), .A2(n7040), .ZN(n5306) );
  NAND2_X1 U6781 ( .A1(n7613), .A2(n7631), .ZN(n8438) );
  INV_X1 U6782 ( .A(n7631), .ZN(n7715) );
  NAND2_X1 U6783 ( .A1(n8570), .A2(n7715), .ZN(n8439) );
  NAND2_X1 U6784 ( .A1(n8570), .A2(n7631), .ZN(n5308) );
  NAND2_X1 U6785 ( .A1(n4486), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5316) );
  INV_X1 U6786 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7029) );
  OR2_X1 U6787 ( .A1(n5637), .A2(n7029), .ZN(n5315) );
  NAND2_X1 U6788 ( .A1(n5310), .A2(n5309), .ZN(n5311) );
  NAND2_X1 U6789 ( .A1(n5329), .A2(n5311), .ZN(n7672) );
  OR2_X1 U6790 ( .A1(n5615), .A2(n7672), .ZN(n5314) );
  INV_X1 U6791 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5312) );
  OR2_X1 U6792 ( .A1(n5229), .A2(n5312), .ZN(n5313) );
  NOR2_X1 U6793 ( .A1(n5317), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5358) );
  OR2_X1 U6794 ( .A1(n5358), .A2(n9022), .ZN(n5325) );
  XNOR2_X1 U6795 ( .A(n5325), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8585) );
  AOI22_X1 U6796 ( .A1(n5222), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5453), .B2(
        n8585), .ZN(n5321) );
  XNOR2_X1 U6797 ( .A(n5319), .B(n5318), .ZN(n6693) );
  NAND2_X1 U6798 ( .A1(n6693), .A2(n8352), .ZN(n5320) );
  NAND2_X1 U6799 ( .A1(n5321), .A2(n5320), .ZN(n7675) );
  NAND2_X1 U6800 ( .A1(n7742), .A2(n7675), .ZN(n8440) );
  INV_X1 U6801 ( .A(n7742), .ZN(n8569) );
  NAND2_X1 U6802 ( .A1(n8569), .A2(n10429), .ZN(n8450) );
  NAND2_X1 U6803 ( .A1(n7670), .A2(n7669), .ZN(n7668) );
  NAND2_X1 U6804 ( .A1(n7742), .A2(n10429), .ZN(n5322) );
  XNOR2_X1 U6805 ( .A(n5324), .B(n5323), .ZN(n6704) );
  NAND2_X1 U6806 ( .A1(n6704), .A2(n8352), .ZN(n5328) );
  NAND2_X1 U6807 ( .A1(n5325), .A2(n5355), .ZN(n5326) );
  NAND2_X1 U6808 ( .A1(n5326), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5337) );
  XNOR2_X1 U6809 ( .A(n5337), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7098) );
  AOI22_X1 U6810 ( .A1(n4481), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5453), .B2(
        n7098), .ZN(n5327) );
  NAND2_X1 U6811 ( .A1(n4487), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6812 ( .A1(n5634), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5333) );
  INV_X1 U6813 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9977) );
  NAND2_X1 U6814 ( .A1(n5329), .A2(n9977), .ZN(n5330) );
  NAND2_X1 U6815 ( .A1(n5343), .A2(n5330), .ZN(n7749) );
  OR2_X1 U6816 ( .A1(n5615), .A2(n7749), .ZN(n5332) );
  INV_X1 U6817 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7028) );
  OR2_X1 U6818 ( .A1(n5637), .A2(n7028), .ZN(n5331) );
  NAND4_X1 U6819 ( .A1(n5334), .A2(n5333), .A3(n5332), .A4(n5331), .ZN(n8568)
         );
  NAND2_X1 U6820 ( .A1(n7748), .A2(n8568), .ZN(n8449) );
  INV_X1 U6821 ( .A(n8568), .ZN(n7761) );
  NAND2_X1 U6822 ( .A1(n7761), .A2(n8981), .ZN(n8448) );
  XNOR2_X1 U6823 ( .A(n5336), .B(n5335), .ZN(n6707) );
  NAND2_X1 U6824 ( .A1(n6707), .A2(n8352), .ZN(n5341) );
  INV_X1 U6825 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6826 ( .A1(n5337), .A2(n5356), .ZN(n5338) );
  NAND2_X1 U6827 ( .A1(n5338), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5339) );
  XNOR2_X1 U6828 ( .A(n5339), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7165) );
  AOI22_X1 U6829 ( .A1(n5222), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5453), .B2(
        n7165), .ZN(n5340) );
  NAND2_X1 U6830 ( .A1(n5634), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5348) );
  INV_X1 U6831 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7764) );
  OR2_X1 U6832 ( .A1(n5476), .A2(n7764), .ZN(n5347) );
  INV_X1 U6833 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7097) );
  OR2_X1 U6834 ( .A1(n5214), .A2(n7097), .ZN(n5346) );
  NAND2_X1 U6835 ( .A1(n5343), .A2(n5342), .ZN(n5344) );
  NAND2_X1 U6836 ( .A1(n5363), .A2(n5344), .ZN(n7763) );
  OR2_X1 U6837 ( .A1(n5615), .A2(n7763), .ZN(n5345) );
  NAND2_X1 U6838 ( .A1(n7766), .A2(n7793), .ZN(n8456) );
  NAND2_X1 U6839 ( .A1(n8460), .A2(n8456), .ZN(n7758) );
  INV_X1 U6840 ( .A(n7758), .ZN(n5349) );
  OR2_X1 U6841 ( .A1(n8444), .A2(n5349), .ZN(n5351) );
  NAND2_X1 U6842 ( .A1(n8981), .A2(n8568), .ZN(n7755) );
  INV_X1 U6843 ( .A(n7793), .ZN(n8567) );
  XNOR2_X1 U6844 ( .A(n5353), .B(n5352), .ZN(n6720) );
  NAND2_X1 U6845 ( .A1(n6720), .A2(n8352), .ZN(n5361) );
  INV_X1 U6846 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5354) );
  AND3_X1 U6847 ( .A1(n5356), .A2(n5355), .A3(n5354), .ZN(n5357) );
  AND2_X1 U6848 ( .A1(n5358), .A2(n5357), .ZN(n5374) );
  OR2_X1 U6849 ( .A1(n5374), .A2(n9022), .ZN(n5359) );
  XNOR2_X1 U6850 ( .A(n5359), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7293) );
  AOI22_X1 U6851 ( .A1(n4481), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5453), .B2(
        n7293), .ZN(n5360) );
  NAND2_X1 U6852 ( .A1(n4486), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5369) );
  INV_X1 U6853 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5362) );
  OR2_X1 U6854 ( .A1(n5637), .A2(n5362), .ZN(n5368) );
  INV_X1 U6855 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9789) );
  NAND2_X1 U6856 ( .A1(n5363), .A2(n9789), .ZN(n5364) );
  NAND2_X1 U6857 ( .A1(n5378), .A2(n5364), .ZN(n7799) );
  OR2_X1 U6858 ( .A1(n5615), .A2(n7799), .ZN(n5367) );
  INV_X1 U6859 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5365) );
  OR2_X1 U6860 ( .A1(n5229), .A2(n5365), .ZN(n5366) );
  NAND2_X1 U6861 ( .A1(n7805), .A2(n7878), .ZN(n8463) );
  INV_X1 U6862 ( .A(n7878), .ZN(n8566) );
  XNOR2_X1 U6863 ( .A(n5372), .B(n5371), .ZN(n6785) );
  NAND2_X1 U6864 ( .A1(n6785), .A2(n8352), .ZN(n5376) );
  NAND2_X1 U6865 ( .A1(n5374), .A2(n5373), .ZN(n5422) );
  NAND2_X1 U6866 ( .A1(n5422), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5387) );
  XNOR2_X1 U6867 ( .A(n5387), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7395) );
  AOI22_X1 U6868 ( .A1(n5222), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5453), .B2(
        n7395), .ZN(n5375) );
  NAND2_X1 U6869 ( .A1(n5634), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5383) );
  INV_X1 U6870 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5377) );
  OR2_X1 U6871 ( .A1(n5637), .A2(n5377), .ZN(n5382) );
  INV_X1 U6872 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7884) );
  OR2_X1 U6873 ( .A1(n5476), .A2(n7884), .ZN(n5381) );
  NAND2_X1 U6874 ( .A1(n5378), .A2(n7282), .ZN(n5379) );
  NAND2_X1 U6875 ( .A1(n5395), .A2(n5379), .ZN(n7883) );
  OR2_X1 U6876 ( .A1(n5615), .A2(n7883), .ZN(n5380) );
  OR2_X1 U6877 ( .A1(n10079), .A2(n8893), .ZN(n8466) );
  NAND2_X1 U6878 ( .A1(n10079), .A2(n8893), .ZN(n8458) );
  INV_X1 U6879 ( .A(n8893), .ZN(n8565) );
  XNOR2_X1 U6880 ( .A(n5386), .B(n5385), .ZN(n6788) );
  NAND2_X1 U6881 ( .A1(n6788), .A2(n8352), .ZN(n5393) );
  INV_X1 U6882 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6883 ( .A1(n5387), .A2(n5420), .ZN(n5388) );
  NAND2_X1 U6884 ( .A1(n5388), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6885 ( .A1(n5390), .A2(n5389), .ZN(n5404) );
  OR2_X1 U6886 ( .A1(n5390), .A2(n5389), .ZN(n5391) );
  AND2_X1 U6887 ( .A1(n5404), .A2(n5391), .ZN(n7649) );
  AOI22_X1 U6888 ( .A1(n4481), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5453), .B2(
        n7649), .ZN(n5392) );
  NAND2_X1 U6889 ( .A1(n5634), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5400) );
  INV_X1 U6890 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5394) );
  OR2_X1 U6891 ( .A1(n5476), .A2(n5394), .ZN(n5399) );
  INV_X1 U6892 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8977) );
  OR2_X1 U6893 ( .A1(n5637), .A2(n8977), .ZN(n5398) );
  NAND2_X1 U6894 ( .A1(n5395), .A2(n9755), .ZN(n5396) );
  NAND2_X1 U6895 ( .A1(n5409), .A2(n5396), .ZN(n8883) );
  OR2_X1 U6896 ( .A1(n5615), .A2(n8883), .ZN(n5397) );
  NAND2_X1 U6897 ( .A1(n8886), .A2(n8860), .ZN(n8471) );
  INV_X1 U6898 ( .A(n8860), .ZN(n8564) );
  OR2_X1 U6899 ( .A1(n8886), .A2(n8564), .ZN(n5401) );
  NAND2_X1 U6900 ( .A1(n5047), .A2(n5401), .ZN(n8866) );
  XNOR2_X1 U6901 ( .A(n5403), .B(n5402), .ZN(n7024) );
  NAND2_X1 U6902 ( .A1(n7024), .A2(n8352), .ZN(n5407) );
  NAND2_X1 U6903 ( .A1(n5404), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5405) );
  XNOR2_X1 U6904 ( .A(n5405), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7772) );
  AOI22_X1 U6905 ( .A1(n4481), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5453), .B2(
        n7772), .ZN(n5406) );
  NAND2_X1 U6906 ( .A1(n5634), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5414) );
  INV_X1 U6907 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5408) );
  OR2_X1 U6908 ( .A1(n5637), .A2(n5408), .ZN(n5413) );
  INV_X1 U6909 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8871) );
  OR2_X1 U6910 ( .A1(n5476), .A2(n8871), .ZN(n5412) );
  INV_X1 U6911 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8340) );
  NAND2_X1 U6912 ( .A1(n5409), .A2(n8340), .ZN(n5410) );
  NAND2_X1 U6913 ( .A1(n5429), .A2(n5410), .ZN(n8870) );
  OR2_X1 U6914 ( .A1(n5615), .A2(n8870), .ZN(n5411) );
  NAND2_X1 U6915 ( .A1(n8967), .A2(n8891), .ZN(n8474) );
  NAND2_X1 U6916 ( .A1(n8475), .A2(n8474), .ZN(n8865) );
  NAND2_X1 U6917 ( .A1(n8866), .A2(n8865), .ZN(n8864) );
  INV_X1 U6918 ( .A(n8891), .ZN(n8563) );
  OR2_X1 U6919 ( .A1(n8967), .A2(n8563), .ZN(n5415) );
  XNOR2_X1 U6920 ( .A(n5417), .B(n5416), .ZN(n7090) );
  NAND2_X1 U6921 ( .A1(n7090), .A2(n8352), .ZN(n5426) );
  INV_X1 U6922 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5419) );
  NAND3_X1 U6923 ( .A1(n5420), .A2(n5389), .A3(n5419), .ZN(n5421) );
  OAI21_X1 U6924 ( .B1(n5422), .B2(n5421), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5423) );
  MUX2_X1 U6925 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5423), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5424) );
  AND2_X1 U6926 ( .A1(n5418), .A2(n5424), .ZN(n7811) );
  AOI22_X1 U6927 ( .A1(n5222), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5453), .B2(
        n7811), .ZN(n5425) );
  NAND2_X1 U6928 ( .A1(n4487), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5435) );
  INV_X1 U6929 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n5427) );
  OR2_X1 U6930 ( .A1(n5214), .A2(n5427), .ZN(n5434) );
  INV_X1 U6931 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U6932 ( .A1(n5429), .A2(n5428), .ZN(n5430) );
  NAND2_X1 U6933 ( .A1(n5442), .A2(n5430), .ZN(n8296) );
  OR2_X1 U6934 ( .A1(n5615), .A2(n8296), .ZN(n5433) );
  INV_X1 U6935 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n5431) );
  OR2_X1 U6936 ( .A1(n5229), .A2(n5431), .ZN(n5432) );
  OR2_X1 U6937 ( .A1(n8850), .A2(n8859), .ZN(n8477) );
  NAND2_X1 U6938 ( .A1(n8850), .A2(n8859), .ZN(n8810) );
  INV_X1 U6939 ( .A(n8859), .ZN(n8817) );
  XNOR2_X1 U6940 ( .A(n5437), .B(n5436), .ZN(n7154) );
  NAND2_X1 U6941 ( .A1(n7154), .A2(n8352), .ZN(n5440) );
  NAND2_X1 U6942 ( .A1(n5418), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5438) );
  XNOR2_X1 U6943 ( .A(n5438), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8594) );
  AOI22_X1 U6944 ( .A1(n4481), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5453), .B2(
        n8594), .ZN(n5439) );
  NAND2_X1 U6945 ( .A1(n5674), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5447) );
  INV_X1 U6946 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8827) );
  OR2_X1 U6947 ( .A1(n5476), .A2(n8827), .ZN(n5446) );
  NAND2_X1 U6948 ( .A1(n5442), .A2(n5441), .ZN(n5443) );
  NAND2_X1 U6949 ( .A1(n5456), .A2(n5443), .ZN(n8826) );
  OR2_X1 U6950 ( .A1(n5615), .A2(n8826), .ZN(n5445) );
  INV_X1 U6951 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9011) );
  OR2_X1 U6952 ( .A1(n5229), .A2(n9011), .ZN(n5444) );
  NAND2_X1 U6953 ( .A1(n8825), .A2(n8842), .ZN(n8481) );
  NAND2_X1 U6954 ( .A1(n8800), .A2(n8481), .ZN(n8821) );
  INV_X1 U6955 ( .A(n8842), .ZN(n8803) );
  XNOR2_X1 U6956 ( .A(n5450), .B(n5449), .ZN(n7247) );
  NAND2_X1 U6957 ( .A1(n7247), .A2(n8352), .ZN(n5455) );
  NAND2_X1 U6958 ( .A1(n5451), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5452) );
  XNOR2_X1 U6959 ( .A(n5452), .B(n5030), .ZN(n8616) );
  INV_X1 U6960 ( .A(n8616), .ZN(n8601) );
  AOI22_X1 U6961 ( .A1(n5222), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5453), .B2(
        n8601), .ZN(n5454) );
  NAND2_X1 U6962 ( .A1(n5634), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5463) );
  INV_X1 U6963 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8615) );
  OR2_X1 U6964 ( .A1(n5637), .A2(n8615), .ZN(n5462) );
  INV_X1 U6965 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9781) );
  NAND2_X1 U6966 ( .A1(n5456), .A2(n9781), .ZN(n5457) );
  NAND2_X1 U6967 ( .A1(n5458), .A2(n5457), .ZN(n8796) );
  OR2_X1 U6968 ( .A1(n5615), .A2(n8796), .ZN(n5461) );
  INV_X1 U6969 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5459) );
  OR2_X1 U6970 ( .A1(n5476), .A2(n5459), .ZN(n5460) );
  NAND4_X1 U6971 ( .A1(n5463), .A2(n5462), .A3(n5461), .A4(n5460), .ZN(n8814)
         );
  NAND2_X1 U6972 ( .A1(n8950), .A2(n8814), .ZN(n5465) );
  INV_X1 U6973 ( .A(n8950), .ZN(n8799) );
  INV_X1 U6974 ( .A(n8814), .ZN(n8304) );
  OAI21_X1 U6975 ( .B1(n8946), .B2(n8804), .A(n8778), .ZN(n5466) );
  INV_X1 U6976 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7495) );
  INV_X1 U6977 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7496) );
  MUX2_X1 U6978 ( .A(n7495), .B(n7496), .S(n7982), .Z(n5470) );
  INV_X1 U6979 ( .A(SI_20_), .ZN(n9718) );
  NAND2_X1 U6980 ( .A1(n5470), .A2(n9718), .ZN(n5487) );
  INV_X1 U6981 ( .A(n5470), .ZN(n5471) );
  NAND2_X1 U6982 ( .A1(n5471), .A2(SI_20_), .ZN(n5472) );
  XNOR2_X1 U6983 ( .A(n5486), .B(n5485), .ZN(n7494) );
  NAND2_X1 U6984 ( .A1(n7494), .A2(n8352), .ZN(n5474) );
  NAND2_X1 U6985 ( .A1(n4481), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U6986 ( .A1(n5674), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5484) );
  INV_X1 U6987 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5475) );
  OR2_X1 U6988 ( .A1(n5476), .A2(n5475), .ZN(n5483) );
  INV_X1 U6989 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9744) );
  NAND2_X1 U6990 ( .A1(n5478), .A2(n9744), .ZN(n5479) );
  NAND2_X1 U6991 ( .A1(n5493), .A2(n5479), .ZN(n8761) );
  OR2_X1 U6992 ( .A1(n5615), .A2(n8761), .ZN(n5482) );
  INV_X1 U6993 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n5480) );
  OR2_X1 U6994 ( .A1(n5229), .A2(n5480), .ZN(n5481) );
  NAND2_X1 U6995 ( .A1(n8940), .A2(n8275), .ZN(n8496) );
  NAND2_X1 U6996 ( .A1(n8493), .A2(n8496), .ZN(n8771) );
  INV_X1 U6997 ( .A(n8275), .ZN(n8788) );
  INV_X1 U6998 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7526) );
  INV_X1 U6999 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n5488) );
  MUX2_X1 U7000 ( .A(n7526), .B(n5488), .S(n7982), .Z(n5499) );
  XNOR2_X1 U7001 ( .A(n5499), .B(SI_21_), .ZN(n5498) );
  XNOR2_X1 U7002 ( .A(n5503), .B(n5498), .ZN(n7525) );
  NAND2_X1 U7003 ( .A1(n7525), .A2(n8352), .ZN(n5490) );
  NAND2_X1 U7004 ( .A1(n5222), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5489) );
  INV_X1 U7005 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U7006 ( .A1(n4486), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5491) );
  OAI21_X1 U7007 ( .B1(n5229), .B2(n5492), .A(n5491), .ZN(n5497) );
  INV_X1 U7008 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9955) );
  NAND2_X1 U7009 ( .A1(n5493), .A2(n9955), .ZN(n5494) );
  NAND2_X1 U7010 ( .A1(n5511), .A2(n5494), .ZN(n8747) );
  NAND2_X1 U7011 ( .A1(n5674), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5495) );
  OAI21_X1 U7012 ( .B1(n8747), .B2(n5615), .A(n5495), .ZN(n5496) );
  INV_X1 U7013 ( .A(n5498), .ZN(n5502) );
  INV_X1 U7014 ( .A(n5499), .ZN(n5500) );
  NAND2_X1 U7015 ( .A1(n5500), .A2(SI_21_), .ZN(n5501) );
  INV_X1 U7016 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7663) );
  INV_X1 U7017 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9929) );
  MUX2_X1 U7018 ( .A(n7663), .B(n9929), .S(n7982), .Z(n5504) );
  INV_X1 U7019 ( .A(SI_22_), .ZN(n9991) );
  NAND2_X1 U7020 ( .A1(n5504), .A2(n9991), .ZN(n5516) );
  INV_X1 U7021 ( .A(n5504), .ZN(n5505) );
  NAND2_X1 U7022 ( .A1(n5505), .A2(SI_22_), .ZN(n5506) );
  NAND2_X1 U7023 ( .A1(n5516), .A2(n5506), .ZN(n5517) );
  XNOR2_X1 U7024 ( .A(n5518), .B(n5517), .ZN(n7660) );
  NAND2_X1 U7025 ( .A1(n7660), .A2(n8352), .ZN(n5508) );
  NAND2_X1 U7026 ( .A1(n4480), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5507) );
  INV_X1 U7027 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U7028 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  NAND2_X1 U7029 ( .A1(n5532), .A2(n5512), .ZN(n8731) );
  OR2_X1 U7030 ( .A1(n8731), .A2(n5615), .ZN(n5515) );
  AOI22_X1 U7031 ( .A1(n5634), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n4486), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U7032 ( .A1(n5674), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U7033 ( .A1(n8930), .A2(n8274), .ZN(n8499) );
  INV_X1 U7034 ( .A(n8274), .ZN(n8753) );
  INV_X1 U7035 ( .A(n5527), .ZN(n5524) );
  INV_X1 U7036 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5520) );
  INV_X1 U7037 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5519) );
  MUX2_X1 U7038 ( .A(n5520), .B(n5519), .S(n7982), .Z(n5521) );
  INV_X1 U7039 ( .A(SI_23_), .ZN(n9817) );
  NAND2_X1 U7040 ( .A1(n5521), .A2(n9817), .ZN(n5537) );
  INV_X1 U7041 ( .A(n5521), .ZN(n5522) );
  NAND2_X1 U7042 ( .A1(n5522), .A2(SI_23_), .ZN(n5523) );
  NAND2_X1 U7043 ( .A1(n5537), .A2(n5523), .ZN(n5525) );
  NAND2_X1 U7044 ( .A1(n5524), .A2(n5525), .ZN(n5528) );
  INV_X1 U7045 ( .A(n5525), .ZN(n5526) );
  NAND2_X1 U7046 ( .A1(n5528), .A2(n5538), .ZN(n7680) );
  NAND2_X1 U7047 ( .A1(n7680), .A2(n8352), .ZN(n5530) );
  NAND2_X1 U7048 ( .A1(n4481), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5529) );
  INV_X1 U7049 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U7050 ( .A1(n5532), .A2(n5531), .ZN(n5533) );
  AND2_X1 U7051 ( .A1(n5542), .A2(n5533), .ZN(n8723) );
  NAND2_X1 U7052 ( .A1(n8723), .A2(n5195), .ZN(n5536) );
  AOI22_X1 U7053 ( .A1(n4487), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n5674), .B2(
        P2_REG1_REG_23__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U7054 ( .A1(n5634), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U7055 ( .A1(n8722), .A2(n8738), .ZN(n8505) );
  INV_X1 U7056 ( .A(n8738), .ZN(n6933) );
  INV_X1 U7057 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7790) );
  INV_X1 U7058 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7821) );
  MUX2_X1 U7059 ( .A(n7790), .B(n7821), .S(n7982), .Z(n5550) );
  XNOR2_X1 U7060 ( .A(n5550), .B(SI_24_), .ZN(n5549) );
  NAND2_X1 U7061 ( .A1(n5222), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5539) );
  INV_X1 U7062 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U7063 ( .A1(n5542), .A2(n9752), .ZN(n5543) );
  NAND2_X1 U7064 ( .A1(n5559), .A2(n5543), .ZN(n8697) );
  OR2_X1 U7065 ( .A1(n8697), .A2(n5615), .ZN(n5546) );
  AOI22_X1 U7066 ( .A1(n4486), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n5674), .B2(
        P2_REG1_REG_24__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7067 ( .A1(n5634), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7068 ( .A1(n8920), .A2(n8257), .ZN(n8506) );
  NAND2_X1 U7069 ( .A1(n8694), .A2(n8701), .ZN(n8693) );
  INV_X1 U7070 ( .A(n5550), .ZN(n5551) );
  INV_X1 U7071 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7829) );
  INV_X1 U7072 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9921) );
  MUX2_X1 U7073 ( .A(n7829), .B(n9921), .S(n7982), .Z(n5553) );
  INV_X1 U7074 ( .A(SI_25_), .ZN(n9765) );
  NAND2_X1 U7075 ( .A1(n5553), .A2(n9765), .ZN(n5566) );
  INV_X1 U7076 ( .A(n5553), .ZN(n5554) );
  NAND2_X1 U7077 ( .A1(n5554), .A2(SI_25_), .ZN(n5555) );
  NAND2_X1 U7078 ( .A1(n5566), .A2(n5555), .ZN(n5567) );
  XNOR2_X1 U7079 ( .A(n5568), .B(n5567), .ZN(n7824) );
  NAND2_X1 U7080 ( .A1(n7824), .A2(n8352), .ZN(n5557) );
  NAND2_X1 U7081 ( .A1(n4480), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5556) );
  INV_X1 U7082 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U7083 ( .A1(n5559), .A2(n5558), .ZN(n5560) );
  NAND2_X1 U7084 ( .A1(n5589), .A2(n5560), .ZN(n8686) );
  OR2_X1 U7085 ( .A1(n8686), .A2(n5615), .ZN(n5565) );
  INV_X1 U7086 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8997) );
  NAND2_X1 U7087 ( .A1(n5674), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U7088 ( .A1(n4486), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5561) );
  OAI211_X1 U7089 ( .C1(n8997), .C2(n5229), .A(n5562), .B(n5561), .ZN(n5563)
         );
  INV_X1 U7090 ( .A(n5563), .ZN(n5564) );
  INV_X1 U7091 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7913) );
  INV_X1 U7092 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9978) );
  MUX2_X1 U7093 ( .A(n7913), .B(n9978), .S(n7982), .Z(n5569) );
  INV_X1 U7094 ( .A(SI_26_), .ZN(n9731) );
  NAND2_X1 U7095 ( .A1(n5569), .A2(n9731), .ZN(n5572) );
  INV_X1 U7096 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U7097 ( .A1(n5570), .A2(SI_26_), .ZN(n5571) );
  INV_X1 U7098 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7929) );
  INV_X1 U7099 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9777) );
  MUX2_X1 U7100 ( .A(n7929), .B(n9777), .S(n7982), .Z(n5575) );
  INV_X1 U7101 ( .A(SI_27_), .ZN(n5574) );
  NAND2_X1 U7102 ( .A1(n5575), .A2(n5574), .ZN(n5607) );
  INV_X1 U7103 ( .A(n5575), .ZN(n5576) );
  NAND2_X1 U7104 ( .A1(n5576), .A2(SI_27_), .ZN(n5577) );
  AND2_X1 U7105 ( .A1(n5607), .A2(n5577), .ZN(n5578) );
  NAND2_X1 U7106 ( .A1(n4481), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5580) );
  INV_X1 U7107 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9779) );
  XNOR2_X1 U7108 ( .A(n5613), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n7960) );
  INV_X1 U7109 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U7110 ( .A1(n5674), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U7111 ( .A1(n4487), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5582) );
  OAI211_X1 U7112 ( .C1(n6567), .C2(n5229), .A(n5583), .B(n5582), .ZN(n5584)
         );
  AOI21_X2 U7113 ( .B1(n7960), .B2(n5195), .A(n5584), .ZN(n8650) );
  INV_X1 U7114 ( .A(n8379), .ZN(n5595) );
  NAND2_X1 U7115 ( .A1(n7912), .A2(n8352), .ZN(n5588) );
  NAND2_X1 U7116 ( .A1(n4481), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5587) );
  INV_X1 U7117 ( .A(n8668), .ZN(n8995) );
  NAND2_X1 U7118 ( .A1(n5589), .A2(n9779), .ZN(n5590) );
  INV_X1 U7119 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8993) );
  NAND2_X1 U7120 ( .A1(n5674), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7121 ( .A1(n4487), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5592) );
  OAI211_X1 U7122 ( .C1(n8993), .C2(n5229), .A(n5593), .B(n5592), .ZN(n5594)
         );
  NAND2_X1 U7123 ( .A1(n8995), .A2(n8284), .ZN(n6556) );
  OR2_X1 U7124 ( .A1(n5595), .A2(n6556), .ZN(n5597) );
  NAND2_X1 U7125 ( .A1(n4840), .A2(n8650), .ZN(n5596) );
  INV_X1 U7126 ( .A(n5602), .ZN(n5599) );
  NAND2_X1 U7127 ( .A1(n8668), .A2(n8284), .ZN(n8515) );
  NAND2_X2 U7128 ( .A1(n8516), .A2(n8515), .ZN(n8659) );
  AND2_X1 U7129 ( .A1(n8659), .A2(n8379), .ZN(n5598) );
  AND2_X1 U7130 ( .A1(n8677), .A2(n5601), .ZN(n5600) );
  NAND2_X1 U7131 ( .A1(n8675), .A2(n5600), .ZN(n5606) );
  INV_X1 U7132 ( .A(n5601), .ZN(n5604) );
  NAND2_X1 U7133 ( .A1(n8999), .A2(n8702), .ZN(n6555) );
  AND2_X1 U7134 ( .A1(n6555), .A2(n5602), .ZN(n5603) );
  NAND2_X1 U7135 ( .A1(n5606), .A2(n5605), .ZN(n8638) );
  MUX2_X1 U7136 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7982), .Z(n5625) );
  INV_X1 U7137 ( .A(SI_28_), .ZN(n5626) );
  XNOR2_X1 U7138 ( .A(n5625), .B(n5626), .ZN(n5623) );
  NAND2_X1 U7139 ( .A1(n7931), .A2(n8352), .ZN(n5610) );
  NAND2_X1 U7140 ( .A1(n5222), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5609) );
  INV_X1 U7141 ( .A(n5613), .ZN(n5612) );
  AND2_X1 U7142 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5611) );
  NAND2_X1 U7143 ( .A1(n5612), .A2(n5611), .ZN(n7949) );
  INV_X1 U7144 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9935) );
  INV_X1 U7145 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6531) );
  OAI21_X1 U7146 ( .B1(n5613), .B2(n9935), .A(n6531), .ZN(n5614) );
  NAND2_X1 U7147 ( .A1(n7949), .A2(n5614), .ZN(n8642) );
  OR2_X1 U7148 ( .A1(n8642), .A2(n5615), .ZN(n5621) );
  INV_X1 U7149 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U7150 ( .A1(n5674), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7151 ( .A1(n4486), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5616) );
  OAI211_X1 U7152 ( .C1(n5618), .C2(n5229), .A(n5617), .B(n5616), .ZN(n5619)
         );
  INV_X1 U7153 ( .A(n5619), .ZN(n5620) );
  NAND2_X1 U7154 ( .A1(n8905), .A2(n8524), .ZN(n8522) );
  INV_X1 U7155 ( .A(n8524), .ZN(n8560) );
  NOR2_X1 U7156 ( .A1(n8905), .A2(n8560), .ZN(n5622) );
  INV_X1 U7157 ( .A(n5625), .ZN(n5627) );
  NAND2_X1 U7158 ( .A1(n5627), .A2(n5626), .ZN(n5628) );
  MUX2_X1 U7159 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n7982), .Z(n7975) );
  INV_X1 U7160 ( .A(SI_29_), .ZN(n5630) );
  XNOR2_X1 U7161 ( .A(n7975), .B(n5630), .ZN(n5631) );
  NAND2_X1 U7162 ( .A1(n9029), .A2(n8352), .ZN(n5633) );
  NAND2_X1 U7163 ( .A1(n4481), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5632) );
  INV_X1 U7164 ( .A(n7949), .ZN(n5639) );
  INV_X1 U7165 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6543) );
  NAND2_X1 U7166 ( .A1(n4487), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U7167 ( .A1(n5634), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5635) );
  OAI211_X1 U7168 ( .C1(n6543), .C2(n5637), .A(n5636), .B(n5635), .ZN(n5638)
         );
  AOI21_X1 U7169 ( .B1(n5639), .B2(n5195), .A(n5638), .ZN(n8649) );
  NAND2_X1 U7170 ( .A1(n7954), .A2(n8649), .ZN(n8533) );
  XNOR2_X1 U7171 ( .A(n5640), .B(n8530), .ZN(n7947) );
  NAND2_X1 U7172 ( .A1(n5641), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5699) );
  XNOR2_X1 U7173 ( .A(n5699), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8554) );
  NAND2_X1 U7174 ( .A1(n4505), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5642) );
  INV_X1 U7175 ( .A(n5643), .ZN(n5644) );
  NAND2_X1 U7176 ( .A1(n5644), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5645) );
  MUX2_X1 U7177 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5645), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5646) );
  NAND2_X1 U7178 ( .A1(n5646), .A2(n4505), .ZN(n8366) );
  NAND2_X1 U7179 ( .A1(n8407), .A2(n8366), .ZN(n7189) );
  XNOR2_X1 U7180 ( .A(n8554), .B(n7189), .ZN(n5647) );
  NAND2_X1 U7181 ( .A1(n5647), .A2(n8622), .ZN(n7882) );
  AND2_X1 U7182 ( .A1(n8366), .A2(n8390), .ZN(n5648) );
  NAND2_X1 U7183 ( .A1(n7661), .A2(n5648), .ZN(n10077) );
  NAND2_X1 U7184 ( .A1(n7882), .A2(n10077), .ZN(n10440) );
  INV_X1 U7185 ( .A(n7194), .ZN(n5651) );
  NAND2_X1 U7186 ( .A1(n5651), .A2(n7193), .ZN(n7195) );
  NAND2_X1 U7187 ( .A1(n7195), .A2(n8421), .ZN(n7345) );
  INV_X1 U7188 ( .A(n8403), .ZN(n5652) );
  AND2_X1 U7189 ( .A1(n8395), .A2(n7403), .ZN(n8398) );
  NAND2_X1 U7190 ( .A1(n7371), .A2(n8404), .ZN(n5654) );
  INV_X1 U7191 ( .A(n8368), .ZN(n5653) );
  NAND2_X1 U7192 ( .A1(n5654), .A2(n5653), .ZN(n7370) );
  INV_X1 U7193 ( .A(n7549), .ZN(n8430) );
  NAND2_X1 U7194 ( .A1(n7624), .A2(n8438), .ZN(n7664) );
  NAND2_X1 U7195 ( .A1(n7664), .A2(n8450), .ZN(n7739) );
  NAND2_X1 U7196 ( .A1(n7739), .A2(n8440), .ZN(n5655) );
  NAND2_X1 U7197 ( .A1(n5655), .A2(n8444), .ZN(n7741) );
  NAND2_X1 U7198 ( .A1(n7741), .A2(n8448), .ZN(n7759) );
  NAND2_X1 U7199 ( .A1(n8895), .A2(n8470), .ZN(n8857) );
  INV_X1 U7200 ( .A(n8865), .ZN(n8473) );
  NAND2_X1 U7201 ( .A1(n8857), .A2(n8473), .ZN(n8862) );
  INV_X1 U7202 ( .A(n8834), .ZN(n8838) );
  INV_X1 U7203 ( .A(n8810), .ZN(n5656) );
  NOR2_X1 U7204 ( .A1(n8821), .A2(n5656), .ZN(n8765) );
  NAND2_X1 U7205 ( .A1(n8950), .A2(n8304), .ZN(n8783) );
  NAND2_X1 U7206 ( .A1(n8946), .A2(n8321), .ZN(n8490) );
  AND2_X1 U7207 ( .A1(n8783), .A2(n8490), .ZN(n8767) );
  AND2_X1 U7208 ( .A1(n8767), .A2(n8496), .ZN(n5657) );
  AND2_X1 U7209 ( .A1(n8765), .A2(n5657), .ZN(n5663) );
  INV_X1 U7210 ( .A(n5657), .ZN(n5658) );
  OR2_X1 U7211 ( .A1(n8950), .A2(n8304), .ZN(n8488) );
  AND2_X1 U7212 ( .A1(n8488), .A2(n8800), .ZN(n8766) );
  OR2_X1 U7213 ( .A1(n5658), .A2(n8766), .ZN(n5662) );
  INV_X1 U7214 ( .A(n8496), .ZN(n5660) );
  INV_X1 U7215 ( .A(n8490), .ZN(n5659) );
  OR2_X1 U7216 ( .A1(n8946), .A2(n8321), .ZN(n8492) );
  OR2_X1 U7217 ( .A1(n5659), .A2(n8787), .ZN(n8768) );
  OR2_X1 U7218 ( .A1(n5660), .A2(n8768), .ZN(n5661) );
  NAND2_X1 U7219 ( .A1(n5664), .A2(n8493), .ZN(n8752) );
  XNOR2_X1 U7220 ( .A(n8935), .B(n8737), .ZN(n8751) );
  NAND2_X1 U7221 ( .A1(n8935), .A2(n8737), .ZN(n8495) );
  OAI21_X1 U7222 ( .B1(n8752), .B2(n8751), .A(n8495), .ZN(n8736) );
  INV_X1 U7223 ( .A(n8736), .ZN(n5665) );
  NAND2_X1 U7224 ( .A1(n5665), .A2(n8377), .ZN(n8712) );
  INV_X1 U7225 ( .A(n8711), .ZN(n8714) );
  INV_X1 U7226 ( .A(n8713), .ZN(n5666) );
  NOR2_X1 U7227 ( .A1(n8714), .A2(n5666), .ZN(n5667) );
  NAND2_X1 U7228 ( .A1(n8712), .A2(n5667), .ZN(n5668) );
  INV_X1 U7229 ( .A(n8701), .ZN(n5669) );
  NAND2_X1 U7230 ( .A1(n5670), .A2(n8508), .ZN(n8657) );
  NOR2_X1 U7231 ( .A1(n8685), .A2(n8702), .ZN(n8512) );
  NOR2_X1 U7232 ( .A1(n8659), .A2(n8512), .ZN(n5671) );
  NOR2_X1 U7233 ( .A1(n8388), .A2(n8650), .ZN(n8393) );
  NOR2_X1 U7234 ( .A1(n8648), .A2(n8647), .ZN(n8646) );
  INV_X1 U7235 ( .A(n8521), .ZN(n5672) );
  XNOR2_X1 U7236 ( .A(n8351), .B(n8530), .ZN(n5682) );
  NAND2_X1 U7237 ( .A1(n8554), .A2(n8390), .ZN(n8384) );
  NAND2_X1 U7238 ( .A1(n8407), .A2(n8546), .ZN(n8361) );
  NAND2_X1 U7239 ( .A1(n8384), .A2(n8361), .ZN(n10357) );
  NAND2_X1 U7240 ( .A1(n8554), .A2(n8407), .ZN(n6696) );
  NOR2_X2 U7241 ( .A1(n5673), .A2(n6696), .ZN(n8816) );
  AND2_X1 U7242 ( .A1(n8560), .A2(n8816), .ZN(n5680) );
  INV_X1 U7243 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7244 ( .A1(n4486), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U7245 ( .A1(n5674), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5675) );
  OAI211_X1 U7246 ( .C1(n5229), .C2(n5677), .A(n5676), .B(n5675), .ZN(n8559)
         );
  INV_X1 U7247 ( .A(n6696), .ZN(n6794) );
  NAND2_X1 U7248 ( .A1(n5673), .A2(n6794), .ZN(n8890) );
  INV_X1 U7249 ( .A(P2_B_REG_SCAN_IN), .ZN(n9956) );
  NOR2_X1 U7250 ( .A1(n8552), .A2(n9956), .ZN(n5678) );
  NOR2_X1 U7251 ( .A1(n8890), .A2(n5678), .ZN(n8630) );
  INV_X1 U7252 ( .A(n7954), .ZN(n5724) );
  NAND2_X1 U7253 ( .A1(n7745), .A2(n7748), .ZN(n7746) );
  INV_X1 U7254 ( .A(n8886), .ZN(n9020) );
  INV_X1 U7255 ( .A(n8825), .ZN(n9013) );
  INV_X1 U7256 ( .A(n8940), .ZN(n8764) );
  INV_X1 U7257 ( .A(n8905), .ZN(n8645) );
  INV_X1 U7258 ( .A(n5683), .ZN(n8641) );
  OR2_X4 U7259 ( .A1(n8385), .A2(n8546), .ZN(n10436) );
  OAI211_X1 U7260 ( .C1(n5724), .C2(n8641), .A(n8634), .B(n8951), .ZN(n7951)
         );
  NAND2_X1 U7261 ( .A1(n7957), .A2(n7951), .ZN(n5684) );
  NOR4_X1 U7262 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5693) );
  INV_X1 U7263 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10400) );
  INV_X1 U7264 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10399) );
  INV_X1 U7265 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n10398) );
  INV_X1 U7266 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10397) );
  NAND4_X1 U7267 ( .A1(n10400), .A2(n10399), .A3(n10398), .A4(n10397), .ZN(
        n5690) );
  NOR4_X1 U7268 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5688) );
  NOR4_X1 U7269 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5687) );
  NOR4_X1 U7270 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5686) );
  NOR4_X1 U7271 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5685) );
  NAND4_X1 U7272 ( .A1(n5688), .A2(n5687), .A3(n5686), .A4(n5685), .ZN(n5689)
         );
  NOR4_X1 U7273 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n5690), .A4(n5689), .ZN(n5692) );
  NOR4_X1 U7274 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5691) );
  NAND3_X1 U7275 ( .A1(n5693), .A2(n5692), .A3(n5691), .ZN(n5709) );
  NAND2_X1 U7276 ( .A1(n5694), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5695) );
  MUX2_X1 U7277 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5695), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5697) );
  NAND2_X1 U7278 ( .A1(n5697), .A2(n5705), .ZN(n7827) );
  INV_X1 U7279 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5698) );
  NAND2_X1 U7280 ( .A1(n5699), .A2(n5698), .ZN(n5700) );
  NAND2_X1 U7281 ( .A1(n5700), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5713) );
  INV_X1 U7282 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U7283 ( .A1(n5713), .A2(n5712), .ZN(n5701) );
  NAND2_X1 U7284 ( .A1(n5701), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5703) );
  INV_X1 U7285 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5702) );
  XNOR2_X1 U7286 ( .A(n7791), .B(P2_B_REG_SCAN_IN), .ZN(n5704) );
  AND2_X1 U7287 ( .A1(n7827), .A2(n5704), .ZN(n5708) );
  NAND2_X1 U7288 ( .A1(n5705), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5706) );
  MUX2_X1 U7289 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5706), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5707) );
  NAND2_X1 U7290 ( .A1(n5707), .A2(n5162), .ZN(n7914) );
  AND2_X1 U7291 ( .A1(n5709), .A2(n10369), .ZN(n7185) );
  INV_X1 U7292 ( .A(n7791), .ZN(n5711) );
  NOR2_X1 U7293 ( .A1(n7914), .A2(n7827), .ZN(n5710) );
  NAND2_X1 U7294 ( .A1(n5711), .A2(n5710), .ZN(n6791) );
  AND2_X1 U7295 ( .A1(n8366), .A2(n8622), .ZN(n6533) );
  XNOR2_X1 U7296 ( .A(n5713), .B(n5712), .ZN(n6695) );
  OAI21_X1 U7297 ( .B1(n6696), .B2(n6533), .A(n6695), .ZN(n5714) );
  INV_X1 U7298 ( .A(n5714), .ZN(n5715) );
  NAND2_X1 U7299 ( .A1(n6791), .A2(n5715), .ZN(n6911) );
  NAND2_X1 U7300 ( .A1(n6527), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5716) );
  OR2_X1 U7301 ( .A1(n6911), .A2(n5716), .ZN(n5717) );
  NOR2_X1 U7302 ( .A1(n7185), .A2(n5717), .ZN(n5719) );
  INV_X1 U7303 ( .A(n10369), .ZN(n5718) );
  NAND2_X1 U7304 ( .A1(n7827), .A2(n7914), .ZN(n10403) );
  OAI21_X1 U7305 ( .B1(P2_D_REG_1__SCAN_IN), .B2(n5718), .A(n10403), .ZN(n6516) );
  INV_X1 U7306 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U7307 ( .A1(n10369), .A2(n5720), .ZN(n5721) );
  NAND2_X1 U7308 ( .A1(n7791), .A2(n7914), .ZN(n10401) );
  NAND2_X1 U7309 ( .A1(n5721), .A2(n10401), .ZN(n7182) );
  NAND2_X1 U7310 ( .A1(n10444), .A2(n8982), .ZN(n9019) );
  INV_X1 U7311 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5722) );
  OR2_X1 U7312 ( .A1(n10444), .A2(n5722), .ZN(n5723) );
  NOR2_X1 U7313 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5732) );
  NOR2_X1 U7314 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5731) );
  INV_X1 U7315 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5735) );
  INV_X2 U7316 ( .A(n5738), .ZN(n9625) );
  NAND2_X1 U7317 ( .A1(n6195), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5743) );
  INV_X1 U7318 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7014) );
  OR2_X1 U7319 ( .A1(n4484), .A2(n7014), .ZN(n5742) );
  NAND2_X4 U7320 ( .A1(n5737), .A2(n9625), .ZN(n8076) );
  INV_X1 U7321 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6631) );
  OR2_X1 U7322 ( .A1(n8076), .A2(n6631), .ZN(n5741) );
  INV_X1 U7323 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6639) );
  INV_X1 U7324 ( .A(n9168), .ZN(n7556) );
  INV_X1 U7325 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5750) );
  AND2_X1 U7326 ( .A1(n5750), .A2(n6128), .ZN(n5744) );
  NAND2_X1 U7327 ( .A1(n9992), .A2(n5744), .ZN(n5745) );
  INV_X1 U7328 ( .A(n6335), .ZN(n6337) );
  XNOR2_X1 U7329 ( .A(n5746), .B(P1_IR_REG_20__SCAN_IN), .ZN(n7074) );
  INV_X1 U7330 ( .A(n7334), .ZN(n5763) );
  NOR2_X1 U7331 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5752) );
  NOR2_X1 U7332 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5751) );
  NAND2_X1 U7333 ( .A1(n5756), .A2(n5757), .ZN(n5754) );
  INV_X1 U7334 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5755) );
  INV_X1 U7335 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5759) );
  OR2_X1 U7336 ( .A1(n5755), .A2(n5759), .ZN(n5760) );
  NAND2_X1 U7337 ( .A1(n5761), .A2(n5760), .ZN(n5762) );
  NAND2_X1 U7338 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  INV_X1 U7339 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U7340 ( .A1(n4503), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5770) );
  XNOR2_X1 U7341 ( .A(n5770), .B(n5769), .ZN(n9322) );
  NAND2_X1 U7342 ( .A1(n5786), .A2(n8242), .ZN(n7059) );
  INV_X1 U7343 ( .A(n5771), .ZN(n5772) );
  XNOR2_X2 U7344 ( .A(n5774), .B(n5734), .ZN(n6955) );
  INV_X1 U7345 ( .A(n6664), .ZN(n5775) );
  NAND2_X1 U7346 ( .A1(n5873), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5782) );
  NOR2_X1 U7347 ( .A1(n5776), .A2(n5755), .ZN(n5777) );
  MUX2_X1 U7348 ( .A(n5755), .B(n5777), .S(P1_IR_REG_2__SCAN_IN), .Z(n5780) );
  INV_X1 U7349 ( .A(n5778), .ZN(n5779) );
  NAND2_X1 U7350 ( .A1(n6629), .A2(n7020), .ZN(n5781) );
  AND3_X2 U7351 ( .A1(n5783), .A2(n5782), .A3(n5781), .ZN(n7333) );
  OAI22_X1 U7352 ( .A1(n7556), .A2(n5882), .B1(n7333), .B2(n5852), .ZN(n5829)
         );
  NAND2_X1 U7353 ( .A1(n9168), .A2(n5814), .ZN(n5785) );
  OR2_X1 U7354 ( .A1(n7333), .A2(n6306), .ZN(n5784) );
  NAND2_X1 U7355 ( .A1(n5785), .A2(n5784), .ZN(n5787) );
  NAND2_X4 U7356 ( .A1(n7058), .A2(n5763), .ZN(n7437) );
  XNOR2_X1 U7357 ( .A(n5787), .B(n7437), .ZN(n5828) );
  NAND2_X1 U7358 ( .A1(n6195), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5793) );
  INV_X1 U7359 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5788) );
  INV_X1 U7360 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5789) );
  INV_X1 U7361 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6743) );
  OR2_X1 U7362 ( .A1(n6376), .A2(n6743), .ZN(n5790) );
  NAND2_X1 U7363 ( .A1(n7982), .A2(SI_0_), .ZN(n5795) );
  INV_X1 U7364 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7365 ( .A1(n5795), .A2(n5794), .ZN(n5797) );
  AND2_X1 U7366 ( .A1(n5797), .A2(n5796), .ZN(n9627) );
  MUX2_X1 U7367 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9627), .S(n5798), .Z(n7480) );
  AOI22_X1 U7368 ( .A1(n5814), .A2(n7480), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n5799), .ZN(n5800) );
  AND2_X1 U7369 ( .A1(n5801), .A2(n5800), .ZN(n6937) );
  NOR2_X1 U7370 ( .A1(n6598), .A2(n6743), .ZN(n5802) );
  AOI21_X1 U7371 ( .B1(n5803), .B2(n7480), .A(n5802), .ZN(n5805) );
  NAND2_X1 U7372 ( .A1(n7063), .A2(n5814), .ZN(n5804) );
  AND2_X1 U7373 ( .A1(n5805), .A2(n5804), .ZN(n5806) );
  INV_X1 U7374 ( .A(n5806), .ZN(n6936) );
  NAND2_X1 U7375 ( .A1(n6937), .A2(n6936), .ZN(n6935) );
  NAND2_X1 U7376 ( .A1(n5806), .A2(n7437), .ZN(n5807) );
  NAND2_X1 U7377 ( .A1(n6935), .A2(n5807), .ZN(n5823) );
  INV_X1 U7378 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U7379 ( .A1(n6195), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5812) );
  INV_X1 U7380 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5809) );
  OR2_X2 U7381 ( .A1(n8076), .A2(n5809), .ZN(n5811) );
  INV_X1 U7382 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7430) );
  OR2_X1 U7383 ( .A1(n5888), .A2(n7430), .ZN(n5810) );
  NAND2_X1 U7384 ( .A1(n7062), .A2(n5814), .ZN(n5821) );
  INV_X1 U7385 ( .A(n6677), .ZN(n5815) );
  NAND2_X1 U7386 ( .A1(n5834), .A2(n5815), .ZN(n5819) );
  NAND2_X1 U7387 ( .A1(n5873), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5818) );
  INV_X1 U7388 ( .A(n5776), .ZN(n5816) );
  NAND2_X1 U7389 ( .A1(n6629), .A2(n7007), .ZN(n5817) );
  NAND2_X1 U7390 ( .A1(n5821), .A2(n5820), .ZN(n5822) );
  INV_X4 U7391 ( .A(n7437), .ZN(n6254) );
  XNOR2_X1 U7392 ( .A(n5822), .B(n6254), .ZN(n5824) );
  NAND2_X1 U7393 ( .A1(n5823), .A2(n5824), .ZN(n7049) );
  INV_X1 U7394 ( .A(n7062), .ZN(n8211) );
  OAI22_X1 U7395 ( .A1(n8211), .A2(n5882), .B1(n7274), .B2(n5852), .ZN(n7052)
         );
  NAND2_X1 U7396 ( .A1(n7049), .A2(n7052), .ZN(n5827) );
  INV_X1 U7397 ( .A(n5823), .ZN(n5826) );
  INV_X1 U7398 ( .A(n5824), .ZN(n5825) );
  NAND2_X1 U7399 ( .A1(n5826), .A2(n5825), .ZN(n7050) );
  NAND2_X1 U7400 ( .A1(n6195), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5833) );
  INV_X1 U7401 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6642) );
  OR2_X1 U7402 ( .A1(n6376), .A2(n6642), .ZN(n5832) );
  INV_X1 U7403 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6632) );
  OR2_X1 U7404 ( .A1(n8076), .A2(n6632), .ZN(n5831) );
  OR2_X1 U7405 ( .A1(n4485), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U7406 ( .A1(n9167), .A2(n6332), .ZN(n5841) );
  INV_X1 U7407 ( .A(n6667), .ZN(n5835) );
  NAND2_X1 U7408 ( .A1(n5873), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U7409 ( .A1(n5778), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5836) );
  XNOR2_X1 U7410 ( .A(n5836), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6775) );
  NAND2_X1 U7411 ( .A1(n6629), .A2(n6775), .ZN(n5837) );
  AND3_X2 U7412 ( .A1(n5839), .A2(n5838), .A3(n5837), .ZN(n10292) );
  OR2_X1 U7413 ( .A1(n10292), .A2(n6306), .ZN(n5840) );
  NAND2_X1 U7414 ( .A1(n5841), .A2(n5840), .ZN(n5842) );
  XNOR2_X1 U7415 ( .A(n5842), .B(n6254), .ZN(n5845) );
  INV_X1 U7416 ( .A(n9167), .ZN(n7303) );
  OAI22_X1 U7417 ( .A1(n7303), .A2(n5882), .B1(n10292), .B2(n5852), .ZN(n5843)
         );
  XNOR2_X1 U7418 ( .A(n5845), .B(n5843), .ZN(n7082) );
  INV_X1 U7419 ( .A(n5843), .ZN(n5844) );
  NAND2_X1 U7420 ( .A1(n5845), .A2(n5844), .ZN(n5846) );
  NAND2_X1 U7421 ( .A1(n6195), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5851) );
  INV_X1 U7422 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5847) );
  OR2_X1 U7423 ( .A1(n6376), .A2(n5847), .ZN(n5850) );
  XNOR2_X1 U7424 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7939) );
  OR2_X1 U7425 ( .A1(n4484), .A2(n7939), .ZN(n5849) );
  INV_X1 U7426 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6633) );
  OR2_X1 U7427 ( .A1(n8076), .A2(n6633), .ZN(n5848) );
  NAND4_X1 U7428 ( .A1(n5851), .A2(n5850), .A3(n5849), .A4(n5848), .ZN(n9166)
         );
  NAND2_X1 U7429 ( .A1(n9166), .A2(n6332), .ZN(n5860) );
  INV_X1 U7430 ( .A(n6680), .ZN(n5853) );
  NAND2_X1 U7431 ( .A1(n6265), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U7432 ( .A1(n5854), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5855) );
  XNOR2_X1 U7433 ( .A(n5855), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6954) );
  NAND2_X1 U7434 ( .A1(n6629), .A2(n6954), .ZN(n5856) );
  AND3_X2 U7435 ( .A1(n5858), .A2(n5857), .A3(n5856), .ZN(n7940) );
  OR2_X1 U7436 ( .A1(n7940), .A2(n6306), .ZN(n5859) );
  INV_X1 U7437 ( .A(n9166), .ZN(n7555) );
  OAI22_X1 U7438 ( .A1(n7555), .A2(n5882), .B1(n7940), .B2(n5852), .ZN(n5862)
         );
  NAND2_X1 U7439 ( .A1(n5863), .A2(n5862), .ZN(n5864) );
  AOI21_X1 U7440 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5865) );
  NOR2_X1 U7441 ( .A1(n5865), .A2(n5889), .ZN(n9085) );
  NAND2_X1 U7442 ( .A1(n6299), .A2(n9085), .ZN(n5871) );
  INV_X1 U7443 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5866) );
  OR2_X1 U7444 ( .A1(n6376), .A2(n5866), .ZN(n5870) );
  INV_X1 U7445 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5867) );
  OR2_X1 U7446 ( .A1(n6134), .A2(n5867), .ZN(n5869) );
  INV_X1 U7447 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6634) );
  OR2_X1 U7448 ( .A1(n8076), .A2(n6634), .ZN(n5868) );
  NAND4_X1 U7449 ( .A1(n5871), .A2(n5870), .A3(n5869), .A4(n5868), .ZN(n9165)
         );
  NAND2_X1 U7450 ( .A1(n9165), .A2(n6332), .ZN(n5880) );
  INV_X1 U7451 ( .A(n6673), .ZN(n5872) );
  NAND2_X1 U7452 ( .A1(n6265), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5877) );
  OR2_X1 U7453 ( .A1(n5874), .A2(n5755), .ZN(n5875) );
  XNOR2_X1 U7454 ( .A(n5875), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U7455 ( .A1(n6629), .A2(n6757), .ZN(n5876) );
  OR2_X1 U7456 ( .A1(n9081), .A2(n6306), .ZN(n5879) );
  NAND2_X1 U7457 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  XNOR2_X1 U7458 ( .A(n5881), .B(n6254), .ZN(n5884) );
  NOR2_X1 U7459 ( .A1(n9081), .A2(n5852), .ZN(n5883) );
  AOI21_X1 U7460 ( .B1(n6308), .B2(n9165), .A(n5883), .ZN(n9078) );
  NAND2_X1 U7461 ( .A1(n9079), .A2(n9078), .ZN(n9077) );
  INV_X1 U7462 ( .A(n5884), .ZN(n5885) );
  OR2_X1 U7463 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  NAND2_X1 U7464 ( .A1(n9077), .A2(n5887), .ZN(n7381) );
  NAND2_X1 U7465 ( .A1(n6195), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5893) );
  INV_X1 U7466 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6644) );
  OR2_X1 U7467 ( .A1(n6376), .A2(n6644), .ZN(n5892) );
  OAI21_X1 U7468 ( .B1(n5889), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5908), .ZN(
        n7514) );
  OR2_X1 U7469 ( .A1(n4485), .A2(n7514), .ZN(n5891) );
  INV_X1 U7470 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7515) );
  OR2_X1 U7471 ( .A1(n8076), .A2(n7515), .ZN(n5890) );
  NAND4_X1 U7472 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), .ZN(n9164)
         );
  NAND2_X1 U7473 ( .A1(n9164), .A2(n6332), .ZN(n5901) );
  INV_X1 U7474 ( .A(n6682), .ZN(n5894) );
  NAND2_X1 U7475 ( .A1(n6265), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5898) );
  OR2_X1 U7476 ( .A1(n5895), .A2(n5755), .ZN(n5896) );
  XNOR2_X1 U7477 ( .A(n5896), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6645) );
  NAND2_X1 U7478 ( .A1(n6629), .A2(n6645), .ZN(n5897) );
  OR2_X1 U7479 ( .A1(n10304), .A2(n6306), .ZN(n5900) );
  NAND2_X1 U7480 ( .A1(n5901), .A2(n5900), .ZN(n5902) );
  XNOR2_X1 U7481 ( .A(n5902), .B(n6254), .ZN(n5905) );
  INV_X1 U7482 ( .A(n9164), .ZN(n9082) );
  OAI22_X1 U7483 ( .A1(n9082), .A2(n5882), .B1(n10304), .B2(n5852), .ZN(n5903)
         );
  XNOR2_X1 U7484 ( .A(n5905), .B(n5903), .ZN(n7382) );
  INV_X1 U7485 ( .A(n5903), .ZN(n5904) );
  NAND2_X1 U7486 ( .A1(n5905), .A2(n5904), .ZN(n5906) );
  NAND2_X1 U7487 ( .A1(n6195), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5914) );
  INV_X1 U7488 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7470) );
  OR2_X1 U7489 ( .A1(n8076), .A2(n7470), .ZN(n5913) );
  AND2_X1 U7490 ( .A1(n5908), .A2(n5907), .ZN(n5909) );
  OR2_X1 U7491 ( .A1(n5909), .A2(n5928), .ZN(n7534) );
  OR2_X1 U7492 ( .A1(n4485), .A2(n7534), .ZN(n5912) );
  INV_X1 U7493 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5910) );
  OR2_X1 U7494 ( .A1(n6376), .A2(n5910), .ZN(n5911) );
  NAND4_X1 U7495 ( .A1(n5914), .A2(n5913), .A3(n5912), .A4(n5911), .ZN(n9163)
         );
  NAND2_X1 U7496 ( .A1(n9163), .A2(n6332), .ZN(n5921) );
  OR2_X1 U7497 ( .A1(n6024), .A2(n6685), .ZN(n5919) );
  NAND2_X1 U7498 ( .A1(n6265), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n5918) );
  INV_X1 U7499 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U7500 ( .A1(n5895), .A2(n5915), .ZN(n5935) );
  NAND2_X1 U7501 ( .A1(n5935), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5916) );
  XNOR2_X1 U7502 ( .A(n5916), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6768) );
  NAND2_X1 U7503 ( .A1(n6629), .A2(n6768), .ZN(n5917) );
  INV_X1 U7504 ( .A(n10312), .ZN(n7476) );
  NAND2_X1 U7505 ( .A1(n7476), .A2(n6317), .ZN(n5920) );
  NAND2_X1 U7506 ( .A1(n5921), .A2(n5920), .ZN(n5922) );
  XNOR2_X1 U7507 ( .A(n5922), .B(n6254), .ZN(n7528) );
  NOR2_X1 U7508 ( .A1(n10312), .A2(n5852), .ZN(n5923) );
  AOI21_X1 U7509 ( .B1(n6308), .B2(n9163), .A(n5923), .ZN(n5924) );
  AND2_X1 U7510 ( .A1(n7528), .A2(n5924), .ZN(n5927) );
  INV_X1 U7511 ( .A(n7528), .ZN(n5925) );
  INV_X1 U7512 ( .A(n5924), .ZN(n7529) );
  NAND2_X1 U7513 ( .A1(n5925), .A2(n7529), .ZN(n5926) );
  NAND2_X1 U7514 ( .A1(n6195), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5934) );
  INV_X1 U7515 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7593) );
  OR2_X1 U7516 ( .A1(n8076), .A2(n7593), .ZN(n5933) );
  NAND2_X1 U7517 ( .A1(n5928), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5950) );
  OR2_X1 U7518 ( .A1(n5928), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7519 ( .A1(n5950), .A2(n5929), .ZN(n7643) );
  OR2_X1 U7520 ( .A1(n4484), .A2(n7643), .ZN(n5932) );
  INV_X1 U7521 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5930) );
  OR2_X1 U7522 ( .A1(n6376), .A2(n5930), .ZN(n5931) );
  NAND4_X1 U7523 ( .A1(n5934), .A2(n5933), .A3(n5932), .A4(n5931), .ZN(n10262)
         );
  NAND2_X1 U7524 ( .A1(n5945), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5936) );
  XNOR2_X1 U7525 ( .A(n5936), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6738) );
  AOI22_X1 U7526 ( .A1(n6265), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6629), .B2(
        n6738), .ZN(n5937) );
  INV_X1 U7527 ( .A(n10316), .ZN(n7685) );
  AOI22_X1 U7528 ( .A1(n6308), .A2(n10262), .B1(n7685), .B2(n6309), .ZN(n7638)
         );
  NAND2_X1 U7529 ( .A1(n10262), .A2(n6332), .ZN(n5940) );
  OR2_X1 U7530 ( .A1(n6306), .A2(n10316), .ZN(n5939) );
  NAND2_X1 U7531 ( .A1(n5940), .A2(n5939), .ZN(n5941) );
  XNOR2_X1 U7532 ( .A(n5941), .B(n6254), .ZN(n7637) );
  INV_X1 U7533 ( .A(n7637), .ZN(n5943) );
  INV_X1 U7534 ( .A(n7638), .ZN(n5942) );
  NAND2_X1 U7535 ( .A1(n5943), .A2(n5942), .ZN(n5944) );
  NAND2_X1 U7536 ( .A1(n5966), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5946) );
  XNOR2_X1 U7537 ( .A(n5946), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6882) );
  AOI22_X1 U7538 ( .A1(n6265), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6629), .B2(
        n6882), .ZN(n5947) );
  NAND2_X1 U7539 ( .A1(n10277), .A2(n6317), .ZN(n5959) );
  NAND2_X1 U7540 ( .A1(n6195), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U7541 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  NAND2_X1 U7542 ( .A1(n5972), .A2(n5951), .ZN(n10273) );
  OR2_X1 U7543 ( .A1(n4485), .A2(n10273), .ZN(n5956) );
  INV_X1 U7544 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n5952) );
  OR2_X1 U7545 ( .A1(n8076), .A2(n5952), .ZN(n5955) );
  INV_X1 U7546 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5953) );
  OR2_X1 U7547 ( .A1(n6376), .A2(n5953), .ZN(n5954) );
  NAND4_X1 U7548 ( .A1(n5957), .A2(n5956), .A3(n5955), .A4(n5954), .ZN(n9162)
         );
  NAND2_X1 U7549 ( .A1(n9162), .A2(n6332), .ZN(n5958) );
  NAND2_X1 U7550 ( .A1(n5959), .A2(n5958), .ZN(n5960) );
  XNOR2_X1 U7551 ( .A(n5960), .B(n6254), .ZN(n5962) );
  AOI22_X1 U7552 ( .A1(n6308), .A2(n9162), .B1(n10277), .B2(n6309), .ZN(n5961)
         );
  NAND2_X1 U7553 ( .A1(n5962), .A2(n5961), .ZN(n5965) );
  OR2_X1 U7554 ( .A1(n5962), .A2(n5961), .ZN(n5963) );
  NAND2_X1 U7555 ( .A1(n5965), .A2(n5963), .ZN(n7707) );
  OAI21_X1 U7556 ( .B1(n5966), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5968) );
  OR2_X1 U7557 ( .A1(n5968), .A2(n5967), .ZN(n5969) );
  NAND2_X1 U7558 ( .A1(n5968), .A2(n5967), .ZN(n5984) );
  AOI22_X1 U7559 ( .A1(n6265), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6629), .B2(
        n6962), .ZN(n5970) );
  NAND2_X1 U7560 ( .A1(n7831), .A2(n6317), .ZN(n5979) );
  NAND2_X1 U7561 ( .A1(n6195), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5977) );
  INV_X1 U7562 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6885) );
  OR2_X1 U7563 ( .A1(n6376), .A2(n6885), .ZN(n5976) );
  NAND2_X1 U7564 ( .A1(n5972), .A2(n6894), .ZN(n5973) );
  NAND2_X1 U7565 ( .A1(n5991), .A2(n5973), .ZN(n7699) );
  OR2_X1 U7566 ( .A1(n4484), .A2(n7699), .ZN(n5975) );
  INV_X1 U7567 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6889) );
  OR2_X1 U7568 ( .A1(n8076), .A2(n6889), .ZN(n5974) );
  OR2_X1 U7569 ( .A1(n10130), .A2(n5852), .ZN(n5978) );
  NAND2_X1 U7570 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  XNOR2_X1 U7571 ( .A(n5980), .B(n6254), .ZN(n5982) );
  AOI22_X1 U7572 ( .A1(n7831), .A2(n6332), .B1(n10265), .B2(n6308), .ZN(n5981)
         );
  OR2_X1 U7573 ( .A1(n5982), .A2(n5981), .ZN(n7726) );
  NAND2_X1 U7574 ( .A1(n7724), .A2(n7726), .ZN(n5983) );
  NAND2_X1 U7575 ( .A1(n5982), .A2(n5981), .ZN(n7725) );
  NAND2_X1 U7576 ( .A1(n5984), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5986) );
  INV_X1 U7577 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5985) );
  XNOR2_X1 U7578 ( .A(n5986), .B(n5985), .ZN(n7123) );
  INV_X1 U7579 ( .A(n7123), .ZN(n5987) );
  AOI22_X1 U7580 ( .A1(n5873), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6629), .B2(
        n5987), .ZN(n5988) );
  NAND2_X1 U7581 ( .A1(n10163), .A2(n6317), .ZN(n5998) );
  NAND2_X1 U7582 ( .A1(n6195), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5996) );
  INV_X1 U7583 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6971) );
  OR2_X1 U7584 ( .A1(n6376), .A2(n6971), .ZN(n5995) );
  INV_X1 U7585 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5990) );
  AND2_X1 U7586 ( .A1(n5991), .A2(n5990), .ZN(n5992) );
  OR2_X1 U7587 ( .A1(n5992), .A2(n6010), .ZN(n10136) );
  OR2_X1 U7588 ( .A1(n4485), .A2(n10136), .ZN(n5994) );
  INV_X1 U7589 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7122) );
  OR2_X1 U7590 ( .A1(n8076), .A2(n7122), .ZN(n5993) );
  NAND4_X1 U7591 ( .A1(n5996), .A2(n5995), .A3(n5994), .A4(n5993), .ZN(n9161)
         );
  NAND2_X1 U7592 ( .A1(n9161), .A2(n6332), .ZN(n5997) );
  NAND2_X1 U7593 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  XNOR2_X1 U7594 ( .A(n5999), .B(n6254), .ZN(n6001) );
  INV_X1 U7595 ( .A(n9161), .ZN(n10060) );
  NOR2_X1 U7596 ( .A1(n10060), .A2(n5882), .ZN(n6000) );
  AOI21_X1 U7597 ( .B1(n10163), .B2(n6309), .A(n6000), .ZN(n6002) );
  XNOR2_X1 U7598 ( .A(n6001), .B(n6002), .ZN(n7860) );
  INV_X1 U7599 ( .A(n6001), .ZN(n6004) );
  INV_X1 U7600 ( .A(n6002), .ZN(n6003) );
  NAND2_X1 U7601 ( .A1(n6004), .A2(n6003), .ZN(n6005) );
  NAND2_X1 U7602 ( .A1(n5747), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6006) );
  XNOR2_X1 U7603 ( .A(n6006), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9179) );
  AOI22_X1 U7604 ( .A1(n6265), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6629), .B2(
        n9179), .ZN(n6007) );
  NAND2_X1 U7605 ( .A1(n7893), .A2(n6317), .ZN(n6017) );
  NAND2_X1 U7606 ( .A1(n6195), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6015) );
  INV_X1 U7607 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7840) );
  OR2_X1 U7608 ( .A1(n8076), .A2(n7840), .ZN(n6014) );
  INV_X1 U7609 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6009) );
  OR2_X1 U7610 ( .A1(n6376), .A2(n6009), .ZN(n6013) );
  NOR2_X1 U7611 ( .A1(n6010), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6011) );
  OR2_X1 U7612 ( .A1(n6029), .A2(n6011), .ZN(n10071) );
  OR2_X1 U7613 ( .A1(n4484), .A2(n10071), .ZN(n6012) );
  OR2_X1 U7614 ( .A1(n10127), .A2(n5852), .ZN(n6016) );
  NAND2_X1 U7615 ( .A1(n6017), .A2(n6016), .ZN(n6018) );
  XNOR2_X1 U7616 ( .A(n6018), .B(n7437), .ZN(n6020) );
  NOR2_X1 U7617 ( .A1(n10127), .A2(n5882), .ZN(n6019) );
  AOI21_X1 U7618 ( .B1(n7893), .B2(n6309), .A(n6019), .ZN(n6021) );
  XNOR2_X1 U7619 ( .A(n6020), .B(n6021), .ZN(n10065) );
  INV_X1 U7620 ( .A(n6020), .ZN(n6022) );
  NAND2_X1 U7621 ( .A1(n6022), .A2(n6021), .ZN(n6023) );
  NAND2_X1 U7622 ( .A1(n6785), .A2(n8072), .ZN(n6028) );
  NAND2_X1 U7623 ( .A1(n6025), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6026) );
  XNOR2_X1 U7624 ( .A(n6026), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U7625 ( .A1(n6265), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6629), .B2(
        n10187), .ZN(n6027) );
  NAND2_X1 U7626 ( .A1(n10122), .A2(n6317), .ZN(n6037) );
  NAND2_X1 U7627 ( .A1(n6195), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6035) );
  INV_X1 U7628 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9182) );
  OR2_X1 U7629 ( .A1(n6376), .A2(n9182), .ZN(n6034) );
  NOR2_X1 U7630 ( .A1(n6029), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6030) );
  OR2_X1 U7631 ( .A1(n6047), .A2(n6030), .ZN(n10117) );
  OR2_X1 U7632 ( .A1(n4485), .A2(n10117), .ZN(n6033) );
  INV_X1 U7633 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6031) );
  OR2_X1 U7634 ( .A1(n8076), .A2(n6031), .ZN(n6032) );
  NAND4_X1 U7635 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(n10089)
         );
  NAND2_X1 U7636 ( .A1(n10089), .A2(n6332), .ZN(n6036) );
  NAND2_X1 U7637 ( .A1(n6037), .A2(n6036), .ZN(n6038) );
  XNOR2_X1 U7638 ( .A(n6038), .B(n6254), .ZN(n7866) );
  INV_X1 U7639 ( .A(n10089), .ZN(n10059) );
  NOR2_X1 U7640 ( .A1(n10059), .A2(n5882), .ZN(n6039) );
  AOI21_X1 U7641 ( .B1(n10122), .B2(n6309), .A(n6039), .ZN(n7865) );
  AND2_X1 U7642 ( .A1(n7866), .A2(n7865), .ZN(n6043) );
  INV_X1 U7643 ( .A(n7866), .ZN(n6041) );
  INV_X1 U7644 ( .A(n7865), .ZN(n6040) );
  NAND2_X1 U7645 ( .A1(n6041), .A2(n6040), .ZN(n6042) );
  NAND2_X1 U7646 ( .A1(n6788), .A2(n8072), .ZN(n6046) );
  OR2_X1 U7647 ( .A1(n6044), .A2(n5755), .ZN(n6063) );
  INV_X1 U7648 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6062) );
  XNOR2_X1 U7649 ( .A(n6063), .B(n6062), .ZN(n9184) );
  INV_X1 U7650 ( .A(n9184), .ZN(n10199) );
  AOI22_X1 U7651 ( .A1(n6265), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6629), .B2(
        n10199), .ZN(n6045) );
  NAND2_X1 U7652 ( .A1(n10096), .A2(n6317), .ZN(n6055) );
  NAND2_X1 U7653 ( .A1(n6195), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6053) );
  INV_X1 U7654 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9183) );
  OR2_X1 U7655 ( .A1(n6376), .A2(n9183), .ZN(n6052) );
  INV_X1 U7656 ( .A(n6047), .ZN(n6048) );
  INV_X1 U7657 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10088) );
  NAND2_X1 U7658 ( .A1(n6048), .A2(n10088), .ZN(n6049) );
  NAND2_X1 U7659 ( .A1(n6070), .A2(n6049), .ZN(n10105) );
  OR2_X1 U7660 ( .A1(n4484), .A2(n10105), .ZN(n6051) );
  INV_X1 U7661 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7906) );
  OR2_X1 U7662 ( .A1(n8076), .A2(n7906), .ZN(n6050) );
  NAND4_X1 U7663 ( .A1(n6053), .A2(n6052), .A3(n6051), .A4(n6050), .ZN(n9217)
         );
  NAND2_X1 U7664 ( .A1(n9217), .A2(n6332), .ZN(n6054) );
  NAND2_X1 U7665 ( .A1(n6055), .A2(n6054), .ZN(n6056) );
  XNOR2_X1 U7666 ( .A(n6056), .B(n6254), .ZN(n10098) );
  INV_X1 U7667 ( .A(n9217), .ZN(n10109) );
  NOR2_X1 U7668 ( .A1(n10109), .A2(n5882), .ZN(n6057) );
  AOI21_X1 U7669 ( .B1(n10096), .B2(n6309), .A(n6057), .ZN(n10097) );
  NAND2_X1 U7670 ( .A1(n10098), .A2(n10097), .ZN(n6058) );
  INV_X1 U7671 ( .A(n10098), .ZN(n6060) );
  INV_X1 U7672 ( .A(n10097), .ZN(n6059) );
  NAND2_X1 U7673 ( .A1(n6060), .A2(n6059), .ZN(n6061) );
  NAND2_X1 U7674 ( .A1(n7024), .A2(n8072), .ZN(n6067) );
  NAND2_X1 U7675 ( .A1(n6063), .A2(n6062), .ZN(n6064) );
  NAND2_X1 U7676 ( .A1(n6064), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6065) );
  XNOR2_X1 U7677 ( .A(n6065), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U7678 ( .A1(n6265), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6629), .B2(
        n10212), .ZN(n6066) );
  NAND2_X1 U7679 ( .A1(n6195), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6075) );
  INV_X1 U7680 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6068) );
  OR2_X1 U7681 ( .A1(n6376), .A2(n6068), .ZN(n6074) );
  INV_X1 U7682 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7683 ( .A1(n6070), .A2(n6069), .ZN(n6071) );
  NAND2_X1 U7684 ( .A1(n6089), .A2(n6071), .ZN(n9506) );
  OR2_X1 U7685 ( .A1(n4485), .A2(n9506), .ZN(n6073) );
  INV_X1 U7686 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9507) );
  OR2_X1 U7687 ( .A1(n8076), .A2(n9507), .ZN(n6072) );
  OAI22_X1 U7688 ( .A1(n9592), .A2(n6306), .B1(n10093), .B2(n5852), .ZN(n6076)
         );
  XNOR2_X1 U7689 ( .A(n6076), .B(n6254), .ZN(n9149) );
  OR2_X1 U7690 ( .A1(n9592), .A2(n5852), .ZN(n6078) );
  INV_X1 U7691 ( .A(n10093), .ZN(n9220) );
  NAND2_X1 U7692 ( .A1(n9220), .A2(n6308), .ZN(n6077) );
  AND2_X1 U7693 ( .A1(n6078), .A2(n6077), .ZN(n6080) );
  NAND2_X1 U7694 ( .A1(n9149), .A2(n6080), .ZN(n6079) );
  NAND2_X1 U7695 ( .A1(n9147), .A2(n6079), .ZN(n6083) );
  INV_X1 U7696 ( .A(n9149), .ZN(n6081) );
  INV_X1 U7697 ( .A(n6080), .ZN(n9148) );
  NAND2_X1 U7698 ( .A1(n6081), .A2(n9148), .ZN(n6082) );
  NAND2_X1 U7699 ( .A1(n7090), .A2(n8072), .ZN(n6086) );
  NAND2_X1 U7700 ( .A1(n6107), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6084) );
  XNOR2_X1 U7701 ( .A(n6084), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10223) );
  AOI22_X1 U7702 ( .A1(n5873), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6629), .B2(
        n10223), .ZN(n6085) );
  NAND2_X1 U7703 ( .A1(n9483), .A2(n6317), .ZN(n6096) );
  NAND2_X1 U7704 ( .A1(n6195), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6094) );
  INV_X1 U7705 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9188) );
  OR2_X1 U7706 ( .A1(n6376), .A2(n9188), .ZN(n6093) );
  INV_X1 U7707 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7708 ( .A1(n6089), .A2(n6088), .ZN(n6090) );
  NAND2_X1 U7709 ( .A1(n6113), .A2(n6090), .ZN(n9486) );
  OR2_X1 U7710 ( .A1(n4485), .A2(n9486), .ZN(n6092) );
  INV_X1 U7711 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9487) );
  OR2_X1 U7712 ( .A1(n8076), .A2(n9487), .ZN(n6091) );
  OR2_X1 U7713 ( .A1(n9496), .A2(n5852), .ZN(n6095) );
  NAND2_X1 U7714 ( .A1(n6096), .A2(n6095), .ZN(n6097) );
  XNOR2_X1 U7715 ( .A(n6097), .B(n6254), .ZN(n6099) );
  NOR2_X1 U7716 ( .A1(n9496), .A2(n5882), .ZN(n6098) );
  AOI21_X1 U7717 ( .B1(n9483), .B2(n6309), .A(n6098), .ZN(n6100) );
  NAND2_X1 U7718 ( .A1(n6099), .A2(n6100), .ZN(n6106) );
  INV_X1 U7719 ( .A(n6099), .ZN(n6102) );
  INV_X1 U7720 ( .A(n6100), .ZN(n6101) );
  NAND2_X1 U7721 ( .A1(n6102), .A2(n6101), .ZN(n6103) );
  NAND2_X1 U7722 ( .A1(n6106), .A2(n6103), .ZN(n9071) );
  INV_X1 U7723 ( .A(n9071), .ZN(n6104) );
  NAND2_X1 U7724 ( .A1(n7154), .A2(n8072), .ZN(n6110) );
  OR2_X1 U7725 ( .A1(n6107), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7726 ( .A1(n6108), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6129) );
  XNOR2_X1 U7727 ( .A(n6129), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10236) );
  AOI22_X1 U7728 ( .A1(n6265), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6629), .B2(
        n10236), .ZN(n6109) );
  NAND2_X1 U7729 ( .A1(n9581), .A2(n6317), .ZN(n6121) );
  INV_X1 U7730 ( .A(n6376), .ZN(n6196) );
  NAND2_X1 U7731 ( .A1(n6196), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6119) );
  INV_X1 U7732 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n6111) );
  OR2_X1 U7733 ( .A1(n6134), .A2(n6111), .ZN(n6118) );
  INV_X1 U7734 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7735 ( .A1(n6113), .A2(n6112), .ZN(n6114) );
  NAND2_X1 U7736 ( .A1(n6137), .A2(n6114), .ZN(n9461) );
  OR2_X1 U7737 ( .A1(n4484), .A2(n9461), .ZN(n6117) );
  INV_X1 U7738 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n6115) );
  OR2_X1 U7739 ( .A1(n8076), .A2(n6115), .ZN(n6116) );
  NAND4_X1 U7740 ( .A1(n6119), .A2(n6118), .A3(n6117), .A4(n6116), .ZN(n9223)
         );
  NAND2_X1 U7741 ( .A1(n9223), .A2(n6332), .ZN(n6120) );
  NAND2_X1 U7742 ( .A1(n6121), .A2(n6120), .ZN(n6122) );
  XNOR2_X1 U7743 ( .A(n6122), .B(n7437), .ZN(n6124) );
  NOR2_X1 U7744 ( .A1(n9478), .A2(n5882), .ZN(n6123) );
  AOI21_X1 U7745 ( .B1(n9581), .B2(n6309), .A(n6123), .ZN(n6125) );
  XNOR2_X1 U7746 ( .A(n6124), .B(n6125), .ZN(n9091) );
  INV_X1 U7747 ( .A(n6124), .ZN(n6126) );
  NAND2_X1 U7748 ( .A1(n6126), .A2(n6125), .ZN(n6127) );
  NAND2_X1 U7749 ( .A1(n7247), .A2(n8072), .ZN(n6133) );
  NAND2_X1 U7750 ( .A1(n6129), .A2(n6128), .ZN(n6130) );
  NAND2_X1 U7751 ( .A1(n6130), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6131) );
  XNOR2_X1 U7752 ( .A(n6131), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U7753 ( .A1(n6265), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6629), .B2(
        n10252), .ZN(n6132) );
  NAND2_X1 U7754 ( .A1(n9578), .A2(n6317), .ZN(n6144) );
  NAND2_X1 U7755 ( .A1(n6195), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6142) );
  INV_X1 U7756 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9192) );
  OR2_X1 U7757 ( .A1(n6376), .A2(n9192), .ZN(n6141) );
  INV_X1 U7758 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7759 ( .A1(n6137), .A2(n6136), .ZN(n6138) );
  NAND2_X1 U7760 ( .A1(n6156), .A2(n6138), .ZN(n9446) );
  OR2_X1 U7761 ( .A1(n4485), .A2(n9446), .ZN(n6140) );
  INV_X1 U7762 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9447) );
  OR2_X1 U7763 ( .A1(n8076), .A2(n9447), .ZN(n6139) );
  OR2_X1 U7764 ( .A1(n9437), .A2(n5852), .ZN(n6143) );
  NAND2_X1 U7765 ( .A1(n6144), .A2(n6143), .ZN(n6145) );
  XNOR2_X1 U7766 ( .A(n6145), .B(n7437), .ZN(n6148) );
  NOR2_X1 U7767 ( .A1(n9437), .A2(n5882), .ZN(n6146) );
  AOI21_X1 U7768 ( .B1(n9578), .B2(n6309), .A(n6146), .ZN(n9128) );
  NAND2_X1 U7769 ( .A1(n9127), .A2(n9128), .ZN(n6151) );
  INV_X1 U7770 ( .A(n6147), .ZN(n6150) );
  INV_X1 U7771 ( .A(n6148), .ZN(n6149) );
  NAND2_X1 U7772 ( .A1(n6150), .A2(n6149), .ZN(n9126) );
  NAND2_X1 U7773 ( .A1(n7320), .A2(n8072), .ZN(n6153) );
  AOI22_X1 U7774 ( .A1(n6265), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9200), .B2(
        n6629), .ZN(n6152) );
  NAND2_X1 U7775 ( .A1(n9573), .A2(n6317), .ZN(n6164) );
  NAND2_X1 U7776 ( .A1(n6195), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6162) );
  INV_X1 U7777 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9431) );
  OR2_X1 U7778 ( .A1(n8076), .A2(n9431), .ZN(n6161) );
  INV_X1 U7779 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7780 ( .A1(n6156), .A2(n6155), .ZN(n6157) );
  NAND2_X1 U7781 ( .A1(n6176), .A2(n6157), .ZN(n9430) );
  OR2_X1 U7782 ( .A1(n9430), .A2(n4484), .ZN(n6160) );
  INV_X1 U7783 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n6158) );
  OR2_X1 U7784 ( .A1(n6376), .A2(n6158), .ZN(n6159) );
  NAND4_X1 U7785 ( .A1(n6162), .A2(n6161), .A3(n6160), .A4(n6159), .ZN(n9421)
         );
  NAND2_X1 U7786 ( .A1(n9421), .A2(n6309), .ZN(n6163) );
  NAND2_X1 U7787 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  XNOR2_X1 U7788 ( .A(n6165), .B(n7437), .ZN(n6168) );
  NAND2_X1 U7789 ( .A1(n9573), .A2(n6309), .ZN(n6167) );
  NAND2_X1 U7790 ( .A1(n6308), .A2(n9421), .ZN(n6166) );
  NAND2_X1 U7791 ( .A1(n6167), .A2(n6166), .ZN(n6169) );
  NAND2_X1 U7792 ( .A1(n6168), .A2(n6169), .ZN(n9046) );
  INV_X1 U7793 ( .A(n6168), .ZN(n6171) );
  INV_X1 U7794 ( .A(n6169), .ZN(n6170) );
  NAND2_X1 U7795 ( .A1(n6171), .A2(n6170), .ZN(n9045) );
  NAND2_X1 U7796 ( .A1(n7494), .A2(n8072), .ZN(n6173) );
  NAND2_X1 U7797 ( .A1(n6265), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7798 ( .A1(n9566), .A2(n6317), .ZN(n6182) );
  INV_X1 U7799 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7800 ( .A1(n6196), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7801 ( .A1(n6195), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6174) );
  AND2_X1 U7802 ( .A1(n6175), .A2(n6174), .ZN(n6179) );
  INV_X1 U7803 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9111) );
  NAND2_X1 U7804 ( .A1(n6176), .A2(n9111), .ZN(n6177) );
  NAND2_X1 U7805 ( .A1(n6193), .A2(n6177), .ZN(n9415) );
  OR2_X1 U7806 ( .A1(n9415), .A2(n4485), .ZN(n6178) );
  OAI211_X1 U7807 ( .C1(n8076), .C2(n6180), .A(n6179), .B(n6178), .ZN(n9226)
         );
  NAND2_X1 U7808 ( .A1(n9226), .A2(n6309), .ZN(n6181) );
  NAND2_X1 U7809 ( .A1(n6182), .A2(n6181), .ZN(n6183) );
  XNOR2_X1 U7810 ( .A(n6183), .B(n7437), .ZN(n6186) );
  NAND2_X1 U7811 ( .A1(n9566), .A2(n6309), .ZN(n6185) );
  NAND2_X1 U7812 ( .A1(n6308), .A2(n9226), .ZN(n6184) );
  NAND2_X1 U7813 ( .A1(n6185), .A2(n6184), .ZN(n6187) );
  NAND2_X1 U7814 ( .A1(n6186), .A2(n6187), .ZN(n9108) );
  INV_X1 U7815 ( .A(n6186), .ZN(n6189) );
  INV_X1 U7816 ( .A(n6187), .ZN(n6188) );
  NAND2_X1 U7817 ( .A1(n6189), .A2(n6188), .ZN(n9109) );
  NAND2_X1 U7818 ( .A1(n7525), .A2(n8072), .ZN(n6191) );
  NAND2_X1 U7819 ( .A1(n6265), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7820 ( .A1(n9563), .A2(n6317), .ZN(n6201) );
  INV_X1 U7821 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7822 ( .A1(n6193), .A2(n6192), .ZN(n6194) );
  AND2_X1 U7823 ( .A1(n6211), .A2(n6194), .ZN(n9406) );
  NAND2_X1 U7824 ( .A1(n9406), .A2(n6299), .ZN(n6199) );
  AOI22_X1 U7825 ( .A1(n6372), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n6195), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7826 ( .A1(n6196), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6197) );
  INV_X1 U7827 ( .A(n9377), .ZN(n9422) );
  NAND2_X1 U7828 ( .A1(n9422), .A2(n6332), .ZN(n6200) );
  NAND2_X1 U7829 ( .A1(n6201), .A2(n6200), .ZN(n6202) );
  XNOR2_X1 U7830 ( .A(n6202), .B(n7437), .ZN(n6204) );
  NOR2_X1 U7831 ( .A1(n9377), .A2(n5882), .ZN(n6203) );
  AOI21_X1 U7832 ( .B1(n9563), .B2(n6309), .A(n6203), .ZN(n6205) );
  XNOR2_X1 U7833 ( .A(n6204), .B(n6205), .ZN(n9054) );
  INV_X1 U7834 ( .A(n6204), .ZN(n6206) );
  NAND2_X1 U7835 ( .A1(n6206), .A2(n6205), .ZN(n6224) );
  NAND2_X1 U7836 ( .A1(n7660), .A2(n8072), .ZN(n6208) );
  NAND2_X1 U7837 ( .A1(n6265), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6207) );
  OR2_X1 U7838 ( .A1(n9230), .A2(n5852), .ZN(n6220) );
  INV_X1 U7839 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7840 ( .A1(n6211), .A2(n6210), .ZN(n6212) );
  NAND2_X1 U7841 ( .A1(n6231), .A2(n6212), .ZN(n9383) );
  OR2_X1 U7842 ( .A1(n9383), .A2(n4484), .ZN(n6218) );
  INV_X1 U7843 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U7844 ( .A1(n6372), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U7845 ( .A1(n6195), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6213) );
  OAI211_X1 U7846 ( .C1(n6376), .C2(n6215), .A(n6214), .B(n6213), .ZN(n6216)
         );
  INV_X1 U7847 ( .A(n6216), .ZN(n6217) );
  NAND2_X1 U7848 ( .A1(n9366), .A2(n6308), .ZN(n6219) );
  INV_X1 U7849 ( .A(n6226), .ZN(n6221) );
  AND2_X1 U7850 ( .A1(n6224), .A2(n6221), .ZN(n6222) );
  OAI22_X1 U7851 ( .A1(n9230), .A2(n6306), .B1(n9402), .B2(n5852), .ZN(n6223)
         );
  XNOR2_X1 U7852 ( .A(n6223), .B(n6254), .ZN(n9119) );
  NAND2_X1 U7853 ( .A1(n7680), .A2(n8072), .ZN(n6228) );
  NAND2_X1 U7854 ( .A1(n6265), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6227) );
  NAND2_X1 U7855 ( .A1(n9550), .A2(n6317), .ZN(n6240) );
  INV_X1 U7856 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U7857 ( .A1(n6231), .A2(n6230), .ZN(n6232) );
  NAND2_X1 U7858 ( .A1(n6246), .A2(n6232), .ZN(n9039) );
  OR2_X1 U7859 ( .A1(n9039), .A2(n4485), .ZN(n6238) );
  INV_X1 U7860 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6235) );
  NAND2_X1 U7861 ( .A1(n6195), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U7862 ( .A1(n6372), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6233) );
  OAI211_X1 U7863 ( .C1(n6376), .C2(n6235), .A(n6234), .B(n6233), .ZN(n6236)
         );
  INV_X1 U7864 ( .A(n6236), .ZN(n6237) );
  NAND2_X1 U7865 ( .A1(n6238), .A2(n6237), .ZN(n9375) );
  NAND2_X1 U7866 ( .A1(n9375), .A2(n6332), .ZN(n6239) );
  NAND2_X1 U7867 ( .A1(n6240), .A2(n6239), .ZN(n6241) );
  XNOR2_X1 U7868 ( .A(n6241), .B(n7437), .ZN(n6243) );
  AND2_X1 U7869 ( .A1(n9375), .A2(n6308), .ZN(n6242) );
  AOI21_X1 U7870 ( .B1(n9550), .B2(n6309), .A(n6242), .ZN(n9035) );
  NAND2_X1 U7871 ( .A1(n7789), .A2(n8072), .ZN(n6245) );
  NAND2_X1 U7872 ( .A1(n6265), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6244) );
  INV_X1 U7873 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9102) );
  NAND2_X1 U7874 ( .A1(n6246), .A2(n9102), .ZN(n6247) );
  AND2_X1 U7875 ( .A1(n6269), .A2(n6247), .ZN(n9353) );
  NAND2_X1 U7876 ( .A1(n9353), .A2(n6299), .ZN(n6253) );
  INV_X1 U7877 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U7878 ( .A1(n6372), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U7879 ( .A1(n6195), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6248) );
  OAI211_X1 U7880 ( .C1(n6376), .C2(n6250), .A(n6249), .B(n6248), .ZN(n6251)
         );
  INV_X1 U7881 ( .A(n6251), .ZN(n6252) );
  OAI22_X1 U7882 ( .A1(n9356), .A2(n6306), .B1(n9234), .B2(n5852), .ZN(n6255)
         );
  XNOR2_X1 U7883 ( .A(n6255), .B(n6254), .ZN(n6258) );
  OR2_X1 U7884 ( .A1(n9356), .A2(n5852), .ZN(n6257) );
  INV_X1 U7885 ( .A(n9234), .ZN(n9367) );
  NAND2_X1 U7886 ( .A1(n9367), .A2(n6308), .ZN(n6256) );
  NAND2_X1 U7887 ( .A1(n6258), .A2(n6259), .ZN(n6263) );
  INV_X1 U7888 ( .A(n6258), .ZN(n6261) );
  INV_X1 U7889 ( .A(n6259), .ZN(n6260) );
  NAND2_X1 U7890 ( .A1(n6261), .A2(n6260), .ZN(n6262) );
  NAND2_X1 U7891 ( .A1(n6263), .A2(n6262), .ZN(n9097) );
  INV_X1 U7892 ( .A(n6263), .ZN(n6264) );
  NAND2_X1 U7893 ( .A1(n7824), .A2(n8072), .ZN(n6267) );
  NAND2_X1 U7894 ( .A1(n6265), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6266) );
  INV_X1 U7895 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9062) );
  NAND2_X1 U7896 ( .A1(n6269), .A2(n9062), .ZN(n6270) );
  NAND2_X1 U7897 ( .A1(n6285), .A2(n6270), .ZN(n9333) );
  OR2_X1 U7898 ( .A1(n9333), .A2(n4484), .ZN(n6276) );
  INV_X1 U7899 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7900 ( .A1(n6195), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7901 ( .A1(n6372), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6271) );
  OAI211_X1 U7902 ( .C1(n6273), .C2(n6376), .A(n6272), .B(n6271), .ZN(n6274)
         );
  INV_X1 U7903 ( .A(n6274), .ZN(n6275) );
  AOI22_X1 U7904 ( .A1(n9540), .A2(n6309), .B1(n6308), .B2(n9316), .ZN(n6280)
         );
  NAND2_X1 U7905 ( .A1(n9540), .A2(n6317), .ZN(n6278) );
  NAND2_X1 U7906 ( .A1(n9316), .A2(n6309), .ZN(n6277) );
  NAND2_X1 U7907 ( .A1(n6278), .A2(n6277), .ZN(n6279) );
  XNOR2_X1 U7908 ( .A(n6279), .B(n7437), .ZN(n6282) );
  XOR2_X1 U7909 ( .A(n6280), .B(n6282), .Z(n9061) );
  INV_X1 U7910 ( .A(n6280), .ZN(n6281) );
  NOR2_X1 U7911 ( .A1(n6282), .A2(n6281), .ZN(n9136) );
  NAND2_X1 U7912 ( .A1(n6265), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6283) );
  INV_X1 U7913 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9140) );
  NAND2_X1 U7914 ( .A1(n6285), .A2(n9140), .ZN(n6286) );
  NAND2_X1 U7915 ( .A1(n9321), .A2(n6299), .ZN(n6292) );
  INV_X1 U7916 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U7917 ( .A1(n6195), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7918 ( .A1(n6372), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6287) );
  OAI211_X1 U7919 ( .C1(n6289), .C2(n6376), .A(n6288), .B(n6287), .ZN(n6290)
         );
  INV_X1 U7920 ( .A(n6290), .ZN(n6291) );
  AND2_X1 U7921 ( .A1(n9339), .A2(n6308), .ZN(n6293) );
  AOI21_X1 U7922 ( .B1(n9536), .B2(n6309), .A(n6293), .ZN(n6312) );
  NAND2_X1 U7923 ( .A1(n9536), .A2(n6317), .ZN(n6295) );
  NAND2_X1 U7924 ( .A1(n9339), .A2(n6309), .ZN(n6294) );
  NAND2_X1 U7925 ( .A1(n6295), .A2(n6294), .ZN(n6296) );
  XNOR2_X1 U7926 ( .A(n6296), .B(n7437), .ZN(n6314) );
  XOR2_X1 U7927 ( .A(n6312), .B(n6314), .Z(n9135) );
  NAND2_X1 U7928 ( .A1(n7927), .A2(n8072), .ZN(n6298) );
  NAND2_X1 U7929 ( .A1(n5873), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6297) );
  XNOR2_X1 U7930 ( .A(n6319), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9302) );
  NAND2_X1 U7931 ( .A1(n9302), .A2(n6299), .ZN(n6305) );
  INV_X1 U7932 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7933 ( .A1(n6372), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7934 ( .A1(n6195), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6300) );
  OAI211_X1 U7935 ( .C1(n6376), .C2(n6302), .A(n6301), .B(n6300), .ZN(n6303)
         );
  INV_X1 U7936 ( .A(n6303), .ZN(n6304) );
  OAI22_X1 U7937 ( .A1(n9304), .A2(n6306), .B1(n9239), .B2(n5852), .ZN(n6307)
         );
  XOR2_X1 U7938 ( .A(n7437), .B(n6307), .Z(n6311) );
  AOI22_X1 U7939 ( .A1(n9531), .A2(n6309), .B1(n6308), .B2(n9317), .ZN(n6310)
         );
  NAND2_X1 U7940 ( .A1(n6311), .A2(n6310), .ZN(n6383) );
  OAI21_X1 U7941 ( .B1(n6311), .B2(n6310), .A(n6383), .ZN(n6583) );
  INV_X1 U7942 ( .A(n6312), .ZN(n6313) );
  NAND2_X1 U7943 ( .A1(n7931), .A2(n8072), .ZN(n6316) );
  NAND2_X1 U7944 ( .A1(n6265), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U7945 ( .A1(n9284), .A2(n6317), .ZN(n6330) );
  INV_X1 U7946 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6587) );
  INV_X1 U7947 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6318) );
  OAI21_X1 U7948 ( .B1(n6319), .B2(n6587), .A(n6318), .ZN(n6322) );
  INV_X1 U7949 ( .A(n6319), .ZN(n6321) );
  AND2_X1 U7950 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6320) );
  NAND2_X1 U7951 ( .A1(n6321), .A2(n6320), .ZN(n9273) );
  NAND2_X1 U7952 ( .A1(n6322), .A2(n9273), .ZN(n6366) );
  OR2_X1 U7953 ( .A1(n6366), .A2(n4485), .ZN(n6328) );
  INV_X1 U7954 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U7955 ( .A1(n6195), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U7956 ( .A1(n6372), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6323) );
  OAI211_X1 U7957 ( .C1(n6376), .C2(n6325), .A(n6324), .B(n6323), .ZN(n6326)
         );
  INV_X1 U7958 ( .A(n6326), .ZN(n6327) );
  NAND2_X1 U7959 ( .A1(n9307), .A2(n6309), .ZN(n6329) );
  NAND2_X1 U7960 ( .A1(n6330), .A2(n6329), .ZN(n6331) );
  XNOR2_X1 U7961 ( .A(n6331), .B(n7437), .ZN(n6334) );
  AOI22_X1 U7962 ( .A1(n9284), .A2(n6332), .B1(n6308), .B2(n9307), .ZN(n6333)
         );
  XNOR2_X1 U7963 ( .A(n6334), .B(n6333), .ZN(n6359) );
  INV_X1 U7964 ( .A(n6359), .ZN(n6384) );
  NAND2_X1 U7965 ( .A1(n5786), .A2(n8253), .ZN(n7329) );
  NAND2_X1 U7966 ( .A1(n6336), .A2(n6337), .ZN(n8204) );
  AND2_X1 U7967 ( .A1(n10323), .A2(n8204), .ZN(n6357) );
  NAND2_X1 U7968 ( .A1(n7823), .A2(P1_B_REG_SCAN_IN), .ZN(n6338) );
  OAI22_X1 U7969 ( .A1(n7825), .A2(n6338), .B1(P1_B_REG_SCAN_IN), .B2(n7823), 
        .ZN(n6340) );
  OAI22_X1 U7970 ( .A1(n10287), .A2(P1_D_REG_0__SCAN_IN), .B1(n6353), .B2(
        n6341), .ZN(n6904) );
  NOR2_X1 U7971 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .ZN(
        n6345) );
  NOR4_X1 U7972 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6344) );
  NOR4_X1 U7973 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6343) );
  NOR4_X1 U7974 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6342) );
  NAND4_X1 U7975 ( .A1(n6345), .A2(n6344), .A3(n6343), .A4(n6342), .ZN(n6351)
         );
  NOR4_X1 U7976 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6349) );
  NOR4_X1 U7977 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6348) );
  NOR4_X1 U7978 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6347) );
  NOR4_X1 U7979 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6346) );
  NAND4_X1 U7980 ( .A1(n6349), .A2(n6348), .A3(n6347), .A4(n6346), .ZN(n6350)
         );
  NOR2_X1 U7981 ( .A1(n6351), .A2(n6350), .ZN(n6352) );
  NOR2_X1 U7982 ( .A1(n10287), .A2(n6352), .ZN(n6903) );
  OR2_X1 U7983 ( .A1(n6904), .A2(n6903), .ZN(n7078) );
  OAI22_X1 U7984 ( .A1(n10287), .A2(P1_D_REG_1__SCAN_IN), .B1(n6353), .B2(
        n7825), .ZN(n7323) );
  OR2_X1 U7985 ( .A1(n7078), .A2(n7323), .ZN(n6938) );
  NAND2_X1 U7986 ( .A1(n6354), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6355) );
  XNOR2_X1 U7987 ( .A(n6355), .B(n4765), .ZN(n7681) );
  AND2_X1 U7988 ( .A1(n7681), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6356) );
  INV_X1 U7989 ( .A(n10288), .ZN(n6700) );
  NOR2_X1 U7990 ( .A1(n6938), .A2(n6700), .ZN(n6364) );
  NAND3_X1 U7991 ( .A1(n6384), .A2(n10101), .A3(n6383), .ZN(n6358) );
  NAND3_X1 U7992 ( .A1(n6586), .A2(n6359), .A3(n10101), .ZN(n6388) );
  NAND2_X1 U7993 ( .A1(n6367), .A2(n10288), .ZN(n7326) );
  INV_X1 U7994 ( .A(n7326), .ZN(n6362) );
  OR2_X1 U7995 ( .A1(n7329), .A2(n8244), .ZN(n7331) );
  INV_X1 U7996 ( .A(n7331), .ZN(n6361) );
  AND2_X1 U7997 ( .A1(n6938), .A2(n10288), .ZN(n6360) );
  NAND2_X1 U7998 ( .A1(n6361), .A2(n6360), .ZN(n6370) );
  INV_X1 U7999 ( .A(n9284), .ZN(n9287) );
  NOR2_X1 U8000 ( .A1(n9287), .A2(n10323), .ZN(n9525) );
  OR2_X1 U8001 ( .A1(n7058), .A2(n5763), .ZN(n8197) );
  INV_X1 U8002 ( .A(n8197), .ZN(n6363) );
  NAND2_X1 U8003 ( .A1(n6364), .A2(n6363), .ZN(n6380) );
  INV_X1 U8004 ( .A(n6366), .ZN(n9285) );
  NAND2_X1 U8005 ( .A1(n6938), .A2(n10323), .ZN(n6368) );
  NAND4_X1 U8006 ( .A1(n6368), .A2(n6598), .A3(n7681), .A4(n6367), .ZN(n6369)
         );
  NAND2_X1 U8007 ( .A1(n6369), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6371) );
  INV_X1 U8008 ( .A(n10106), .ZN(n9143) );
  AOI22_X1 U8009 ( .A1(n9285), .A2(n9143), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6382) );
  OR2_X1 U8010 ( .A1(n9273), .A2(n4484), .ZN(n6379) );
  INV_X1 U8011 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6375) );
  NAND2_X1 U8012 ( .A1(n6372), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U8013 ( .A1(n6195), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6373) );
  OAI211_X1 U8014 ( .C1(n6376), .C2(n6375), .A(n6374), .B(n6373), .ZN(n6377)
         );
  INV_X1 U8015 ( .A(n6377), .ZN(n6378) );
  NAND2_X1 U8016 ( .A1(n6379), .A2(n6378), .ZN(n9294) );
  NAND2_X1 U8017 ( .A1(n9294), .A2(n9152), .ZN(n6381) );
  OAI211_X1 U8018 ( .C1(n9239), .C2(n10061), .A(n6382), .B(n6381), .ZN(n6386)
         );
  NOR3_X1 U8019 ( .A1(n6384), .A2(n6383), .A3(n9156), .ZN(n6385) );
  AOI211_X1 U8020 ( .C1(n10067), .C2(n9525), .A(n6386), .B(n6385), .ZN(n6387)
         );
  NAND3_X1 U8021 ( .A1(n6389), .A2(n6388), .A3(n6387), .ZN(P1_U3218) );
  NAND3_X1 U8022 ( .A1(n8384), .A2(n8385), .A3(n8355), .ZN(n6390) );
  NAND2_X2 U8023 ( .A1(n6390), .A2(n7189), .ZN(n6513) );
  XNOR2_X1 U8024 ( .A(n6391), .B(n6513), .ZN(n6393) );
  INV_X1 U8025 ( .A(n6393), .ZN(n6394) );
  NAND2_X1 U8026 ( .A1(n6395), .A2(n6394), .ZN(n6398) );
  NAND2_X1 U8027 ( .A1(n8579), .A2(n10436), .ZN(n6397) );
  INV_X1 U8028 ( .A(n10408), .ZN(n10361) );
  MUX2_X1 U8029 ( .A(n6397), .B(n6513), .S(n10361), .Z(n7112) );
  NAND2_X1 U8030 ( .A1(n7111), .A2(n6398), .ZN(n7137) );
  OR2_X1 U8031 ( .A1(n6399), .A2(n8951), .ZN(n6400) );
  XNOR2_X1 U8032 ( .A(n7231), .B(n6488), .ZN(n6401) );
  XNOR2_X1 U8033 ( .A(n6400), .B(n6401), .ZN(n7138) );
  OR2_X1 U8034 ( .A1(n7198), .A2(n8951), .ZN(n6402) );
  XNOR2_X1 U8035 ( .A(n7351), .B(n6513), .ZN(n6403) );
  XNOR2_X1 U8036 ( .A(n6402), .B(n6403), .ZN(n7147) );
  INV_X1 U8037 ( .A(n6402), .ZN(n6404) );
  NAND2_X1 U8038 ( .A1(n6404), .A2(n6403), .ZN(n6405) );
  OR2_X1 U8039 ( .A1(n7407), .A2(n8951), .ZN(n6407) );
  XNOR2_X1 U8040 ( .A(n7362), .B(n6488), .ZN(n6406) );
  NAND2_X1 U8041 ( .A1(n6407), .A2(n6406), .ZN(n6409) );
  OAI21_X1 U8042 ( .B1(n6407), .B2(n6406), .A(n6409), .ZN(n7175) );
  NAND2_X1 U8043 ( .A1(n7173), .A2(n6409), .ZN(n7209) );
  OR2_X1 U8044 ( .A1(n7489), .A2(n8951), .ZN(n6410) );
  XNOR2_X1 U8045 ( .A(n7576), .B(n6488), .ZN(n6411) );
  XNOR2_X1 U8046 ( .A(n6410), .B(n6411), .ZN(n7208) );
  INV_X1 U8047 ( .A(n6410), .ZN(n6413) );
  INV_X1 U8048 ( .A(n6411), .ZN(n6412) );
  NOR2_X1 U8049 ( .A1(n7423), .A2(n8951), .ZN(n6415) );
  XNOR2_X1 U8050 ( .A(n7603), .B(n6513), .ZN(n6416) );
  NAND2_X1 U8051 ( .A1(n6415), .A2(n6416), .ZN(n6419) );
  INV_X1 U8052 ( .A(n6415), .ZN(n6418) );
  INV_X1 U8053 ( .A(n6416), .ZN(n6417) );
  NAND2_X1 U8054 ( .A1(n6418), .A2(n6417), .ZN(n7419) );
  AND2_X1 U8055 ( .A1(n6419), .A2(n7419), .ZN(n7485) );
  INV_X1 U8056 ( .A(n6424), .ZN(n6421) );
  XNOR2_X1 U8057 ( .A(n4482), .B(n6488), .ZN(n6423) );
  INV_X1 U8058 ( .A(n6423), .ZN(n6420) );
  NAND2_X1 U8059 ( .A1(n6421), .A2(n6420), .ZN(n6422) );
  XNOR2_X1 U8060 ( .A(n6424), .B(n6423), .ZN(n7420) );
  OR2_X1 U8061 ( .A1(n7613), .A2(n8951), .ZN(n6427) );
  XNOR2_X1 U8062 ( .A(n7631), .B(n6513), .ZN(n6425) );
  XNOR2_X1 U8063 ( .A(n6427), .B(n6425), .ZN(n7499) );
  INV_X1 U8064 ( .A(n6425), .ZN(n6426) );
  NOR2_X1 U8065 ( .A1(n7742), .A2(n8951), .ZN(n6428) );
  XNOR2_X1 U8066 ( .A(n7675), .B(n6513), .ZN(n6429) );
  NAND2_X1 U8067 ( .A1(n6428), .A2(n6429), .ZN(n6432) );
  INV_X1 U8068 ( .A(n6428), .ZN(n6431) );
  INV_X1 U8069 ( .A(n6429), .ZN(n6430) );
  NAND2_X1 U8070 ( .A1(n6431), .A2(n6430), .ZN(n6433) );
  AND2_X1 U8071 ( .A1(n6432), .A2(n6433), .ZN(n7611) );
  XNOR2_X1 U8072 ( .A(n7748), .B(n6513), .ZN(n6434) );
  NAND2_X1 U8073 ( .A1(n8568), .A2(n10436), .ZN(n6435) );
  XNOR2_X1 U8074 ( .A(n6434), .B(n6435), .ZN(n6613) );
  INV_X1 U8075 ( .A(n6434), .ZN(n6437) );
  INV_X1 U8076 ( .A(n6435), .ZN(n6436) );
  NAND2_X1 U8077 ( .A1(n6437), .A2(n6436), .ZN(n6438) );
  XNOR2_X1 U8078 ( .A(n7766), .B(n6488), .ZN(n6439) );
  NOR2_X1 U8079 ( .A1(n7793), .A2(n8951), .ZN(n6440) );
  XNOR2_X1 U8080 ( .A(n6439), .B(n6440), .ZN(n6621) );
  INV_X1 U8081 ( .A(n6439), .ZN(n6441) );
  NAND2_X1 U8082 ( .A1(n6441), .A2(n6440), .ZN(n6442) );
  XNOR2_X1 U8083 ( .A(n7805), .B(n6488), .ZN(n6443) );
  NOR2_X1 U8084 ( .A1(n7878), .A2(n8951), .ZN(n6444) );
  XNOR2_X1 U8085 ( .A(n6443), .B(n6444), .ZN(n6600) );
  INV_X1 U8086 ( .A(n6443), .ZN(n6445) );
  XNOR2_X1 U8087 ( .A(n10079), .B(n6488), .ZN(n6446) );
  NOR2_X1 U8088 ( .A1(n8893), .A2(n8951), .ZN(n6447) );
  XNOR2_X1 U8089 ( .A(n6446), .B(n6447), .ZN(n6607) );
  NAND2_X1 U8090 ( .A1(n6606), .A2(n6607), .ZN(n6450) );
  INV_X1 U8091 ( .A(n6446), .ZN(n6448) );
  NAND2_X1 U8092 ( .A1(n6448), .A2(n6447), .ZN(n6449) );
  XNOR2_X1 U8093 ( .A(n8886), .B(n6488), .ZN(n6451) );
  OR2_X1 U8094 ( .A1(n8860), .A2(n8951), .ZN(n6452) );
  NAND2_X1 U8095 ( .A1(n6451), .A2(n6452), .ZN(n6457) );
  INV_X1 U8096 ( .A(n6451), .ZN(n6454) );
  INV_X1 U8097 ( .A(n6452), .ZN(n6453) );
  NAND2_X1 U8098 ( .A1(n6454), .A2(n6453), .ZN(n6455) );
  NAND2_X1 U8099 ( .A1(n6457), .A2(n6455), .ZN(n7848) );
  XNOR2_X1 U8100 ( .A(n8967), .B(n6488), .ZN(n6459) );
  INV_X1 U8101 ( .A(n6459), .ZN(n6458) );
  OR2_X1 U8102 ( .A1(n8891), .A2(n8951), .ZN(n8338) );
  NAND2_X1 U8103 ( .A1(n6460), .A2(n6459), .ZN(n8336) );
  XNOR2_X1 U8104 ( .A(n8850), .B(n6488), .ZN(n6462) );
  OR2_X1 U8105 ( .A1(n8859), .A2(n8951), .ZN(n6463) );
  NAND2_X1 U8106 ( .A1(n6462), .A2(n6463), .ZN(n6467) );
  INV_X1 U8107 ( .A(n6462), .ZN(n6465) );
  INV_X1 U8108 ( .A(n6463), .ZN(n6464) );
  NAND2_X1 U8109 ( .A1(n6465), .A2(n6464), .ZN(n6466) );
  AND2_X1 U8110 ( .A1(n6467), .A2(n6466), .ZN(n8294) );
  XNOR2_X1 U8111 ( .A(n8825), .B(n6513), .ZN(n6469) );
  NOR2_X1 U8112 ( .A1(n8842), .A2(n8951), .ZN(n6468) );
  XNOR2_X1 U8113 ( .A(n6469), .B(n6468), .ZN(n8302) );
  XNOR2_X1 U8114 ( .A(n8950), .B(n6513), .ZN(n6472) );
  NAND2_X1 U8115 ( .A1(n8814), .A2(n10436), .ZN(n6470) );
  XNOR2_X1 U8116 ( .A(n6472), .B(n6470), .ZN(n7967) );
  INV_X1 U8117 ( .A(n6470), .ZN(n6471) );
  AND2_X1 U8118 ( .A1(n6472), .A2(n6471), .ZN(n6473) );
  XNOR2_X1 U8119 ( .A(n8946), .B(n6488), .ZN(n6474) );
  NAND2_X1 U8120 ( .A1(n8804), .A2(n10436), .ZN(n6475) );
  NAND2_X1 U8121 ( .A1(n6474), .A2(n6475), .ZN(n6479) );
  INV_X1 U8122 ( .A(n6474), .ZN(n6477) );
  INV_X1 U8123 ( .A(n6475), .ZN(n6476) );
  NAND2_X1 U8124 ( .A1(n6477), .A2(n6476), .ZN(n6478) );
  NAND2_X1 U8125 ( .A1(n8265), .A2(n8264), .ZN(n8263) );
  NAND2_X1 U8126 ( .A1(n8263), .A2(n6479), .ZN(n8320) );
  XNOR2_X1 U8127 ( .A(n8940), .B(n6513), .ZN(n6481) );
  NOR2_X1 U8128 ( .A1(n8275), .A2(n8951), .ZN(n6480) );
  XNOR2_X1 U8129 ( .A(n6481), .B(n6480), .ZN(n8319) );
  NAND2_X1 U8130 ( .A1(n6481), .A2(n6480), .ZN(n8271) );
  XNOR2_X1 U8131 ( .A(n8935), .B(n6513), .ZN(n6485) );
  NAND2_X1 U8132 ( .A1(n8772), .A2(n10436), .ZN(n6484) );
  INV_X1 U8133 ( .A(n6484), .ZN(n6482) );
  NAND2_X1 U8134 ( .A1(n6485), .A2(n6482), .ZN(n6483) );
  AND2_X1 U8135 ( .A1(n8271), .A2(n6483), .ZN(n6487) );
  INV_X1 U8136 ( .A(n6483), .ZN(n6486) );
  XNOR2_X1 U8137 ( .A(n6485), .B(n6484), .ZN(n8272) );
  XNOR2_X1 U8138 ( .A(n8930), .B(n6488), .ZN(n6489) );
  XNOR2_X1 U8139 ( .A(n6491), .B(n6489), .ZN(n8328) );
  OR2_X1 U8140 ( .A1(n8274), .A2(n8951), .ZN(n8327) );
  NAND2_X1 U8141 ( .A1(n8328), .A2(n8327), .ZN(n8326) );
  INV_X1 U8142 ( .A(n6489), .ZN(n6490) );
  XNOR2_X1 U8143 ( .A(n8722), .B(n6513), .ZN(n6495) );
  INV_X1 U8144 ( .A(n6495), .ZN(n6493) );
  NOR2_X1 U8145 ( .A1(n6496), .A2(n6493), .ZN(n8309) );
  NOR2_X1 U8146 ( .A1(n8257), .A2(n8951), .ZN(n8311) );
  XNOR2_X1 U8147 ( .A(n6496), .B(n6495), .ZN(n8255) );
  NOR2_X1 U8148 ( .A1(n8738), .A2(n8951), .ZN(n8310) );
  NAND2_X1 U8149 ( .A1(n8255), .A2(n6498), .ZN(n6499) );
  NAND2_X1 U8150 ( .A1(n6500), .A2(n6499), .ZN(n8280) );
  XNOR2_X1 U8151 ( .A(n8999), .B(n6513), .ZN(n8282) );
  INV_X1 U8152 ( .A(n8282), .ZN(n6501) );
  NAND2_X1 U8153 ( .A1(n8280), .A2(n6501), .ZN(n6503) );
  NOR2_X1 U8154 ( .A1(n8702), .A2(n8951), .ZN(n8281) );
  INV_X1 U8155 ( .A(n8281), .ZN(n6502) );
  NAND2_X1 U8156 ( .A1(n6504), .A2(n8282), .ZN(n6505) );
  XNOR2_X1 U8157 ( .A(n8668), .B(n6513), .ZN(n6508) );
  NOR2_X1 U8158 ( .A1(n8284), .A2(n8951), .ZN(n6507) );
  NAND2_X1 U8159 ( .A1(n6508), .A2(n6507), .ZN(n6509) );
  OAI21_X1 U8160 ( .B1(n6508), .B2(n6507), .A(n6509), .ZN(n6548) );
  INV_X1 U8161 ( .A(n6509), .ZN(n6510) );
  XNOR2_X1 U8162 ( .A(n8388), .B(n6513), .ZN(n6512) );
  NOR2_X1 U8163 ( .A1(n8650), .A2(n8951), .ZN(n6511) );
  NAND2_X1 U8164 ( .A1(n6512), .A2(n6511), .ZN(n6522) );
  INV_X1 U8165 ( .A(n6521), .ZN(n6574) );
  NOR2_X1 U8166 ( .A1(n8524), .A2(n8951), .ZN(n6514) );
  XNOR2_X1 U8167 ( .A(n6514), .B(n6513), .ZN(n6515) );
  XNOR2_X1 U8168 ( .A(n8905), .B(n6515), .ZN(n6524) );
  INV_X1 U8169 ( .A(n6524), .ZN(n6520) );
  INV_X1 U8170 ( .A(n6516), .ZN(n7187) );
  NOR2_X1 U8171 ( .A1(n7185), .A2(n7182), .ZN(n6517) );
  NAND2_X1 U8172 ( .A1(n7187), .A2(n6517), .ZN(n6528) );
  NAND2_X1 U8173 ( .A1(n6695), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10404) );
  INV_X1 U8174 ( .A(n10404), .ZN(n6518) );
  NAND2_X1 U8175 ( .A1(n6791), .A2(n6518), .ZN(n10368) );
  NAND2_X1 U8176 ( .A1(n10434), .A2(n6696), .ZN(n6519) );
  NAND2_X1 U8177 ( .A1(n6574), .A2(n5054), .ZN(n6540) );
  NAND3_X1 U8178 ( .A1(n6521), .A2(n8329), .A3(n6524), .ZN(n6539) );
  INV_X1 U8179 ( .A(n6522), .ZN(n6523) );
  NAND3_X1 U8180 ( .A1(n6524), .A2(n6523), .A3(n8329), .ZN(n6538) );
  OR2_X1 U8181 ( .A1(n8385), .A2(n8366), .ZN(n7199) );
  OR2_X1 U8182 ( .A1(n10368), .A2(n7199), .ZN(n6525) );
  OR2_X1 U8183 ( .A1(n6528), .A2(n6525), .ZN(n6526) );
  NAND2_X1 U8184 ( .A1(n6528), .A2(n6527), .ZN(n6912) );
  INV_X1 U8185 ( .A(n6911), .ZN(n6529) );
  NAND2_X1 U8186 ( .A1(n6912), .A2(n6529), .ZN(n6530) );
  OAI22_X1 U8187 ( .A1(n8642), .A2(n8341), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6531), .ZN(n6536) );
  INV_X1 U8188 ( .A(n6532), .ZN(n6534) );
  NAND2_X1 U8189 ( .A1(n6534), .A2(n6533), .ZN(n6919) );
  OAI22_X1 U8190 ( .A1(n8650), .A2(n8343), .B1(n8649), .B2(n8342), .ZN(n6535)
         );
  AOI211_X1 U8191 ( .C1(n8905), .C2(n8346), .A(n6536), .B(n6535), .ZN(n6537)
         );
  NAND3_X1 U8192 ( .A1(n6540), .A2(n6539), .A3(n5049), .ZN(P2_U3222) );
  INV_X1 U8193 ( .A(n7182), .ZN(n6541) );
  NOR2_X1 U8194 ( .A1(n10452), .A2(n6543), .ZN(n6544) );
  NAND2_X1 U8195 ( .A1(n8668), .A2(n8346), .ZN(n6554) );
  OR2_X1 U8196 ( .A1(n8650), .A2(n8890), .ZN(n6550) );
  INV_X1 U8197 ( .A(n8702), .ZN(n8561) );
  NAND2_X1 U8198 ( .A1(n8561), .A2(n8816), .ZN(n6549) );
  AND2_X1 U8199 ( .A1(n6550), .A2(n6549), .ZN(n8664) );
  INV_X1 U8200 ( .A(n8341), .ZN(n8299) );
  AOI22_X1 U8201 ( .A1(n8299), .A2(n8669), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n6551) );
  OAI21_X1 U8202 ( .B1(n8664), .B2(n6919), .A(n6551), .ZN(n6552) );
  NAND2_X1 U8203 ( .A1(n8656), .A2(n8659), .ZN(n6557) );
  NAND2_X1 U8204 ( .A1(n6557), .A2(n6556), .ZN(n6558) );
  XNOR2_X1 U8205 ( .A(n6558), .B(n8379), .ZN(n7958) );
  NAND2_X1 U8206 ( .A1(n6559), .A2(n8379), .ZN(n6560) );
  NAND2_X1 U8207 ( .A1(n6560), .A2(n10357), .ZN(n6561) );
  OR2_X1 U8208 ( .A1(n4553), .A2(n6561), .ZN(n6563) );
  OAI22_X1 U8209 ( .A1(n8524), .A2(n8890), .B1(n8284), .B2(n8892), .ZN(n6577)
         );
  INV_X1 U8210 ( .A(n6577), .ZN(n6562) );
  NAND2_X1 U8211 ( .A1(n6563), .A2(n6562), .ZN(n7964) );
  AOI211_X1 U8212 ( .C1(n8388), .C2(n8666), .A(n10436), .B(n8640), .ZN(n7959)
         );
  AOI21_X1 U8213 ( .B1(n7958), .B2(n10440), .A(n6566), .ZN(n6594) );
  MUX2_X1 U8214 ( .A(n6567), .B(n6594), .S(n10444), .Z(n6570) );
  INV_X1 U8215 ( .A(n9019), .ZN(n6568) );
  NAND2_X1 U8216 ( .A1(n8388), .A2(n6568), .ZN(n6569) );
  NAND2_X1 U8217 ( .A1(n6570), .A2(n6569), .ZN(P2_U3515) );
  NAND2_X1 U8218 ( .A1(n6571), .A2(n6572), .ZN(n6573) );
  NAND3_X1 U8219 ( .A1(n6574), .A2(n6573), .A3(n8329), .ZN(n6581) );
  INV_X1 U8220 ( .A(n6919), .ZN(n8287) );
  INV_X1 U8221 ( .A(n7960), .ZN(n6575) );
  OAI22_X1 U8222 ( .A1(n6575), .A2(n8341), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9935), .ZN(n6576) );
  AOI21_X1 U8223 ( .B1(n6577), .B2(n8287), .A(n6576), .ZN(n6578) );
  INV_X1 U8224 ( .A(n6579), .ZN(n6580) );
  NAND2_X1 U8225 ( .A1(n6581), .A2(n6580), .ZN(P2_U3216) );
  INV_X1 U8226 ( .A(n6582), .ZN(n6585) );
  INV_X1 U8227 ( .A(n6583), .ZN(n6584) );
  NAND2_X1 U8228 ( .A1(n10067), .A2(n10164), .ZN(n9146) );
  INV_X1 U8229 ( .A(n9339), .ZN(n8093) );
  OAI22_X1 U8230 ( .A1(n8093), .A2(n10061), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6587), .ZN(n6589) );
  NOR2_X1 U8231 ( .A1(n9269), .A2(n10092), .ZN(n6588) );
  AOI211_X1 U8232 ( .C1(n9302), .C2(n9143), .A(n6589), .B(n6588), .ZN(n6590)
         );
  OAI21_X1 U8233 ( .B1(n9304), .B2(n9146), .A(n6590), .ZN(n6591) );
  INV_X1 U8234 ( .A(n6591), .ZN(n6592) );
  NAND2_X1 U8235 ( .A1(n6593), .A2(n6592), .ZN(P1_U3212) );
  INV_X1 U8236 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6595) );
  MUX2_X1 U8237 ( .A(n6595), .B(n6594), .S(n10452), .Z(n6597) );
  NAND2_X1 U8238 ( .A1(n8388), .A2(n7604), .ZN(n6596) );
  NAND2_X1 U8239 ( .A1(n6597), .A2(n6596), .ZN(P2_U3547) );
  INV_X1 U8240 ( .A(n7681), .ZN(n6627) );
  OR2_X2 U8241 ( .A1(n6655), .A2(P1_U3084), .ZN(n9159) );
  XNOR2_X1 U8242 ( .A(n6599), .B(n6600), .ZN(n6601) );
  NOR2_X1 U8243 ( .A1(n6601), .A2(n8348), .ZN(n6605) );
  AND2_X1 U8244 ( .A1(n7805), .A2(n8346), .ZN(n6604) );
  OAI22_X1 U8245 ( .A1(n8341), .A2(n7799), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9789), .ZN(n6603) );
  OAI22_X1 U8246 ( .A1(n7793), .A2(n8343), .B1(n8342), .B2(n8893), .ZN(n6602)
         );
  OR4_X1 U8247 ( .A1(n6605), .A2(n6604), .A3(n6603), .A4(n6602), .ZN(P2_U3226)
         );
  XNOR2_X1 U8248 ( .A(n6606), .B(n6607), .ZN(n6608) );
  NOR2_X1 U8249 ( .A1(n6608), .A2(n8348), .ZN(n6612) );
  AND2_X1 U8250 ( .A1(n10079), .A2(n8346), .ZN(n6611) );
  OAI22_X1 U8251 ( .A1(n8341), .A2(n7883), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7282), .ZN(n6610) );
  OAI22_X1 U8252 ( .A1(n7878), .A2(n8343), .B1(n8342), .B2(n8860), .ZN(n6609)
         );
  OR4_X1 U8253 ( .A1(n6612), .A2(n6611), .A3(n6610), .A4(n6609), .ZN(P2_U3236)
         );
  NOR2_X2 U8254 ( .A1(n6791), .A2(n10404), .ZN(P2_U3966) );
  XNOR2_X1 U8255 ( .A(n6614), .B(n6613), .ZN(n6615) );
  NOR2_X1 U8256 ( .A1(n6615), .A2(n8348), .ZN(n6619) );
  AND2_X1 U8257 ( .A1(n8346), .A2(n8981), .ZN(n6618) );
  OAI22_X1 U8258 ( .A1(n8341), .A2(n7749), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9977), .ZN(n6617) );
  OAI22_X1 U8259 ( .A1(n7742), .A2(n8343), .B1(n8342), .B2(n7793), .ZN(n6616)
         );
  OR4_X1 U8260 ( .A1(n6619), .A2(n6618), .A3(n6617), .A4(n6616), .ZN(P2_U3219)
         );
  XNOR2_X1 U8261 ( .A(n6620), .B(n6621), .ZN(n6622) );
  NOR2_X1 U8262 ( .A1(n6622), .A2(n8348), .ZN(n6626) );
  AND2_X1 U8263 ( .A1(n8346), .A2(n7766), .ZN(n6625) );
  OAI22_X1 U8264 ( .A1(n8341), .A2(n7763), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5342), .ZN(n6624) );
  OAI22_X1 U8265 ( .A1(n7761), .A2(n8343), .B1(n8342), .B2(n7878), .ZN(n6623)
         );
  OR4_X1 U8266 ( .A1(n6626), .A2(n6625), .A3(n6624), .A4(n6623), .ZN(P2_U3238)
         );
  OR2_X1 U8267 ( .A1(n8204), .A2(n6627), .ZN(n6628) );
  NAND2_X1 U8268 ( .A1(n6628), .A2(n6655), .ZN(n6650) );
  OR2_X1 U8269 ( .A1(n6650), .A2(n6629), .ZN(n6747) );
  NAND2_X1 U8270 ( .A1(n6747), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U8271 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7709) );
  INV_X1 U8272 ( .A(n6645), .ZN(n6924) );
  INV_X1 U8273 ( .A(n6954), .ZN(n6679) );
  INV_X1 U8274 ( .A(n6775), .ZN(n6666) );
  INV_X1 U8275 ( .A(n7020), .ZN(n6663) );
  XNOR2_X1 U8276 ( .A(n7007), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n7003) );
  NAND2_X1 U8277 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n7004) );
  NOR2_X1 U8278 ( .A1(n7003), .A2(n7004), .ZN(n7002) );
  AOI21_X1 U8279 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n7007), .A(n7002), .ZN(
        n7017) );
  XNOR2_X1 U8280 ( .A(n7020), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n7016) );
  INV_X1 U8281 ( .A(n7015), .ZN(n6630) );
  OAI21_X1 U8282 ( .B1(n6631), .B2(n6663), .A(n6630), .ZN(n6773) );
  XOR2_X1 U8283 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6775), .Z(n6774) );
  NAND2_X1 U8284 ( .A1(n6773), .A2(n6774), .ZN(n6772) );
  OAI21_X1 U8285 ( .B1(n6632), .B2(n6666), .A(n6772), .ZN(n6949) );
  MUX2_X1 U8286 ( .A(n6633), .B(P1_REG2_REG_4__SCAN_IN), .S(n6954), .Z(n6950)
         );
  NOR2_X1 U8287 ( .A1(n6949), .A2(n6950), .ZN(n6948) );
  INV_X1 U8288 ( .A(n6752), .ZN(n6635) );
  XNOR2_X1 U8289 ( .A(n6757), .B(n6634), .ZN(n6751) );
  INV_X1 U8290 ( .A(n6757), .ZN(n6672) );
  AOI22_X1 U8291 ( .A1(n6635), .A2(n6751), .B1(n6672), .B2(n6634), .ZN(n6928)
         );
  XNOR2_X1 U8292 ( .A(n6645), .B(n7515), .ZN(n6929) );
  NAND2_X1 U8293 ( .A1(n6928), .A2(n6929), .ZN(n6927) );
  XNOR2_X1 U8294 ( .A(n6768), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n6763) );
  NOR2_X1 U8295 ( .A1(n6738), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6636) );
  AOI21_X1 U8296 ( .B1(n6738), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6636), .ZN(
        n6730) );
  NAND2_X1 U8297 ( .A1(n6729), .A2(n6730), .ZN(n6728) );
  OAI21_X1 U8298 ( .B1(n6738), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6728), .ZN(
        n6638) );
  NAND2_X1 U8299 ( .A1(n6882), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6891) );
  OAI21_X1 U8300 ( .B1(n6882), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6891), .ZN(
        n6637) );
  OR2_X1 U8301 ( .A1(n6955), .A2(P1_U3084), .ZN(n7924) );
  NOR2_X1 U8302 ( .A1(n6654), .A2(n6958), .ZN(n9195) );
  AOI211_X1 U8303 ( .C1(n6638), .C2(n6637), .A(n6890), .B(n10245), .ZN(n6659)
         );
  XNOR2_X1 U8304 ( .A(n7020), .B(n6639), .ZN(n7012) );
  XNOR2_X1 U8305 ( .A(n6676), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n7000) );
  AND2_X1 U8306 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6999) );
  NAND2_X1 U8307 ( .A1(n7000), .A2(n6999), .ZN(n6998) );
  NAND2_X1 U8308 ( .A1(n7007), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U8309 ( .A1(n6998), .A2(n6640), .ZN(n7011) );
  NAND2_X1 U8310 ( .A1(n7012), .A2(n7011), .ZN(n7010) );
  NAND2_X1 U8311 ( .A1(n7020), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U8312 ( .A1(n7010), .A2(n6641), .ZN(n6777) );
  XNOR2_X1 U8313 ( .A(n6775), .B(n6642), .ZN(n6778) );
  NAND2_X1 U8314 ( .A1(n6777), .A2(n6778), .ZN(n6776) );
  OAI21_X1 U8315 ( .B1(n6642), .B2(n6666), .A(n6776), .ZN(n6944) );
  MUX2_X1 U8316 ( .A(n5847), .B(P1_REG1_REG_4__SCAN_IN), .S(n6954), .Z(n6945)
         );
  NOR2_X1 U8317 ( .A1(n6944), .A2(n6945), .ZN(n6943) );
  INV_X1 U8318 ( .A(n6943), .ZN(n6643) );
  OAI21_X1 U8319 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n6954), .A(n6643), .ZN(
        n6754) );
  XNOR2_X1 U8320 ( .A(n6757), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n6755) );
  NOR2_X1 U8321 ( .A1(n6754), .A2(n6755), .ZN(n6753) );
  AOI21_X1 U8322 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n6757), .A(n6753), .ZN(
        n6921) );
  XNOR2_X1 U8323 ( .A(n6645), .B(n6644), .ZN(n6922) );
  NAND2_X1 U8324 ( .A1(n6921), .A2(n6922), .ZN(n6920) );
  OAI21_X1 U8325 ( .B1(n6645), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6920), .ZN(
        n6765) );
  INV_X1 U8326 ( .A(n6765), .ZN(n6646) );
  XNOR2_X1 U8327 ( .A(n6768), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n6764) );
  OAI22_X1 U8328 ( .A1(n6646), .A2(n6764), .B1(n6768), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n6734) );
  AND2_X1 U8329 ( .A1(n6738), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6731) );
  INV_X1 U8330 ( .A(n6731), .ZN(n6647) );
  NOR2_X1 U8331 ( .A1(n6738), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6732) );
  AOI21_X1 U8332 ( .B1(n6734), .B2(n6647), .A(n6732), .ZN(n6649) );
  INV_X1 U8333 ( .A(n6882), .ZN(n6701) );
  AOI22_X1 U8334 ( .A1(n6882), .A2(n5953), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6701), .ZN(n6648) );
  NOR2_X1 U8335 ( .A1(n6649), .A2(n6648), .ZN(n6883) );
  AOI21_X1 U8336 ( .B1(n6649), .B2(n6648), .A(n6883), .ZN(n6653) );
  INV_X1 U8337 ( .A(n6650), .ZN(n6652) );
  NOR2_X1 U8338 ( .A1(n6958), .A2(P1_U3084), .ZN(n7932) );
  AND2_X1 U8339 ( .A1(n7932), .A2(n6955), .ZN(n6651) );
  NOR2_X1 U8340 ( .A1(n6653), .A2(n10257), .ZN(n6658) );
  NOR2_X2 U8341 ( .A1(n6654), .A2(n8195), .ZN(n10251) );
  INV_X1 U8342 ( .A(n10251), .ZN(n6967) );
  INV_X1 U8343 ( .A(n6655), .ZN(n6656) );
  INV_X1 U8344 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10482) );
  OAI22_X1 U8345 ( .A1(n6967), .A2(n6701), .B1(n10260), .B2(n10482), .ZN(n6657) );
  OR4_X1 U8346 ( .A1(n7709), .A2(n6659), .A3(n6658), .A4(n6657), .ZN(P1_U3250)
         );
  XNOR2_X1 U8347 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NOR2_X2 U8348 ( .A1(n6660), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9030) );
  AOI22_X1 U8349 ( .A1(n9030), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n10041), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6661) );
  OAI21_X1 U8350 ( .B1(n6664), .B2(n6706), .A(n6661), .ZN(P2_U3356) );
  AOI22_X1 U8351 ( .A1(n9030), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n6853), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6662) );
  OAI21_X1 U8352 ( .B1(n6667), .B2(n6706), .A(n6662), .ZN(P2_U3355) );
  OR2_X1 U8353 ( .A1(n7982), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9622) );
  INV_X1 U8354 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6665) );
  AND2_X1 U8355 ( .A1(n7982), .A2(P1_U3084), .ZN(n7923) );
  INV_X2 U8356 ( .A(n7923), .ZN(n9624) );
  OAI222_X1 U8357 ( .A1(n9622), .A2(n6665), .B1(n9624), .B2(n6664), .C1(
        P1_U3084), .C2(n6663), .ZN(P1_U3351) );
  INV_X1 U8358 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6668) );
  AOI22_X1 U8359 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n9030), .B1(n6840), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6669) );
  OAI21_X1 U8360 ( .B1(n6680), .B2(n6706), .A(n6669), .ZN(P2_U3354) );
  AOI22_X1 U8361 ( .A1(n9030), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n10023), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6670) );
  OAI21_X1 U8362 ( .B1(n6677), .B2(n6706), .A(n6670), .ZN(P2_U3357) );
  AOI22_X1 U8363 ( .A1(n6880), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n9030), .ZN(n6671) );
  OAI21_X1 U8364 ( .B1(n6673), .B2(n6706), .A(n6671), .ZN(P2_U3353) );
  INV_X1 U8365 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6674) );
  OAI222_X1 U8366 ( .A1(n9622), .A2(n6674), .B1(n9624), .B2(n6673), .C1(
        P1_U3084), .C2(n6672), .ZN(P1_U3348) );
  AOI22_X1 U8367 ( .A1(n6864), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n9030), .ZN(n6675) );
  OAI21_X1 U8368 ( .B1(n6682), .B2(n6706), .A(n6675), .ZN(P2_U3352) );
  INV_X1 U8369 ( .A(n9622), .ZN(n9617) );
  INV_X1 U8370 ( .A(n9617), .ZN(n9626) );
  INV_X1 U8371 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6678) );
  OAI222_X1 U8372 ( .A1(n9626), .A2(n6678), .B1(n9624), .B2(n6677), .C1(
        P1_U3084), .C2(n6676), .ZN(P1_U3352) );
  INV_X1 U8373 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6681) );
  OAI222_X1 U8374 ( .A1(n9626), .A2(n6681), .B1(n9624), .B2(n6680), .C1(
        P1_U3084), .C2(n6679), .ZN(P1_U3349) );
  INV_X1 U8375 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9802) );
  OAI222_X1 U8376 ( .A1(n9626), .A2(n9802), .B1(n9624), .B2(n6682), .C1(
        P1_U3084), .C2(n6924), .ZN(P1_U3347) );
  AOI22_X1 U8377 ( .A1(n6983), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n9030), .ZN(n6683) );
  OAI21_X1 U8378 ( .B1(n6685), .B2(n6706), .A(n6683), .ZN(P2_U3351) );
  AOI22_X1 U8379 ( .A1(n6768), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9617), .ZN(n6684) );
  OAI21_X1 U8380 ( .B1(n6685), .B2(n9624), .A(n6684), .ZN(P1_U3346) );
  INV_X1 U8381 ( .A(n9030), .ZN(n7930) );
  INV_X1 U8382 ( .A(n6686), .ZN(n6689) );
  INV_X1 U8383 ( .A(n7040), .ZN(n7031) );
  OAI222_X1 U8384 ( .A1(n7930), .A2(n6687), .B1(n6706), .B2(n6689), .C1(
        P2_U3152), .C2(n7031), .ZN(P2_U3350) );
  INV_X1 U8385 ( .A(n6738), .ZN(n6688) );
  OAI222_X1 U8386 ( .A1(n9622), .A2(n9987), .B1(n9624), .B2(n6689), .C1(
        P1_U3084), .C2(n6688), .ZN(P1_U3345) );
  INV_X1 U8387 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6692) );
  INV_X1 U8388 ( .A(n7323), .ZN(n6690) );
  NAND2_X1 U8389 ( .A1(n6690), .A2(n10288), .ZN(n6691) );
  OAI21_X1 U8390 ( .B1(n10288), .B2(n6692), .A(n6691), .ZN(P1_U3441) );
  INV_X1 U8391 ( .A(n6693), .ZN(n6702) );
  AOI22_X1 U8392 ( .A1(n8585), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n9030), .ZN(n6694) );
  OAI21_X1 U8393 ( .B1(n6702), .B2(n6706), .A(n6694), .ZN(P2_U3349) );
  OR2_X1 U8394 ( .A1(n6695), .A2(P2_U3152), .ZN(n8557) );
  OAI21_X1 U8395 ( .B1(n5210), .B2(n8557), .A(n10368), .ZN(n6698) );
  NAND2_X1 U8396 ( .A1(n5210), .A2(n6696), .ZN(n6697) );
  NAND2_X1 U8397 ( .A1(n6698), .A2(n6697), .ZN(n10026) );
  NOR2_X1 U8398 ( .A1(n10350), .A2(P2_U3966), .ZN(P2_U3151) );
  NAND2_X1 U8399 ( .A1(n6700), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6699) );
  OAI21_X1 U8400 ( .B1(n6904), .B2(n6700), .A(n6699), .ZN(P1_U3440) );
  OAI222_X1 U8401 ( .A1(n9626), .A2(n6703), .B1(n9624), .B2(n6702), .C1(n6701), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U8402 ( .A(n6704), .ZN(n6710) );
  AOI22_X1 U8403 ( .A1(n7098), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n9030), .ZN(n6705) );
  OAI21_X1 U8404 ( .B1(n6710), .B2(n6706), .A(n6705), .ZN(P2_U3348) );
  INV_X1 U8405 ( .A(n6707), .ZN(n6711) );
  AOI22_X1 U8406 ( .A1(n7165), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n9030), .ZN(n6708) );
  OAI21_X1 U8407 ( .B1(n6711), .B2(n6706), .A(n6708), .ZN(P2_U3347) );
  INV_X1 U8408 ( .A(n6962), .ZN(n6970) );
  OAI222_X1 U8409 ( .A1(P1_U3084), .A2(n6970), .B1(n9624), .B2(n6710), .C1(
        n6709), .C2(n9626), .ZN(P1_U3343) );
  OAI222_X1 U8410 ( .A1(P1_U3084), .A2(n7123), .B1(n9624), .B2(n6711), .C1(
        n9805), .C2(n9626), .ZN(P1_U3342) );
  INV_X1 U8411 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6713) );
  NAND2_X1 U8412 ( .A1(n7063), .A2(P1_U4006), .ZN(n6712) );
  OAI21_X1 U8413 ( .B1(P1_U4006), .B2(n6713), .A(n6712), .ZN(P1_U3555) );
  INV_X1 U8414 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6719) );
  NAND2_X1 U8415 ( .A1(n6195), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6717) );
  INV_X1 U8416 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6714) );
  OR2_X1 U8417 ( .A1(n6376), .A2(n6714), .ZN(n6716) );
  INV_X1 U8418 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9210) );
  OR2_X1 U8419 ( .A1(n8076), .A2(n9210), .ZN(n6715) );
  AND3_X1 U8420 ( .A1(n6717), .A2(n6716), .A3(n6715), .ZN(n9209) );
  INV_X1 U8421 ( .A(n9209), .ZN(n8086) );
  NAND2_X1 U8422 ( .A1(n8086), .A2(P1_U4006), .ZN(n6718) );
  OAI21_X1 U8423 ( .B1(P1_U4006), .B2(n6719), .A(n6718), .ZN(P1_U3586) );
  INV_X1 U8424 ( .A(n6720), .ZN(n6725) );
  AOI22_X1 U8425 ( .A1(n7293), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n9030), .ZN(n6721) );
  OAI21_X1 U8426 ( .B1(n6725), .B2(n6706), .A(n6721), .ZN(P2_U3346) );
  INV_X1 U8427 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9740) );
  INV_X1 U8428 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8988) );
  NAND2_X1 U8429 ( .A1(n4487), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6723) );
  INV_X1 U8430 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8903) );
  OR2_X1 U8431 ( .A1(n5637), .A2(n8903), .ZN(n6722) );
  OAI211_X1 U8432 ( .C1(n5229), .C2(n8988), .A(n6723), .B(n6722), .ZN(n8631)
         );
  NAND2_X1 U8433 ( .A1(n8631), .A2(P2_U3966), .ZN(n6724) );
  OAI21_X1 U8434 ( .B1(P2_U3966), .B2(n9740), .A(n6724), .ZN(P2_U3583) );
  INV_X1 U8435 ( .A(n9179), .ZN(n7119) );
  OAI222_X1 U8436 ( .A1(n9622), .A2(n6726), .B1(n9624), .B2(n6725), .C1(
        P1_U3084), .C2(n7119), .ZN(P1_U3341) );
  NAND2_X1 U8437 ( .A1(n8772), .A2(P2_U3966), .ZN(n6727) );
  OAI21_X1 U8438 ( .B1(P2_U3966), .B2(n5488), .A(n6727), .ZN(P2_U3573) );
  INV_X1 U8439 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6741) );
  OAI21_X1 U8440 ( .B1(n6730), .B2(n6729), .A(n6728), .ZN(n6736) );
  NOR2_X1 U8441 ( .A1(n6732), .A2(n6731), .ZN(n6733) );
  XNOR2_X1 U8442 ( .A(n6734), .B(n6733), .ZN(n6735) );
  AOI22_X1 U8443 ( .A1(n6736), .A2(n9195), .B1(n10238), .B2(n6735), .ZN(n6740)
         );
  INV_X1 U8444 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6737) );
  NOR2_X1 U8445 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6737), .ZN(n7640) );
  AOI21_X1 U8446 ( .B1(n10251), .B2(n6738), .A(n7640), .ZN(n6739) );
  OAI211_X1 U8447 ( .C1(n10260), .C2(n6741), .A(n6740), .B(n6739), .ZN(
        P1_U3249) );
  INV_X1 U8448 ( .A(n10260), .ZN(n6899) );
  INV_X1 U8449 ( .A(n6955), .ZN(n9207) );
  NAND2_X1 U8450 ( .A1(n9207), .A2(n5789), .ZN(n6742) );
  NAND2_X1 U8451 ( .A1(n8195), .A2(n6742), .ZN(n6745) );
  AOI21_X1 U8452 ( .B1(n6955), .B2(n6743), .A(P1_IR_REG_0__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U8453 ( .A1(n6745), .A2(n4756), .ZN(n6957) );
  OAI211_X1 U8454 ( .C1(n6745), .C2(n6744), .A(n6957), .B(P1_STATE_REG_SCAN_IN), .ZN(n6746) );
  OAI22_X1 U8455 ( .A1(n6747), .A2(n6746), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5788), .ZN(n6749) );
  NOR3_X1 U8456 ( .A1(n10257), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n4756), .ZN(
        n6748) );
  AOI211_X1 U8457 ( .C1(P1_ADDR_REG_0__SCAN_IN), .C2(n6899), .A(n6749), .B(
        n6748), .ZN(n6750) );
  INV_X1 U8458 ( .A(n6750), .ZN(P1_U3241) );
  XNOR2_X1 U8459 ( .A(n6752), .B(n6751), .ZN(n6760) );
  AND2_X1 U8460 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9084) );
  AOI211_X1 U8461 ( .C1(n6755), .C2(n6754), .A(n6753), .B(n10257), .ZN(n6756)
         );
  AOI211_X1 U8462 ( .C1(n10251), .C2(n6757), .A(n9084), .B(n6756), .ZN(n6759)
         );
  NAND2_X1 U8463 ( .A1(n6899), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n6758) );
  OAI211_X1 U8464 ( .C1(n10245), .C2(n6760), .A(n6759), .B(n6758), .ZN(
        P1_U3246) );
  AOI21_X1 U8465 ( .B1(n6763), .B2(n6762), .A(n6761), .ZN(n6771) );
  AND2_X1 U8466 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7531) );
  XNOR2_X1 U8467 ( .A(n6765), .B(n6764), .ZN(n6766) );
  NOR2_X1 U8468 ( .A1(n10257), .A2(n6766), .ZN(n6767) );
  AOI211_X1 U8469 ( .C1(n10251), .C2(n6768), .A(n7531), .B(n6767), .ZN(n6770)
         );
  NAND2_X1 U8470 ( .A1(n6899), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6769) );
  OAI211_X1 U8471 ( .C1(n6771), .C2(n10245), .A(n6770), .B(n6769), .ZN(
        P1_U3248) );
  INV_X1 U8472 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6784) );
  OAI211_X1 U8473 ( .C1(n6774), .C2(n6773), .A(n9195), .B(n6772), .ZN(n6782)
         );
  INV_X1 U8474 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7564) );
  NOR2_X1 U8475 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7564), .ZN(n7083) );
  INV_X1 U8476 ( .A(n7083), .ZN(n6781) );
  NAND2_X1 U8477 ( .A1(n10251), .A2(n6775), .ZN(n6780) );
  OAI211_X1 U8478 ( .C1(n6778), .C2(n6777), .A(n10238), .B(n6776), .ZN(n6779)
         );
  AND4_X1 U8479 ( .A1(n6782), .A2(n6781), .A3(n6780), .A4(n6779), .ZN(n6783)
         );
  OAI21_X1 U8480 ( .B1(n6784), .B2(n10260), .A(n6783), .ZN(P1_U3244) );
  INV_X1 U8481 ( .A(n6785), .ZN(n6787) );
  INV_X1 U8482 ( .A(n7395), .ZN(n7391) );
  OAI222_X1 U8483 ( .A1(n7930), .A2(n6786), .B1(n6706), .B2(n6787), .C1(n7391), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  OAI222_X1 U8484 ( .A1(n9622), .A2(n9792), .B1(n9624), .B2(n6787), .C1(n4633), 
        .C2(P1_U3084), .ZN(P1_U3340) );
  INV_X1 U8485 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6789) );
  INV_X1 U8486 ( .A(n6788), .ZN(n6790) );
  INV_X1 U8487 ( .A(n7649), .ZN(n7652) );
  OAI222_X1 U8488 ( .A1(n7930), .A2(n6789), .B1(n6706), .B2(n6790), .C1(n7652), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8489 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9914) );
  OAI222_X1 U8490 ( .A1(P1_U3084), .A2(n9184), .B1(n9624), .B2(n6790), .C1(
        n9914), .C2(n9626), .ZN(P1_U3339) );
  NOR2_X1 U8491 ( .A1(n5673), .A2(P2_U3152), .ZN(n7934) );
  INV_X1 U8492 ( .A(n6791), .ZN(n6792) );
  NAND2_X1 U8493 ( .A1(n7934), .A2(n6792), .ZN(n6793) );
  OAI211_X1 U8494 ( .C1(n6794), .C2(n10368), .A(n6793), .B(n8557), .ZN(n6797)
         );
  NAND2_X1 U8495 ( .A1(n6797), .A2(n5210), .ZN(n6795) );
  INV_X2 U8496 ( .A(P2_U3966), .ZN(n8578) );
  NAND2_X1 U8497 ( .A1(n6795), .A2(n8578), .ZN(n6823) );
  AND2_X1 U8498 ( .A1(n6823), .A2(n5673), .ZN(n10042) );
  AND2_X1 U8499 ( .A1(n5210), .A2(n8552), .ZN(n6796) );
  NAND2_X1 U8500 ( .A1(n6797), .A2(n6796), .ZN(n10344) );
  NAND2_X1 U8501 ( .A1(n6880), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U8502 ( .A1(n6853), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6803) );
  MUX2_X1 U8503 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6798), .S(n6853), .Z(n6843)
         );
  NAND2_X1 U8504 ( .A1(n10041), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6802) );
  MUX2_X1 U8505 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6799), .S(n10041), .Z(n10044) );
  NAND2_X1 U8506 ( .A1(n10023), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6801) );
  MUX2_X1 U8507 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6800), .S(n10023), .Z(n10033) );
  NAND3_X1 U8508 ( .A1(n10355), .A2(P2_REG1_REG_0__SCAN_IN), .A3(n10033), .ZN(
        n10032) );
  NAND2_X1 U8509 ( .A1(n6801), .A2(n10032), .ZN(n10045) );
  NAND2_X1 U8510 ( .A1(n10044), .A2(n10045), .ZN(n10043) );
  NAND2_X1 U8511 ( .A1(n6802), .A2(n10043), .ZN(n6844) );
  NAND2_X1 U8512 ( .A1(n6843), .A2(n6844), .ZN(n6842) );
  NAND2_X1 U8513 ( .A1(n6803), .A2(n6842), .ZN(n6831) );
  INV_X1 U8514 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6804) );
  MUX2_X1 U8515 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6804), .S(n6840), .Z(n6830)
         );
  NAND2_X1 U8516 ( .A1(n6831), .A2(n6830), .ZN(n6829) );
  NAND2_X1 U8517 ( .A1(n6840), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6805) );
  NAND2_X1 U8518 ( .A1(n6829), .A2(n6805), .ZN(n6872) );
  MUX2_X1 U8519 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6806), .S(n6880), .Z(n6871)
         );
  NAND2_X1 U8520 ( .A1(n6872), .A2(n6871), .ZN(n6807) );
  NAND2_X1 U8521 ( .A1(n6808), .A2(n6807), .ZN(n6811) );
  MUX2_X1 U8522 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6809), .S(n6864), .Z(n6810)
         );
  NAND2_X1 U8523 ( .A1(n6810), .A2(n6811), .ZN(n6855) );
  OAI21_X1 U8524 ( .B1(n6811), .B2(n6810), .A(n6855), .ZN(n6814) );
  NAND2_X1 U8525 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7487) );
  INV_X1 U8526 ( .A(n7487), .ZN(n6812) );
  AOI21_X1 U8527 ( .B1(n10350), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6812), .ZN(
        n6813) );
  OAI21_X1 U8528 ( .B1(n10344), .B2(n6814), .A(n6813), .ZN(n6827) );
  MUX2_X1 U8529 ( .A(n6815), .B(P2_REG2_REG_4__SCAN_IN), .S(n6840), .Z(n6836)
         );
  INV_X1 U8530 ( .A(n10355), .ZN(n10353) );
  INV_X1 U8531 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10360) );
  OR2_X1 U8532 ( .A1(n10023), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6817) );
  NAND2_X1 U8533 ( .A1(n10023), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6816) );
  NAND2_X1 U8534 ( .A1(n6817), .A2(n6816), .ZN(n10019) );
  NAND2_X1 U8535 ( .A1(n10041), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6818) );
  OAI21_X1 U8536 ( .B1(n10041), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6818), .ZN(
        n10038) );
  NAND2_X1 U8537 ( .A1(n6853), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6819) );
  OAI21_X1 U8538 ( .B1(n6853), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6819), .ZN(
        n6849) );
  NOR2_X1 U8539 ( .A1(n6850), .A2(n6849), .ZN(n6848) );
  NAND2_X1 U8540 ( .A1(n6880), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6820) );
  OAI21_X1 U8541 ( .B1(n6880), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6820), .ZN(
        n6876) );
  NAND2_X1 U8542 ( .A1(n6864), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6821) );
  OAI21_X1 U8543 ( .B1(n6864), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6821), .ZN(
        n6824) );
  NOR2_X1 U8544 ( .A1(n6825), .A2(n6824), .ZN(n6863) );
  NOR2_X1 U8545 ( .A1(n5673), .A2(n8552), .ZN(n6822) );
  NAND2_X1 U8546 ( .A1(n6823), .A2(n6822), .ZN(n10347) );
  AOI211_X1 U8547 ( .C1(n6825), .C2(n6824), .A(n6863), .B(n10347), .ZN(n6826)
         );
  AOI211_X1 U8548 ( .C1(n10042), .C2(n6864), .A(n6827), .B(n6826), .ZN(n6828)
         );
  INV_X1 U8549 ( .A(n6828), .ZN(P2_U3251) );
  OAI21_X1 U8550 ( .B1(n6831), .B2(n6830), .A(n6829), .ZN(n6834) );
  NAND2_X1 U8551 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7176) );
  INV_X1 U8552 ( .A(n7176), .ZN(n6832) );
  AOI21_X1 U8553 ( .B1(n10350), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6832), .ZN(
        n6833) );
  OAI21_X1 U8554 ( .B1(n10344), .B2(n6834), .A(n6833), .ZN(n6839) );
  AOI211_X1 U8555 ( .C1(n6837), .C2(n6836), .A(n6835), .B(n10347), .ZN(n6838)
         );
  AOI211_X1 U8556 ( .C1(n10042), .C2(n6840), .A(n6839), .B(n6838), .ZN(n6841)
         );
  INV_X1 U8557 ( .A(n6841), .ZN(P2_U3249) );
  OAI21_X1 U8558 ( .B1(n6844), .B2(n6843), .A(n6842), .ZN(n6847) );
  INV_X1 U8559 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9801) );
  NOR2_X1 U8560 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9801), .ZN(n6845) );
  AOI21_X1 U8561 ( .B1(n10350), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6845), .ZN(
        n6846) );
  OAI21_X1 U8562 ( .B1(n10344), .B2(n6847), .A(n6846), .ZN(n6852) );
  AOI211_X1 U8563 ( .C1(n6850), .C2(n6849), .A(n6848), .B(n10347), .ZN(n6851)
         );
  AOI211_X1 U8564 ( .C1(n10042), .C2(n6853), .A(n6852), .B(n6851), .ZN(n6854)
         );
  INV_X1 U8565 ( .A(n6854), .ZN(P2_U3248) );
  NAND2_X1 U8566 ( .A1(n6864), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6856) );
  NAND2_X1 U8567 ( .A1(n6856), .A2(n6855), .ZN(n6859) );
  MUX2_X1 U8568 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6857), .S(n6983), .Z(n6858)
         );
  NAND2_X1 U8569 ( .A1(n6858), .A2(n6859), .ZN(n6984) );
  OAI21_X1 U8570 ( .B1(n6859), .B2(n6858), .A(n6984), .ZN(n6862) );
  NOR2_X1 U8571 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5275), .ZN(n6860) );
  AOI21_X1 U8572 ( .B1(n10350), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6860), .ZN(
        n6861) );
  OAI21_X1 U8573 ( .B1(n10344), .B2(n6862), .A(n6861), .ZN(n6869) );
  AOI21_X1 U8574 ( .B1(n6864), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6863), .ZN(
        n6867) );
  NAND2_X1 U8575 ( .A1(n6983), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6865) );
  OAI21_X1 U8576 ( .B1(n6983), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6865), .ZN(
        n6866) );
  NOR2_X1 U8577 ( .A1(n6867), .A2(n6866), .ZN(n6979) );
  AOI211_X1 U8578 ( .C1(n6867), .C2(n6866), .A(n6979), .B(n10347), .ZN(n6868)
         );
  AOI211_X1 U8579 ( .C1(n10042), .C2(n6983), .A(n6869), .B(n6868), .ZN(n6870)
         );
  INV_X1 U8580 ( .A(n6870), .ZN(P2_U3252) );
  XNOR2_X1 U8581 ( .A(n6872), .B(n6871), .ZN(n6875) );
  NOR2_X1 U8582 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9924), .ZN(n6873) );
  AOI21_X1 U8583 ( .B1(n10350), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6873), .ZN(
        n6874) );
  OAI21_X1 U8584 ( .B1(n10344), .B2(n6875), .A(n6874), .ZN(n6879) );
  AOI211_X1 U8585 ( .C1(n6877), .C2(n6876), .A(n4515), .B(n10347), .ZN(n6878)
         );
  AOI211_X1 U8586 ( .C1(n10042), .C2(n6880), .A(n6879), .B(n6878), .ZN(n6881)
         );
  INV_X1 U8587 ( .A(n6881), .ZN(P2_U3250) );
  NOR2_X1 U8588 ( .A1(n6882), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6884) );
  NOR2_X1 U8589 ( .A1(n6884), .A2(n6883), .ZN(n6888) );
  MUX2_X1 U8590 ( .A(n6885), .B(P1_REG1_REG_10__SCAN_IN), .S(n6962), .Z(n6887)
         );
  INV_X1 U8591 ( .A(n6974), .ZN(n6886) );
  AOI21_X1 U8592 ( .B1(n6888), .B2(n6887), .A(n6886), .ZN(n6901) );
  XNOR2_X1 U8593 ( .A(n6962), .B(n6889), .ZN(n6893) );
  OAI211_X1 U8594 ( .C1(n6893), .C2(n6892), .A(n9195), .B(n6964), .ZN(n6897)
         );
  NOR2_X1 U8595 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6894), .ZN(n7729) );
  INV_X1 U8596 ( .A(n7729), .ZN(n6896) );
  NAND2_X1 U8597 ( .A1(n10251), .A2(n6962), .ZN(n6895) );
  NAND3_X1 U8598 ( .A1(n6897), .A2(n6896), .A3(n6895), .ZN(n6898) );
  AOI21_X1 U8599 ( .B1(n6899), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n6898), .ZN(
        n6900) );
  OAI21_X1 U8600 ( .B1(n6901), .B2(n10257), .A(n6900), .ZN(P1_U3251) );
  OR2_X2 U8601 ( .A1(n7329), .A2(n7074), .ZN(n10325) );
  OAI21_X1 U8602 ( .B1(n10325), .B2(n9322), .A(n7323), .ZN(n6902) );
  INV_X1 U8603 ( .A(n6903), .ZN(n6905) );
  NAND2_X1 U8604 ( .A1(n6905), .A2(n6904), .ZN(n7324) );
  INV_X1 U8605 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6909) );
  INV_X1 U8606 ( .A(n7480), .ZN(n7273) );
  INV_X1 U8607 ( .A(n7063), .ZN(n7070) );
  NOR2_X1 U8608 ( .A1(n7070), .A2(n7480), .ZN(n8208) );
  NOR2_X1 U8609 ( .A1(n8208), .A2(n7065), .ZN(n8102) );
  NAND2_X1 U8610 ( .A1(n8197), .A2(n7329), .ZN(n6906) );
  INV_X1 U8611 ( .A(n8204), .ZN(n7069) );
  OAI22_X1 U8612 ( .A1(n8102), .A2(n6906), .B1(n8211), .B2(n10128), .ZN(n7479)
         );
  INV_X1 U8613 ( .A(n7479), .ZN(n6907) );
  OAI21_X1 U8614 ( .B1(n7273), .B2(n7329), .A(n6907), .ZN(n9598) );
  NAND2_X1 U8615 ( .A1(n9598), .A2(n10333), .ZN(n6908) );
  OAI21_X1 U8616 ( .B1(n10333), .B2(n6909), .A(n6908), .ZN(P1_U3454) );
  NOR2_X1 U8617 ( .A1(n6910), .A2(n8890), .ZN(n10356) );
  INV_X1 U8618 ( .A(n10356), .ZN(n6918) );
  OR2_X1 U8619 ( .A1(n6911), .A2(P2_U3152), .ZN(n8553) );
  INV_X1 U8620 ( .A(n8553), .ZN(n7183) );
  NAND2_X1 U8621 ( .A1(n6912), .A2(n7183), .ZN(n7139) );
  AOI22_X1 U8622 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n7139), .B1(n8346), .B2(
        n10408), .ZN(n6917) );
  INV_X1 U8623 ( .A(n8363), .ZN(n6915) );
  NAND2_X1 U8624 ( .A1(n8579), .A2(n10361), .ZN(n8408) );
  INV_X1 U8625 ( .A(n8408), .ZN(n6913) );
  MUX2_X1 U8626 ( .A(n6913), .B(n10408), .S(n8951), .Z(n6914) );
  OAI21_X1 U8627 ( .B1(n6915), .B2(n6914), .A(n8329), .ZN(n6916) );
  OAI211_X1 U8628 ( .C1(n6919), .C2(n6918), .A(n6917), .B(n6916), .ZN(P2_U3234) );
  INV_X1 U8629 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6932) );
  OAI21_X1 U8630 ( .B1(n6922), .B2(n6921), .A(n6920), .ZN(n6926) );
  INV_X1 U8631 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6923) );
  NOR2_X1 U8632 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6923), .ZN(n7383) );
  NOR2_X1 U8633 ( .A1(n6967), .A2(n6924), .ZN(n6925) );
  AOI211_X1 U8634 ( .C1(n10238), .C2(n6926), .A(n7383), .B(n6925), .ZN(n6931)
         );
  OAI211_X1 U8635 ( .C1(n6929), .C2(n6928), .A(n9195), .B(n6927), .ZN(n6930)
         );
  OAI211_X1 U8636 ( .C1(n6932), .C2(n10260), .A(n6931), .B(n6930), .ZN(
        P1_U3247) );
  NAND2_X1 U8637 ( .A1(n6933), .A2(P2_U3966), .ZN(n6934) );
  OAI21_X1 U8638 ( .B1(P2_U3966), .B2(n5519), .A(n6934), .ZN(P2_U3575) );
  OAI21_X1 U8639 ( .B1(n6937), .B2(n6936), .A(n6935), .ZN(n6956) );
  AOI22_X1 U8640 ( .A1(n6956), .A2(n10101), .B1(n9152), .B2(n7062), .ZN(n6942)
         );
  INV_X1 U8641 ( .A(n6938), .ZN(n6939) );
  NAND2_X1 U8642 ( .A1(n10067), .A2(n6939), .ZN(n6940) );
  NAND2_X1 U8643 ( .A1(n9146), .A2(n6940), .ZN(n7053) );
  INV_X1 U8644 ( .A(n7053), .ZN(n6994) );
  NAND2_X1 U8645 ( .A1(n6994), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6941) );
  OAI211_X1 U8646 ( .C1(n9146), .C2(n7273), .A(n6942), .B(n6941), .ZN(P1_U3230) );
  INV_X1 U8647 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6961) );
  AOI21_X1 U8648 ( .B1(n6945), .B2(n6944), .A(n6943), .ZN(n6947) );
  AND2_X1 U8649 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7250) );
  INV_X1 U8650 ( .A(n7250), .ZN(n6946) );
  OAI21_X1 U8651 ( .B1(n10257), .B2(n6947), .A(n6946), .ZN(n6953) );
  AOI21_X1 U8652 ( .B1(n6950), .B2(n6949), .A(n6948), .ZN(n6951) );
  NOR2_X1 U8653 ( .A1(n10245), .A2(n6951), .ZN(n6952) );
  AOI211_X1 U8654 ( .C1(n10251), .C2(n6954), .A(n6953), .B(n6952), .ZN(n6960)
         );
  MUX2_X1 U8655 ( .A(n7004), .B(n6956), .S(n6955), .Z(n6959) );
  OAI211_X1 U8656 ( .C1(n6959), .C2(n6958), .A(P1_U4006), .B(n6957), .ZN(n7021) );
  OAI211_X1 U8657 ( .C1(n6961), .C2(n10260), .A(n6960), .B(n7021), .ZN(
        P1_U3245) );
  INV_X1 U8658 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6978) );
  NAND2_X1 U8659 ( .A1(n6962), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6963) );
  MUX2_X1 U8660 ( .A(n7122), .B(P1_REG2_REG_11__SCAN_IN), .S(n7123), .Z(n6965)
         );
  NAND2_X1 U8661 ( .A1(n6965), .A2(n6966), .ZN(n7125) );
  OAI21_X1 U8662 ( .B1(n6966), .B2(n6965), .A(n7125), .ZN(n6969) );
  AND2_X1 U8663 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7854) );
  NOR2_X1 U8664 ( .A1(n6967), .A2(n7123), .ZN(n6968) );
  AOI211_X1 U8665 ( .C1(n9195), .C2(n6969), .A(n7854), .B(n6968), .ZN(n6977)
         );
  NAND2_X1 U8666 ( .A1(n6970), .A2(n6885), .ZN(n6972) );
  MUX2_X1 U8667 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6971), .S(n7123), .Z(n6973)
         );
  AOI21_X1 U8668 ( .B1(n6974), .B2(n6972), .A(n6973), .ZN(n7118) );
  AND3_X1 U8669 ( .A1(n6974), .A2(n6973), .A3(n6972), .ZN(n6975) );
  OAI21_X1 U8670 ( .B1(n7118), .B2(n6975), .A(n10238), .ZN(n6976) );
  OAI211_X1 U8671 ( .C1(n10260), .C2(n6978), .A(n6977), .B(n6976), .ZN(
        P1_U3252) );
  XNOR2_X1 U8672 ( .A(n7040), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n6980) );
  NOR2_X1 U8673 ( .A1(n6981), .A2(n6980), .ZN(n7039) );
  AOI211_X1 U8674 ( .C1(n6981), .C2(n6980), .A(n7039), .B(n10347), .ZN(n6991)
         );
  INV_X1 U8675 ( .A(n10042), .ZN(n10346) );
  NOR2_X1 U8676 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7502), .ZN(n6982) );
  AOI21_X1 U8677 ( .B1(n10350), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6982), .ZN(
        n6989) );
  NAND2_X1 U8678 ( .A1(n6983), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6985) );
  NAND2_X1 U8679 ( .A1(n6985), .A2(n6984), .ZN(n6987) );
  MUX2_X1 U8680 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7032), .S(n7040), .Z(n6986)
         );
  INV_X1 U8681 ( .A(n10344), .ZN(n10342) );
  NAND2_X1 U8682 ( .A1(n6987), .A2(n6986), .ZN(n7030) );
  OAI211_X1 U8683 ( .C1(n6987), .C2(n6986), .A(n10342), .B(n7030), .ZN(n6988)
         );
  OAI211_X1 U8684 ( .C1(n10346), .C2(n7031), .A(n6989), .B(n6988), .ZN(n6990)
         );
  OR2_X1 U8685 ( .A1(n6991), .A2(n6990), .ZN(P2_U3253) );
  NOR2_X1 U8686 ( .A1(n10323), .A2(n7333), .ZN(n7276) );
  OAI22_X1 U8687 ( .A1(n7303), .A2(n10092), .B1(n10061), .B2(n8211), .ZN(n6993) );
  AOI21_X1 U8688 ( .B1(n7276), .B2(n7053), .A(n6993), .ZN(n6996) );
  NAND2_X1 U8689 ( .A1(n6994), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6995) );
  OAI211_X1 U8690 ( .C1(n6997), .C2(n9156), .A(n6996), .B(n6995), .ZN(P1_U3235) );
  INV_X1 U8691 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7009) );
  OAI211_X1 U8692 ( .C1(n7000), .C2(n6999), .A(n10238), .B(n6998), .ZN(n7001)
         );
  OAI21_X1 U8693 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7430), .A(n7001), .ZN(n7006) );
  AOI211_X1 U8694 ( .C1(n7004), .C2(n7003), .A(n7002), .B(n10245), .ZN(n7005)
         );
  AOI211_X1 U8695 ( .C1(n10251), .C2(n7007), .A(n7006), .B(n7005), .ZN(n7008)
         );
  OAI21_X1 U8696 ( .B1(n10260), .B2(n7009), .A(n7008), .ZN(P1_U3242) );
  INV_X1 U8697 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7023) );
  OAI211_X1 U8698 ( .C1(n7012), .C2(n7011), .A(n10238), .B(n7010), .ZN(n7013)
         );
  OAI21_X1 U8699 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7014), .A(n7013), .ZN(n7019) );
  AOI211_X1 U8700 ( .C1(n7017), .C2(n7016), .A(n7015), .B(n10245), .ZN(n7018)
         );
  AOI211_X1 U8701 ( .C1(n10251), .C2(n7020), .A(n7019), .B(n7018), .ZN(n7022)
         );
  OAI211_X1 U8702 ( .C1(n7023), .C2(n10260), .A(n7022), .B(n7021), .ZN(
        P1_U3243) );
  INV_X1 U8703 ( .A(n7024), .ZN(n7026) );
  INV_X1 U8704 ( .A(n10212), .ZN(n9186) );
  OAI222_X1 U8705 ( .A1(n9622), .A2(n7025), .B1(n9624), .B2(n7026), .C1(
        P1_U3084), .C2(n9186), .ZN(P1_U3338) );
  INV_X1 U8706 ( .A(n7772), .ZN(n7780) );
  OAI222_X1 U8707 ( .A1(n7930), .A2(n7027), .B1(n6706), .B2(n7026), .C1(
        P2_U3152), .C2(n7780), .ZN(P2_U3343) );
  MUX2_X1 U8708 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7028), .S(n7098), .Z(n7035)
         );
  NAND2_X1 U8709 ( .A1(n8585), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7033) );
  MUX2_X1 U8710 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7029), .S(n8585), .Z(n8587)
         );
  OAI21_X1 U8711 ( .B1(n7032), .B2(n7031), .A(n7030), .ZN(n8588) );
  NAND2_X1 U8712 ( .A1(n8587), .A2(n8588), .ZN(n8586) );
  NAND2_X1 U8713 ( .A1(n7033), .A2(n8586), .ZN(n7034) );
  NAND2_X1 U8714 ( .A1(n7035), .A2(n7034), .ZN(n7099) );
  OAI21_X1 U8715 ( .B1(n7035), .B2(n7034), .A(n7099), .ZN(n7038) );
  NOR2_X1 U8716 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9977), .ZN(n7036) );
  AOI21_X1 U8717 ( .B1(n10350), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7036), .ZN(
        n7037) );
  OAI21_X1 U8718 ( .B1(n10344), .B2(n7038), .A(n7037), .ZN(n7047) );
  OR2_X1 U8719 ( .A1(n8585), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7042) );
  NAND2_X1 U8720 ( .A1(n8585), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7041) );
  NAND2_X1 U8721 ( .A1(n7042), .A2(n7041), .ZN(n8581) );
  NOR2_X1 U8722 ( .A1(n8582), .A2(n8581), .ZN(n8580) );
  AOI21_X1 U8723 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n8585), .A(n8580), .ZN(
        n7045) );
  NAND2_X1 U8724 ( .A1(n7098), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7043) );
  OAI21_X1 U8725 ( .B1(n7098), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7043), .ZN(
        n7044) );
  AOI211_X1 U8726 ( .C1(n7045), .C2(n7044), .A(n7094), .B(n10347), .ZN(n7046)
         );
  AOI211_X1 U8727 ( .C1(n10042), .C2(n7098), .A(n7047), .B(n7046), .ZN(n7048)
         );
  INV_X1 U8728 ( .A(n7048), .ZN(P2_U3255) );
  NAND2_X1 U8729 ( .A1(n7050), .A2(n7049), .ZN(n7051) );
  XOR2_X1 U8730 ( .A(n7052), .B(n7051), .Z(n7057) );
  NOR2_X1 U8731 ( .A1(n10323), .A2(n7274), .ZN(n7076) );
  OAI22_X1 U8732 ( .A1(n7070), .A2(n10061), .B1(n10092), .B2(n7556), .ZN(n7055) );
  NOR2_X1 U8733 ( .A1(n7053), .A2(n7430), .ZN(n7054) );
  AOI211_X1 U8734 ( .C1(n10067), .C2(n7076), .A(n7055), .B(n7054), .ZN(n7056)
         );
  OAI21_X1 U8735 ( .B1(n7057), .B2(n9156), .A(n7056), .ZN(P1_U3220) );
  OR2_X1 U8736 ( .A1(n7058), .A2(n7334), .ZN(n7061) );
  OR2_X1 U8737 ( .A1(n7059), .A2(n8253), .ZN(n7060) );
  AND2_X1 U8738 ( .A1(n7063), .A2(n7480), .ZN(n7064) );
  OAI21_X1 U8739 ( .B1(n8105), .B2(n7064), .A(n7261), .ZN(n7436) );
  NAND2_X1 U8740 ( .A1(n7066), .A2(n7065), .ZN(n7267) );
  OAI21_X1 U8741 ( .B1(n7066), .B2(n7065), .A(n7267), .ZN(n7072) );
  NAND2_X1 U8742 ( .A1(n6336), .A2(n9200), .ZN(n7068) );
  NAND2_X1 U8743 ( .A1(n6337), .A2(n7074), .ZN(n7067) );
  OAI22_X1 U8744 ( .A1(n7070), .A2(n10129), .B1(n10128), .B2(n7556), .ZN(n7071) );
  AOI21_X1 U8745 ( .B1(n7072), .B2(n10266), .A(n7071), .ZN(n7073) );
  OAI21_X1 U8746 ( .B1(n10272), .B2(n7436), .A(n7073), .ZN(n7433) );
  NAND2_X1 U8747 ( .A1(n5786), .A2(n9200), .ZN(n8061) );
  OR2_X1 U8748 ( .A1(n8061), .A2(n7074), .ZN(n10170) );
  NOR2_X1 U8749 ( .A1(n7436), .A2(n10170), .ZN(n7077) );
  XNOR2_X1 U8750 ( .A(n7274), .B(n7273), .ZN(n7075) );
  NOR2_X1 U8751 ( .A1(n7075), .A2(n10325), .ZN(n7429) );
  NOR4_X1 U8752 ( .A1(n7433), .A2(n7077), .A3(n7076), .A4(n7429), .ZN(n10291)
         );
  NAND2_X1 U8753 ( .A1(n10339), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7080) );
  OAI21_X1 U8754 ( .B1(n10291), .B2(n10339), .A(n7080), .ZN(P1_U3524) );
  XNOR2_X1 U8755 ( .A(n7081), .B(n7082), .ZN(n7088) );
  NOR2_X1 U8756 ( .A1(n9146), .A2(n10292), .ZN(n7087) );
  AOI21_X1 U8757 ( .B1(n9152), .B2(n9166), .A(n7083), .ZN(n7085) );
  NAND2_X1 U8758 ( .A1(n10090), .A2(n9168), .ZN(n7084) );
  OAI211_X1 U8759 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n10106), .A(n7085), .B(
        n7084), .ZN(n7086) );
  AOI211_X1 U8760 ( .C1(n7088), .C2(n10101), .A(n7087), .B(n7086), .ZN(n7089)
         );
  INV_X1 U8761 ( .A(n7089), .ZN(P1_U3216) );
  INV_X1 U8762 ( .A(n7090), .ZN(n7145) );
  AOI22_X1 U8763 ( .A1(n7811), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n9030), .ZN(n7091) );
  OAI21_X1 U8764 ( .B1(n7145), .B2(n6706), .A(n7091), .ZN(P2_U3342) );
  NAND2_X1 U8765 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n8578), .ZN(n7092) );
  OAI21_X1 U8766 ( .B1(n8284), .B2(n8578), .A(n7092), .ZN(P2_U3578) );
  NAND2_X1 U8767 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8578), .ZN(n7093) );
  OAI21_X1 U8768 ( .B1(n8649), .B2(n8578), .A(n7093), .ZN(P2_U3581) );
  INV_X1 U8769 ( .A(n10347), .ZN(n10343) );
  MUX2_X1 U8770 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n7764), .S(n7165), .Z(n7096)
         );
  OAI21_X1 U8771 ( .B1(n7096), .B2(n7095), .A(n7166), .ZN(n7108) );
  MUX2_X1 U8772 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7097), .S(n7165), .Z(n7102)
         );
  NAND2_X1 U8773 ( .A1(n7098), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7100) );
  NAND2_X1 U8774 ( .A1(n7100), .A2(n7099), .ZN(n7101) );
  NAND2_X1 U8775 ( .A1(n7102), .A2(n7101), .ZN(n7157) );
  OAI21_X1 U8776 ( .B1(n7102), .B2(n7101), .A(n7157), .ZN(n7106) );
  NAND2_X1 U8777 ( .A1(n10042), .A2(n7165), .ZN(n7105) );
  NOR2_X1 U8778 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5342), .ZN(n7103) );
  AOI21_X1 U8779 ( .B1(n10350), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7103), .ZN(
        n7104) );
  OAI211_X1 U8780 ( .C1(n10344), .C2(n7106), .A(n7105), .B(n7104), .ZN(n7107)
         );
  AOI21_X1 U8781 ( .B1(n10343), .B2(n7108), .A(n7107), .ZN(n7109) );
  INV_X1 U8782 ( .A(n7109), .ZN(P2_U3256) );
  OAI21_X1 U8783 ( .B1(n7110), .B2(n7112), .A(n7111), .ZN(n7116) );
  NOR2_X1 U8784 ( .A1(n8343), .A2(n8418), .ZN(n7115) );
  AOI22_X1 U8785 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(n7139), .B1(n8346), .B2(
        n6391), .ZN(n7113) );
  OAI21_X1 U8786 ( .B1(n8342), .B2(n6399), .A(n7113), .ZN(n7114) );
  AOI211_X1 U8787 ( .C1(n8329), .C2(n7116), .A(n7115), .B(n7114), .ZN(n7117)
         );
  INV_X1 U8788 ( .A(n7117), .ZN(P2_U3224) );
  AOI21_X1 U8789 ( .B1(n6971), .B2(n7123), .A(n7118), .ZN(n7121) );
  AOI22_X1 U8790 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n7119), .B1(n9179), .B2(
        n6009), .ZN(n7120) );
  NOR2_X1 U8791 ( .A1(n7121), .A2(n7120), .ZN(n9181) );
  AOI21_X1 U8792 ( .B1(n7121), .B2(n7120), .A(n9181), .ZN(n7136) );
  INV_X1 U8793 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7133) );
  AND2_X1 U8794 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10057) );
  AOI21_X1 U8795 ( .B1(n10251), .B2(n9179), .A(n10057), .ZN(n7132) );
  NAND2_X1 U8796 ( .A1(n7123), .A2(n7122), .ZN(n7124) );
  NAND2_X1 U8797 ( .A1(n7125), .A2(n7124), .ZN(n7129) );
  OR2_X1 U8798 ( .A1(n9179), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7127) );
  NAND2_X1 U8799 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9179), .ZN(n7126) );
  NAND2_X1 U8800 ( .A1(n7127), .A2(n7126), .ZN(n7128) );
  AOI21_X1 U8801 ( .B1(n7129), .B2(n7128), .A(n9169), .ZN(n7130) );
  NAND2_X1 U8802 ( .A1(n9195), .A2(n7130), .ZN(n7131) );
  OAI211_X1 U8803 ( .C1(n7133), .C2(n10260), .A(n7132), .B(n7131), .ZN(n7134)
         );
  INV_X1 U8804 ( .A(n7134), .ZN(n7135) );
  OAI21_X1 U8805 ( .B1(n7136), .B2(n10257), .A(n7135), .ZN(P1_U3253) );
  XOR2_X1 U8806 ( .A(n7138), .B(n7137), .Z(n7143) );
  NOR2_X1 U8807 ( .A1(n8343), .A2(n6910), .ZN(n7142) );
  AOI22_X1 U8808 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(n7139), .B1(n8346), .B2(
        n7231), .ZN(n7140) );
  OAI21_X1 U8809 ( .B1(n8342), .B2(n7198), .A(n7140), .ZN(n7141) );
  AOI211_X1 U8810 ( .C1(n7143), .C2(n8329), .A(n7142), .B(n7141), .ZN(n7144)
         );
  INV_X1 U8811 ( .A(n7144), .ZN(P2_U3239) );
  INV_X1 U8812 ( .A(n10223), .ZN(n9189) );
  OAI222_X1 U8813 ( .A1(n9626), .A2(n9804), .B1(n9624), .B2(n7145), .C1(n9189), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  NAND2_X1 U8814 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n8578), .ZN(n7146) );
  OAI21_X1 U8815 ( .B1(n8650), .B2(n8578), .A(n7146), .ZN(P2_U3579) );
  XNOR2_X1 U8816 ( .A(n7148), .B(n7147), .ZN(n7153) );
  NAND2_X1 U8817 ( .A1(n8346), .A2(n7351), .ZN(n7149) );
  OAI21_X1 U8818 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n9801), .A(n7149), .ZN(n7151) );
  OAI22_X1 U8819 ( .A1(n6399), .A2(n8343), .B1(n8342), .B2(n7407), .ZN(n7150)
         );
  AOI211_X1 U8820 ( .C1(n8299), .C2(n9801), .A(n7151), .B(n7150), .ZN(n7152)
         );
  OAI21_X1 U8821 ( .B1(n7153), .B2(n8348), .A(n7152), .ZN(P2_U3220) );
  INV_X1 U8822 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7155) );
  INV_X1 U8823 ( .A(n7154), .ZN(n7156) );
  INV_X1 U8824 ( .A(n8594), .ZN(n8600) );
  OAI222_X1 U8825 ( .A1(n7930), .A2(n7155), .B1(n6706), .B2(n7156), .C1(n8600), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8826 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9937) );
  INV_X1 U8827 ( .A(n10236), .ZN(n9191) );
  OAI222_X1 U8828 ( .A1(n9626), .A2(n9937), .B1(n9624), .B2(n7156), .C1(n9191), 
        .C2(P1_U3084), .ZN(P1_U3336) );
  INV_X1 U8829 ( .A(n7293), .ZN(n7284) );
  INV_X1 U8830 ( .A(n7157), .ZN(n7158) );
  AOI21_X1 U8831 ( .B1(n7165), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7158), .ZN(
        n7160) );
  MUX2_X1 U8832 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n5362), .S(n7293), .Z(n7159)
         );
  NAND2_X1 U8833 ( .A1(n7160), .A2(n7159), .ZN(n7286) );
  OAI21_X1 U8834 ( .B1(n7160), .B2(n7159), .A(n7286), .ZN(n7164) );
  NOR2_X1 U8835 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9789), .ZN(n7163) );
  INV_X1 U8836 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7161) );
  NOR2_X1 U8837 ( .A1(n10026), .A2(n7161), .ZN(n7162) );
  AOI211_X1 U8838 ( .C1(n10342), .C2(n7164), .A(n7163), .B(n7162), .ZN(n7171)
         );
  INV_X1 U8839 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7800) );
  XNOR2_X1 U8840 ( .A(n7293), .B(n7800), .ZN(n7169) );
  OR2_X1 U8841 ( .A1(n7165), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7167) );
  NAND2_X1 U8842 ( .A1(n7168), .A2(n7169), .ZN(n7295) );
  OAI211_X1 U8843 ( .C1(n7169), .C2(n7168), .A(n10343), .B(n7295), .ZN(n7170)
         );
  OAI211_X1 U8844 ( .C1(n10346), .C2(n7284), .A(n7171), .B(n7170), .ZN(
        P2_U3257) );
  AOI21_X1 U8845 ( .B1(n7172), .B2(n7175), .A(n7174), .ZN(n7181) );
  INV_X1 U8846 ( .A(n7240), .ZN(n7179) );
  OAI21_X1 U8847 ( .B1(n8335), .B2(n7239), .A(n7176), .ZN(n7178) );
  OAI22_X1 U8848 ( .A1(n7198), .A2(n8343), .B1(n8342), .B2(n7489), .ZN(n7177)
         );
  AOI211_X1 U8849 ( .C1(n7179), .C2(n8299), .A(n7178), .B(n7177), .ZN(n7180)
         );
  OAI21_X1 U8850 ( .B1(n7181), .B2(n8348), .A(n7180), .ZN(P2_U3232) );
  NAND2_X1 U8851 ( .A1(n7183), .A2(n7182), .ZN(n7184) );
  NOR2_X1 U8852 ( .A1(n7185), .A2(n7184), .ZN(n7186) );
  NAND2_X1 U8853 ( .A1(n7187), .A2(n7186), .ZN(n7202) );
  INV_X1 U8854 ( .A(n8877), .ZN(n7188) );
  OR2_X1 U8855 ( .A1(n7189), .A2(n8622), .ZN(n7350) );
  AND2_X1 U8856 ( .A1(n7882), .A2(n7350), .ZN(n7190) );
  XNOR2_X1 U8857 ( .A(n7191), .B(n7193), .ZN(n7230) );
  INV_X1 U8858 ( .A(n7230), .ZN(n7207) );
  INV_X1 U8859 ( .A(n7195), .ZN(n7196) );
  AOI21_X1 U8860 ( .B1(n7192), .B2(n7194), .A(n7196), .ZN(n7197) );
  OAI222_X1 U8861 ( .A1(n8890), .A2(n7198), .B1(n8892), .B2(n6910), .C1(n8889), 
        .C2(n7197), .ZN(n7228) );
  INV_X1 U8862 ( .A(n7200), .ZN(n8417) );
  INV_X1 U8863 ( .A(n7352), .ZN(n7201) );
  AOI211_X1 U8864 ( .C1(n7231), .C2(n8417), .A(n10436), .B(n7201), .ZN(n7229)
         );
  OR2_X1 U8865 ( .A1(n7202), .A2(n8390), .ZN(n7950) );
  INV_X1 U8866 ( .A(n7950), .ZN(n8830) );
  NAND2_X1 U8867 ( .A1(n7229), .A2(n8830), .ZN(n7204) );
  INV_X1 U8868 ( .A(n10358), .ZN(n8848) );
  AOI22_X1 U8869 ( .A1(n8877), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n8848), .ZN(n7203) );
  OAI211_X1 U8870 ( .C1(n7233), .C2(n10362), .A(n7204), .B(n7203), .ZN(n7205)
         );
  AOI21_X1 U8871 ( .B1(n7228), .B2(n7188), .A(n7205), .ZN(n7206) );
  OAI21_X1 U8872 ( .B1(n8809), .B2(n7207), .A(n7206), .ZN(P2_U3294) );
  XNOR2_X1 U8873 ( .A(n7209), .B(n7208), .ZN(n7214) );
  INV_X1 U8874 ( .A(n7210), .ZN(n7413) );
  OAI22_X1 U8875 ( .A1(n8335), .A2(n7573), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9924), .ZN(n7212) );
  OAI22_X1 U8876 ( .A1(n7407), .A2(n8343), .B1(n8342), .B2(n7423), .ZN(n7211)
         );
  AOI211_X1 U8877 ( .C1(n7413), .C2(n8299), .A(n7212), .B(n7211), .ZN(n7213)
         );
  OAI21_X1 U8878 ( .B1(n7214), .B2(n8348), .A(n7213), .ZN(P2_U3229) );
  XNOR2_X1 U8879 ( .A(n7215), .B(n8363), .ZN(n7218) );
  NAND2_X1 U8880 ( .A1(n8579), .A2(n8816), .ZN(n7216) );
  OAI21_X1 U8881 ( .B1(n6399), .B2(n8890), .A(n7216), .ZN(n7217) );
  AOI21_X1 U8882 ( .B1(n7218), .B2(n10357), .A(n7217), .ZN(n10416) );
  OR2_X1 U8883 ( .A1(n7219), .A2(n7215), .ZN(n7220) );
  AND2_X1 U8884 ( .A1(n7221), .A2(n7220), .ZN(n10415) );
  NAND2_X1 U8885 ( .A1(n10408), .A2(n6391), .ZN(n8420) );
  AND2_X1 U8886 ( .A1(n8420), .A2(n8951), .ZN(n7222) );
  NAND2_X1 U8887 ( .A1(n8417), .A2(n7222), .ZN(n10412) );
  INV_X1 U8888 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10024) );
  OAI22_X1 U8889 ( .A1(n7950), .A2(n10412), .B1(n10024), .B2(n10358), .ZN(
        n7223) );
  INV_X1 U8890 ( .A(n7223), .ZN(n7225) );
  NAND2_X1 U8891 ( .A1(n8877), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7224) );
  OAI211_X1 U8892 ( .C1(n10362), .C2(n10413), .A(n7225), .B(n7224), .ZN(n7226)
         );
  AOI21_X1 U8893 ( .B1(n10366), .B2(n10415), .A(n7226), .ZN(n7227) );
  OAI21_X1 U8894 ( .B1(n8897), .B2(n10416), .A(n7227), .ZN(P2_U3295) );
  AOI211_X1 U8895 ( .C1(n7230), .C2(n10440), .A(n7229), .B(n7228), .ZN(n7236)
         );
  AOI22_X1 U8896 ( .A1(n7604), .A2(n7231), .B1(n10450), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n7232) );
  OAI21_X1 U8897 ( .B1(n7236), .B2(n10450), .A(n7232), .ZN(P2_U3522) );
  OAI22_X1 U8898 ( .A1(n9019), .A2(n7233), .B1(n10444), .B2(n5213), .ZN(n7234)
         );
  INV_X1 U8899 ( .A(n7234), .ZN(n7235) );
  OAI21_X1 U8900 ( .B1(n7236), .B2(n10442), .A(n7235), .ZN(P2_U3457) );
  XOR2_X1 U8901 ( .A(n7237), .B(n8364), .Z(n7238) );
  AOI222_X1 U8902 ( .A1(n10357), .A2(n7238), .B1(n8573), .B2(n8815), .C1(n8575), .C2(n8816), .ZN(n7365) );
  AOI21_X1 U8903 ( .B1(n7362), .B2(n7353), .A(n7410), .ZN(n7363) );
  NOR2_X1 U8904 ( .A1(n7950), .A2(n10436), .ZN(n8874) );
  NOR2_X1 U8905 ( .A1(n10362), .A2(n7239), .ZN(n7242) );
  OAI22_X1 U8906 ( .A1(n7188), .A2(n6815), .B1(n7240), .B2(n10358), .ZN(n7241)
         );
  AOI211_X1 U8907 ( .C1(n7363), .C2(n8874), .A(n7242), .B(n7241), .ZN(n7246)
         );
  OAI21_X1 U8908 ( .B1(n7244), .B2(n8364), .A(n7243), .ZN(n7361) );
  NAND2_X1 U8909 ( .A1(n7361), .A2(n10366), .ZN(n7245) );
  OAI211_X1 U8910 ( .C1(n7365), .C2(n8877), .A(n7246), .B(n7245), .ZN(P2_U3292) );
  INV_X1 U8911 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7248) );
  INV_X1 U8912 ( .A(n7247), .ZN(n7249) );
  OAI222_X1 U8913 ( .A1(n7930), .A2(n7248), .B1(n6706), .B2(n7249), .C1(
        P2_U3152), .C2(n8616), .ZN(P2_U3340) );
  INV_X1 U8914 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9920) );
  INV_X1 U8915 ( .A(n10252), .ZN(n9193) );
  OAI222_X1 U8916 ( .A1(n9626), .A2(n9920), .B1(n9624), .B2(n7249), .C1(
        P1_U3084), .C2(n9193), .ZN(P1_U3335) );
  INV_X1 U8917 ( .A(n7940), .ZN(n7307) );
  AOI21_X1 U8918 ( .B1(n9152), .B2(n9165), .A(n7250), .ZN(n7252) );
  NAND2_X1 U8919 ( .A1(n10090), .A2(n9167), .ZN(n7251) );
  OAI211_X1 U8920 ( .C1(n10106), .C2(n7939), .A(n7252), .B(n7251), .ZN(n7258)
         );
  INV_X1 U8921 ( .A(n7254), .ZN(n7255) );
  AOI211_X1 U8922 ( .C1(n7256), .C2(n7253), .A(n9156), .B(n7255), .ZN(n7257)
         );
  AOI211_X1 U8923 ( .C1(n10095), .C2(n7307), .A(n7258), .B(n7257), .ZN(n7259)
         );
  INV_X1 U8924 ( .A(n7259), .ZN(P1_U3228) );
  INV_X1 U8925 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7279) );
  NAND2_X1 U8926 ( .A1(n9168), .A2(n7333), .ZN(n8217) );
  INV_X1 U8927 ( .A(n7274), .ZN(n8210) );
  NAND2_X1 U8928 ( .A1(n7062), .A2(n8210), .ZN(n7260) );
  NAND2_X1 U8929 ( .A1(n7261), .A2(n7260), .ZN(n7265) );
  INV_X1 U8930 ( .A(n7265), .ZN(n7263) );
  NAND2_X1 U8931 ( .A1(n7263), .A2(n7262), .ZN(n7302) );
  INV_X1 U8932 ( .A(n7302), .ZN(n7264) );
  AOI21_X1 U8933 ( .B1(n8100), .B2(n7265), .A(n7264), .ZN(n7336) );
  NAND2_X1 U8934 ( .A1(n8211), .A2(n8210), .ZN(n7266) );
  AOI22_X1 U8935 ( .A1(n10264), .A2(n9167), .B1(n10263), .B2(n7062), .ZN(n7268) );
  OAI21_X1 U8936 ( .B1(n7336), .B2(n10272), .A(n7268), .ZN(n7269) );
  AOI21_X1 U8937 ( .B1(n7270), .B2(n10266), .A(n7269), .ZN(n7341) );
  INV_X1 U8938 ( .A(n10325), .ZN(n10165) );
  INV_X1 U8939 ( .A(n7333), .ZN(n7272) );
  NAND2_X1 U8940 ( .A1(n7274), .A2(n7273), .ZN(n7271) );
  NAND2_X1 U8941 ( .A1(n7272), .A2(n7271), .ZN(n7275) );
  NAND3_X1 U8942 ( .A1(n7333), .A2(n7274), .A3(n7273), .ZN(n7560) );
  AND2_X1 U8943 ( .A1(n7275), .A2(n7560), .ZN(n7339) );
  AOI21_X1 U8944 ( .B1(n10165), .B2(n7339), .A(n7276), .ZN(n7277) );
  OAI211_X1 U8945 ( .C1(n7336), .C2(n10170), .A(n7341), .B(n7277), .ZN(n7280)
         );
  NAND2_X1 U8946 ( .A1(n7280), .A2(n10333), .ZN(n7278) );
  OAI21_X1 U8947 ( .B1(n10333), .B2(n7279), .A(n7278), .ZN(P1_U3460) );
  NAND2_X1 U8948 ( .A1(n7280), .A2(n10341), .ZN(n7281) );
  OAI21_X1 U8949 ( .B1(n10341), .B2(n6639), .A(n7281), .ZN(P1_U3525) );
  INV_X1 U8950 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7283) );
  OAI22_X1 U8951 ( .A1(n10026), .A2(n7283), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7282), .ZN(n7291) );
  AOI22_X1 U8952 ( .A1(n7395), .A2(n5377), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7391), .ZN(n7288) );
  NAND2_X1 U8953 ( .A1(n7284), .A2(n5362), .ZN(n7285) );
  AND2_X1 U8954 ( .A1(n7286), .A2(n7285), .ZN(n7287) );
  NOR2_X1 U8955 ( .A1(n7287), .A2(n7288), .ZN(n7390) );
  AOI21_X1 U8956 ( .B1(n7288), .B2(n7287), .A(n7390), .ZN(n7289) );
  NOR2_X1 U8957 ( .A1(n10344), .A2(n7289), .ZN(n7290) );
  AOI211_X1 U8958 ( .C1(n10042), .C2(n7395), .A(n7291), .B(n7290), .ZN(n7300)
         );
  NOR2_X1 U8959 ( .A1(n7395), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7292) );
  AOI21_X1 U8960 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7395), .A(n7292), .ZN(
        n7297) );
  NAND2_X1 U8961 ( .A1(n7293), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7294) );
  OAI21_X1 U8962 ( .B1(n7297), .B2(n7296), .A(n7394), .ZN(n7298) );
  NAND2_X1 U8963 ( .A1(n10343), .A2(n7298), .ZN(n7299) );
  NAND2_X1 U8964 ( .A1(n7300), .A2(n7299), .ZN(P2_U3258) );
  INV_X1 U8965 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7317) );
  INV_X1 U8966 ( .A(n10170), .ZN(n10330) );
  NAND2_X1 U8967 ( .A1(n7556), .A2(n7333), .ZN(n7301) );
  NAND2_X1 U8968 ( .A1(n7302), .A2(n7301), .ZN(n7554) );
  OR2_X1 U8969 ( .A1(n9167), .A2(n10292), .ZN(n8215) );
  NAND2_X1 U8970 ( .A1(n9167), .A2(n10292), .ZN(n8219) );
  NAND2_X1 U8971 ( .A1(n8215), .A2(n8219), .ZN(n8103) );
  NAND2_X1 U8972 ( .A1(n7554), .A2(n8103), .ZN(n7553) );
  NAND2_X1 U8973 ( .A1(n7303), .A2(n10292), .ZN(n7304) );
  NAND2_X1 U8974 ( .A1(n7553), .A2(n7304), .ZN(n7305) );
  NAND2_X1 U8975 ( .A1(n9166), .A2(n7940), .ZN(n7999) );
  NAND2_X1 U8976 ( .A1(n8157), .A2(n7999), .ZN(n8104) );
  OR2_X1 U8977 ( .A1(n7305), .A2(n8104), .ZN(n7306) );
  NAND2_X1 U8978 ( .A1(n7440), .A2(n7306), .ZN(n7938) );
  INV_X1 U8979 ( .A(n10292), .ZN(n7563) );
  OR2_X1 U8980 ( .A1(n7560), .A2(n7563), .ZN(n7562) );
  INV_X1 U8981 ( .A(n7449), .ZN(n7450) );
  NAND2_X1 U8982 ( .A1(n7562), .A2(n7307), .ZN(n7308) );
  NAND2_X1 U8983 ( .A1(n7450), .A2(n7308), .ZN(n7944) );
  OAI22_X1 U8984 ( .A1(n7944), .A2(n10325), .B1(n7940), .B2(n10323), .ZN(n7315) );
  NAND2_X1 U8985 ( .A1(n7309), .A2(n8213), .ZN(n8159) );
  INV_X1 U8986 ( .A(n8103), .ZN(n7310) );
  NAND2_X1 U8987 ( .A1(n8159), .A2(n7310), .ZN(n7311) );
  XNOR2_X1 U8988 ( .A(n8000), .B(n8104), .ZN(n7314) );
  INV_X1 U8989 ( .A(n10272), .ZN(n7697) );
  NAND2_X1 U8990 ( .A1(n7938), .A2(n7697), .ZN(n7313) );
  AOI22_X1 U8991 ( .A1(n10264), .A2(n9165), .B1(n10263), .B2(n9167), .ZN(n7312) );
  OAI211_X1 U8992 ( .C1(n9477), .C2(n7314), .A(n7313), .B(n7312), .ZN(n7937)
         );
  AOI211_X1 U8993 ( .C1(n10330), .C2(n7938), .A(n7315), .B(n7937), .ZN(n7318)
         );
  OR2_X1 U8994 ( .A1(n7318), .A2(n10331), .ZN(n7316) );
  OAI21_X1 U8995 ( .B1(n10333), .B2(n7317), .A(n7316), .ZN(P1_U3466) );
  OR2_X1 U8996 ( .A1(n7318), .A2(n10339), .ZN(n7319) );
  OAI21_X1 U8997 ( .B1(n10341), .B2(n5847), .A(n7319), .ZN(P1_U3527) );
  INV_X1 U8998 ( .A(n7320), .ZN(n7322) );
  OAI222_X1 U8999 ( .A1(n7930), .A2(n7321), .B1(n6706), .B2(n7322), .C1(
        P2_U3152), .C2(n8622), .ZN(P2_U3339) );
  OAI222_X1 U9000 ( .A1(n9626), .A2(n9950), .B1(n9624), .B2(n7322), .C1(n9322), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OR2_X1 U9001 ( .A1(n7324), .A2(n7323), .ZN(n7325) );
  NAND2_X1 U9002 ( .A1(n10288), .A2(n9200), .ZN(n7327) );
  INV_X1 U9003 ( .A(n8242), .ZN(n7328) );
  OR2_X1 U9004 ( .A1(n7329), .A2(n7328), .ZN(n7330) );
  INV_X1 U9005 ( .A(n9512), .ZN(n10282) );
  INV_X1 U9006 ( .A(n9505), .ZN(n10275) );
  AOI22_X1 U9007 ( .A1(n4483), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10275), .ZN(n7332) );
  OAI21_X1 U9008 ( .B1(n9484), .B2(n7333), .A(n7332), .ZN(n7338) );
  NAND2_X1 U9009 ( .A1(n7334), .A2(n9200), .ZN(n7335) );
  OR2_X1 U9010 ( .A1(n4483), .A2(n7335), .ZN(n7845) );
  NOR2_X1 U9011 ( .A1(n7336), .A2(n7845), .ZN(n7337) );
  AOI211_X1 U9012 ( .C1(n7339), .C2(n10282), .A(n7338), .B(n7337), .ZN(n7340)
         );
  OAI21_X1 U9013 ( .B1(n4483), .B2(n7341), .A(n7340), .ZN(P1_U3289) );
  OAI21_X1 U9014 ( .B1(n7343), .B2(n8367), .A(n7342), .ZN(n10422) );
  INV_X1 U9015 ( .A(n10422), .ZN(n7349) );
  OAI21_X1 U9016 ( .B1(n8413), .B2(n7345), .A(n7344), .ZN(n7347) );
  OAI22_X1 U9017 ( .A1(n6399), .A2(n8892), .B1(n7407), .B2(n8890), .ZN(n7346)
         );
  AOI21_X1 U9018 ( .B1(n7347), .B2(n10357), .A(n7346), .ZN(n7348) );
  OAI21_X1 U9019 ( .B1(n7349), .B2(n7882), .A(n7348), .ZN(n10420) );
  INV_X1 U9020 ( .A(n10420), .ZN(n7360) );
  NOR2_X1 U9021 ( .A1(n8897), .A2(n7350), .ZN(n8854) );
  AOI21_X1 U9022 ( .B1(n7352), .B2(n7351), .A(n10436), .ZN(n7354) );
  NAND2_X1 U9023 ( .A1(n7354), .A2(n7353), .ZN(n10418) );
  NOR2_X1 U9024 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(n10358), .ZN(n7356) );
  NOR2_X1 U9025 ( .A1(n10362), .A2(n10419), .ZN(n7355) );
  AOI211_X1 U9026 ( .C1(n8877), .C2(P2_REG2_REG_3__SCAN_IN), .A(n7356), .B(
        n7355), .ZN(n7357) );
  OAI21_X1 U9027 ( .B1(n7950), .B2(n10418), .A(n7357), .ZN(n7358) );
  AOI21_X1 U9028 ( .B1(n8854), .B2(n10422), .A(n7358), .ZN(n7359) );
  OAI21_X1 U9029 ( .B1(n7360), .B2(n8897), .A(n7359), .ZN(P2_U3293) );
  INV_X1 U9030 ( .A(n10440), .ZN(n8971) );
  INV_X1 U9031 ( .A(n7361), .ZN(n7366) );
  AOI22_X1 U9032 ( .A1(n7363), .A2(n8951), .B1(n8982), .B2(n7362), .ZN(n7364)
         );
  OAI211_X1 U9033 ( .C1(n8971), .C2(n7366), .A(n7365), .B(n7364), .ZN(n7368)
         );
  NAND2_X1 U9034 ( .A1(n7368), .A2(n10452), .ZN(n7367) );
  OAI21_X1 U9035 ( .B1(n10452), .B2(n6804), .A(n7367), .ZN(P2_U3524) );
  NAND2_X1 U9036 ( .A1(n7368), .A2(n10444), .ZN(n7369) );
  OAI21_X1 U9037 ( .B1(n10444), .B2(n5240), .A(n7369), .ZN(P2_U3463) );
  NAND3_X1 U9038 ( .A1(n7371), .A2(n8368), .A3(n8404), .ZN(n7372) );
  NAND2_X1 U9039 ( .A1(n7370), .A2(n7372), .ZN(n7373) );
  AOI222_X1 U9040 ( .A1(n10357), .A2(n7373), .B1(n8571), .B2(n8815), .C1(n8573), .C2(n8816), .ZN(n7600) );
  INV_X1 U9041 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7374) );
  OAI22_X1 U9042 ( .A1(n7188), .A2(n7374), .B1(n7488), .B2(n10358), .ZN(n7376)
         );
  OAI211_X1 U9043 ( .C1(n7411), .C2(n7606), .A(n8951), .B(n7543), .ZN(n7599)
         );
  NOR2_X1 U9044 ( .A1(n7599), .A2(n7950), .ZN(n7375) );
  AOI211_X1 U9045 ( .C1(n8885), .C2(n7603), .A(n7376), .B(n7375), .ZN(n7380)
         );
  OAI21_X1 U9046 ( .B1(n7378), .B2(n8368), .A(n7377), .ZN(n7602) );
  NAND2_X1 U9047 ( .A1(n7602), .A2(n10366), .ZN(n7379) );
  OAI211_X1 U9048 ( .C1(n7600), .C2(n8877), .A(n7380), .B(n7379), .ZN(P2_U3290) );
  XNOR2_X1 U9049 ( .A(n7381), .B(n7382), .ZN(n7388) );
  NOR2_X1 U9050 ( .A1(n9146), .A2(n10304), .ZN(n7387) );
  AOI21_X1 U9051 ( .B1(n9152), .B2(n9163), .A(n7383), .ZN(n7385) );
  NAND2_X1 U9052 ( .A1(n10090), .A2(n9165), .ZN(n7384) );
  OAI211_X1 U9053 ( .C1(n10106), .C2(n7514), .A(n7385), .B(n7384), .ZN(n7386)
         );
  AOI211_X1 U9054 ( .C1(n7388), .C2(n10101), .A(n7387), .B(n7386), .ZN(n7389)
         );
  INV_X1 U9055 ( .A(n7389), .ZN(P1_U3237) );
  AOI21_X1 U9056 ( .B1(n7391), .B2(n5377), .A(n7390), .ZN(n7393) );
  AOI22_X1 U9057 ( .A1(n7649), .A2(n8977), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7652), .ZN(n7392) );
  NOR2_X1 U9058 ( .A1(n7393), .A2(n7392), .ZN(n7651) );
  AOI21_X1 U9059 ( .B1(n7393), .B2(n7392), .A(n7651), .ZN(n7402) );
  AOI22_X1 U9060 ( .A1(n7649), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n5394), .B2(
        n7652), .ZN(n7397) );
  OAI21_X1 U9061 ( .B1(n7397), .B2(n7396), .A(n7648), .ZN(n7400) );
  NAND2_X1 U9062 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7849) );
  NAND2_X1 U9063 ( .A1(n10350), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7398) );
  OAI211_X1 U9064 ( .C1(n10346), .C2(n7652), .A(n7849), .B(n7398), .ZN(n7399)
         );
  AOI21_X1 U9065 ( .B1(n7400), .B2(n10343), .A(n7399), .ZN(n7401) );
  OAI21_X1 U9066 ( .B1(n7402), .B2(n10344), .A(n7401), .ZN(P2_U3259) );
  NAND2_X1 U9067 ( .A1(n7404), .A2(n7403), .ZN(n7405) );
  XOR2_X1 U9068 ( .A(n8365), .B(n7405), .Z(n7406) );
  OAI222_X1 U9069 ( .A1(n8890), .A2(n7423), .B1(n8892), .B2(n7407), .C1(n8889), 
        .C2(n7406), .ZN(n7570) );
  INV_X1 U9070 ( .A(n7570), .ZN(n7418) );
  OAI21_X1 U9071 ( .B1(n7409), .B2(n8365), .A(n7408), .ZN(n7572) );
  INV_X1 U9072 ( .A(n7410), .ZN(n7412) );
  AOI211_X1 U9073 ( .C1(n7576), .C2(n7412), .A(n10436), .B(n7411), .ZN(n7571)
         );
  NAND2_X1 U9074 ( .A1(n7571), .A2(n8830), .ZN(n7415) );
  AOI22_X1 U9075 ( .A1(n8877), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n7413), .B2(
        n8848), .ZN(n7414) );
  OAI211_X1 U9076 ( .C1(n7573), .C2(n10362), .A(n7415), .B(n7414), .ZN(n7416)
         );
  AOI21_X1 U9077 ( .B1(n10366), .B2(n7572), .A(n7416), .ZN(n7417) );
  OAI21_X1 U9078 ( .B1(n7418), .B2(n8897), .A(n7417), .ZN(P2_U3291) );
  NAND2_X1 U9079 ( .A1(n7484), .A2(n7485), .ZN(n7483) );
  NAND2_X1 U9080 ( .A1(n7483), .A2(n7419), .ZN(n7421) );
  XNOR2_X1 U9081 ( .A(n7421), .B(n7420), .ZN(n7428) );
  INV_X1 U9082 ( .A(n7541), .ZN(n7426) );
  NAND2_X1 U9083 ( .A1(n8346), .A2(n4482), .ZN(n7422) );
  OAI21_X1 U9084 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n5275), .A(n7422), .ZN(n7425) );
  OAI22_X1 U9085 ( .A1(n7423), .A2(n8343), .B1(n8342), .B2(n7613), .ZN(n7424)
         );
  AOI211_X1 U9086 ( .C1(n7426), .C2(n8299), .A(n7425), .B(n7424), .ZN(n7427)
         );
  OAI21_X1 U9087 ( .B1(n7428), .B2(n8348), .A(n7427), .ZN(P2_U3215) );
  INV_X1 U9088 ( .A(n7429), .ZN(n7431) );
  OAI22_X1 U9089 ( .A1(n7431), .A2(n9200), .B1(n9505), .B2(n7430), .ZN(n7432)
         );
  OAI21_X1 U9090 ( .B1(n7433), .B2(n7432), .A(n9508), .ZN(n7435) );
  AOI22_X1 U9091 ( .A1(n10276), .A2(n8210), .B1(n4483), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7434) );
  OAI211_X1 U9092 ( .C1(n7436), .C2(n7845), .A(n7435), .B(n7434), .ZN(P1_U3290) );
  NAND2_X1 U9093 ( .A1(n8197), .A2(n7437), .ZN(n7438) );
  NAND2_X1 U9094 ( .A1(n7555), .A2(n7940), .ZN(n7439) );
  NAND2_X1 U9095 ( .A1(n9165), .A2(n9081), .ZN(n7457) );
  OAI21_X1 U9096 ( .B1(n7441), .B2(n7444), .A(n7467), .ZN(n10299) );
  INV_X1 U9097 ( .A(n8157), .ZN(n7442) );
  OR2_X1 U9098 ( .A1(n8000), .A2(n7442), .ZN(n7443) );
  NAND2_X1 U9099 ( .A1(n7443), .A2(n7999), .ZN(n7445) );
  NOR2_X1 U9100 ( .A1(n7445), .A2(n7444), .ZN(n7509) );
  AND2_X1 U9101 ( .A1(n7445), .A2(n7444), .ZN(n7446) );
  OAI21_X1 U9102 ( .B1(n7509), .B2(n7446), .A(n10266), .ZN(n7448) );
  AOI22_X1 U9103 ( .A1(n10263), .A2(n9166), .B1(n10264), .B2(n9164), .ZN(n7447) );
  NAND2_X1 U9104 ( .A1(n7448), .A2(n7447), .ZN(n10302) );
  INV_X1 U9105 ( .A(n9081), .ZN(n7465) );
  AOI211_X1 U9106 ( .C1(n7465), .C2(n7450), .A(n10325), .B(n4888), .ZN(n10300)
         );
  INV_X1 U9107 ( .A(n10300), .ZN(n7452) );
  INV_X1 U9108 ( .A(n9085), .ZN(n7451) );
  OAI22_X1 U9109 ( .A1(n7452), .A2(n9200), .B1(n9505), .B2(n7451), .ZN(n7453)
         );
  OAI21_X1 U9110 ( .B1(n10302), .B2(n7453), .A(n9508), .ZN(n7455) );
  AOI22_X1 U9111 ( .A1(n10276), .A2(n7465), .B1(n4483), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n7454) );
  OAI211_X1 U9112 ( .C1(n9481), .C2(n10299), .A(n7455), .B(n7454), .ZN(
        P1_U3286) );
  NAND2_X1 U9113 ( .A1(n9163), .A2(n10312), .ZN(n8225) );
  NAND2_X1 U9114 ( .A1(n8006), .A2(n8225), .ZN(n8003) );
  INV_X1 U9115 ( .A(n8003), .ZN(n7463) );
  NAND2_X1 U9116 ( .A1(n7999), .A2(n7457), .ZN(n8220) );
  NAND2_X1 U9117 ( .A1(n9164), .A2(n10304), .ZN(n8005) );
  INV_X1 U9118 ( .A(n8005), .ZN(n8222) );
  NOR2_X1 U9119 ( .A1(n8220), .A2(n8222), .ZN(n7456) );
  NAND2_X1 U9120 ( .A1(n8000), .A2(n7456), .ZN(n7461) );
  NAND2_X1 U9121 ( .A1(n8157), .A2(n8160), .ZN(n7458) );
  NAND2_X1 U9122 ( .A1(n7458), .A2(n7457), .ZN(n8001) );
  INV_X1 U9123 ( .A(n8001), .ZN(n7460) );
  INV_X1 U9124 ( .A(n8161), .ZN(n7459) );
  AOI21_X1 U9125 ( .B1(n7460), .B2(n8005), .A(n7459), .ZN(n8224) );
  NAND2_X1 U9126 ( .A1(n7461), .A2(n8224), .ZN(n7462) );
  OAI21_X1 U9127 ( .B1(n7463), .B2(n7462), .A(n7587), .ZN(n7464) );
  AOI222_X1 U9128 ( .A1(n10266), .A2(n7464), .B1(n10262), .B2(n10264), .C1(
        n9164), .C2(n10263), .ZN(n10311) );
  NAND2_X1 U9129 ( .A1(n9165), .A2(n7465), .ZN(n7466) );
  NAND2_X1 U9130 ( .A1(n8161), .A2(n8005), .ZN(n8002) );
  NAND2_X1 U9131 ( .A1(n7508), .A2(n8002), .ZN(n7507) );
  NAND2_X1 U9132 ( .A1(n9082), .A2(n10304), .ZN(n7468) );
  NAND2_X1 U9133 ( .A1(n7469), .A2(n8003), .ZN(n7581) );
  OAI21_X1 U9134 ( .B1(n7469), .B2(n8003), .A(n7581), .ZN(n10314) );
  INV_X1 U9135 ( .A(n9481), .ZN(n9382) );
  NAND2_X1 U9136 ( .A1(n10314), .A2(n9382), .ZN(n7478) );
  OAI22_X1 U9137 ( .A1(n9508), .A2(n7470), .B1(n7534), .B2(n9505), .ZN(n7475)
         );
  INV_X1 U9138 ( .A(n10304), .ZN(n7521) );
  INV_X1 U9139 ( .A(n7518), .ZN(n7472) );
  INV_X1 U9140 ( .A(n7592), .ZN(n7471) );
  OAI211_X1 U9141 ( .C1(n10312), .C2(n7472), .A(n7471), .B(n10165), .ZN(n10310) );
  NOR2_X1 U9142 ( .A1(n7473), .A2(n9200), .ZN(n9490) );
  INV_X1 U9143 ( .A(n9490), .ZN(n9387) );
  NOR2_X1 U9144 ( .A1(n10310), .A2(n9387), .ZN(n7474) );
  AOI211_X1 U9145 ( .C1(n10276), .C2(n7476), .A(n7475), .B(n7474), .ZN(n7477)
         );
  OAI211_X1 U9146 ( .C1(n4483), .C2(n10311), .A(n7478), .B(n7477), .ZN(
        P1_U3284) );
  AOI22_X1 U9147 ( .A1(n7479), .A2(n9508), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n10275), .ZN(n7482) );
  OAI21_X1 U9148 ( .B1(n10282), .B2(n10276), .A(n7480), .ZN(n7481) );
  OAI211_X1 U9149 ( .C1(n5789), .C2(n9508), .A(n7482), .B(n7481), .ZN(P1_U3291) );
  OAI21_X1 U9150 ( .B1(n7485), .B2(n7484), .A(n7483), .ZN(n7492) );
  NAND2_X1 U9151 ( .A1(n8346), .A2(n7603), .ZN(n7486) );
  OAI211_X1 U9152 ( .C1(n8341), .C2(n7488), .A(n7487), .B(n7486), .ZN(n7491)
         );
  OAI22_X1 U9153 ( .A1(n7489), .A2(n8343), .B1(n8342), .B2(n7625), .ZN(n7490)
         );
  AOI211_X1 U9154 ( .C1(n7492), .C2(n8329), .A(n7491), .B(n7490), .ZN(n7493)
         );
  INV_X1 U9155 ( .A(n7493), .ZN(P2_U3241) );
  INV_X1 U9156 ( .A(n7494), .ZN(n7497) );
  OAI222_X1 U9157 ( .A1(P2_U3152), .A2(n8366), .B1(n6706), .B2(n7497), .C1(
        n7495), .C2(n7930), .ZN(P2_U3338) );
  OAI222_X1 U9158 ( .A1(P1_U3084), .A2(n8244), .B1(n9624), .B2(n7497), .C1(
        n7496), .C2(n9622), .ZN(P1_U3333) );
  XNOR2_X1 U9159 ( .A(n7498), .B(n7499), .ZN(n7506) );
  INV_X1 U9160 ( .A(n7500), .ZN(n7630) );
  NAND2_X1 U9161 ( .A1(n8346), .A2(n7631), .ZN(n7501) );
  OAI21_X1 U9162 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7502), .A(n7501), .ZN(n7504) );
  OAI22_X1 U9163 ( .A1(n7625), .A2(n8343), .B1(n8342), .B2(n7742), .ZN(n7503)
         );
  AOI211_X1 U9164 ( .C1(n7630), .C2(n8299), .A(n7504), .B(n7503), .ZN(n7505)
         );
  OAI21_X1 U9165 ( .B1(n7506), .B2(n8348), .A(n7505), .ZN(P2_U3223) );
  OAI21_X1 U9166 ( .B1(n7508), .B2(n8002), .A(n7507), .ZN(n10308) );
  INV_X1 U9167 ( .A(n10308), .ZN(n7524) );
  INV_X1 U9168 ( .A(n8160), .ZN(n7997) );
  NOR2_X1 U9169 ( .A1(n7509), .A2(n7997), .ZN(n7510) );
  XOR2_X1 U9170 ( .A(n8002), .B(n7510), .Z(n7513) );
  AOI22_X1 U9171 ( .A1(n10263), .A2(n9165), .B1(n10264), .B2(n9163), .ZN(n7512) );
  NAND2_X1 U9172 ( .A1(n10308), .A2(n7697), .ZN(n7511) );
  OAI211_X1 U9173 ( .C1(n7513), .C2(n9477), .A(n7512), .B(n7511), .ZN(n10306)
         );
  NAND2_X1 U9174 ( .A1(n10306), .A2(n9508), .ZN(n7523) );
  OAI22_X1 U9175 ( .A1(n9508), .A2(n7515), .B1(n7514), .B2(n9505), .ZN(n7520)
         );
  NAND2_X1 U9176 ( .A1(n7516), .A2(n7521), .ZN(n7517) );
  NAND2_X1 U9177 ( .A1(n7518), .A2(n7517), .ZN(n10305) );
  NOR2_X1 U9178 ( .A1(n10305), .A2(n9512), .ZN(n7519) );
  AOI211_X1 U9179 ( .C1(n10276), .C2(n7521), .A(n7520), .B(n7519), .ZN(n7522)
         );
  OAI211_X1 U9180 ( .C1(n7524), .C2(n7845), .A(n7523), .B(n7522), .ZN(P1_U3285) );
  INV_X1 U9181 ( .A(n7525), .ZN(n8254) );
  OAI222_X1 U9182 ( .A1(P2_U3152), .A2(n8355), .B1(n6706), .B2(n8254), .C1(
        n7526), .C2(n7930), .ZN(P2_U3337) );
  XNOR2_X1 U9183 ( .A(n7529), .B(n7528), .ZN(n7530) );
  XNOR2_X1 U9184 ( .A(n7527), .B(n7530), .ZN(n7537) );
  NOR2_X1 U9185 ( .A1(n9146), .A2(n10312), .ZN(n7536) );
  AOI21_X1 U9186 ( .B1(n9152), .B2(n10262), .A(n7531), .ZN(n7533) );
  NAND2_X1 U9187 ( .A1(n10090), .A2(n9164), .ZN(n7532) );
  OAI211_X1 U9188 ( .C1(n10106), .C2(n7534), .A(n7533), .B(n7532), .ZN(n7535)
         );
  AOI211_X1 U9189 ( .C1(n7537), .C2(n10101), .A(n7536), .B(n7535), .ZN(n7538)
         );
  INV_X1 U9190 ( .A(n7538), .ZN(P1_U3211) );
  OAI21_X1 U9191 ( .B1(n8430), .B2(n7539), .A(n7622), .ZN(n7540) );
  AOI222_X1 U9192 ( .A1(n10357), .A2(n7540), .B1(n8570), .B2(n8815), .C1(n8572), .C2(n8816), .ZN(n10425) );
  INV_X1 U9193 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7542) );
  OAI22_X1 U9194 ( .A1(n7188), .A2(n7542), .B1(n7541), .B2(n10358), .ZN(n7546)
         );
  AOI21_X1 U9195 ( .B1(n7543), .B2(n4482), .A(n10436), .ZN(n7544) );
  NAND2_X1 U9196 ( .A1(n7544), .A2(n7628), .ZN(n10424) );
  NOR2_X1 U9197 ( .A1(n10424), .A2(n7950), .ZN(n7545) );
  AOI211_X1 U9198 ( .C1(n8885), .C2(n4482), .A(n7546), .B(n7545), .ZN(n7552)
         );
  OAI21_X1 U9199 ( .B1(n7550), .B2(n7549), .A(n7548), .ZN(n10428) );
  NAND2_X1 U9200 ( .A1(n10428), .A2(n10366), .ZN(n7551) );
  OAI211_X1 U9201 ( .C1(n10425), .C2(n8877), .A(n7552), .B(n7551), .ZN(
        P2_U3289) );
  XNOR2_X1 U9202 ( .A(n8159), .B(n8103), .ZN(n7559) );
  OAI21_X1 U9203 ( .B1(n7554), .B2(n8103), .A(n7553), .ZN(n10296) );
  OAI22_X1 U9204 ( .A1(n7556), .A2(n10129), .B1(n10128), .B2(n7555), .ZN(n7557) );
  AOI21_X1 U9205 ( .B1(n10296), .B2(n7697), .A(n7557), .ZN(n7558) );
  OAI21_X1 U9206 ( .B1(n9477), .B2(n7559), .A(n7558), .ZN(n10294) );
  INV_X1 U9207 ( .A(n10294), .ZN(n7569) );
  NAND2_X1 U9208 ( .A1(n7560), .A2(n7563), .ZN(n7561) );
  NAND2_X1 U9209 ( .A1(n7562), .A2(n7561), .ZN(n10293) );
  NAND2_X1 U9210 ( .A1(n10276), .A2(n7563), .ZN(n7566) );
  AOI22_X1 U9211 ( .A1(n4483), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10275), .B2(
        n7564), .ZN(n7565) );
  OAI211_X1 U9212 ( .C1(n10293), .C2(n9512), .A(n7566), .B(n7565), .ZN(n7567)
         );
  AOI21_X1 U9213 ( .B1(n10296), .B2(n10283), .A(n7567), .ZN(n7568) );
  OAI21_X1 U9214 ( .B1(n7569), .B2(n4483), .A(n7568), .ZN(P1_U3288) );
  AOI211_X1 U9215 ( .C1(n10440), .C2(n7572), .A(n7571), .B(n7570), .ZN(n7578)
         );
  OAI22_X1 U9216 ( .A1(n9019), .A2(n7573), .B1(n10444), .B2(n5251), .ZN(n7574)
         );
  INV_X1 U9217 ( .A(n7574), .ZN(n7575) );
  OAI21_X1 U9218 ( .B1(n7578), .B2(n10442), .A(n7575), .ZN(P2_U3466) );
  AOI22_X1 U9219 ( .A1(n7604), .A2(n7576), .B1(n10450), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n7577) );
  OAI21_X1 U9220 ( .B1(n7578), .B2(n10450), .A(n7577), .ZN(P2_U3525) );
  OR2_X1 U9221 ( .A1(n10262), .A2(n10316), .ZN(n8146) );
  NAND2_X1 U9222 ( .A1(n10262), .A2(n10316), .ZN(n8167) );
  NAND2_X1 U9223 ( .A1(n8146), .A2(n8167), .ZN(n7585) );
  INV_X1 U9224 ( .A(n7585), .ZN(n8108) );
  INV_X1 U9225 ( .A(n9163), .ZN(n7579) );
  NAND2_X1 U9226 ( .A1(n7579), .A2(n10312), .ZN(n7580) );
  NAND2_X1 U9227 ( .A1(n7581), .A2(n7580), .ZN(n7584) );
  INV_X1 U9228 ( .A(n7584), .ZN(n7582) );
  NAND2_X1 U9229 ( .A1(n7582), .A2(n7585), .ZN(n7687) );
  INV_X1 U9230 ( .A(n7687), .ZN(n7583) );
  AOI21_X1 U9231 ( .B1(n8108), .B2(n7584), .A(n7583), .ZN(n10321) );
  INV_X1 U9232 ( .A(n10321), .ZN(n7598) );
  INV_X1 U9233 ( .A(n8006), .ZN(n8154) );
  NOR2_X1 U9234 ( .A1(n8154), .A2(n7585), .ZN(n7586) );
  NAND2_X1 U9235 ( .A1(n7587), .A2(n7586), .ZN(n7690) );
  NAND2_X1 U9236 ( .A1(n7690), .A2(n10266), .ZN(n7590) );
  AOI21_X1 U9237 ( .B1(n7587), .B2(n8006), .A(n8108), .ZN(n7589) );
  AOI22_X1 U9238 ( .A1(n10263), .A2(n9163), .B1(n10264), .B2(n9162), .ZN(n7588) );
  OAI21_X1 U9239 ( .B1(n7590), .B2(n7589), .A(n7588), .ZN(n10319) );
  INV_X1 U9240 ( .A(n10280), .ZN(n7591) );
  OAI21_X1 U9241 ( .B1(n10316), .B2(n7592), .A(n7591), .ZN(n10317) );
  OAI22_X1 U9242 ( .A1(n9508), .A2(n7593), .B1(n7643), .B2(n9505), .ZN(n7594)
         );
  AOI21_X1 U9243 ( .B1(n10276), .B2(n7685), .A(n7594), .ZN(n7595) );
  OAI21_X1 U9244 ( .B1(n10317), .B2(n9512), .A(n7595), .ZN(n7596) );
  AOI21_X1 U9245 ( .B1(n10319), .B2(n9508), .A(n7596), .ZN(n7597) );
  OAI21_X1 U9246 ( .B1(n7598), .B2(n9481), .A(n7597), .ZN(P1_U3283) );
  NAND2_X1 U9247 ( .A1(n7600), .A2(n7599), .ZN(n7601) );
  AOI21_X1 U9248 ( .B1(n10440), .B2(n7602), .A(n7601), .ZN(n7609) );
  AOI22_X1 U9249 ( .A1(n7604), .A2(n7603), .B1(n10450), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n7605) );
  OAI21_X1 U9250 ( .B1(n7609), .B2(n10450), .A(n7605), .ZN(P2_U3526) );
  OAI22_X1 U9251 ( .A1(n9019), .A2(n7606), .B1(n10444), .B2(n5263), .ZN(n7607)
         );
  INV_X1 U9252 ( .A(n7607), .ZN(n7608) );
  OAI21_X1 U9253 ( .B1(n7609), .B2(n10442), .A(n7608), .ZN(P2_U3469) );
  OAI21_X1 U9254 ( .B1(n4575), .B2(n7611), .A(n7610), .ZN(n7612) );
  NAND2_X1 U9255 ( .A1(n7612), .A2(n8329), .ZN(n7618) );
  OR2_X1 U9256 ( .A1(n7613), .A2(n8892), .ZN(n7615) );
  NAND2_X1 U9257 ( .A1(n8568), .A2(n8815), .ZN(n7614) );
  NAND2_X1 U9258 ( .A1(n7615), .A2(n7614), .ZN(n7665) );
  NOR2_X1 U9259 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5309), .ZN(n8584) );
  NOR2_X1 U9260 ( .A1(n8341), .A2(n7672), .ZN(n7616) );
  AOI211_X1 U9261 ( .C1(n8287), .C2(n7665), .A(n8584), .B(n7616), .ZN(n7617)
         );
  OAI211_X1 U9262 ( .C1(n10429), .C2(n8335), .A(n7618), .B(n7617), .ZN(
        P2_U3233) );
  NAND2_X1 U9263 ( .A1(n7619), .A2(n8436), .ZN(n7620) );
  AND2_X1 U9264 ( .A1(n7621), .A2(n7620), .ZN(n7714) );
  INV_X1 U9265 ( .A(n7882), .ZN(n8845) );
  NAND3_X1 U9266 ( .A1(n7622), .A2(n4942), .A3(n8433), .ZN(n7623) );
  AOI21_X1 U9267 ( .B1(n7624), .B2(n7623), .A(n8889), .ZN(n7627) );
  OAI22_X1 U9268 ( .A1(n7625), .A2(n8892), .B1(n7742), .B2(n8890), .ZN(n7626)
         );
  AOI211_X1 U9269 ( .C1(n7714), .C2(n8845), .A(n7627), .B(n7626), .ZN(n7719)
         );
  AND2_X1 U9270 ( .A1(n7628), .A2(n7631), .ZN(n7629) );
  OR2_X1 U9271 ( .A1(n7629), .A2(n4573), .ZN(n7716) );
  INV_X1 U9272 ( .A(n8874), .ZN(n10363) );
  AOI22_X1 U9273 ( .A1(n8897), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7630), .B2(
        n8848), .ZN(n7633) );
  NAND2_X1 U9274 ( .A1(n8885), .A2(n7631), .ZN(n7632) );
  OAI211_X1 U9275 ( .C1(n7716), .C2(n10363), .A(n7633), .B(n7632), .ZN(n7634)
         );
  AOI21_X1 U9276 ( .B1(n7714), .B2(n8854), .A(n7634), .ZN(n7635) );
  OAI21_X1 U9277 ( .B1(n7719), .B2(n8897), .A(n7635), .ZN(P2_U3288) );
  XNOR2_X1 U9278 ( .A(n7638), .B(n7637), .ZN(n7639) );
  XNOR2_X1 U9279 ( .A(n7636), .B(n7639), .ZN(n7646) );
  NOR2_X1 U9280 ( .A1(n9146), .A2(n10316), .ZN(n7645) );
  AOI21_X1 U9281 ( .B1(n9152), .B2(n9162), .A(n7640), .ZN(n7642) );
  NAND2_X1 U9282 ( .A1(n10090), .A2(n9163), .ZN(n7641) );
  OAI211_X1 U9283 ( .C1(n10106), .C2(n7643), .A(n7642), .B(n7641), .ZN(n7644)
         );
  AOI211_X1 U9284 ( .C1(n7646), .C2(n10101), .A(n7645), .B(n7644), .ZN(n7647)
         );
  INV_X1 U9285 ( .A(n7647), .ZN(P1_U3219) );
  XNOR2_X1 U9286 ( .A(n7779), .B(n7772), .ZN(n7650) );
  OAI21_X1 U9287 ( .B1(n7650), .B2(n8871), .A(n7781), .ZN(n7658) );
  AOI21_X1 U9288 ( .B1(n7652), .B2(n8977), .A(n7651), .ZN(n7771) );
  XNOR2_X1 U9289 ( .A(n7771), .B(n7780), .ZN(n7653) );
  NAND2_X1 U9290 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7653), .ZN(n7773) );
  OAI211_X1 U9291 ( .C1(n7653), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10342), .B(
        n7773), .ZN(n7656) );
  NOR2_X1 U9292 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8340), .ZN(n7654) );
  AOI21_X1 U9293 ( .B1(n10350), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7654), .ZN(
        n7655) );
  OAI211_X1 U9294 ( .C1(n10346), .C2(n7780), .A(n7656), .B(n7655), .ZN(n7657)
         );
  AOI21_X1 U9295 ( .B1(n10343), .B2(n7658), .A(n7657), .ZN(n7659) );
  INV_X1 U9296 ( .A(n7659), .ZN(P2_U3260) );
  INV_X1 U9297 ( .A(n7660), .ZN(n7662) );
  OAI222_X1 U9298 ( .A1(n9626), .A2(n9929), .B1(n9624), .B2(n7662), .C1(
        P1_U3084), .C2(n5786), .ZN(P1_U3331) );
  OAI222_X1 U9299 ( .A1(n7930), .A2(n7663), .B1(n6706), .B2(n7662), .C1(
        P2_U3152), .C2(n7661), .ZN(P2_U3336) );
  XOR2_X1 U9300 ( .A(n7664), .B(n8443), .Z(n7667) );
  INV_X1 U9301 ( .A(n7665), .ZN(n7666) );
  OAI21_X1 U9302 ( .B1(n7667), .B2(n8889), .A(n7666), .ZN(n10431) );
  INV_X1 U9303 ( .A(n10431), .ZN(n7679) );
  INV_X1 U9304 ( .A(n8443), .ZN(n7669) );
  OAI21_X1 U9305 ( .B1(n7670), .B2(n7669), .A(n7668), .ZN(n10433) );
  NOR2_X1 U9306 ( .A1(n4573), .A2(n10429), .ZN(n7671) );
  OR2_X1 U9307 ( .A1(n7745), .A2(n7671), .ZN(n10430) );
  INV_X1 U9308 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7673) );
  OAI22_X1 U9309 ( .A1(n7188), .A2(n7673), .B1(n7672), .B2(n10358), .ZN(n7674)
         );
  AOI21_X1 U9310 ( .B1(n8885), .B2(n7675), .A(n7674), .ZN(n7676) );
  OAI21_X1 U9311 ( .B1(n10430), .B2(n10363), .A(n7676), .ZN(n7677) );
  AOI21_X1 U9312 ( .B1(n10433), .B2(n10366), .A(n7677), .ZN(n7678) );
  OAI21_X1 U9313 ( .B1(n7679), .B2(n8897), .A(n7678), .ZN(P2_U3287) );
  INV_X1 U9314 ( .A(n7680), .ZN(n7684) );
  NOR2_X1 U9315 ( .A1(n7681), .A2(P1_U3084), .ZN(n8250) );
  AOI21_X1 U9316 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9617), .A(n8250), .ZN(
        n7682) );
  OAI21_X1 U9317 ( .B1(n7684), .B2(n9624), .A(n7682), .ZN(P1_U3330) );
  NAND2_X1 U9318 ( .A1(n9030), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7683) );
  OAI211_X1 U9319 ( .C1(n7684), .C2(n6706), .A(n7683), .B(n8557), .ZN(P2_U3335) );
  NAND2_X1 U9320 ( .A1(n10262), .A2(n7685), .ZN(n7686) );
  NAND2_X1 U9321 ( .A1(n7687), .A2(n7686), .ZN(n10261) );
  AND2_X1 U9322 ( .A1(n10277), .A2(n9162), .ZN(n7689) );
  OR2_X1 U9323 ( .A1(n10277), .A2(n9162), .ZN(n7688) );
  NAND2_X1 U9324 ( .A1(n7831), .A2(n10130), .ZN(n8015) );
  NAND2_X1 U9325 ( .A1(n8147), .A2(n8015), .ZN(n8110) );
  XNOR2_X1 U9326 ( .A(n7830), .B(n8110), .ZN(n10052) );
  NAND2_X1 U9327 ( .A1(n7690), .A2(n8167), .ZN(n10269) );
  INV_X1 U9328 ( .A(n9162), .ZN(n7691) );
  OR2_X1 U9329 ( .A1(n7691), .A2(n10277), .ZN(n8014) );
  NAND2_X1 U9330 ( .A1(n7691), .A2(n10277), .ZN(n8012) );
  NAND2_X1 U9331 ( .A1(n10269), .A2(n10268), .ZN(n10267) );
  NAND2_X1 U9332 ( .A1(n10267), .A2(n8014), .ZN(n7693) );
  INV_X1 U9333 ( .A(n8110), .ZN(n7692) );
  NAND2_X1 U9334 ( .A1(n7693), .A2(n7692), .ZN(n7834) );
  OAI211_X1 U9335 ( .C1(n7693), .C2(n7692), .A(n7834), .B(n10266), .ZN(n7695)
         );
  AOI22_X1 U9336 ( .A1(n10263), .A2(n9162), .B1(n10264), .B2(n9161), .ZN(n7694) );
  NAND2_X1 U9337 ( .A1(n7695), .A2(n7694), .ZN(n7696) );
  AOI21_X1 U9338 ( .B1(n10052), .B2(n7697), .A(n7696), .ZN(n10054) );
  INV_X1 U9339 ( .A(n10277), .ZN(n10324) );
  NAND2_X1 U9340 ( .A1(n10280), .A2(n10324), .ZN(n10279) );
  AOI21_X1 U9341 ( .B1(n10279), .B2(n7831), .A(n10325), .ZN(n7698) );
  NAND2_X1 U9342 ( .A1(n7698), .A2(n10139), .ZN(n10050) );
  INV_X1 U9343 ( .A(n7699), .ZN(n7733) );
  AOI22_X1 U9344 ( .A1(n4483), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7733), .B2(
        n10275), .ZN(n7701) );
  NAND2_X1 U9345 ( .A1(n10276), .A2(n7831), .ZN(n7700) );
  OAI211_X1 U9346 ( .C1(n10050), .C2(n9387), .A(n7701), .B(n7700), .ZN(n7702)
         );
  AOI21_X1 U9347 ( .B1(n10052), .B2(n10283), .A(n7702), .ZN(n7703) );
  OAI21_X1 U9348 ( .B1(n10054), .B2(n4483), .A(n7703), .ZN(P1_U3281) );
  INV_X1 U9349 ( .A(n7704), .ZN(n7705) );
  AOI21_X1 U9350 ( .B1(n7707), .B2(n7706), .A(n7705), .ZN(n7713) );
  NOR2_X1 U9351 ( .A1(n10092), .A2(n10130), .ZN(n7708) );
  AOI211_X1 U9352 ( .C1(n10090), .C2(n10262), .A(n7709), .B(n7708), .ZN(n7710)
         );
  OAI21_X1 U9353 ( .B1(n10106), .B2(n10273), .A(n7710), .ZN(n7711) );
  AOI21_X1 U9354 ( .B1(n10095), .B2(n10277), .A(n7711), .ZN(n7712) );
  OAI21_X1 U9355 ( .B1(n7713), .B2(n9156), .A(n7712), .ZN(P1_U3229) );
  INV_X1 U9356 ( .A(n7714), .ZN(n7720) );
  OAI22_X1 U9357 ( .A1(n7716), .A2(n10436), .B1(n7715), .B2(n10434), .ZN(n7717) );
  INV_X1 U9358 ( .A(n7717), .ZN(n7718) );
  OAI211_X1 U9359 ( .C1(n10077), .C2(n7720), .A(n7719), .B(n7718), .ZN(n7722)
         );
  NAND2_X1 U9360 ( .A1(n7722), .A2(n10452), .ZN(n7721) );
  OAI21_X1 U9361 ( .B1(n10452), .B2(n7032), .A(n7721), .ZN(P2_U3528) );
  NAND2_X1 U9362 ( .A1(n7722), .A2(n10444), .ZN(n7723) );
  OAI21_X1 U9363 ( .B1(n10444), .B2(n5293), .A(n7723), .ZN(P2_U3475) );
  NAND2_X1 U9364 ( .A1(n7726), .A2(n7725), .ZN(n7727) );
  XNOR2_X1 U9365 ( .A(n7724), .B(n7727), .ZN(n7735) );
  INV_X1 U9366 ( .A(n10067), .ZN(n7728) );
  NAND2_X1 U9367 ( .A1(n7831), .A2(n10164), .ZN(n10049) );
  NOR2_X1 U9368 ( .A1(n7728), .A2(n10049), .ZN(n7732) );
  AOI21_X1 U9369 ( .B1(n10090), .B2(n9162), .A(n7729), .ZN(n7730) );
  OAI21_X1 U9370 ( .B1(n10060), .B2(n10092), .A(n7730), .ZN(n7731) );
  AOI211_X1 U9371 ( .C1(n7733), .C2(n9143), .A(n7732), .B(n7731), .ZN(n7734)
         );
  OAI21_X1 U9372 ( .B1(n7735), .B2(n9156), .A(n7734), .ZN(P1_U3215) );
  NAND2_X1 U9373 ( .A1(n7736), .A2(n8444), .ZN(n7737) );
  INV_X1 U9374 ( .A(n8444), .ZN(n7738) );
  NAND3_X1 U9375 ( .A1(n7739), .A2(n7738), .A3(n8440), .ZN(n7740) );
  AOI21_X1 U9376 ( .B1(n7741), .B2(n7740), .A(n8889), .ZN(n7744) );
  OAI22_X1 U9377 ( .A1(n7742), .A2(n8892), .B1(n7793), .B2(n8890), .ZN(n7743)
         );
  AOI211_X1 U9378 ( .C1(n8980), .C2(n8845), .A(n7744), .B(n7743), .ZN(n8985)
         );
  INV_X1 U9379 ( .A(n7745), .ZN(n7747) );
  INV_X1 U9380 ( .A(n7746), .ZN(n7762) );
  AOI21_X1 U9381 ( .B1(n8981), .B2(n7747), .A(n7762), .ZN(n8983) );
  NOR2_X1 U9382 ( .A1(n10362), .A2(n7748), .ZN(n7752) );
  INV_X1 U9383 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7750) );
  OAI22_X1 U9384 ( .A1(n7188), .A2(n7750), .B1(n7749), .B2(n10358), .ZN(n7751)
         );
  AOI211_X1 U9385 ( .C1(n8983), .C2(n8874), .A(n7752), .B(n7751), .ZN(n7754)
         );
  NAND2_X1 U9386 ( .A1(n8980), .A2(n8854), .ZN(n7753) );
  OAI211_X1 U9387 ( .C1(n8985), .C2(n8877), .A(n7754), .B(n7753), .ZN(P2_U3286) );
  NAND2_X1 U9388 ( .A1(n7756), .A2(n7755), .ZN(n7757) );
  XNOR2_X1 U9389 ( .A(n7757), .B(n5349), .ZN(n10441) );
  INV_X1 U9390 ( .A(n10441), .ZN(n7770) );
  XNOR2_X1 U9391 ( .A(n7759), .B(n7758), .ZN(n7760) );
  OAI222_X1 U9392 ( .A1(n8890), .A2(n7878), .B1(n8892), .B2(n7761), .C1(n7760), 
        .C2(n8889), .ZN(n10438) );
  INV_X1 U9393 ( .A(n7766), .ZN(n10435) );
  OAI21_X1 U9394 ( .B1(n7762), .B2(n10435), .A(n7801), .ZN(n10437) );
  OAI22_X1 U9395 ( .A1(n7188), .A2(n7764), .B1(n7763), .B2(n10358), .ZN(n7765)
         );
  AOI21_X1 U9396 ( .B1(n8885), .B2(n7766), .A(n7765), .ZN(n7767) );
  OAI21_X1 U9397 ( .B1(n10437), .B2(n10363), .A(n7767), .ZN(n7768) );
  AOI21_X1 U9398 ( .B1(n10438), .B2(n7188), .A(n7768), .ZN(n7769) );
  OAI21_X1 U9399 ( .B1(n8809), .B2(n7770), .A(n7769), .ZN(P2_U3285) );
  NAND2_X1 U9400 ( .A1(n7772), .A2(n7771), .ZN(n7774) );
  NAND2_X1 U9401 ( .A1(n7774), .A2(n7773), .ZN(n7777) );
  XNOR2_X1 U9402 ( .A(n7811), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7776) );
  INV_X1 U9403 ( .A(n7813), .ZN(n7775) );
  AOI21_X1 U9404 ( .B1(n7777), .B2(n7776), .A(n7775), .ZN(n7788) );
  AND2_X1 U9405 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8298) );
  AOI21_X1 U9406 ( .B1(n10350), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8298), .ZN(
        n7778) );
  INV_X1 U9407 ( .A(n7778), .ZN(n7786) );
  NAND2_X1 U9408 ( .A1(n7780), .A2(n7779), .ZN(n7782) );
  XNOR2_X1 U9409 ( .A(n7811), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n7783) );
  AOI211_X1 U9410 ( .C1(n7784), .C2(n7783), .A(n10347), .B(n4529), .ZN(n7785)
         );
  AOI211_X1 U9411 ( .C1(n10042), .C2(n7811), .A(n7786), .B(n7785), .ZN(n7787)
         );
  OAI21_X1 U9412 ( .B1(n7788), .B2(n10344), .A(n7787), .ZN(P2_U3261) );
  INV_X1 U9413 ( .A(n7789), .ZN(n7822) );
  OAI222_X1 U9414 ( .A1(P2_U3152), .A2(n7791), .B1(n6706), .B2(n7822), .C1(
        n7790), .C2(n7930), .ZN(P2_U3334) );
  AOI21_X1 U9415 ( .B1(n7792), .B2(n8372), .A(n8889), .ZN(n7796) );
  OAI22_X1 U9416 ( .A1(n7793), .A2(n8892), .B1(n8893), .B2(n8890), .ZN(n7794)
         );
  AOI21_X1 U9417 ( .B1(n7796), .B2(n7795), .A(n7794), .ZN(n7915) );
  XNOR2_X1 U9418 ( .A(n7798), .B(n7797), .ZN(n7918) );
  NAND2_X1 U9419 ( .A1(n7918), .A2(n10366), .ZN(n7807) );
  OAI22_X1 U9420 ( .A1(n7188), .A2(n7800), .B1(n7799), .B2(n10358), .ZN(n7804)
         );
  INV_X1 U9421 ( .A(n7801), .ZN(n7802) );
  INV_X1 U9422 ( .A(n7805), .ZN(n7922) );
  NOR2_X1 U9423 ( .A1(n7916), .A2(n10363), .ZN(n7803) );
  AOI211_X1 U9424 ( .C1(n8885), .C2(n7805), .A(n7804), .B(n7803), .ZN(n7806)
         );
  OAI211_X1 U9425 ( .C1(n8897), .C2(n7915), .A(n7807), .B(n7806), .ZN(P2_U3284) );
  NAND2_X1 U9426 ( .A1(n8594), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7808) );
  OAI21_X1 U9427 ( .B1(n8594), .B2(P2_REG2_REG_17__SCAN_IN), .A(n7808), .ZN(
        n7809) );
  NOR2_X1 U9428 ( .A1(n7810), .A2(n7809), .ZN(n8593) );
  AOI211_X1 U9429 ( .C1(n7810), .C2(n7809), .A(n10347), .B(n8593), .ZN(n7820)
         );
  OR2_X1 U9430 ( .A1(n7811), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7812) );
  AND2_X1 U9431 ( .A1(n7813), .A2(n7812), .ZN(n7815) );
  INV_X1 U9432 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8959) );
  XNOR2_X1 U9433 ( .A(n8594), .B(n8959), .ZN(n7814) );
  NAND3_X1 U9434 ( .A1(n7813), .A2(n7814), .A3(n7812), .ZN(n8599) );
  OAI211_X1 U9435 ( .C1(n7815), .C2(n7814), .A(n10342), .B(n8599), .ZN(n7818)
         );
  NOR2_X1 U9436 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5441), .ZN(n7816) );
  AOI21_X1 U9437 ( .B1(n10350), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n7816), .ZN(
        n7817) );
  OAI211_X1 U9438 ( .C1(n10346), .C2(n8600), .A(n7818), .B(n7817), .ZN(n7819)
         );
  OR2_X1 U9439 ( .A1(n7820), .A2(n7819), .ZN(P2_U3262) );
  OAI222_X1 U9440 ( .A1(P1_U3084), .A2(n7823), .B1(n9624), .B2(n7822), .C1(
        n7821), .C2(n9626), .ZN(P1_U3329) );
  INV_X1 U9441 ( .A(n7824), .ZN(n7828) );
  INV_X1 U9442 ( .A(n7825), .ZN(n7826) );
  OAI222_X1 U9443 ( .A1(n9626), .A2(n9921), .B1(n9624), .B2(n7828), .C1(
        P1_U3084), .C2(n7826), .ZN(P1_U3328) );
  OAI222_X1 U9444 ( .A1(n7930), .A2(n7829), .B1(n6706), .B2(n7828), .C1(
        P2_U3152), .C2(n7827), .ZN(P2_U3333) );
  XNOR2_X1 U9445 ( .A(n10163), .B(n9161), .ZN(n10131) );
  OR2_X1 U9446 ( .A1(n7893), .A2(n10127), .ZN(n8017) );
  NAND2_X1 U9447 ( .A1(n7893), .A2(n10127), .ZN(n8020) );
  NAND2_X1 U9448 ( .A1(n8017), .A2(n8020), .ZN(n8111) );
  OR2_X1 U9449 ( .A1(n7832), .A2(n8111), .ZN(n7833) );
  NAND2_X1 U9450 ( .A1(n10111), .A2(n7833), .ZN(n10158) );
  NAND2_X1 U9451 ( .A1(n10163), .A2(n10060), .ZN(n8016) );
  NAND2_X1 U9452 ( .A1(n10126), .A2(n8016), .ZN(n7897) );
  OR2_X1 U9453 ( .A1(n10163), .A2(n10060), .ZN(n7896) );
  NAND2_X1 U9454 ( .A1(n7897), .A2(n7896), .ZN(n7835) );
  XNOR2_X1 U9455 ( .A(n7835), .B(n8111), .ZN(n7837) );
  OAI22_X1 U9456 ( .A1(n10060), .A2(n10129), .B1(n10128), .B2(n10059), .ZN(
        n7836) );
  AOI21_X1 U9457 ( .B1(n7837), .B2(n10266), .A(n7836), .ZN(n7838) );
  OAI21_X1 U9458 ( .B1(n10158), .B2(n10272), .A(n7838), .ZN(n10162) );
  NAND2_X1 U9459 ( .A1(n10162), .A2(n9508), .ZN(n7844) );
  NOR2_X1 U9460 ( .A1(n10139), .A2(n10163), .ZN(n10138) );
  INV_X1 U9461 ( .A(n10138), .ZN(n7839) );
  INV_X1 U9462 ( .A(n7893), .ZN(n10066) );
  AOI211_X1 U9463 ( .C1(n7893), .C2(n7839), .A(n10325), .B(n10119), .ZN(n10159) );
  NOR2_X1 U9464 ( .A1(n10066), .A2(n9484), .ZN(n7842) );
  OAI22_X1 U9465 ( .A1(n9508), .A2(n7840), .B1(n10071), .B2(n9505), .ZN(n7841)
         );
  AOI211_X1 U9466 ( .C1(n10159), .C2(n9490), .A(n7842), .B(n7841), .ZN(n7843)
         );
  OAI211_X1 U9467 ( .C1(n10158), .C2(n7845), .A(n7844), .B(n7843), .ZN(
        P1_U3279) );
  AOI21_X1 U9468 ( .B1(n7848), .B2(n7847), .A(n6456), .ZN(n7853) );
  OAI21_X1 U9469 ( .B1(n8341), .B2(n8883), .A(n7849), .ZN(n7851) );
  OAI22_X1 U9470 ( .A1(n8893), .A2(n8343), .B1(n8342), .B2(n8891), .ZN(n7850)
         );
  AOI211_X1 U9471 ( .C1(n8886), .C2(n8346), .A(n7851), .B(n7850), .ZN(n7852)
         );
  OAI21_X1 U9472 ( .B1(n7853), .B2(n8348), .A(n7852), .ZN(P2_U3217) );
  INV_X1 U9473 ( .A(n10127), .ZN(n9160) );
  AOI21_X1 U9474 ( .B1(n9152), .B2(n9160), .A(n7854), .ZN(n7856) );
  NAND2_X1 U9475 ( .A1(n10090), .A2(n10265), .ZN(n7855) );
  OAI211_X1 U9476 ( .C1(n10106), .C2(n10136), .A(n7856), .B(n7855), .ZN(n7862)
         );
  INV_X1 U9477 ( .A(n7857), .ZN(n7858) );
  AOI211_X1 U9478 ( .C1(n7860), .C2(n7859), .A(n9156), .B(n7858), .ZN(n7861)
         );
  AOI211_X1 U9479 ( .C1(n10095), .C2(n10163), .A(n7862), .B(n7861), .ZN(n7863)
         );
  INV_X1 U9480 ( .A(n7863), .ZN(P1_U3234) );
  XNOR2_X1 U9481 ( .A(n7866), .B(n7865), .ZN(n7867) );
  XNOR2_X1 U9482 ( .A(n7864), .B(n7867), .ZN(n7872) );
  AND2_X1 U9483 ( .A1(n10122), .A2(n10164), .ZN(n10152) );
  AND2_X1 U9484 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10186) );
  NOR2_X1 U9485 ( .A1(n10061), .A2(n10127), .ZN(n7868) );
  AOI211_X1 U9486 ( .C1(n9152), .C2(n9217), .A(n10186), .B(n7868), .ZN(n7869)
         );
  OAI21_X1 U9487 ( .B1(n10106), .B2(n10117), .A(n7869), .ZN(n7870) );
  AOI21_X1 U9488 ( .B1(n10067), .B2(n10152), .A(n7870), .ZN(n7871) );
  OAI21_X1 U9489 ( .B1(n7872), .B2(n9156), .A(n7871), .ZN(P1_U3232) );
  NAND2_X1 U9490 ( .A1(n7873), .A2(n8464), .ZN(n7874) );
  NAND2_X1 U9491 ( .A1(n7875), .A2(n7874), .ZN(n10078) );
  INV_X1 U9492 ( .A(n8854), .ZN(n7892) );
  OAI21_X1 U9493 ( .B1(n7877), .B2(n8464), .A(n7876), .ZN(n7880) );
  OAI22_X1 U9494 ( .A1(n7878), .A2(n8892), .B1(n8860), .B2(n8890), .ZN(n7879)
         );
  AOI21_X1 U9495 ( .B1(n7880), .B2(n10357), .A(n7879), .ZN(n7881) );
  OAI21_X1 U9496 ( .B1(n10078), .B2(n7882), .A(n7881), .ZN(n10082) );
  NAND2_X1 U9497 ( .A1(n10082), .A2(n7188), .ZN(n7891) );
  OAI22_X1 U9498 ( .A1(n7188), .A2(n7884), .B1(n7883), .B2(n10358), .ZN(n7889)
         );
  INV_X1 U9499 ( .A(n8881), .ZN(n7887) );
  NAND2_X1 U9500 ( .A1(n7885), .A2(n10079), .ZN(n7886) );
  NAND2_X1 U9501 ( .A1(n7887), .A2(n7886), .ZN(n10081) );
  NOR2_X1 U9502 ( .A1(n10081), .A2(n10363), .ZN(n7888) );
  AOI211_X1 U9503 ( .C1(n8885), .C2(n10079), .A(n7889), .B(n7888), .ZN(n7890)
         );
  OAI211_X1 U9504 ( .C1(n10078), .C2(n7892), .A(n7891), .B(n7890), .ZN(
        P2_U3283) );
  NAND2_X1 U9505 ( .A1(n7893), .A2(n9160), .ZN(n10110) );
  NAND2_X1 U9506 ( .A1(n10122), .A2(n10089), .ZN(n7894) );
  AND2_X1 U9507 ( .A1(n10110), .A2(n7894), .ZN(n7895) );
  AOI21_X1 U9508 ( .B1(n10111), .B2(n7895), .A(n4492), .ZN(n9219) );
  OR2_X1 U9509 ( .A1(n10096), .A2(n10109), .ZN(n9241) );
  NAND2_X1 U9510 ( .A1(n10096), .A2(n10109), .ZN(n8145) );
  NAND2_X1 U9511 ( .A1(n9241), .A2(n8145), .ZN(n7899) );
  INV_X1 U9512 ( .A(n7899), .ZN(n8114) );
  XNOR2_X1 U9513 ( .A(n9219), .B(n8114), .ZN(n10151) );
  INV_X1 U9514 ( .A(n10151), .ZN(n7911) );
  AND2_X1 U9515 ( .A1(n8017), .A2(n7896), .ZN(n8022) );
  NAND2_X1 U9516 ( .A1(n7897), .A2(n8022), .ZN(n7898) );
  NAND2_X1 U9517 ( .A1(n7898), .A2(n8020), .ZN(n10108) );
  OR2_X1 U9518 ( .A1(n10122), .A2(n10059), .ZN(n8019) );
  NAND2_X1 U9519 ( .A1(n10122), .A2(n10059), .ZN(n8151) );
  INV_X1 U9520 ( .A(n8151), .ZN(n8171) );
  NOR2_X1 U9521 ( .A1(n7899), .A2(n8171), .ZN(n7900) );
  NAND2_X1 U9522 ( .A1(n10107), .A2(n7900), .ZN(n9242) );
  NAND2_X1 U9523 ( .A1(n9242), .A2(n10266), .ZN(n7903) );
  AOI21_X1 U9524 ( .B1(n10107), .B2(n8151), .A(n8114), .ZN(n7902) );
  AOI22_X1 U9525 ( .A1(n9220), .A2(n10264), .B1(n10263), .B2(n10089), .ZN(
        n7901) );
  OAI21_X1 U9526 ( .B1(n7903), .B2(n7902), .A(n7901), .ZN(n10150) );
  INV_X1 U9527 ( .A(n10122), .ZN(n7904) );
  NAND2_X1 U9528 ( .A1(n10119), .A2(n7904), .ZN(n7905) );
  INV_X1 U9529 ( .A(n7905), .ZN(n10120) );
  INV_X1 U9530 ( .A(n10096), .ZN(n10148) );
  OAI211_X1 U9531 ( .C1(n10120), .C2(n10148), .A(n10165), .B(n9502), .ZN(
        n10147) );
  OAI22_X1 U9532 ( .A1(n9508), .A2(n7906), .B1(n10105), .B2(n9505), .ZN(n7907)
         );
  AOI21_X1 U9533 ( .B1(n10096), .B2(n10276), .A(n7907), .ZN(n7908) );
  OAI21_X1 U9534 ( .B1(n10147), .B2(n9387), .A(n7908), .ZN(n7909) );
  AOI21_X1 U9535 ( .B1(n10150), .B2(n9508), .A(n7909), .ZN(n7910) );
  OAI21_X1 U9536 ( .B1(n7911), .B2(n9481), .A(n7910), .ZN(P1_U3277) );
  INV_X1 U9537 ( .A(n7912), .ZN(n7926) );
  OAI222_X1 U9538 ( .A1(P2_U3152), .A2(n7914), .B1(n6706), .B2(n7926), .C1(
        n7913), .C2(n7930), .ZN(P2_U3332) );
  OAI21_X1 U9539 ( .B1(n10436), .B2(n7916), .A(n7915), .ZN(n7917) );
  AOI21_X1 U9540 ( .B1(n7918), .B2(n10440), .A(n7917), .ZN(n7920) );
  MUX2_X1 U9541 ( .A(n5362), .B(n7920), .S(n10452), .Z(n7919) );
  OAI21_X1 U9542 ( .B1(n7922), .B2(n8979), .A(n7919), .ZN(P2_U3532) );
  MUX2_X1 U9543 ( .A(n5365), .B(n7920), .S(n10444), .Z(n7921) );
  OAI21_X1 U9544 ( .B1(n7922), .B2(n9019), .A(n7921), .ZN(P2_U3487) );
  NAND2_X1 U9545 ( .A1(n7927), .A2(n7923), .ZN(n7925) );
  OAI211_X1 U9546 ( .C1(n9622), .C2(n9777), .A(n7925), .B(n7924), .ZN(P1_U3326) );
  OAI222_X1 U9547 ( .A1(P1_U3084), .A2(n6339), .B1(n9624), .B2(n7926), .C1(
        n9978), .C2(n9622), .ZN(P1_U3327) );
  INV_X1 U9548 ( .A(n7927), .ZN(n7928) );
  OAI222_X1 U9549 ( .A1(n7930), .A2(n7929), .B1(n6706), .B2(n7928), .C1(
        P2_U3152), .C2(n8552), .ZN(P2_U3331) );
  INV_X1 U9550 ( .A(n7931), .ZN(n7936) );
  AOI21_X1 U9551 ( .B1(n9617), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n7932), .ZN(
        n7933) );
  OAI21_X1 U9552 ( .B1(n7936), .B2(n9624), .A(n7933), .ZN(P1_U3325) );
  AOI21_X1 U9553 ( .B1(n9030), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n7934), .ZN(
        n7935) );
  OAI21_X1 U9554 ( .B1(n7936), .B2(n6706), .A(n7935), .ZN(P2_U3330) );
  MUX2_X1 U9555 ( .A(n7937), .B(P1_REG2_REG_4__SCAN_IN), .S(n4483), .Z(n7946)
         );
  NAND2_X1 U9556 ( .A1(n7938), .A2(n10283), .ZN(n7943) );
  OAI22_X1 U9557 ( .A1(n9484), .A2(n7940), .B1(n7939), .B2(n9505), .ZN(n7941)
         );
  INV_X1 U9558 ( .A(n7941), .ZN(n7942) );
  OAI211_X1 U9559 ( .C1(n9512), .C2(n7944), .A(n7943), .B(n7942), .ZN(n7945)
         );
  OR2_X1 U9560 ( .A1(n7946), .A2(n7945), .ZN(P1_U3287) );
  NAND2_X1 U9561 ( .A1(n7947), .A2(n10366), .ZN(n7956) );
  INV_X1 U9562 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n7948) );
  OAI22_X1 U9563 ( .A1(n7949), .A2(n10358), .B1(n7948), .B2(n7188), .ZN(n7953)
         );
  NOR2_X1 U9564 ( .A1(n7951), .A2(n7950), .ZN(n7952) );
  AOI211_X1 U9565 ( .C1(n8885), .C2(n7954), .A(n7953), .B(n7952), .ZN(n7955)
         );
  OAI211_X1 U9566 ( .C1(n7957), .C2(n8877), .A(n7956), .B(n7955), .ZN(P2_U3267) );
  INV_X1 U9567 ( .A(n7958), .ZN(n7966) );
  NAND2_X1 U9568 ( .A1(n7959), .A2(n8830), .ZN(n7962) );
  AOI22_X1 U9569 ( .A1(n7960), .A2(n8848), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n8897), .ZN(n7961) );
  OAI211_X1 U9570 ( .C1(n4840), .C2(n10362), .A(n7962), .B(n7961), .ZN(n7963)
         );
  AOI21_X1 U9571 ( .B1(n7964), .B2(n7188), .A(n7963), .ZN(n7965) );
  OAI21_X1 U9572 ( .B1(n7966), .B2(n8809), .A(n7965), .ZN(P2_U3269) );
  XNOR2_X1 U9573 ( .A(n7968), .B(n7967), .ZN(n7972) );
  OAI22_X1 U9574 ( .A1(n8341), .A2(n8796), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9781), .ZN(n7970) );
  OAI22_X1 U9575 ( .A1(n8842), .A2(n8343), .B1(n8342), .B2(n8321), .ZN(n7969)
         );
  AOI211_X1 U9576 ( .C1(n8950), .C2(n8346), .A(n7970), .B(n7969), .ZN(n7971)
         );
  OAI21_X1 U9577 ( .B1(n7972), .B2(n8348), .A(n7971), .ZN(P2_U3240) );
  NOR2_X1 U9578 ( .A1(n7975), .A2(SI_29_), .ZN(n7973) );
  NAND2_X1 U9579 ( .A1(n7975), .A2(SI_29_), .ZN(n7976) );
  MUX2_X1 U9580 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7982), .Z(n7978) );
  NAND2_X1 U9581 ( .A1(n7977), .A2(SI_30_), .ZN(n7981) );
  NAND2_X1 U9582 ( .A1(n7979), .A2(n7978), .ZN(n7980) );
  NAND2_X1 U9583 ( .A1(n7981), .A2(n7980), .ZN(n7986) );
  MUX2_X1 U9584 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7982), .Z(n7984) );
  INV_X1 U9585 ( .A(SI_31_), .ZN(n7983) );
  XNOR2_X1 U9586 ( .A(n7984), .B(n7983), .ZN(n7985) );
  NAND2_X1 U9587 ( .A1(n6265), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7987) );
  NAND2_X1 U9588 ( .A1(n9516), .A2(n9209), .ZN(n8239) );
  INV_X1 U9589 ( .A(n8239), .ZN(n8123) );
  NOR2_X1 U9590 ( .A1(n8123), .A2(n8039), .ZN(n8085) );
  NAND2_X1 U9591 ( .A1(n9029), .A2(n8072), .ZN(n7990) );
  NAND2_X1 U9592 ( .A1(n6265), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7989) );
  INV_X1 U9593 ( .A(n9294), .ZN(n8092) );
  INV_X1 U9594 ( .A(n8127), .ZN(n8070) );
  INV_X1 U9595 ( .A(n9375), .ZN(n9349) );
  OR2_X1 U9596 ( .A1(n9550), .A2(n9349), .ZN(n9257) );
  NAND2_X1 U9597 ( .A1(n8094), .A2(n9257), .ZN(n8142) );
  NAND2_X1 U9598 ( .A1(n8142), .A2(n9258), .ZN(n7992) );
  NAND2_X1 U9599 ( .A1(n9540), .A2(n9350), .ZN(n9262) );
  NAND2_X1 U9600 ( .A1(n9550), .A2(n9349), .ZN(n8095) );
  NAND2_X1 U9601 ( .A1(n9258), .A2(n8095), .ZN(n8043) );
  NAND2_X1 U9602 ( .A1(n8043), .A2(n8094), .ZN(n7993) );
  AND2_X1 U9603 ( .A1(n9262), .A2(n7993), .ZN(n8133) );
  NAND2_X1 U9604 ( .A1(n8133), .A2(n8039), .ZN(n7994) );
  NAND2_X1 U9605 ( .A1(n7995), .A2(n7994), .ZN(n8048) );
  INV_X1 U9606 ( .A(n9421), .ZN(n9454) );
  OR2_X1 U9607 ( .A1(n9573), .A2(n9454), .ZN(n8135) );
  OR2_X1 U9608 ( .A1(n9578), .A2(n9437), .ZN(n8099) );
  AND2_X1 U9609 ( .A1(n8135), .A2(n8099), .ZN(n8035) );
  NAND2_X1 U9610 ( .A1(n9578), .A2(n9437), .ZN(n9249) );
  AND2_X1 U9611 ( .A1(n9581), .A2(n9478), .ZN(n9247) );
  INV_X1 U9612 ( .A(n9247), .ZN(n8030) );
  AND2_X1 U9613 ( .A1(n9249), .A2(n8030), .ZN(n7996) );
  OR2_X1 U9614 ( .A1(n9581), .A2(n9478), .ZN(n9450) );
  AND2_X1 U9615 ( .A1(n8099), .A2(n9450), .ZN(n9248) );
  MUX2_X1 U9616 ( .A(n7996), .B(n9248), .S(n8061), .Z(n8033) );
  NAND2_X1 U9617 ( .A1(n8101), .A2(n8157), .ZN(n7998) );
  NOR2_X1 U9618 ( .A1(n8003), .A2(n8002), .ZN(n8107) );
  NAND2_X1 U9619 ( .A1(n8006), .A2(n8161), .ZN(n8004) );
  NAND2_X1 U9620 ( .A1(n8004), .A2(n8225), .ZN(n8008) );
  NAND2_X1 U9621 ( .A1(n8225), .A2(n8005), .ZN(n8163) );
  NAND2_X1 U9622 ( .A1(n8163), .A2(n8006), .ZN(n8007) );
  MUX2_X1 U9623 ( .A(n8008), .B(n8007), .S(n8039), .Z(n8009) );
  NAND2_X1 U9624 ( .A1(n8010), .A2(n8009), .ZN(n8013) );
  NAND2_X1 U9625 ( .A1(n8014), .A2(n8167), .ZN(n8011) );
  NAND2_X1 U9626 ( .A1(n8015), .A2(n8012), .ZN(n8148) );
  NAND2_X1 U9627 ( .A1(n8147), .A2(n8014), .ZN(n8169) );
  NAND2_X1 U9628 ( .A1(n8020), .A2(n8016), .ZN(n8149) );
  AND2_X1 U9629 ( .A1(n8149), .A2(n8017), .ZN(n8018) );
  INV_X1 U9630 ( .A(n8020), .ZN(n8021) );
  NOR2_X1 U9631 ( .A1(n8022), .A2(n8021), .ZN(n8170) );
  OR2_X1 U9632 ( .A1(n9510), .A2(n10093), .ZN(n9473) );
  NAND2_X1 U9633 ( .A1(n9510), .A2(n10093), .ZN(n9243) );
  NAND2_X1 U9634 ( .A1(n8023), .A2(n9241), .ZN(n8025) );
  NAND2_X1 U9635 ( .A1(n8176), .A2(n8145), .ZN(n8024) );
  MUX2_X1 U9636 ( .A(n8025), .B(n8024), .S(n8039), .Z(n8026) );
  NAND3_X1 U9637 ( .A1(n8027), .A2(n9497), .A3(n8026), .ZN(n8029) );
  OR2_X1 U9638 ( .A1(n9483), .A2(n9496), .ZN(n8178) );
  NAND2_X1 U9639 ( .A1(n9483), .A2(n9496), .ZN(n9245) );
  MUX2_X1 U9640 ( .A(n9243), .B(n9473), .S(n8061), .Z(n8028) );
  NAND3_X1 U9641 ( .A1(n8029), .A2(n9479), .A3(n8028), .ZN(n8032) );
  MUX2_X1 U9642 ( .A(n8178), .B(n9245), .S(n8061), .Z(n8031) );
  INV_X1 U9643 ( .A(n9226), .ZN(n9438) );
  AND2_X1 U9644 ( .A1(n9566), .A2(n9438), .ZN(n9252) );
  NAND2_X1 U9645 ( .A1(n9573), .A2(n9454), .ZN(n9250) );
  INV_X1 U9646 ( .A(n9250), .ZN(n8185) );
  OR2_X1 U9647 ( .A1(n9252), .A2(n8185), .ZN(n8034) );
  AND2_X1 U9648 ( .A1(n9250), .A2(n9249), .ZN(n8134) );
  AND2_X1 U9649 ( .A1(n9418), .A2(n9226), .ZN(n9253) );
  INV_X1 U9650 ( .A(n8135), .ZN(n8036) );
  OR2_X1 U9651 ( .A1(n9253), .A2(n8036), .ZN(n8037) );
  INV_X1 U9652 ( .A(n9253), .ZN(n9395) );
  OR2_X1 U9653 ( .A1(n9563), .A2(n9377), .ZN(n8098) );
  NAND2_X1 U9654 ( .A1(n9395), .A2(n8098), .ZN(n8138) );
  NAND2_X1 U9655 ( .A1(n9390), .A2(n9402), .ZN(n8096) );
  NAND2_X1 U9656 ( .A1(n9563), .A2(n9377), .ZN(n9372) );
  AND2_X1 U9657 ( .A1(n8096), .A2(n9372), .ZN(n9256) );
  OAI21_X1 U9658 ( .B1(n8042), .B2(n8138), .A(n9256), .ZN(n8038) );
  AND2_X1 U9659 ( .A1(n9230), .A2(n9366), .ZN(n9255) );
  INV_X1 U9660 ( .A(n9255), .ZN(n8139) );
  NAND2_X1 U9661 ( .A1(n8038), .A2(n8139), .ZN(n8040) );
  NAND2_X1 U9662 ( .A1(n8098), .A2(n9252), .ZN(n8041) );
  NAND2_X1 U9663 ( .A1(n9256), .A2(n8041), .ZN(n8184) );
  AOI21_X1 U9664 ( .B1(n8042), .B2(n8098), .A(n8184), .ZN(n8045) );
  INV_X1 U9665 ( .A(n8043), .ZN(n8044) );
  OAI21_X1 U9666 ( .B1(n8045), .B2(n9255), .A(n8044), .ZN(n8046) );
  NAND2_X1 U9667 ( .A1(n8058), .A2(n9260), .ZN(n8049) );
  INV_X1 U9668 ( .A(n9536), .ZN(n9313) );
  AOI21_X1 U9669 ( .B1(n8049), .B2(n9313), .A(n9339), .ZN(n8052) );
  NAND2_X1 U9670 ( .A1(n8058), .A2(n9262), .ZN(n8050) );
  AOI21_X1 U9671 ( .B1(n8050), .B2(n8093), .A(n9536), .ZN(n8051) );
  MUX2_X1 U9672 ( .A(n8052), .B(n8051), .S(n8061), .Z(n8064) );
  NAND2_X1 U9673 ( .A1(n9536), .A2(n9260), .ZN(n8053) );
  NAND2_X1 U9674 ( .A1(n8128), .A2(n8053), .ZN(n8056) );
  NAND2_X1 U9675 ( .A1(n9262), .A2(n9339), .ZN(n8054) );
  NAND2_X1 U9676 ( .A1(n9264), .A2(n8054), .ZN(n8055) );
  MUX2_X1 U9677 ( .A(n8056), .B(n8055), .S(n8061), .Z(n8057) );
  INV_X1 U9678 ( .A(n8057), .ZN(n8060) );
  NOR2_X1 U9679 ( .A1(n8058), .A2(n9305), .ZN(n8059) );
  MUX2_X1 U9680 ( .A(n9264), .B(n8128), .S(n8061), .Z(n8062) );
  OAI21_X1 U9681 ( .B1(n8064), .B2(n8063), .A(n8062), .ZN(n8065) );
  NAND2_X1 U9682 ( .A1(n9284), .A2(n9269), .ZN(n9266) );
  INV_X1 U9683 ( .A(n9289), .ZN(n9265) );
  NAND2_X1 U9684 ( .A1(n8065), .A2(n9265), .ZN(n8067) );
  MUX2_X1 U9685 ( .A(n9266), .B(n8126), .S(n8039), .Z(n8066) );
  NOR2_X1 U9686 ( .A1(n8081), .A2(n9294), .ZN(n8069) );
  AOI21_X1 U9687 ( .B1(n8081), .B2(n9294), .A(n8039), .ZN(n8068) );
  NAND2_X1 U9688 ( .A1(n9026), .A2(n8072), .ZN(n8074) );
  NAND2_X1 U9689 ( .A1(n6265), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U9690 ( .A1(n6195), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8079) );
  INV_X1 U9691 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8075) );
  OR2_X1 U9692 ( .A1(n6376), .A2(n8075), .ZN(n8078) );
  INV_X1 U9693 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9214) );
  OR2_X1 U9694 ( .A1(n8076), .A2(n9214), .ZN(n8077) );
  AND3_X1 U9695 ( .A1(n8079), .A2(n8078), .A3(n8077), .ZN(n9270) );
  NOR2_X1 U9696 ( .A1(n10146), .A2(n9270), .ZN(n8236) );
  NAND2_X1 U9697 ( .A1(n8236), .A2(n9516), .ZN(n8080) );
  NAND2_X1 U9698 ( .A1(n8080), .A2(n8239), .ZN(n8125) );
  INV_X1 U9699 ( .A(n8081), .ZN(n8082) );
  NAND3_X1 U9700 ( .A1(n8082), .A2(n8039), .A3(n9294), .ZN(n8083) );
  INV_X1 U9701 ( .A(n9270), .ZN(n9158) );
  NAND2_X1 U9702 ( .A1(n9158), .A2(n8086), .ZN(n8084) );
  NAND2_X1 U9703 ( .A1(n10146), .A2(n8084), .ZN(n8190) );
  NOR2_X1 U9704 ( .A1(n6336), .A2(n8253), .ZN(n8089) );
  INV_X1 U9705 ( .A(n8191), .ZN(n8091) );
  NAND2_X1 U9706 ( .A1(n10146), .A2(n9270), .ZN(n8090) );
  NAND2_X1 U9707 ( .A1(n8091), .A2(n8090), .ZN(n8240) );
  NAND2_X1 U9708 ( .A1(n9523), .A2(n8092), .ZN(n8131) );
  NAND2_X1 U9709 ( .A1(n8094), .A2(n9258), .ZN(n9347) );
  NAND2_X1 U9710 ( .A1(n9257), .A2(n8095), .ZN(n9365) );
  INV_X1 U9711 ( .A(n8096), .ZN(n8097) );
  NAND2_X1 U9712 ( .A1(n8098), .A2(n9372), .ZN(n9400) );
  NOR2_X1 U9713 ( .A1(n9253), .A2(n9252), .ZN(n9419) );
  NAND2_X1 U9714 ( .A1(n8099), .A2(n9249), .ZN(n9441) );
  INV_X1 U9715 ( .A(n9465), .ZN(n8117) );
  INV_X1 U9716 ( .A(n9479), .ZN(n8116) );
  INV_X1 U9717 ( .A(n9497), .ZN(n9494) );
  NAND3_X1 U9718 ( .A1(n8102), .A2(n8101), .A3(n8100), .ZN(n8106) );
  NOR4_X1 U9719 ( .A1(n8106), .A2(n8105), .A3(n8104), .A4(n8103), .ZN(n8109)
         );
  NAND4_X1 U9720 ( .A1(n8109), .A2(n10268), .A3(n8108), .A4(n8107), .ZN(n8112)
         );
  NOR3_X1 U9721 ( .A1(n8112), .A2(n8111), .A3(n8110), .ZN(n8113) );
  NAND4_X1 U9722 ( .A1(n8114), .A2(n10113), .A3(n8113), .A4(n10131), .ZN(n8115) );
  NOR4_X1 U9723 ( .A1(n8117), .A2(n8116), .A3(n9494), .A4(n8115), .ZN(n8118)
         );
  NAND4_X1 U9724 ( .A1(n9419), .A2(n9435), .A3(n4879), .A4(n8118), .ZN(n8119)
         );
  OR4_X1 U9725 ( .A1(n9365), .A2(n9380), .A3(n9400), .A4(n8119), .ZN(n8120) );
  NOR4_X1 U9726 ( .A1(n9305), .A2(n9337), .A3(n9347), .A4(n8120), .ZN(n8121)
         );
  NAND4_X1 U9727 ( .A1(n9267), .A2(n9265), .A3(n9314), .A4(n8121), .ZN(n8122)
         );
  NOR4_X1 U9728 ( .A1(n8240), .A2(n8123), .A3(n8236), .A4(n8122), .ZN(n8124)
         );
  NOR2_X1 U9729 ( .A1(n8124), .A2(n6337), .ZN(n8202) );
  INV_X1 U9730 ( .A(n8125), .ZN(n8193) );
  NAND2_X1 U9731 ( .A1(n8127), .A2(n8126), .ZN(n8235) );
  INV_X1 U9732 ( .A(n9264), .ZN(n9290) );
  OAI211_X1 U9733 ( .C1(n9290), .C2(n4510), .A(n9266), .B(n8128), .ZN(n8129)
         );
  INV_X1 U9734 ( .A(n8129), .ZN(n8130) );
  OR2_X1 U9735 ( .A1(n8235), .A2(n8130), .ZN(n8132) );
  AND2_X1 U9736 ( .A1(n8132), .A2(n8131), .ZN(n8238) );
  INV_X1 U9737 ( .A(n8133), .ZN(n8186) );
  INV_X1 U9738 ( .A(n8134), .ZN(n8136) );
  OAI21_X1 U9739 ( .B1(n8136), .B2(n9248), .A(n8135), .ZN(n8137) );
  NOR2_X1 U9740 ( .A1(n8138), .A2(n8137), .ZN(n8140) );
  OAI21_X1 U9741 ( .B1(n8184), .B2(n8140), .A(n8139), .ZN(n8141) );
  NOR2_X1 U9742 ( .A1(n8142), .A2(n8141), .ZN(n8143) );
  OAI211_X1 U9743 ( .C1(n8186), .C2(n8143), .A(n9263), .B(n9260), .ZN(n8233)
         );
  NOR2_X1 U9744 ( .A1(n9247), .A2(n4778), .ZN(n8144) );
  NAND2_X1 U9745 ( .A1(n8144), .A2(n9249), .ZN(n8166) );
  NAND2_X1 U9746 ( .A1(n9243), .A2(n8145), .ZN(n8179) );
  INV_X1 U9747 ( .A(n8146), .ZN(n8155) );
  INV_X1 U9748 ( .A(n8147), .ZN(n8153) );
  INV_X1 U9749 ( .A(n8148), .ZN(n8152) );
  INV_X1 U9750 ( .A(n8149), .ZN(n8150) );
  OAI211_X1 U9751 ( .C1(n8153), .C2(n8152), .A(n8151), .B(n8150), .ZN(n8175)
         );
  OR4_X1 U9752 ( .A1(n8179), .A2(n8155), .A3(n8154), .A4(n8175), .ZN(n8156) );
  NOR2_X1 U9753 ( .A1(n8166), .A2(n8156), .ZN(n8229) );
  NAND2_X1 U9754 ( .A1(n8157), .A2(n8215), .ZN(n8158) );
  AOI21_X1 U9755 ( .B1(n8159), .B2(n8219), .A(n8158), .ZN(n8162) );
  OAI211_X1 U9756 ( .C1(n8162), .C2(n8220), .A(n8161), .B(n8160), .ZN(n8165)
         );
  INV_X1 U9757 ( .A(n8163), .ZN(n8164) );
  NAND2_X1 U9758 ( .A1(n8165), .A2(n8164), .ZN(n8183) );
  INV_X1 U9759 ( .A(n8166), .ZN(n8182) );
  INV_X1 U9760 ( .A(n8167), .ZN(n8168) );
  NOR2_X1 U9761 ( .A1(n8169), .A2(n8168), .ZN(n8174) );
  INV_X1 U9762 ( .A(n8170), .ZN(n8172) );
  OR2_X1 U9763 ( .A1(n8172), .A2(n8171), .ZN(n8173) );
  OAI21_X1 U9764 ( .B1(n8175), .B2(n8174), .A(n8173), .ZN(n8177) );
  NOR2_X1 U9765 ( .A1(n8177), .A2(n8176), .ZN(n8180) );
  AND2_X1 U9766 ( .A1(n8178), .A2(n9473), .ZN(n9244) );
  OAI21_X1 U9767 ( .B1(n8180), .B2(n8179), .A(n9244), .ZN(n8181) );
  AND2_X1 U9768 ( .A1(n8182), .A2(n8181), .ZN(n8207) );
  AOI21_X1 U9769 ( .B1(n8229), .B2(n8183), .A(n8207), .ZN(n8187) );
  OR3_X1 U9770 ( .A1(n8186), .A2(n8185), .A3(n8184), .ZN(n8230) );
  OAI21_X1 U9771 ( .B1(n8187), .B2(n8230), .A(n9264), .ZN(n8188) );
  OR3_X1 U9772 ( .A1(n8235), .A2(n8233), .A3(n8188), .ZN(n8189) );
  NAND3_X1 U9773 ( .A1(n8190), .A2(n8238), .A3(n8189), .ZN(n8192) );
  AOI211_X1 U9774 ( .C1(n8193), .C2(n8192), .A(n8253), .B(n8191), .ZN(n8194)
         );
  NOR3_X1 U9775 ( .A1(n8202), .A2(n9200), .A3(n8194), .ZN(n8201) );
  NAND3_X1 U9776 ( .A1(n10288), .A2(n8195), .A3(n9207), .ZN(n8196) );
  OR2_X1 U9777 ( .A1(n8197), .A2(n8196), .ZN(n8200) );
  INV_X1 U9778 ( .A(P1_B_REG_SCAN_IN), .ZN(n8198) );
  AOI21_X1 U9779 ( .B1(n5786), .B2(n8250), .A(n8198), .ZN(n8199) );
  AND2_X1 U9780 ( .A1(n8200), .A2(n8199), .ZN(n8249) );
  INV_X1 U9781 ( .A(n8202), .ZN(n8203) );
  OAI21_X1 U9782 ( .B1(n8205), .B2(n8204), .A(n8203), .ZN(n8206) );
  NAND2_X1 U9783 ( .A1(n8206), .A2(n9200), .ZN(n8252) );
  INV_X1 U9784 ( .A(n8207), .ZN(n8232) );
  INV_X1 U9785 ( .A(n8208), .ZN(n8209) );
  OAI211_X1 U9786 ( .C1(n8211), .C2(n8210), .A(n6337), .B(n8209), .ZN(n8212)
         );
  NAND3_X1 U9787 ( .A1(n8214), .A2(n8213), .A3(n8212), .ZN(n8218) );
  INV_X1 U9788 ( .A(n8215), .ZN(n8216) );
  AOI21_X1 U9789 ( .B1(n8218), .B2(n8217), .A(n8216), .ZN(n8223) );
  INV_X1 U9790 ( .A(n8219), .ZN(n8221) );
  NOR4_X1 U9791 ( .A1(n8223), .A2(n8222), .A3(n8221), .A4(n8220), .ZN(n8227)
         );
  INV_X1 U9792 ( .A(n8224), .ZN(n8226) );
  OAI21_X1 U9793 ( .B1(n8227), .B2(n8226), .A(n8225), .ZN(n8228) );
  NAND2_X1 U9794 ( .A1(n8229), .A2(n8228), .ZN(n8231) );
  AOI21_X1 U9795 ( .B1(n8232), .B2(n8231), .A(n8230), .ZN(n8234) );
  OR4_X1 U9796 ( .A1(n8235), .A2(n9305), .A3(n8234), .A4(n8233), .ZN(n8237) );
  AOI21_X1 U9797 ( .B1(n8238), .B2(n8237), .A(n8236), .ZN(n8241) );
  OAI21_X1 U9798 ( .B1(n8241), .B2(n8240), .A(n8239), .ZN(n8243) );
  INV_X1 U9799 ( .A(n8249), .ZN(n8245) );
  NAND3_X1 U9800 ( .A1(n8243), .A2(n8242), .A3(n8245), .ZN(n8248) );
  INV_X1 U9801 ( .A(n8243), .ZN(n8246) );
  NAND4_X1 U9802 ( .A1(n8246), .A2(n9200), .A3(n8245), .A4(n8244), .ZN(n8247)
         );
  OAI211_X1 U9803 ( .C1(n8250), .C2(n8249), .A(n8248), .B(n8247), .ZN(n8251)
         );
  OAI222_X1 U9804 ( .A1(n9624), .A2(n8254), .B1(n9622), .B2(n5488), .C1(n8253), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  XNOR2_X1 U9805 ( .A(n8256), .B(n8310), .ZN(n8262) );
  INV_X1 U9806 ( .A(n8723), .ZN(n8259) );
  OAI22_X1 U9807 ( .A1(n8257), .A2(n8890), .B1(n8274), .B2(n8892), .ZN(n8717)
         );
  AOI22_X1 U9808 ( .A1(n8717), .A2(n8287), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8258) );
  OAI21_X1 U9809 ( .B1(n8259), .B2(n8341), .A(n8258), .ZN(n8260) );
  AOI21_X1 U9810 ( .B1(n8722), .B2(n8346), .A(n8260), .ZN(n8261) );
  OAI21_X1 U9811 ( .B1(n8262), .B2(n8348), .A(n8261), .ZN(P2_U3218) );
  OAI21_X1 U9812 ( .B1(n8265), .B2(n8264), .A(n8263), .ZN(n8266) );
  NAND2_X1 U9813 ( .A1(n8266), .A2(n8329), .ZN(n8270) );
  INV_X1 U9814 ( .A(n8267), .ZN(n8780) );
  AND2_X1 U9815 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8623) );
  OAI22_X1 U9816 ( .A1(n8304), .A2(n8343), .B1(n8342), .B2(n8275), .ZN(n8268)
         );
  AOI211_X1 U9817 ( .C1(n8299), .C2(n8780), .A(n8623), .B(n8268), .ZN(n8269)
         );
  OAI211_X1 U9818 ( .C1(n8782), .C2(n8335), .A(n8270), .B(n8269), .ZN(P2_U3221) );
  NAND2_X1 U9819 ( .A1(n4506), .A2(n8271), .ZN(n8273) );
  XNOR2_X1 U9820 ( .A(n8273), .B(n8272), .ZN(n8279) );
  OAI22_X1 U9821 ( .A1(n8341), .A2(n8747), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9955), .ZN(n8277) );
  OAI22_X1 U9822 ( .A1(n8275), .A2(n8343), .B1(n8342), .B2(n8274), .ZN(n8276)
         );
  AOI211_X1 U9823 ( .C1(n8935), .C2(n8346), .A(n8277), .B(n8276), .ZN(n8278)
         );
  OAI21_X1 U9824 ( .B1(n8279), .B2(n8348), .A(n8278), .ZN(P2_U3225) );
  XNOR2_X1 U9825 ( .A(n8282), .B(n8281), .ZN(n8283) );
  XNOR2_X1 U9826 ( .A(n8280), .B(n8283), .ZN(n8291) );
  OR2_X1 U9827 ( .A1(n8284), .A2(n8890), .ZN(n8286) );
  NAND2_X1 U9828 ( .A1(n8562), .A2(n8816), .ZN(n8285) );
  NAND2_X1 U9829 ( .A1(n8286), .A2(n8285), .ZN(n8679) );
  AOI22_X1 U9830 ( .A1(n8679), .A2(n8287), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8288) );
  OAI21_X1 U9831 ( .B1(n8686), .B2(n8341), .A(n8288), .ZN(n8289) );
  AOI21_X1 U9832 ( .B1(n8685), .B2(n8346), .A(n8289), .ZN(n8290) );
  OAI21_X1 U9833 ( .B1(n8291), .B2(n8348), .A(n8290), .ZN(P2_U3227) );
  OAI21_X1 U9834 ( .B1(n8294), .B2(n8293), .A(n8292), .ZN(n8295) );
  NAND2_X1 U9835 ( .A1(n8295), .A2(n8329), .ZN(n8301) );
  INV_X1 U9836 ( .A(n8296), .ZN(n8849) );
  OAI22_X1 U9837 ( .A1(n8891), .A2(n8343), .B1(n8342), .B2(n8842), .ZN(n8297)
         );
  AOI211_X1 U9838 ( .C1(n8849), .C2(n8299), .A(n8298), .B(n8297), .ZN(n8300)
         );
  OAI211_X1 U9839 ( .C1(n4834), .C2(n8335), .A(n8301), .B(n8300), .ZN(P2_U3228) );
  XNOR2_X1 U9840 ( .A(n8303), .B(n8302), .ZN(n8308) );
  OAI22_X1 U9841 ( .A1(n8341), .A2(n8826), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5441), .ZN(n8306) );
  OAI22_X1 U9842 ( .A1(n8304), .A2(n8342), .B1(n8343), .B2(n8859), .ZN(n8305)
         );
  AOI211_X1 U9843 ( .C1(n8825), .C2(n8346), .A(n8306), .B(n8305), .ZN(n8307)
         );
  OAI21_X1 U9844 ( .B1(n8308), .B2(n8348), .A(n8307), .ZN(P2_U3230) );
  AOI21_X1 U9845 ( .B1(n8310), .B2(n8256), .A(n8309), .ZN(n8314) );
  XNOR2_X1 U9846 ( .A(n8312), .B(n8311), .ZN(n8313) );
  XNOR2_X1 U9847 ( .A(n8314), .B(n8313), .ZN(n8318) );
  OAI22_X1 U9848 ( .A1(n8341), .A2(n8697), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9752), .ZN(n8316) );
  OAI22_X1 U9849 ( .A1(n8702), .A2(n8342), .B1(n8343), .B2(n8738), .ZN(n8315)
         );
  AOI211_X1 U9850 ( .C1(n8920), .C2(n8346), .A(n8316), .B(n8315), .ZN(n8317)
         );
  OAI21_X1 U9851 ( .B1(n8318), .B2(n8348), .A(n8317), .ZN(P2_U3231) );
  XNOR2_X1 U9852 ( .A(n8320), .B(n8319), .ZN(n8325) );
  OAI22_X1 U9853 ( .A1(n8341), .A2(n8761), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9744), .ZN(n8323) );
  OAI22_X1 U9854 ( .A1(n8321), .A2(n8343), .B1(n8342), .B2(n8737), .ZN(n8322)
         );
  AOI211_X1 U9855 ( .C1(n8940), .C2(n8346), .A(n8323), .B(n8322), .ZN(n8324)
         );
  OAI21_X1 U9856 ( .B1(n8325), .B2(n8348), .A(n8324), .ZN(P2_U3235) );
  INV_X1 U9857 ( .A(n8930), .ZN(n8734) );
  OAI21_X1 U9858 ( .B1(n8328), .B2(n8327), .A(n8326), .ZN(n8330) );
  NAND2_X1 U9859 ( .A1(n8330), .A2(n8329), .ZN(n8334) );
  NOR2_X1 U9860 ( .A1(n8341), .A2(n8731), .ZN(n8332) );
  OAI22_X1 U9861 ( .A1(n8737), .A2(n8343), .B1(n8342), .B2(n8738), .ZN(n8331)
         );
  AOI211_X1 U9862 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3152), .A(n8332), 
        .B(n8331), .ZN(n8333) );
  OAI211_X1 U9863 ( .C1(n8734), .C2(n8335), .A(n8334), .B(n8333), .ZN(P2_U3237) );
  NAND2_X1 U9864 ( .A1(n8337), .A2(n8336), .ZN(n8339) );
  XNOR2_X1 U9865 ( .A(n8339), .B(n8338), .ZN(n8349) );
  OAI22_X1 U9866 ( .A1(n8341), .A2(n8870), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8340), .ZN(n8345) );
  OAI22_X1 U9867 ( .A1(n8860), .A2(n8343), .B1(n8342), .B2(n8859), .ZN(n8344)
         );
  AOI211_X1 U9868 ( .C1(n8967), .C2(n8346), .A(n8345), .B(n8344), .ZN(n8347)
         );
  OAI21_X1 U9869 ( .B1(n8349), .B2(n8348), .A(n8347), .ZN(P2_U3243) );
  INV_X1 U9870 ( .A(n8533), .ZN(n8350) );
  NAND2_X1 U9871 ( .A1(n9026), .A2(n8352), .ZN(n8354) );
  NAND2_X1 U9872 ( .A1(n4480), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8353) );
  INV_X1 U9873 ( .A(n8559), .ZN(n8358) );
  NOR2_X1 U9874 ( .A1(n8627), .A2(n8358), .ZN(n8541) );
  INV_X1 U9875 ( .A(n8631), .ZN(n8360) );
  NOR2_X1 U9876 ( .A1(n8628), .A2(n8360), .ZN(n8542) );
  AND2_X1 U9877 ( .A1(n8627), .A2(n8358), .ZN(n8387) );
  INV_X1 U9878 ( .A(n8541), .ZN(n8362) );
  INV_X1 U9879 ( .A(n8787), .ZN(n8777) );
  NAND2_X1 U9880 ( .A1(n8488), .A2(n8783), .ZN(n8801) );
  INV_X1 U9881 ( .A(n8821), .ZN(n8479) );
  NAND2_X1 U9882 ( .A1(n8363), .A2(n8408), .ZN(n10409) );
  NOR4_X1 U9883 ( .A1(n8365), .A2(n8364), .A3(n10409), .A4(n7215), .ZN(n8370)
         );
  NOR4_X1 U9884 ( .A1(n7192), .A2(n8368), .A3(n8367), .A4(n8366), .ZN(n8369)
         );
  AND4_X1 U9885 ( .A1(n8370), .A2(n8369), .A3(n8436), .A4(n8430), .ZN(n8371)
         );
  NAND4_X1 U9886 ( .A1(n8371), .A2(n5349), .A3(n8444), .A4(n8443), .ZN(n8373)
         );
  NOR4_X1 U9887 ( .A1(n5040), .A2(n8373), .A3(n5384), .A4(n8372), .ZN(n8374)
         );
  NAND4_X1 U9888 ( .A1(n8479), .A2(n8834), .A3(n8473), .A4(n8374), .ZN(n8375)
         );
  NOR4_X1 U9889 ( .A1(n8771), .A2(n8777), .A3(n8801), .A4(n8375), .ZN(n8376)
         );
  NAND3_X1 U9890 ( .A1(n8711), .A2(n8377), .A3(n8376), .ZN(n8378) );
  NOR4_X1 U9891 ( .A1(n8659), .A2(n8751), .A3(n8701), .A4(n8378), .ZN(n8380)
         );
  NAND4_X1 U9892 ( .A1(n8639), .A2(n8380), .A3(n8508), .A4(n5595), .ZN(n8381)
         );
  OAI22_X1 U9893 ( .A1(n8383), .A2(n8407), .B1(n8546), .B2(n8384), .ZN(n8550)
         );
  INV_X1 U9894 ( .A(n8384), .ZN(n8386) );
  INV_X1 U9895 ( .A(n8385), .ZN(n10407) );
  INV_X1 U9896 ( .A(n8387), .ZN(n8537) );
  NAND2_X1 U9897 ( .A1(n8388), .A2(n8650), .ZN(n8389) );
  NAND2_X1 U9898 ( .A1(n8522), .A2(n8389), .ZN(n8392) );
  NAND2_X1 U9899 ( .A1(n8407), .A2(n8390), .ZN(n8391) );
  OR2_X1 U9900 ( .A1(n8554), .A2(n8391), .ZN(n8543) );
  MUX2_X1 U9901 ( .A(n8393), .B(n8392), .S(n8543), .Z(n8529) );
  INV_X1 U9902 ( .A(n8543), .ZN(n8523) );
  AND2_X1 U9903 ( .A1(n8404), .A2(n8403), .ZN(n8394) );
  MUX2_X1 U9904 ( .A(n8394), .B(n8398), .S(n8543), .Z(n8414) );
  INV_X1 U9905 ( .A(n8414), .ZN(n8396) );
  NAND2_X1 U9906 ( .A1(n8396), .A2(n8395), .ZN(n8401) );
  NAND2_X1 U9907 ( .A1(n8398), .A2(n8397), .ZN(n8400) );
  INV_X1 U9908 ( .A(n8426), .ZN(n8399) );
  AOI21_X1 U9909 ( .B1(n8401), .B2(n8400), .A(n8399), .ZN(n8429) );
  NAND2_X1 U9910 ( .A1(n8403), .A2(n8402), .ZN(n8406) );
  NAND2_X1 U9911 ( .A1(n8432), .A2(n8404), .ZN(n8405) );
  AOI21_X1 U9912 ( .B1(n8414), .B2(n8406), .A(n8405), .ZN(n8416) );
  AND2_X1 U9913 ( .A1(n8408), .A2(n8407), .ZN(n8409) );
  OAI211_X1 U9914 ( .C1(n8410), .C2(n8409), .A(n8423), .B(n5650), .ZN(n8411)
         );
  NAND3_X1 U9915 ( .A1(n8411), .A2(n8421), .A3(n8543), .ZN(n8412) );
  NAND3_X1 U9916 ( .A1(n8414), .A2(n8413), .A3(n8412), .ZN(n8415) );
  OAI21_X1 U9917 ( .B1(n8416), .B2(n8523), .A(n8415), .ZN(n8427) );
  NAND2_X1 U9918 ( .A1(n8417), .A2(n6910), .ZN(n8422) );
  NAND2_X1 U9919 ( .A1(n5650), .A2(n8418), .ZN(n8419) );
  NAND4_X1 U9920 ( .A1(n8422), .A2(n8421), .A3(n8420), .A4(n8419), .ZN(n8424)
         );
  NAND3_X1 U9921 ( .A1(n8424), .A2(n8523), .A3(n8423), .ZN(n8425) );
  NAND3_X1 U9922 ( .A1(n8427), .A2(n8426), .A3(n8425), .ZN(n8428) );
  OAI21_X1 U9923 ( .B1(n8429), .B2(n8543), .A(n8428), .ZN(n8431) );
  OAI211_X1 U9924 ( .C1(n8432), .C2(n8543), .A(n8431), .B(n8430), .ZN(n8437)
         );
  MUX2_X1 U9925 ( .A(n8434), .B(n8433), .S(n8543), .Z(n8435) );
  NAND3_X1 U9926 ( .A1(n8437), .A2(n8436), .A3(n8435), .ZN(n8447) );
  MUX2_X1 U9927 ( .A(n8439), .B(n8438), .S(n8523), .Z(n8441) );
  AND2_X1 U9928 ( .A1(n8441), .A2(n8440), .ZN(n8446) );
  AND2_X1 U9929 ( .A1(n8450), .A2(n8523), .ZN(n8442) );
  AOI22_X1 U9930 ( .A1(n8444), .A2(n8443), .B1(n8442), .B2(n8449), .ZN(n8445)
         );
  AOI21_X1 U9931 ( .B1(n8447), .B2(n8446), .A(n8445), .ZN(n8455) );
  NAND2_X1 U9932 ( .A1(n8456), .A2(n8448), .ZN(n8453) );
  INV_X1 U9933 ( .A(n8448), .ZN(n8451) );
  OAI211_X1 U9934 ( .C1(n8451), .C2(n8450), .A(n8460), .B(n8449), .ZN(n8452)
         );
  MUX2_X1 U9935 ( .A(n8453), .B(n8452), .S(n8543), .Z(n8454) );
  OR2_X1 U9936 ( .A1(n8455), .A2(n8454), .ZN(n8462) );
  NAND3_X1 U9937 ( .A1(n8462), .A2(n8463), .A3(n8456), .ZN(n8457) );
  NAND3_X1 U9938 ( .A1(n8457), .A2(n8464), .A3(n8461), .ZN(n8459) );
  NAND2_X1 U9939 ( .A1(n8459), .A2(n8458), .ZN(n8469) );
  NAND3_X1 U9940 ( .A1(n8462), .A2(n8461), .A3(n8460), .ZN(n8465) );
  NAND3_X1 U9941 ( .A1(n8465), .A2(n8464), .A3(n8463), .ZN(n8467) );
  NAND2_X1 U9942 ( .A1(n8467), .A2(n8466), .ZN(n8468) );
  MUX2_X1 U9943 ( .A(n8471), .B(n8470), .S(n8543), .Z(n8472) );
  MUX2_X1 U9944 ( .A(n8475), .B(n8474), .S(n8543), .Z(n8476) );
  MUX2_X1 U9945 ( .A(n8810), .B(n8477), .S(n8543), .Z(n8478) );
  NAND2_X1 U9946 ( .A1(n8480), .A2(n8479), .ZN(n8484) );
  AND2_X1 U9947 ( .A1(n8783), .A2(n8481), .ZN(n8482) );
  MUX2_X1 U9948 ( .A(n8766), .B(n8482), .S(n8523), .Z(n8483) );
  NAND2_X1 U9949 ( .A1(n8484), .A2(n8483), .ZN(n8489) );
  NAND2_X1 U9950 ( .A1(n8489), .A2(n8783), .ZN(n8485) );
  NAND2_X1 U9951 ( .A1(n8485), .A2(n8492), .ZN(n8486) );
  NAND3_X1 U9952 ( .A1(n8486), .A2(n8496), .A3(n8490), .ZN(n8487) );
  OR2_X1 U9953 ( .A1(n8935), .A2(n8737), .ZN(n8498) );
  NAND2_X1 U9954 ( .A1(n8489), .A2(n8488), .ZN(n8491) );
  NAND2_X1 U9955 ( .A1(n8491), .A2(n8490), .ZN(n8494) );
  NAND3_X1 U9956 ( .A1(n8494), .A2(n8493), .A3(n8492), .ZN(n8497) );
  INV_X1 U9957 ( .A(n8500), .ZN(n8501) );
  OAI21_X1 U9958 ( .B1(n8701), .B2(n8501), .A(n8523), .ZN(n8503) );
  INV_X1 U9959 ( .A(n8506), .ZN(n8502) );
  AOI21_X1 U9960 ( .B1(n8504), .B2(n8503), .A(n8502), .ZN(n8511) );
  AOI21_X1 U9961 ( .B1(n8506), .B2(n8505), .A(n8523), .ZN(n8510) );
  NOR2_X1 U9962 ( .A1(n8676), .A2(n8523), .ZN(n8507) );
  NOR2_X1 U9963 ( .A1(n8659), .A2(n8507), .ZN(n8509) );
  INV_X1 U9964 ( .A(n8512), .ZN(n8658) );
  NAND2_X1 U9965 ( .A1(n8658), .A2(n8516), .ZN(n8513) );
  NAND2_X1 U9966 ( .A1(n8513), .A2(n8515), .ZN(n8519) );
  NAND2_X1 U9967 ( .A1(n8685), .A2(n8702), .ZN(n8514) );
  NAND2_X1 U9968 ( .A1(n8515), .A2(n8514), .ZN(n8517) );
  NAND2_X1 U9969 ( .A1(n8517), .A2(n8516), .ZN(n8518) );
  MUX2_X1 U9970 ( .A(n8519), .B(n8518), .S(n8543), .Z(n8520) );
  OAI21_X1 U9971 ( .B1(n8523), .B2(n8905), .A(n8522), .ZN(n8526) );
  NAND2_X1 U9972 ( .A1(n8524), .A2(n8543), .ZN(n8525) );
  NAND2_X1 U9973 ( .A1(n8526), .A2(n8525), .ZN(n8527) );
  OAI21_X1 U9974 ( .B1(n8529), .B2(n8528), .A(n8527), .ZN(n8531) );
  NAND2_X1 U9975 ( .A1(n8531), .A2(n8530), .ZN(n8535) );
  MUX2_X1 U9976 ( .A(n8533), .B(n8532), .S(n8543), .Z(n8534) );
  NAND2_X1 U9977 ( .A1(n8535), .A2(n8534), .ZN(n8536) );
  NAND2_X1 U9978 ( .A1(n8537), .A2(n8536), .ZN(n8540) );
  MUX2_X1 U9979 ( .A(n8538), .B(n4560), .S(n8543), .Z(n8539) );
  OAI21_X1 U9980 ( .B1(n8541), .B2(n8540), .A(n8539), .ZN(n8548) );
  INV_X1 U9981 ( .A(n8542), .ZN(n8544) );
  MUX2_X1 U9982 ( .A(n8545), .B(n8544), .S(n8543), .Z(n8547) );
  AOI21_X1 U9983 ( .B1(n8548), .B2(n8547), .A(n8546), .ZN(n8549) );
  NOR3_X1 U9984 ( .A1(n8892), .A2(n8553), .A3(n8552), .ZN(n8556) );
  OAI21_X1 U9985 ( .B1(n8557), .B2(n8554), .A(P2_B_REG_SCAN_IN), .ZN(n8555) );
  OAI22_X1 U9986 ( .A1(n8558), .A2(n8557), .B1(n8556), .B2(n8555), .ZN(
        P2_U3244) );
  MUX2_X1 U9987 ( .A(n8559), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8578), .Z(
        P2_U3582) );
  MUX2_X1 U9988 ( .A(n8560), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8578), .Z(
        P2_U3580) );
  MUX2_X1 U9989 ( .A(n8561), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8578), .Z(
        P2_U3577) );
  MUX2_X1 U9990 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8562), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U9991 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8753), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9992 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8788), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9993 ( .A(n8804), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8578), .Z(
        P2_U3571) );
  MUX2_X1 U9994 ( .A(n8814), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8578), .Z(
        P2_U3570) );
  MUX2_X1 U9995 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8803), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9996 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8817), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9997 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8563), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9998 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8564), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9999 ( .A(n8565), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8578), .Z(
        P2_U3565) );
  MUX2_X1 U10000 ( .A(n8566), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8578), .Z(
        P2_U3564) );
  MUX2_X1 U10001 ( .A(n8567), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8578), .Z(
        P2_U3563) );
  MUX2_X1 U10002 ( .A(n8568), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8578), .Z(
        P2_U3562) );
  MUX2_X1 U10003 ( .A(n8569), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8578), .Z(
        P2_U3561) );
  MUX2_X1 U10004 ( .A(n8570), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8578), .Z(
        P2_U3560) );
  MUX2_X1 U10005 ( .A(n8571), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8578), .Z(
        P2_U3559) );
  MUX2_X1 U10006 ( .A(n8572), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8578), .Z(
        P2_U3558) );
  MUX2_X1 U10007 ( .A(n8573), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8578), .Z(
        P2_U3557) );
  MUX2_X1 U10008 ( .A(n8574), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8578), .Z(
        P2_U3556) );
  MUX2_X1 U10009 ( .A(n8575), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8578), .Z(
        P2_U3555) );
  MUX2_X1 U10010 ( .A(n8576), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8578), .Z(
        P2_U3554) );
  MUX2_X1 U10011 ( .A(n8577), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8578), .Z(
        P2_U3553) );
  MUX2_X1 U10012 ( .A(n8579), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8578), .Z(
        P2_U3552) );
  AOI211_X1 U10013 ( .C1(n8582), .C2(n8581), .A(n8580), .B(n10347), .ZN(n8583)
         );
  INV_X1 U10014 ( .A(n8583), .ZN(n8592) );
  AOI21_X1 U10015 ( .B1(n10350), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8584), .ZN(
        n8591) );
  NAND2_X1 U10016 ( .A1(n10042), .A2(n8585), .ZN(n8590) );
  OAI211_X1 U10017 ( .C1(n8588), .C2(n8587), .A(n10342), .B(n8586), .ZN(n8589)
         );
  NAND4_X1 U10018 ( .A1(n8592), .A2(n8591), .A3(n8590), .A4(n8589), .ZN(
        P2_U3254) );
  XNOR2_X1 U10019 ( .A(n8616), .B(n8609), .ZN(n8595) );
  NOR2_X1 U10020 ( .A1(n5459), .A2(n8595), .ZN(n8610) );
  AOI21_X1 U10021 ( .B1(n8595), .B2(n5459), .A(n8610), .ZN(n8607) );
  NAND2_X1 U10022 ( .A1(n10042), .A2(n8601), .ZN(n8598) );
  NOR2_X1 U10023 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9781), .ZN(n8596) );
  AOI21_X1 U10024 ( .B1(n10350), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8596), .ZN(
        n8597) );
  NAND2_X1 U10025 ( .A1(n8598), .A2(n8597), .ZN(n8606) );
  OAI21_X1 U10026 ( .B1(n8600), .B2(n8959), .A(n8599), .ZN(n8603) );
  XNOR2_X1 U10027 ( .A(n8601), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8602) );
  NOR2_X1 U10028 ( .A1(n8603), .A2(n8602), .ZN(n8614) );
  AOI21_X1 U10029 ( .B1(n8603), .B2(n8602), .A(n8614), .ZN(n8604) );
  NOR2_X1 U10030 ( .A1(n8604), .A2(n10344), .ZN(n8605) );
  AOI211_X1 U10031 ( .C1(n10343), .C2(n8607), .A(n8606), .B(n8605), .ZN(n8608)
         );
  INV_X1 U10032 ( .A(n8608), .ZN(P2_U3263) );
  NOR2_X1 U10033 ( .A1(n8609), .A2(n8616), .ZN(n8611) );
  NOR2_X1 U10034 ( .A1(n8611), .A2(n8610), .ZN(n8613) );
  XNOR2_X1 U10035 ( .A(n8613), .B(n8612), .ZN(n8621) );
  NAND2_X1 U10036 ( .A1(n8621), .A2(n10343), .ZN(n8619) );
  AOI21_X1 U10037 ( .B1(n8616), .B2(n8615), .A(n8614), .ZN(n8617) );
  XNOR2_X1 U10038 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8617), .ZN(n8620) );
  AOI21_X1 U10039 ( .B1(n8620), .B2(n10342), .A(n10042), .ZN(n8618) );
  INV_X1 U10040 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8625) );
  INV_X1 U10041 ( .A(n8623), .ZN(n8624) );
  OAI21_X1 U10042 ( .B1(n10026), .B2(n8625), .A(n8624), .ZN(n8626) );
  INV_X1 U10043 ( .A(n8628), .ZN(n8990) );
  NOR2_X1 U10044 ( .A1(n8627), .A2(n8634), .ZN(n8629) );
  XNOR2_X1 U10045 ( .A(n8629), .B(n8628), .ZN(n8902) );
  NAND2_X1 U10046 ( .A1(n8902), .A2(n8874), .ZN(n8633) );
  AND2_X1 U10047 ( .A1(n8631), .A2(n8630), .ZN(n8901) );
  INV_X1 U10048 ( .A(n8901), .ZN(n10072) );
  NOR2_X1 U10049 ( .A1(n8877), .A2(n10072), .ZN(n8635) );
  AOI21_X1 U10050 ( .B1(n8897), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8635), .ZN(
        n8632) );
  OAI211_X1 U10051 ( .C1(n8990), .C2(n10362), .A(n8633), .B(n8632), .ZN(
        P2_U3265) );
  XNOR2_X1 U10052 ( .A(n10073), .B(n8634), .ZN(n10075) );
  NAND2_X1 U10053 ( .A1(n10075), .A2(n8874), .ZN(n8637) );
  AOI21_X1 U10054 ( .B1(n8877), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8635), .ZN(
        n8636) );
  OAI211_X1 U10055 ( .C1(n10073), .C2(n10362), .A(n8637), .B(n8636), .ZN(
        P2_U3266) );
  AOI21_X1 U10056 ( .B1(n8905), .B2(n4842), .A(n8641), .ZN(n8906) );
  INV_X1 U10057 ( .A(n8642), .ZN(n8643) );
  AOI22_X1 U10058 ( .A1(n8643), .A2(n8848), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n8897), .ZN(n8644) );
  OAI21_X1 U10059 ( .B1(n8645), .B2(n10362), .A(n8644), .ZN(n8654) );
  AOI211_X1 U10060 ( .C1(n8648), .C2(n8647), .A(n8889), .B(n8646), .ZN(n8652)
         );
  OAI22_X1 U10061 ( .A1(n8650), .A2(n8892), .B1(n8649), .B2(n8890), .ZN(n8651)
         );
  NOR2_X1 U10062 ( .A1(n8652), .A2(n8651), .ZN(n8908) );
  INV_X1 U10063 ( .A(n7188), .ZN(n8897) );
  NOR2_X1 U10064 ( .A1(n8908), .A2(n8897), .ZN(n8653) );
  AOI211_X1 U10065 ( .C1(n8906), .C2(n8874), .A(n8654), .B(n8653), .ZN(n8655)
         );
  OAI21_X1 U10066 ( .B1(n8909), .B2(n8809), .A(n8655), .ZN(P2_U3268) );
  INV_X1 U10067 ( .A(n8912), .ZN(n8674) );
  NAND2_X1 U10068 ( .A1(n8657), .A2(n8658), .ZN(n8660) );
  NAND2_X1 U10069 ( .A1(n8660), .A2(n8659), .ZN(n8662) );
  NAND2_X1 U10070 ( .A1(n8662), .A2(n8661), .ZN(n8663) );
  NAND2_X1 U10071 ( .A1(n8663), .A2(n10357), .ZN(n8665) );
  NAND2_X1 U10072 ( .A1(n8665), .A2(n8664), .ZN(n8910) );
  INV_X1 U10073 ( .A(n8666), .ZN(n8667) );
  AOI211_X1 U10074 ( .C1(n8668), .C2(n8682), .A(n10436), .B(n8667), .ZN(n8911)
         );
  NAND2_X1 U10075 ( .A1(n8911), .A2(n8830), .ZN(n8671) );
  AOI22_X1 U10076 ( .A1(n8669), .A2(n8848), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n8897), .ZN(n8670) );
  OAI211_X1 U10077 ( .C1(n8995), .C2(n10362), .A(n8671), .B(n8670), .ZN(n8672)
         );
  AOI21_X1 U10078 ( .B1(n8910), .B2(n7188), .A(n8672), .ZN(n8673) );
  OAI21_X1 U10079 ( .B1(n8674), .B2(n8809), .A(n8673), .ZN(P2_U3270) );
  XNOR2_X1 U10080 ( .A(n8675), .B(n8677), .ZN(n8917) );
  INV_X1 U10081 ( .A(n8917), .ZN(n8692) );
  NAND3_X1 U10082 ( .A1(n8704), .A2(n8677), .A3(n8676), .ZN(n8678) );
  NAND3_X1 U10083 ( .A1(n8657), .A2(n10357), .A3(n8678), .ZN(n8681) );
  INV_X1 U10084 ( .A(n8679), .ZN(n8680) );
  NAND2_X1 U10085 ( .A1(n8681), .A2(n8680), .ZN(n8915) );
  INV_X1 U10086 ( .A(n8696), .ZN(n8684) );
  INV_X1 U10087 ( .A(n8682), .ZN(n8683) );
  AOI211_X1 U10088 ( .C1(n8685), .C2(n8684), .A(n10436), .B(n8683), .ZN(n8916)
         );
  NAND2_X1 U10089 ( .A1(n8916), .A2(n8830), .ZN(n8689) );
  INV_X1 U10090 ( .A(n8686), .ZN(n8687) );
  AOI22_X1 U10091 ( .A1(n8687), .A2(n8848), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8897), .ZN(n8688) );
  OAI211_X1 U10092 ( .C1(n8999), .C2(n10362), .A(n8689), .B(n8688), .ZN(n8690)
         );
  AOI21_X1 U10093 ( .B1(n8915), .B2(n7188), .A(n8690), .ZN(n8691) );
  OAI21_X1 U10094 ( .B1(n8692), .B2(n8809), .A(n8691), .ZN(P2_U3271) );
  OAI21_X1 U10095 ( .B1(n8694), .B2(n8701), .A(n8693), .ZN(n8695) );
  INV_X1 U10096 ( .A(n8695), .ZN(n8924) );
  AOI21_X1 U10097 ( .B1(n8920), .B2(n8720), .A(n8696), .ZN(n8921) );
  INV_X1 U10098 ( .A(n8697), .ZN(n8698) );
  AOI22_X1 U10099 ( .A1(P2_REG2_REG_24__SCAN_IN), .A2(n8897), .B1(n8698), .B2(
        n8848), .ZN(n8699) );
  OAI21_X1 U10100 ( .B1(n5547), .B2(n10362), .A(n8699), .ZN(n8707) );
  AOI21_X1 U10101 ( .B1(n8700), .B2(n8701), .A(n8889), .ZN(n8705) );
  OAI22_X1 U10102 ( .A1(n8702), .A2(n8890), .B1(n8738), .B2(n8892), .ZN(n8703)
         );
  AOI21_X1 U10103 ( .B1(n8705), .B2(n8704), .A(n8703), .ZN(n8923) );
  NOR2_X1 U10104 ( .A1(n8923), .A2(n8897), .ZN(n8706) );
  AOI211_X1 U10105 ( .C1(n8921), .C2(n8874), .A(n8707), .B(n8706), .ZN(n8708)
         );
  OAI21_X1 U10106 ( .B1(n8924), .B2(n8809), .A(n8708), .ZN(P2_U3272) );
  AOI21_X1 U10107 ( .B1(n8711), .B2(n8710), .A(n8709), .ZN(n8927) );
  INV_X1 U10108 ( .A(n8927), .ZN(n8728) );
  NAND2_X1 U10109 ( .A1(n8712), .A2(n8713), .ZN(n8715) );
  XNOR2_X1 U10110 ( .A(n8715), .B(n8714), .ZN(n8716) );
  NAND2_X1 U10111 ( .A1(n8716), .A2(n10357), .ZN(n8719) );
  INV_X1 U10112 ( .A(n8717), .ZN(n8718) );
  NAND2_X1 U10113 ( .A1(n8719), .A2(n8718), .ZN(n8925) );
  INV_X1 U10114 ( .A(n8722), .ZN(n9004) );
  INV_X1 U10115 ( .A(n8720), .ZN(n8721) );
  AOI211_X1 U10116 ( .C1(n8722), .C2(n8730), .A(n10436), .B(n8721), .ZN(n8926)
         );
  NAND2_X1 U10117 ( .A1(n8926), .A2(n8830), .ZN(n8725) );
  AOI22_X1 U10118 ( .A1(n8877), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8723), .B2(
        n8848), .ZN(n8724) );
  OAI211_X1 U10119 ( .C1(n9004), .C2(n10362), .A(n8725), .B(n8724), .ZN(n8726)
         );
  AOI21_X1 U10120 ( .B1(n8925), .B2(n7188), .A(n8726), .ZN(n8727) );
  OAI21_X1 U10121 ( .B1(n8728), .B2(n8809), .A(n8727), .ZN(P2_U3273) );
  XNOR2_X1 U10122 ( .A(n8729), .B(n8735), .ZN(n8934) );
  AOI21_X1 U10123 ( .B1(n8930), .B2(n8745), .A(n4846), .ZN(n8931) );
  INV_X1 U10124 ( .A(n8731), .ZN(n8732) );
  AOI22_X1 U10125 ( .A1(n8877), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8732), .B2(
        n8848), .ZN(n8733) );
  OAI21_X1 U10126 ( .B1(n8734), .B2(n10362), .A(n8733), .ZN(n8742) );
  AOI21_X1 U10127 ( .B1(n8736), .B2(n8735), .A(n8889), .ZN(n8740) );
  OAI22_X1 U10128 ( .A1(n8738), .A2(n8890), .B1(n8737), .B2(n8892), .ZN(n8739)
         );
  AOI21_X1 U10129 ( .B1(n8740), .B2(n8712), .A(n8739), .ZN(n8933) );
  NOR2_X1 U10130 ( .A1(n8933), .A2(n8897), .ZN(n8741) );
  AOI211_X1 U10131 ( .C1(n8931), .C2(n8874), .A(n8742), .B(n8741), .ZN(n8743)
         );
  OAI21_X1 U10132 ( .B1(n8934), .B2(n8809), .A(n8743), .ZN(P2_U3274) );
  XOR2_X1 U10133 ( .A(n8751), .B(n8744), .Z(n8939) );
  INV_X1 U10134 ( .A(n8759), .ZN(n8746) );
  AOI21_X1 U10135 ( .B1(n8935), .B2(n8746), .A(n4847), .ZN(n8936) );
  INV_X1 U10136 ( .A(n8747), .ZN(n8748) );
  AOI22_X1 U10137 ( .A1(n8877), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8748), .B2(
        n8848), .ZN(n8749) );
  OAI21_X1 U10138 ( .B1(n8750), .B2(n10362), .A(n8749), .ZN(n8756) );
  XNOR2_X1 U10139 ( .A(n8752), .B(n8751), .ZN(n8754) );
  AOI222_X1 U10140 ( .A1(n10357), .A2(n8754), .B1(n8753), .B2(n8815), .C1(
        n8788), .C2(n8816), .ZN(n8938) );
  NOR2_X1 U10141 ( .A1(n8938), .A2(n8897), .ZN(n8755) );
  AOI211_X1 U10142 ( .C1(n8936), .C2(n8874), .A(n8756), .B(n8755), .ZN(n8757)
         );
  OAI21_X1 U10143 ( .B1(n8939), .B2(n8809), .A(n8757), .ZN(P2_U3275) );
  XNOR2_X1 U10144 ( .A(n8758), .B(n8771), .ZN(n8944) );
  INV_X1 U10145 ( .A(n8779), .ZN(n8760) );
  AOI21_X1 U10146 ( .B1(n8940), .B2(n8760), .A(n8759), .ZN(n8941) );
  INV_X1 U10147 ( .A(n8761), .ZN(n8762) );
  AOI22_X1 U10148 ( .A1(n8877), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8762), .B2(
        n8848), .ZN(n8763) );
  OAI21_X1 U10149 ( .B1(n8764), .B2(n10362), .A(n8763), .ZN(n8775) );
  NAND2_X1 U10150 ( .A1(n8841), .A2(n8765), .ZN(n8812) );
  NAND2_X1 U10151 ( .A1(n8812), .A2(n8766), .ZN(n8784) );
  NAND2_X1 U10152 ( .A1(n8784), .A2(n8767), .ZN(n8769) );
  AND2_X1 U10153 ( .A1(n8769), .A2(n8768), .ZN(n8770) );
  XOR2_X1 U10154 ( .A(n8771), .B(n8770), .Z(n8773) );
  AOI222_X1 U10155 ( .A1(n10357), .A2(n8773), .B1(n8772), .B2(n8815), .C1(
        n8804), .C2(n8816), .ZN(n8943) );
  NOR2_X1 U10156 ( .A1(n8943), .A2(n8897), .ZN(n8774) );
  AOI211_X1 U10157 ( .C1(n8941), .C2(n8874), .A(n8775), .B(n8774), .ZN(n8776)
         );
  OAI21_X1 U10158 ( .B1(n8809), .B2(n8944), .A(n8776), .ZN(P2_U3276) );
  XNOR2_X1 U10159 ( .A(n8778), .B(n8777), .ZN(n8949) );
  AOI211_X1 U10160 ( .C1(n8946), .C2(n8794), .A(n10436), .B(n8779), .ZN(n8945)
         );
  AOI22_X1 U10161 ( .A1(n8877), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8780), .B2(
        n8848), .ZN(n8781) );
  OAI21_X1 U10162 ( .B1(n8782), .B2(n10362), .A(n8781), .ZN(n8791) );
  NAND2_X1 U10163 ( .A1(n8784), .A2(n8783), .ZN(n8786) );
  NAND2_X1 U10164 ( .A1(n8786), .A2(n8787), .ZN(n8785) );
  OAI21_X1 U10165 ( .B1(n8787), .B2(n8786), .A(n8785), .ZN(n8789) );
  AOI222_X1 U10166 ( .A1(n10357), .A2(n8789), .B1(n8788), .B2(n8815), .C1(
        n8814), .C2(n8816), .ZN(n8948) );
  NOR2_X1 U10167 ( .A1(n8948), .A2(n8897), .ZN(n8790) );
  AOI211_X1 U10168 ( .C1(n8945), .C2(n8830), .A(n8791), .B(n8790), .ZN(n8792)
         );
  OAI21_X1 U10169 ( .B1(n8949), .B2(n8809), .A(n8792), .ZN(P2_U3277) );
  XOR2_X1 U10170 ( .A(n8801), .B(n8793), .Z(n8955) );
  INV_X1 U10171 ( .A(n8794), .ZN(n8795) );
  AOI21_X1 U10172 ( .B1(n8950), .B2(n8823), .A(n8795), .ZN(n8952) );
  INV_X1 U10173 ( .A(n8796), .ZN(n8797) );
  AOI22_X1 U10174 ( .A1(n8877), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8797), .B2(
        n8848), .ZN(n8798) );
  OAI21_X1 U10175 ( .B1(n8799), .B2(n10362), .A(n8798), .ZN(n8807) );
  NAND2_X1 U10176 ( .A1(n8812), .A2(n8800), .ZN(n8802) );
  XNOR2_X1 U10177 ( .A(n8802), .B(n8801), .ZN(n8805) );
  AOI222_X1 U10178 ( .A1(n10357), .A2(n8805), .B1(n8804), .B2(n8815), .C1(
        n8803), .C2(n8816), .ZN(n8954) );
  NOR2_X1 U10179 ( .A1(n8954), .A2(n8897), .ZN(n8806) );
  AOI211_X1 U10180 ( .C1(n8952), .C2(n8874), .A(n8807), .B(n8806), .ZN(n8808)
         );
  OAI21_X1 U10181 ( .B1(n8955), .B2(n8809), .A(n8808), .ZN(P2_U3278) );
  NAND2_X1 U10182 ( .A1(n8841), .A2(n8810), .ZN(n8811) );
  NAND2_X1 U10183 ( .A1(n8811), .A2(n8821), .ZN(n8813) );
  NAND3_X1 U10184 ( .A1(n8813), .A2(n10357), .A3(n8812), .ZN(n8819) );
  AOI22_X1 U10185 ( .A1(n8817), .A2(n8816), .B1(n8815), .B2(n8814), .ZN(n8818)
         );
  NAND2_X1 U10186 ( .A1(n8819), .A2(n8818), .ZN(n8956) );
  INV_X1 U10187 ( .A(n8956), .ZN(n8833) );
  OAI21_X1 U10188 ( .B1(n8822), .B2(n8821), .A(n8820), .ZN(n8958) );
  NAND2_X1 U10189 ( .A1(n8958), .A2(n10366), .ZN(n8832) );
  INV_X1 U10190 ( .A(n8823), .ZN(n8824) );
  AOI211_X1 U10191 ( .C1(n8825), .C2(n4836), .A(n10436), .B(n8824), .ZN(n8957)
         );
  NOR2_X1 U10192 ( .A1(n9013), .A2(n10362), .ZN(n8829) );
  OAI22_X1 U10193 ( .A1(n7188), .A2(n8827), .B1(n8826), .B2(n10358), .ZN(n8828) );
  AOI211_X1 U10194 ( .C1(n8957), .C2(n8830), .A(n8829), .B(n8828), .ZN(n8831)
         );
  OAI211_X1 U10195 ( .C1(n8877), .C2(n8833), .A(n8832), .B(n8831), .ZN(
        P2_U3279) );
  AND2_X1 U10196 ( .A1(n8835), .A2(n8834), .ZN(n8836) );
  OR2_X1 U10197 ( .A1(n8837), .A2(n8836), .ZN(n8965) );
  INV_X1 U10198 ( .A(n8965), .ZN(n8855) );
  NAND2_X1 U10199 ( .A1(n8839), .A2(n8838), .ZN(n8840) );
  AOI21_X1 U10200 ( .B1(n8841), .B2(n8840), .A(n8889), .ZN(n8844) );
  OAI22_X1 U10201 ( .A1(n8891), .A2(n8892), .B1(n8842), .B2(n8890), .ZN(n8843)
         );
  AOI211_X1 U10202 ( .C1(n8855), .C2(n8845), .A(n8844), .B(n8843), .ZN(n8964)
         );
  AND2_X1 U10203 ( .A1(n8867), .A2(n8850), .ZN(n8847) );
  OR2_X1 U10204 ( .A1(n8847), .A2(n8846), .ZN(n8961) );
  AOI22_X1 U10205 ( .A1(n8877), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8849), .B2(
        n8848), .ZN(n8852) );
  NAND2_X1 U10206 ( .A1(n8850), .A2(n8885), .ZN(n8851) );
  OAI211_X1 U10207 ( .C1(n8961), .C2(n10363), .A(n8852), .B(n8851), .ZN(n8853)
         );
  AOI21_X1 U10208 ( .B1(n8855), .B2(n8854), .A(n8853), .ZN(n8856) );
  OAI21_X1 U10209 ( .B1(n8964), .B2(n8897), .A(n8856), .ZN(P2_U3280) );
  INV_X1 U10210 ( .A(n8857), .ZN(n8858) );
  AOI21_X1 U10211 ( .B1(n8858), .B2(n8865), .A(n8889), .ZN(n8863) );
  OAI22_X1 U10212 ( .A1(n8860), .A2(n8892), .B1(n8859), .B2(n8890), .ZN(n8861)
         );
  AOI21_X1 U10213 ( .B1(n8863), .B2(n8862), .A(n8861), .ZN(n8970) );
  OAI21_X1 U10214 ( .B1(n8866), .B2(n8865), .A(n8864), .ZN(n8966) );
  NAND2_X1 U10215 ( .A1(n8966), .A2(n10366), .ZN(n8876) );
  INV_X1 U10216 ( .A(n8867), .ZN(n8868) );
  AOI21_X1 U10217 ( .B1(n8967), .B2(n8880), .A(n8868), .ZN(n8968) );
  INV_X1 U10218 ( .A(n8967), .ZN(n8869) );
  NOR2_X1 U10219 ( .A1(n8869), .A2(n10362), .ZN(n8873) );
  OAI22_X1 U10220 ( .A1(n7188), .A2(n8871), .B1(n8870), .B2(n10358), .ZN(n8872) );
  AOI211_X1 U10221 ( .C1(n8968), .C2(n8874), .A(n8873), .B(n8872), .ZN(n8875)
         );
  OAI211_X1 U10222 ( .C1(n8970), .C2(n8877), .A(n8876), .B(n8875), .ZN(
        P2_U3281) );
  XNOR2_X1 U10223 ( .A(n8879), .B(n8878), .ZN(n8976) );
  OAI21_X1 U10224 ( .B1(n8881), .B2(n9020), .A(n8880), .ZN(n8974) );
  NAND2_X1 U10225 ( .A1(n8877), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8882) );
  OAI21_X1 U10226 ( .B1(n10358), .B2(n8883), .A(n8882), .ZN(n8884) );
  AOI21_X1 U10227 ( .B1(n8886), .B2(n8885), .A(n8884), .ZN(n8887) );
  OAI21_X1 U10228 ( .B1(n8974), .B2(n10363), .A(n8887), .ZN(n8899) );
  AOI21_X1 U10229 ( .B1(n8888), .B2(n5040), .A(n8889), .ZN(n8896) );
  OAI22_X1 U10230 ( .A1(n8893), .A2(n8892), .B1(n8891), .B2(n8890), .ZN(n8894)
         );
  AOI21_X1 U10231 ( .B1(n8896), .B2(n8895), .A(n8894), .ZN(n8973) );
  NOR2_X1 U10232 ( .A1(n8973), .A2(n8897), .ZN(n8898) );
  AOI211_X1 U10233 ( .C1(n8976), .C2(n10366), .A(n8899), .B(n8898), .ZN(n8900)
         );
  INV_X1 U10234 ( .A(n8900), .ZN(P2_U3282) );
  AOI21_X1 U10235 ( .B1(n8902), .B2(n8951), .A(n8901), .ZN(n8987) );
  MUX2_X1 U10236 ( .A(n8903), .B(n8987), .S(n10452), .Z(n8904) );
  OAI21_X1 U10237 ( .B1(n8990), .B2(n8979), .A(n8904), .ZN(P2_U3551) );
  AOI22_X1 U10238 ( .A1(n8906), .A2(n8951), .B1(n8982), .B2(n8905), .ZN(n8907)
         );
  OAI211_X1 U10239 ( .C1(n8909), .C2(n8971), .A(n8908), .B(n8907), .ZN(n8991)
         );
  MUX2_X1 U10240 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8991), .S(n10452), .Z(
        P2_U3548) );
  INV_X1 U10241 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8913) );
  AOI211_X1 U10242 ( .C1(n8912), .C2(n10440), .A(n8911), .B(n8910), .ZN(n8992)
         );
  MUX2_X1 U10243 ( .A(n8913), .B(n8992), .S(n10452), .Z(n8914) );
  OAI21_X1 U10244 ( .B1(n8995), .B2(n8979), .A(n8914), .ZN(P2_U3546) );
  INV_X1 U10245 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8918) );
  AOI211_X1 U10246 ( .C1(n8917), .C2(n10440), .A(n8916), .B(n8915), .ZN(n8996)
         );
  MUX2_X1 U10247 ( .A(n8918), .B(n8996), .S(n10452), .Z(n8919) );
  OAI21_X1 U10248 ( .B1(n8999), .B2(n8979), .A(n8919), .ZN(P2_U3545) );
  AOI22_X1 U10249 ( .A1(n8921), .A2(n8951), .B1(n8982), .B2(n8920), .ZN(n8922)
         );
  OAI211_X1 U10250 ( .C1(n8924), .C2(n8971), .A(n8923), .B(n8922), .ZN(n9000)
         );
  MUX2_X1 U10251 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9000), .S(n10452), .Z(
        P2_U3544) );
  INV_X1 U10252 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8928) );
  AOI211_X1 U10253 ( .C1(n8927), .C2(n10440), .A(n8926), .B(n8925), .ZN(n9001)
         );
  MUX2_X1 U10254 ( .A(n8928), .B(n9001), .S(n10452), .Z(n8929) );
  OAI21_X1 U10255 ( .B1(n9004), .B2(n8979), .A(n8929), .ZN(P2_U3543) );
  AOI22_X1 U10256 ( .A1(n8931), .A2(n8951), .B1(n8982), .B2(n8930), .ZN(n8932)
         );
  OAI211_X1 U10257 ( .C1(n8934), .C2(n8971), .A(n8933), .B(n8932), .ZN(n9005)
         );
  MUX2_X1 U10258 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9005), .S(n10452), .Z(
        P2_U3542) );
  AOI22_X1 U10259 ( .A1(n8936), .A2(n8951), .B1(n8982), .B2(n8935), .ZN(n8937)
         );
  OAI211_X1 U10260 ( .C1(n8939), .C2(n8971), .A(n8938), .B(n8937), .ZN(n9006)
         );
  MUX2_X1 U10261 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9006), .S(n10452), .Z(
        P2_U3541) );
  AOI22_X1 U10262 ( .A1(n8941), .A2(n8951), .B1(n8982), .B2(n8940), .ZN(n8942)
         );
  OAI211_X1 U10263 ( .C1(n8944), .C2(n8971), .A(n8943), .B(n8942), .ZN(n9007)
         );
  MUX2_X1 U10264 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9007), .S(n10452), .Z(
        P2_U3540) );
  AOI21_X1 U10265 ( .B1(n8982), .B2(n8946), .A(n8945), .ZN(n8947) );
  OAI211_X1 U10266 ( .C1(n8949), .C2(n8971), .A(n8948), .B(n8947), .ZN(n9008)
         );
  MUX2_X1 U10267 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9008), .S(n10452), .Z(
        P2_U3539) );
  AOI22_X1 U10268 ( .A1(n8952), .A2(n8951), .B1(n8982), .B2(n8950), .ZN(n8953)
         );
  OAI211_X1 U10269 ( .C1(n8955), .C2(n8971), .A(n8954), .B(n8953), .ZN(n9009)
         );
  MUX2_X1 U10270 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9009), .S(n10452), .Z(
        P2_U3538) );
  AOI211_X1 U10271 ( .C1(n8958), .C2(n10440), .A(n8957), .B(n8956), .ZN(n9010)
         );
  MUX2_X1 U10272 ( .A(n8959), .B(n9010), .S(n10452), .Z(n8960) );
  OAI21_X1 U10273 ( .B1(n9013), .B2(n8979), .A(n8960), .ZN(P2_U3537) );
  OAI22_X1 U10274 ( .A1(n8961), .A2(n10436), .B1(n4834), .B2(n10434), .ZN(
        n8962) );
  INV_X1 U10275 ( .A(n8962), .ZN(n8963) );
  OAI211_X1 U10276 ( .C1(n10077), .C2(n8965), .A(n8964), .B(n8963), .ZN(n9014)
         );
  MUX2_X1 U10277 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9014), .S(n10452), .Z(
        P2_U3536) );
  INV_X1 U10278 ( .A(n8966), .ZN(n8972) );
  AOI22_X1 U10279 ( .A1(n8968), .A2(n8951), .B1(n8982), .B2(n8967), .ZN(n8969)
         );
  OAI211_X1 U10280 ( .C1(n8972), .C2(n8971), .A(n8970), .B(n8969), .ZN(n9015)
         );
  MUX2_X1 U10281 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9015), .S(n10452), .Z(
        P2_U3535) );
  OAI21_X1 U10282 ( .B1(n10436), .B2(n8974), .A(n8973), .ZN(n8975) );
  AOI21_X1 U10283 ( .B1(n8976), .B2(n10440), .A(n8975), .ZN(n9016) );
  MUX2_X1 U10284 ( .A(n8977), .B(n9016), .S(n10452), .Z(n8978) );
  OAI21_X1 U10285 ( .B1(n9020), .B2(n8979), .A(n8978), .ZN(P2_U3534) );
  INV_X1 U10286 ( .A(n8980), .ZN(n8986) );
  AOI22_X1 U10287 ( .A1(n8983), .A2(n8951), .B1(n8982), .B2(n8981), .ZN(n8984)
         );
  OAI211_X1 U10288 ( .C1(n10077), .C2(n8986), .A(n8985), .B(n8984), .ZN(n9021)
         );
  MUX2_X1 U10289 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9021), .S(n10452), .Z(
        P2_U3530) );
  MUX2_X1 U10290 ( .A(n8988), .B(n8987), .S(n10444), .Z(n8989) );
  OAI21_X1 U10291 ( .B1(n8990), .B2(n9019), .A(n8989), .ZN(P2_U3519) );
  MUX2_X1 U10292 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8991), .S(n10444), .Z(
        P2_U3516) );
  MUX2_X1 U10293 ( .A(n8993), .B(n8992), .S(n10444), .Z(n8994) );
  OAI21_X1 U10294 ( .B1(n8995), .B2(n9019), .A(n8994), .ZN(P2_U3514) );
  MUX2_X1 U10295 ( .A(n8997), .B(n8996), .S(n10444), .Z(n8998) );
  OAI21_X1 U10296 ( .B1(n8999), .B2(n9019), .A(n8998), .ZN(P2_U3513) );
  MUX2_X1 U10297 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9000), .S(n10444), .Z(
        P2_U3512) );
  INV_X1 U10298 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9002) );
  MUX2_X1 U10299 ( .A(n9002), .B(n9001), .S(n10444), .Z(n9003) );
  OAI21_X1 U10300 ( .B1(n9004), .B2(n9019), .A(n9003), .ZN(P2_U3511) );
  MUX2_X1 U10301 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9005), .S(n10444), .Z(
        P2_U3510) );
  MUX2_X1 U10302 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9006), .S(n10444), .Z(
        P2_U3509) );
  MUX2_X1 U10303 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9007), .S(n10444), .Z(
        P2_U3508) );
  MUX2_X1 U10304 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9008), .S(n10444), .Z(
        P2_U3507) );
  MUX2_X1 U10305 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9009), .S(n10444), .Z(
        P2_U3505) );
  MUX2_X1 U10306 ( .A(n9011), .B(n9010), .S(n10444), .Z(n9012) );
  OAI21_X1 U10307 ( .B1(n9013), .B2(n9019), .A(n9012), .ZN(P2_U3502) );
  MUX2_X1 U10308 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9014), .S(n10444), .Z(
        P2_U3499) );
  MUX2_X1 U10309 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9015), .S(n10444), .Z(
        P2_U3496) );
  INV_X1 U10310 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9017) );
  MUX2_X1 U10311 ( .A(n9017), .B(n9016), .S(n10444), .Z(n9018) );
  OAI21_X1 U10312 ( .B1(n9020), .B2(n9019), .A(n9018), .ZN(P2_U3493) );
  MUX2_X1 U10313 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n9021), .S(n10444), .Z(
        P2_U3481) );
  NOR4_X1 U10314 ( .A1(n9023), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9022), .A4(
        P2_U3152), .ZN(n9024) );
  AOI21_X1 U10315 ( .B1(n9030), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9024), .ZN(
        n9025) );
  OAI21_X1 U10316 ( .B1(n9619), .B2(n6706), .A(n9025), .ZN(P2_U3327) );
  INV_X1 U10317 ( .A(n9026), .ZN(n9620) );
  AOI22_X1 U10318 ( .A1(n9027), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9030), .ZN(n9028) );
  OAI21_X1 U10319 ( .B1(n9620), .B2(n6706), .A(n9028), .ZN(P2_U3328) );
  INV_X1 U10320 ( .A(n9029), .ZN(n9623) );
  AOI22_X1 U10321 ( .A1(n9031), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9030), .ZN(n9032) );
  OAI21_X1 U10322 ( .B1(n9623), .B2(n6706), .A(n9032), .ZN(P2_U3329) );
  MUX2_X1 U10323 ( .A(n9033), .B(n10355), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3358) );
  INV_X1 U10324 ( .A(n9550), .ZN(n9363) );
  INV_X1 U10325 ( .A(n9034), .ZN(n9038) );
  OAI21_X1 U10326 ( .B1(n9036), .B2(n9098), .A(n9035), .ZN(n9037) );
  OAI211_X1 U10327 ( .C1(n9038), .C2(n9098), .A(n10101), .B(n9037), .ZN(n9043)
         );
  INV_X1 U10328 ( .A(n9039), .ZN(n9361) );
  AOI22_X1 U10329 ( .A1(n9366), .A2(n10090), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9040) );
  OAI21_X1 U10330 ( .B1(n9234), .B2(n10092), .A(n9040), .ZN(n9041) );
  AOI21_X1 U10331 ( .B1(n9361), .B2(n9143), .A(n9041), .ZN(n9042) );
  OAI211_X1 U10332 ( .C1(n9363), .C2(n9146), .A(n9043), .B(n9042), .ZN(
        P1_U3214) );
  NAND2_X1 U10333 ( .A1(n9046), .A2(n9045), .ZN(n9047) );
  XNOR2_X1 U10334 ( .A(n9044), .B(n9047), .ZN(n9052) );
  INV_X1 U10335 ( .A(n9437), .ZN(n9468) );
  NAND2_X1 U10336 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9202) );
  OAI21_X1 U10337 ( .B1(n10092), .B2(n9438), .A(n9202), .ZN(n9048) );
  AOI21_X1 U10338 ( .B1(n10090), .B2(n9468), .A(n9048), .ZN(n9049) );
  OAI21_X1 U10339 ( .B1(n10106), .B2(n9430), .A(n9049), .ZN(n9050) );
  AOI21_X1 U10340 ( .B1(n9573), .B2(n10095), .A(n9050), .ZN(n9051) );
  OAI21_X1 U10341 ( .B1(n9052), .B2(n9156), .A(n9051), .ZN(P1_U3217) );
  XOR2_X1 U10342 ( .A(n9054), .B(n9053), .Z(n9059) );
  AOI22_X1 U10343 ( .A1(n9366), .A2(n9152), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9056) );
  NAND2_X1 U10344 ( .A1(n9143), .A2(n9406), .ZN(n9055) );
  OAI211_X1 U10345 ( .C1(n9438), .C2(n10061), .A(n9056), .B(n9055), .ZN(n9057)
         );
  AOI21_X1 U10346 ( .B1(n9563), .B2(n10095), .A(n9057), .ZN(n9058) );
  OAI21_X1 U10347 ( .B1(n9059), .B2(n9156), .A(n9058), .ZN(P1_U3221) );
  AOI21_X1 U10348 ( .B1(n4494), .B2(n9061), .A(n9137), .ZN(n9067) );
  NOR2_X1 U10349 ( .A1(n9333), .A2(n10106), .ZN(n9064) );
  OAI22_X1 U10350 ( .A1(n9234), .A2(n10061), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9062), .ZN(n9063) );
  AOI211_X1 U10351 ( .C1(n9152), .C2(n9339), .A(n9064), .B(n9063), .ZN(n9066)
         );
  NAND2_X1 U10352 ( .A1(n9540), .A2(n10095), .ZN(n9065) );
  OAI211_X1 U10353 ( .C1(n9067), .C2(n9156), .A(n9066), .B(n9065), .ZN(
        P1_U3223) );
  INV_X1 U10354 ( .A(n9069), .ZN(n9070) );
  AOI21_X1 U10355 ( .B1(n9068), .B2(n9071), .A(n9070), .ZN(n9076) );
  INV_X1 U10356 ( .A(n9483), .ZN(n9485) );
  NOR2_X1 U10357 ( .A1(n9485), .A2(n10323), .ZN(n9590) );
  NOR2_X1 U10358 ( .A1(n10106), .A2(n9486), .ZN(n9074) );
  NAND2_X1 U10359 ( .A1(n10090), .A2(n9220), .ZN(n9072) );
  NAND2_X1 U10360 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10218)
         );
  OAI211_X1 U10361 ( .C1(n9478), .C2(n10092), .A(n9072), .B(n10218), .ZN(n9073) );
  AOI211_X1 U10362 ( .C1(n9590), .C2(n10067), .A(n9074), .B(n9073), .ZN(n9075)
         );
  OAI21_X1 U10363 ( .B1(n9076), .B2(n9156), .A(n9075), .ZN(P1_U3224) );
  OAI21_X1 U10364 ( .B1(n9079), .B2(n9078), .A(n9077), .ZN(n9080) );
  NAND2_X1 U10365 ( .A1(n9080), .A2(n10101), .ZN(n9088) );
  NOR2_X1 U10366 ( .A1(n10323), .A2(n9081), .ZN(n10301) );
  AOI22_X1 U10367 ( .A1(n10090), .A2(n9166), .B1(n10301), .B2(n10067), .ZN(
        n9087) );
  NOR2_X1 U10368 ( .A1(n10092), .A2(n9082), .ZN(n9083) );
  AOI211_X1 U10369 ( .C1(n9085), .C2(n9143), .A(n9084), .B(n9083), .ZN(n9086)
         );
  NAND3_X1 U10370 ( .A1(n9088), .A2(n9087), .A3(n9086), .ZN(P1_U3225) );
  OAI21_X1 U10371 ( .B1(n9091), .B2(n9090), .A(n9089), .ZN(n9092) );
  NAND2_X1 U10372 ( .A1(n9092), .A2(n10101), .ZN(n9096) );
  INV_X1 U10373 ( .A(n9496), .ZN(n9467) );
  NAND2_X1 U10374 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10230)
         );
  OAI21_X1 U10375 ( .B1(n10092), .B2(n9437), .A(n10230), .ZN(n9094) );
  NOR2_X1 U10376 ( .A1(n10106), .A2(n9461), .ZN(n9093) );
  AOI211_X1 U10377 ( .C1(n10090), .C2(n9467), .A(n9094), .B(n9093), .ZN(n9095)
         );
  OAI211_X1 U10378 ( .C1(n9464), .C2(n9146), .A(n9096), .B(n9095), .ZN(
        P1_U3226) );
  OAI21_X1 U10379 ( .B1(n9034), .B2(n9098), .A(n9097), .ZN(n9099) );
  INV_X1 U10380 ( .A(n9099), .ZN(n9100) );
  OAI21_X1 U10381 ( .B1(n9101), .B2(n9100), .A(n10101), .ZN(n9106) );
  OAI22_X1 U10382 ( .A1(n9349), .A2(n10061), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9102), .ZN(n9104) );
  NOR2_X1 U10383 ( .A1(n9350), .A2(n10092), .ZN(n9103) );
  AOI211_X1 U10384 ( .C1(n9353), .C2(n9143), .A(n9104), .B(n9103), .ZN(n9105)
         );
  OAI211_X1 U10385 ( .C1(n9356), .C2(n9146), .A(n9106), .B(n9105), .ZN(
        P1_U3227) );
  NAND2_X1 U10386 ( .A1(n9109), .A2(n9108), .ZN(n9110) );
  XNOR2_X1 U10387 ( .A(n9107), .B(n9110), .ZN(n9116) );
  OAI22_X1 U10388 ( .A1(n10092), .A2(n9377), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9111), .ZN(n9112) );
  AOI21_X1 U10389 ( .B1(n10090), .B2(n9421), .A(n9112), .ZN(n9113) );
  OAI21_X1 U10390 ( .B1(n10106), .B2(n9415), .A(n9113), .ZN(n9114) );
  AOI21_X1 U10391 ( .B1(n9566), .B2(n10095), .A(n9114), .ZN(n9115) );
  OAI21_X1 U10392 ( .B1(n9116), .B2(n9156), .A(n9115), .ZN(P1_U3231) );
  NAND2_X1 U10393 ( .A1(n9118), .A2(n9117), .ZN(n9120) );
  XNOR2_X1 U10394 ( .A(n9120), .B(n9119), .ZN(n9125) );
  NOR2_X1 U10395 ( .A1(n9230), .A2(n10323), .ZN(n9556) );
  AOI22_X1 U10396 ( .A1(n10090), .A2(n9422), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9122) );
  NAND2_X1 U10397 ( .A1(n9375), .A2(n9152), .ZN(n9121) );
  OAI211_X1 U10398 ( .C1(n10106), .C2(n9383), .A(n9122), .B(n9121), .ZN(n9123)
         );
  AOI21_X1 U10399 ( .B1(n9556), .B2(n10067), .A(n9123), .ZN(n9124) );
  OAI21_X1 U10400 ( .B1(n9125), .B2(n9156), .A(n9124), .ZN(P1_U3233) );
  NAND2_X1 U10401 ( .A1(n9127), .A2(n9126), .ZN(n9129) );
  XNOR2_X1 U10402 ( .A(n9129), .B(n9128), .ZN(n9134) );
  NAND2_X1 U10403 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10244)
         );
  OAI21_X1 U10404 ( .B1(n10092), .B2(n9454), .A(n10244), .ZN(n9130) );
  AOI21_X1 U10405 ( .B1(n10090), .B2(n9223), .A(n9130), .ZN(n9131) );
  OAI21_X1 U10406 ( .B1(n10106), .B2(n9446), .A(n9131), .ZN(n9132) );
  AOI21_X1 U10407 ( .B1(n9578), .B2(n10095), .A(n9132), .ZN(n9133) );
  OAI21_X1 U10408 ( .B1(n9134), .B2(n9156), .A(n9133), .ZN(P1_U3236) );
  OAI21_X1 U10409 ( .B1(n9137), .B2(n9136), .A(n9135), .ZN(n9138) );
  NAND3_X1 U10410 ( .A1(n9139), .A2(n10101), .A3(n9138), .ZN(n9145) );
  OAI22_X1 U10411 ( .A1(n9350), .A2(n10061), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9140), .ZN(n9142) );
  NOR2_X1 U10412 ( .A1(n9239), .A2(n10092), .ZN(n9141) );
  AOI211_X1 U10413 ( .C1(n9321), .C2(n9143), .A(n9142), .B(n9141), .ZN(n9144)
         );
  OAI211_X1 U10414 ( .C1(n9313), .C2(n9146), .A(n9145), .B(n9144), .ZN(
        P1_U3238) );
  XNOR2_X1 U10415 ( .A(n9149), .B(n9148), .ZN(n9150) );
  XNOR2_X1 U10416 ( .A(n9147), .B(n9150), .ZN(n9157) );
  NAND2_X1 U10417 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10207)
         );
  OAI21_X1 U10418 ( .B1(n10061), .B2(n10109), .A(n10207), .ZN(n9151) );
  AOI21_X1 U10419 ( .B1(n9152), .B2(n9467), .A(n9151), .ZN(n9153) );
  OAI21_X1 U10420 ( .B1(n10106), .B2(n9506), .A(n9153), .ZN(n9154) );
  AOI21_X1 U10421 ( .B1(n9510), .B2(n10095), .A(n9154), .ZN(n9155) );
  OAI21_X1 U10422 ( .B1(n9157), .B2(n9156), .A(n9155), .ZN(P1_U3239) );
  MUX2_X1 U10423 ( .A(n9158), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9159), .Z(
        P1_U3585) );
  MUX2_X1 U10424 ( .A(n9294), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9159), .Z(
        P1_U3584) );
  MUX2_X1 U10425 ( .A(n9307), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9159), .Z(
        P1_U3583) );
  MUX2_X1 U10426 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9317), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10427 ( .A(n9339), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9159), .Z(
        P1_U3581) );
  MUX2_X1 U10428 ( .A(n9316), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9159), .Z(
        P1_U3580) );
  MUX2_X1 U10429 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9367), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10430 ( .A(n9375), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9159), .Z(
        P1_U3578) );
  MUX2_X1 U10431 ( .A(n9366), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9159), .Z(
        P1_U3577) );
  MUX2_X1 U10432 ( .A(n9422), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9159), .Z(
        P1_U3576) );
  MUX2_X1 U10433 ( .A(n9226), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9159), .Z(
        P1_U3575) );
  MUX2_X1 U10434 ( .A(n9421), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9159), .Z(
        P1_U3574) );
  MUX2_X1 U10435 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9468), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10436 ( .A(n9223), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9159), .Z(
        P1_U3572) );
  MUX2_X1 U10437 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9467), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10438 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9220), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10439 ( .A(n9217), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9159), .Z(
        P1_U3569) );
  MUX2_X1 U10440 ( .A(n10089), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9159), .Z(
        P1_U3568) );
  MUX2_X1 U10441 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9160), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10442 ( .A(n9161), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9159), .Z(
        P1_U3566) );
  MUX2_X1 U10443 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n10265), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10444 ( .A(n9162), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9159), .Z(
        P1_U3564) );
  MUX2_X1 U10445 ( .A(n10262), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9159), .Z(
        P1_U3563) );
  MUX2_X1 U10446 ( .A(n9163), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9159), .Z(
        P1_U3562) );
  MUX2_X1 U10447 ( .A(n9164), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9159), .Z(
        P1_U3561) );
  MUX2_X1 U10448 ( .A(n9165), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9159), .Z(
        P1_U3560) );
  MUX2_X1 U10449 ( .A(n9166), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9159), .Z(
        P1_U3559) );
  MUX2_X1 U10450 ( .A(n9167), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9159), .Z(
        P1_U3558) );
  MUX2_X1 U10451 ( .A(n9168), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9159), .Z(
        P1_U3557) );
  MUX2_X1 U10452 ( .A(n7062), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9159), .Z(
        P1_U3556) );
  NAND2_X1 U10453 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n10187), .ZN(n9170) );
  OAI21_X1 U10454 ( .B1(n10187), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9170), .ZN(
        n10183) );
  NOR2_X1 U10455 ( .A1(n9171), .A2(n9184), .ZN(n9172) );
  NOR2_X1 U10456 ( .A1(n7906), .A2(n10196), .ZN(n10195) );
  NOR2_X1 U10457 ( .A1(n9172), .A2(n10195), .ZN(n9173) );
  NOR2_X1 U10458 ( .A1(n9173), .A2(n9186), .ZN(n9174) );
  NAND2_X1 U10459 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n10223), .ZN(n9175) );
  OAI21_X1 U10460 ( .B1(n10223), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9175), .ZN(
        n10220) );
  AOI21_X1 U10461 ( .B1(n10223), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10219), 
        .ZN(n10233) );
  NAND2_X1 U10462 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n10236), .ZN(n9176) );
  OAI21_X1 U10463 ( .B1(n10236), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9176), .ZN(
        n10232) );
  NOR2_X1 U10464 ( .A1(n10233), .A2(n10232), .ZN(n10231) );
  MUX2_X1 U10465 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n9447), .S(n10252), .Z(
        n9177) );
  INV_X1 U10466 ( .A(n9177), .ZN(n10247) );
  NOR2_X1 U10467 ( .A1(n10248), .A2(n10247), .ZN(n10246) );
  AOI21_X1 U10468 ( .B1(n10252), .B2(P1_REG2_REG_18__SCAN_IN), .A(n10246), 
        .ZN(n9178) );
  XNOR2_X1 U10469 ( .A(n10252), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n10255) );
  INV_X1 U10470 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9190) );
  XNOR2_X1 U10471 ( .A(n9191), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10240) );
  XOR2_X1 U10472 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10223), .Z(n10225) );
  NOR2_X1 U10473 ( .A1(n9179), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9180) );
  NOR2_X1 U10474 ( .A1(n9181), .A2(n9180), .ZN(n10190) );
  MUX2_X1 U10475 ( .A(n9182), .B(P1_REG1_REG_13__SCAN_IN), .S(n10187), .Z(
        n10189) );
  NOR2_X1 U10476 ( .A1(n10190), .A2(n10189), .ZN(n10188) );
  AOI21_X1 U10477 ( .B1(n4633), .B2(n9182), .A(n10188), .ZN(n10201) );
  MUX2_X1 U10478 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9183), .S(n9184), .Z(
        n10202) );
  NOR2_X1 U10479 ( .A1(n10201), .A2(n10202), .ZN(n10200) );
  AOI21_X1 U10480 ( .B1(n9184), .B2(n9183), .A(n10200), .ZN(n9185) );
  NAND2_X1 U10481 ( .A1(n10212), .A2(n9185), .ZN(n9187) );
  XNOR2_X1 U10482 ( .A(n9186), .B(n9185), .ZN(n10214) );
  NAND2_X1 U10483 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n10214), .ZN(n10213) );
  NAND2_X1 U10484 ( .A1(n9187), .A2(n10213), .ZN(n10226) );
  NAND2_X1 U10485 ( .A1(n10225), .A2(n10226), .ZN(n10224) );
  OAI21_X1 U10486 ( .B1(n9189), .B2(n9188), .A(n10224), .ZN(n10239) );
  NAND2_X1 U10487 ( .A1(n10240), .A2(n10239), .ZN(n10237) );
  OAI21_X1 U10488 ( .B1(n9191), .B2(n9190), .A(n10237), .ZN(n10254) );
  NOR2_X1 U10489 ( .A1(n10255), .A2(n10254), .ZN(n10253) );
  AOI21_X1 U10490 ( .B1(n9193), .B2(n9192), .A(n10253), .ZN(n9194) );
  XNOR2_X1 U10491 ( .A(n9194), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9197) );
  NAND2_X1 U10492 ( .A1(n9196), .A2(n9195), .ZN(n9199) );
  AOI21_X1 U10493 ( .B1(n9197), .B2(n10238), .A(n10251), .ZN(n9198) );
  NAND2_X1 U10494 ( .A1(n9199), .A2(n9198), .ZN(n9201) );
  INV_X1 U10495 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9203) );
  OAI21_X1 U10496 ( .B1(n10260), .B2(n9203), .A(n9202), .ZN(n9204) );
  INV_X1 U10497 ( .A(n9523), .ZN(n9276) );
  OR2_X2 U10498 ( .A1(n9458), .A2(n9578), .ZN(n9443) );
  NOR2_X1 U10499 ( .A1(n9443), .A2(n9573), .ZN(n9428) );
  AND2_X2 U10500 ( .A1(n9360), .A2(n9356), .ZN(n9351) );
  INV_X1 U10501 ( .A(n9540), .ZN(n9336) );
  NAND2_X1 U10502 ( .A1(n9276), .A2(n9283), .ZN(n9272) );
  NOR2_X1 U10503 ( .A1(n10146), .A2(n9272), .ZN(n9205) );
  XNOR2_X1 U10504 ( .A(n9206), .B(n9205), .ZN(n9518) );
  NAND2_X1 U10505 ( .A1(n9207), .A2(P1_B_REG_SCAN_IN), .ZN(n9208) );
  NAND2_X1 U10506 ( .A1(n10264), .A2(n9208), .ZN(n9271) );
  NOR2_X1 U10507 ( .A1(n9271), .A2(n9209), .ZN(n10145) );
  NAND2_X1 U10508 ( .A1(n9508), .A2(n10145), .ZN(n9213) );
  OAI21_X1 U10509 ( .B1(n9508), .B2(n9210), .A(n9213), .ZN(n9211) );
  AOI21_X1 U10510 ( .B1(n9516), .B2(n10276), .A(n9211), .ZN(n9212) );
  OAI21_X1 U10511 ( .B1(n9518), .B2(n9512), .A(n9212), .ZN(P1_U3261) );
  XNOR2_X1 U10512 ( .A(n10146), .B(n9272), .ZN(n10143) );
  OAI21_X1 U10513 ( .B1(n9508), .B2(n9214), .A(n9213), .ZN(n9215) );
  AOI21_X1 U10514 ( .B1(n10146), .B2(n10276), .A(n9215), .ZN(n9216) );
  OAI21_X1 U10515 ( .B1(n10143), .B2(n9512), .A(n9216), .ZN(P1_U3262) );
  AND2_X1 U10516 ( .A1(n10096), .A2(n9217), .ZN(n9218) );
  OAI22_X2 U10517 ( .A1(n9219), .A2(n9218), .B1(n9217), .B2(n10096), .ZN(n9498) );
  OAI21_X1 U10518 ( .B1(n9592), .B2(n10093), .A(n9498), .ZN(n9222) );
  NAND2_X1 U10519 ( .A1(n9222), .A2(n9221), .ZN(n9480) );
  NOR2_X1 U10520 ( .A1(n9581), .A2(n9223), .ZN(n9224) );
  NOR2_X1 U10521 ( .A1(n9573), .A2(n9421), .ZN(n9225) );
  INV_X1 U10522 ( .A(n9573), .ZN(n9429) );
  INV_X1 U10523 ( .A(n9412), .ZN(n9229) );
  NAND2_X1 U10524 ( .A1(n9566), .A2(n9226), .ZN(n9228) );
  AOI21_X1 U10525 ( .B1(n9229), .B2(n9228), .A(n9227), .ZN(n9394) );
  NAND2_X1 U10526 ( .A1(n9394), .A2(n9400), .ZN(n9393) );
  OAI21_X1 U10527 ( .B1(n9377), .B2(n9409), .A(n9393), .ZN(n9381) );
  NAND2_X1 U10528 ( .A1(n9230), .A2(n9402), .ZN(n9231) );
  NAND2_X1 U10529 ( .A1(n9550), .A2(n9375), .ZN(n9233) );
  NOR2_X1 U10530 ( .A1(n9550), .A2(n9375), .ZN(n9232) );
  NAND2_X1 U10531 ( .A1(n9356), .A2(n9234), .ZN(n9236) );
  NOR2_X1 U10532 ( .A1(n9356), .A2(n9234), .ZN(n9235) );
  NAND2_X1 U10533 ( .A1(n9328), .A2(n9337), .ZN(n9327) );
  NAND2_X1 U10534 ( .A1(n9327), .A2(n9237), .ZN(n9312) );
  INV_X1 U10535 ( .A(n9312), .ZN(n9238) );
  XNOR2_X1 U10536 ( .A(n9240), .B(n9267), .ZN(n9519) );
  INV_X1 U10537 ( .A(n9519), .ZN(n9280) );
  NAND2_X1 U10538 ( .A1(n9242), .A2(n9241), .ZN(n9495) );
  NAND2_X1 U10539 ( .A1(n9495), .A2(n9243), .ZN(n9474) );
  NAND2_X1 U10540 ( .A1(n9474), .A2(n9244), .ZN(n9246) );
  NAND2_X1 U10541 ( .A1(n9434), .A2(n9435), .ZN(n9251) );
  NOR2_X1 U10542 ( .A1(n9400), .A2(n9253), .ZN(n9254) );
  INV_X1 U10543 ( .A(n9258), .ZN(n9259) );
  INV_X1 U10544 ( .A(n9260), .ZN(n9261) );
  NAND2_X1 U10545 ( .A1(n9306), .A2(n9299), .ZN(n9288) );
  NAND3_X1 U10546 ( .A1(n9288), .A2(n9265), .A3(n9264), .ZN(n9293) );
  NAND2_X1 U10547 ( .A1(n9293), .A2(n9266), .ZN(n9268) );
  OAI21_X1 U10548 ( .B1(n9276), .B2(n9283), .A(n9272), .ZN(n9520) );
  NOR2_X1 U10549 ( .A1(n9520), .A2(n9512), .ZN(n9278) );
  INV_X1 U10550 ( .A(n9273), .ZN(n9274) );
  AOI22_X1 U10551 ( .A1(n9274), .A2(n10275), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n4483), .ZN(n9275) );
  OAI21_X1 U10552 ( .B1(n9276), .B2(n9484), .A(n9275), .ZN(n9277) );
  AOI211_X1 U10553 ( .C1(n9521), .C2(n9508), .A(n9278), .B(n9277), .ZN(n9279)
         );
  OAI21_X1 U10554 ( .B1(n9280), .B2(n9481), .A(n9279), .ZN(P1_U3355) );
  OAI21_X1 U10555 ( .B1(n9282), .B2(n9289), .A(n9281), .ZN(n9529) );
  AOI211_X1 U10556 ( .C1(n9284), .C2(n4895), .A(n10325), .B(n9283), .ZN(n9526)
         );
  AOI22_X1 U10557 ( .A1(n9285), .A2(n10275), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n4483), .ZN(n9286) );
  OAI21_X1 U10558 ( .B1(n9287), .B2(n9484), .A(n9286), .ZN(n9297) );
  INV_X1 U10559 ( .A(n9288), .ZN(n9291) );
  OAI21_X1 U10560 ( .B1(n9291), .B2(n9290), .A(n9289), .ZN(n9292) );
  NAND2_X1 U10561 ( .A1(n9293), .A2(n9292), .ZN(n9295) );
  AOI222_X1 U10562 ( .A1(n10266), .A2(n9295), .B1(n9294), .B2(n10264), .C1(
        n9317), .C2(n10263), .ZN(n9528) );
  NOR2_X1 U10563 ( .A1(n9528), .A2(n4483), .ZN(n9296) );
  AOI211_X1 U10564 ( .C1(n9490), .C2(n9526), .A(n9297), .B(n9296), .ZN(n9298)
         );
  OAI21_X1 U10565 ( .B1(n9529), .B2(n9481), .A(n9298), .ZN(P1_U3263) );
  XNOR2_X2 U10566 ( .A(n9300), .B(n9299), .ZN(n9534) );
  AOI211_X1 U10567 ( .C1(n9531), .C2(n9319), .A(n10325), .B(n9301), .ZN(n9530)
         );
  AOI22_X1 U10568 ( .A1(n9302), .A2(n10275), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n4483), .ZN(n9303) );
  OAI21_X1 U10569 ( .B1(n9304), .B2(n9484), .A(n9303), .ZN(n9310) );
  XNOR2_X1 U10570 ( .A(n9306), .B(n9305), .ZN(n9308) );
  AOI222_X1 U10571 ( .A1(n10266), .A2(n9308), .B1(n9307), .B2(n10264), .C1(
        n9339), .C2(n10263), .ZN(n9533) );
  NOR2_X1 U10572 ( .A1(n9533), .A2(n4483), .ZN(n9309) );
  AOI211_X1 U10573 ( .C1(n9530), .C2(n9490), .A(n9310), .B(n9309), .ZN(n9311)
         );
  OAI21_X1 U10574 ( .B1(n9534), .B2(n9481), .A(n9311), .ZN(P1_U3264) );
  XNOR2_X1 U10575 ( .A(n9312), .B(n9314), .ZN(n9539) );
  NOR2_X1 U10576 ( .A1(n9313), .A2(n9484), .ZN(n9325) );
  XNOR2_X1 U10577 ( .A(n9315), .B(n9314), .ZN(n9318) );
  AOI222_X1 U10578 ( .A1(n10266), .A2(n9318), .B1(n9317), .B2(n10264), .C1(
        n9316), .C2(n10263), .ZN(n9538) );
  INV_X1 U10579 ( .A(n9319), .ZN(n9320) );
  AOI211_X1 U10580 ( .C1(n9536), .C2(n9330), .A(n10325), .B(n9320), .ZN(n9535)
         );
  AOI22_X1 U10581 ( .A1(n9535), .A2(n9322), .B1(n10275), .B2(n9321), .ZN(n9323) );
  AOI21_X1 U10582 ( .B1(n9538), .B2(n9323), .A(n4483), .ZN(n9324) );
  AOI211_X1 U10583 ( .C1(n4483), .C2(P1_REG2_REG_26__SCAN_IN), .A(n9325), .B(
        n9324), .ZN(n9326) );
  OAI21_X1 U10584 ( .B1(n9539), .B2(n9481), .A(n9326), .ZN(P1_U3265) );
  OAI21_X1 U10585 ( .B1(n9328), .B2(n9337), .A(n9327), .ZN(n9329) );
  INV_X1 U10586 ( .A(n9329), .ZN(n9544) );
  INV_X1 U10587 ( .A(n9351), .ZN(n9332) );
  INV_X1 U10588 ( .A(n9330), .ZN(n9331) );
  AOI21_X1 U10589 ( .B1(n9540), .B2(n9332), .A(n9331), .ZN(n9541) );
  INV_X1 U10590 ( .A(n9333), .ZN(n9334) );
  AOI22_X1 U10591 ( .A1(n9334), .A2(n10275), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n4483), .ZN(n9335) );
  OAI21_X1 U10592 ( .B1(n9336), .B2(n9484), .A(n9335), .ZN(n9342) );
  XNOR2_X1 U10593 ( .A(n9338), .B(n9337), .ZN(n9340) );
  AOI222_X1 U10594 ( .A1(n10266), .A2(n9340), .B1(n9339), .B2(n10264), .C1(
        n9367), .C2(n10263), .ZN(n9543) );
  NOR2_X1 U10595 ( .A1(n9543), .A2(n4483), .ZN(n9341) );
  AOI211_X1 U10596 ( .C1(n9541), .C2(n10282), .A(n9342), .B(n9341), .ZN(n9343)
         );
  OAI21_X1 U10597 ( .B1(n9544), .B2(n9481), .A(n9343), .ZN(P1_U3266) );
  XNOR2_X1 U10598 ( .A(n9344), .B(n9347), .ZN(n9549) );
  AOI21_X1 U10599 ( .B1(n9347), .B2(n9346), .A(n9345), .ZN(n9348) );
  OAI222_X1 U10600 ( .A1(n10128), .A2(n9350), .B1(n10129), .B2(n9349), .C1(
        n9477), .C2(n9348), .ZN(n9545) );
  INV_X1 U10601 ( .A(n9360), .ZN(n9352) );
  AOI211_X1 U10602 ( .C1(n9547), .C2(n9352), .A(n10325), .B(n9351), .ZN(n9546)
         );
  NAND2_X1 U10603 ( .A1(n9546), .A2(n9490), .ZN(n9355) );
  AOI22_X1 U10604 ( .A1(n9353), .A2(n10275), .B1(n4483), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n9354) );
  OAI211_X1 U10605 ( .C1(n9356), .C2(n9484), .A(n9355), .B(n9354), .ZN(n9357)
         );
  AOI21_X1 U10606 ( .B1(n9545), .B2(n9508), .A(n9357), .ZN(n9358) );
  OAI21_X1 U10607 ( .B1(n9549), .B2(n9481), .A(n9358), .ZN(P1_U3267) );
  XOR2_X1 U10608 ( .A(n9365), .B(n9359), .Z(n9554) );
  AOI21_X1 U10609 ( .B1(n9550), .B2(n9385), .A(n9360), .ZN(n9551) );
  AOI22_X1 U10610 ( .A1(P1_REG2_REG_23__SCAN_IN), .A2(n4483), .B1(n9361), .B2(
        n10275), .ZN(n9362) );
  OAI21_X1 U10611 ( .B1(n9363), .B2(n9484), .A(n9362), .ZN(n9370) );
  XOR2_X1 U10612 ( .A(n9365), .B(n9364), .Z(n9368) );
  AOI222_X1 U10613 ( .A1(n10266), .A2(n9368), .B1(n9367), .B2(n10264), .C1(
        n9366), .C2(n10263), .ZN(n9553) );
  NOR2_X1 U10614 ( .A1(n9553), .A2(n4483), .ZN(n9369) );
  AOI211_X1 U10615 ( .C1(n9551), .C2(n10282), .A(n9370), .B(n9369), .ZN(n9371)
         );
  OAI21_X1 U10616 ( .B1(n9554), .B2(n9481), .A(n9371), .ZN(P1_U3268) );
  NAND2_X1 U10617 ( .A1(n9397), .A2(n9372), .ZN(n9374) );
  INV_X1 U10618 ( .A(n9380), .ZN(n9373) );
  XNOR2_X1 U10619 ( .A(n9374), .B(n9373), .ZN(n9379) );
  NAND2_X1 U10620 ( .A1(n9375), .A2(n10264), .ZN(n9376) );
  OAI21_X1 U10621 ( .B1(n9377), .B2(n10129), .A(n9376), .ZN(n9378) );
  AOI21_X1 U10622 ( .B1(n9379), .B2(n10266), .A(n9378), .ZN(n9559) );
  XOR2_X1 U10623 ( .A(n9381), .B(n9380), .Z(n9555) );
  NAND2_X1 U10624 ( .A1(n9555), .A2(n9382), .ZN(n9392) );
  INV_X1 U10625 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9384) );
  OAI22_X1 U10626 ( .A1(n9508), .A2(n9384), .B1(n9383), .B2(n9505), .ZN(n9389)
         );
  AOI21_X1 U10627 ( .B1(n9403), .B2(n9390), .A(n10325), .ZN(n9386) );
  NAND2_X1 U10628 ( .A1(n9386), .A2(n9385), .ZN(n9557) );
  NOR2_X1 U10629 ( .A1(n9557), .A2(n9387), .ZN(n9388) );
  AOI211_X1 U10630 ( .C1(n10276), .C2(n9390), .A(n9389), .B(n9388), .ZN(n9391)
         );
  OAI211_X1 U10631 ( .C1(n4483), .C2(n9559), .A(n9392), .B(n9391), .ZN(
        P1_U3269) );
  OAI21_X1 U10632 ( .B1(n9394), .B2(n9400), .A(n9393), .ZN(n9565) );
  NAND2_X1 U10633 ( .A1(n9396), .A2(n9395), .ZN(n9399) );
  INV_X1 U10634 ( .A(n9397), .ZN(n9398) );
  AOI21_X1 U10635 ( .B1(n9400), .B2(n9399), .A(n9398), .ZN(n9401) );
  OAI222_X1 U10636 ( .A1(n10128), .A2(n9402), .B1(n10129), .B2(n9438), .C1(
        n9477), .C2(n9401), .ZN(n9561) );
  INV_X1 U10637 ( .A(n9413), .ZN(n9405) );
  INV_X1 U10638 ( .A(n9403), .ZN(n9404) );
  AOI211_X1 U10639 ( .C1(n9563), .C2(n9405), .A(n10325), .B(n9404), .ZN(n9562)
         );
  NAND2_X1 U10640 ( .A1(n9562), .A2(n9490), .ZN(n9408) );
  AOI22_X1 U10641 ( .A1(n4483), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9406), .B2(
        n10275), .ZN(n9407) );
  OAI211_X1 U10642 ( .C1(n9409), .C2(n9484), .A(n9408), .B(n9407), .ZN(n9410)
         );
  AOI21_X1 U10643 ( .B1(n9561), .B2(n9508), .A(n9410), .ZN(n9411) );
  OAI21_X1 U10644 ( .B1(n9565), .B2(n9481), .A(n9411), .ZN(P1_U3270) );
  XOR2_X1 U10645 ( .A(n9412), .B(n9419), .Z(n9570) );
  INV_X1 U10646 ( .A(n9428), .ZN(n9414) );
  AOI21_X1 U10647 ( .B1(n9566), .B2(n9414), .A(n9413), .ZN(n9567) );
  INV_X1 U10648 ( .A(n9415), .ZN(n9416) );
  AOI22_X1 U10649 ( .A1(n4483), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9416), .B2(
        n10275), .ZN(n9417) );
  OAI21_X1 U10650 ( .B1(n9418), .B2(n9484), .A(n9417), .ZN(n9425) );
  XNOR2_X1 U10651 ( .A(n9420), .B(n9419), .ZN(n9423) );
  AOI222_X1 U10652 ( .A1(n10266), .A2(n9423), .B1(n9422), .B2(n10264), .C1(
        n9421), .C2(n10263), .ZN(n9569) );
  NOR2_X1 U10653 ( .A1(n9569), .A2(n4483), .ZN(n9424) );
  AOI211_X1 U10654 ( .C1(n9567), .C2(n10282), .A(n9425), .B(n9424), .ZN(n9426)
         );
  OAI21_X1 U10655 ( .B1(n9570), .B2(n9481), .A(n9426), .ZN(P1_U3271) );
  XNOR2_X1 U10656 ( .A(n9427), .B(n9435), .ZN(n9575) );
  AOI211_X1 U10657 ( .C1(n9573), .C2(n9443), .A(n10325), .B(n9428), .ZN(n9572)
         );
  NOR2_X1 U10658 ( .A1(n9429), .A2(n9484), .ZN(n9433) );
  OAI22_X1 U10659 ( .A1(n9508), .A2(n9431), .B1(n9430), .B2(n9505), .ZN(n9432)
         );
  AOI211_X1 U10660 ( .C1(n9572), .C2(n9490), .A(n9433), .B(n9432), .ZN(n9440)
         );
  XOR2_X1 U10661 ( .A(n9435), .B(n9434), .Z(n9436) );
  OAI222_X1 U10662 ( .A1(n10128), .A2(n9438), .B1(n10129), .B2(n9437), .C1(
        n9436), .C2(n9477), .ZN(n9571) );
  NAND2_X1 U10663 ( .A1(n9571), .A2(n9508), .ZN(n9439) );
  OAI211_X1 U10664 ( .C1(n9575), .C2(n9481), .A(n9440), .B(n9439), .ZN(
        P1_U3272) );
  XNOR2_X1 U10665 ( .A(n9442), .B(n9441), .ZN(n9580) );
  INV_X1 U10666 ( .A(n9443), .ZN(n9444) );
  AOI211_X1 U10667 ( .C1(n9578), .C2(n9458), .A(n10325), .B(n9444), .ZN(n9577)
         );
  INV_X1 U10668 ( .A(n9578), .ZN(n9445) );
  NOR2_X1 U10669 ( .A1(n9445), .A2(n9484), .ZN(n9449) );
  OAI22_X1 U10670 ( .A1(n9508), .A2(n9447), .B1(n9446), .B2(n9505), .ZN(n9448)
         );
  AOI211_X1 U10671 ( .C1(n9577), .C2(n9490), .A(n9449), .B(n9448), .ZN(n9456)
         );
  NAND2_X1 U10672 ( .A1(n9451), .A2(n9450), .ZN(n9452) );
  XNOR2_X1 U10673 ( .A(n9452), .B(n4879), .ZN(n9453) );
  OAI222_X1 U10674 ( .A1(n10128), .A2(n9454), .B1(n10129), .B2(n9478), .C1(
        n9477), .C2(n9453), .ZN(n9576) );
  NAND2_X1 U10675 ( .A1(n9576), .A2(n9508), .ZN(n9455) );
  OAI211_X1 U10676 ( .C1(n9580), .C2(n9481), .A(n9456), .B(n9455), .ZN(
        P1_U3273) );
  XNOR2_X1 U10677 ( .A(n9457), .B(n9465), .ZN(n9585) );
  INV_X1 U10678 ( .A(n9482), .ZN(n9460) );
  INV_X1 U10679 ( .A(n9458), .ZN(n9459) );
  AOI21_X1 U10680 ( .B1(n9581), .B2(n9460), .A(n9459), .ZN(n9582) );
  INV_X1 U10681 ( .A(n9461), .ZN(n9462) );
  AOI22_X1 U10682 ( .A1(n4483), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9462), .B2(
        n10275), .ZN(n9463) );
  OAI21_X1 U10683 ( .B1(n9464), .B2(n9484), .A(n9463), .ZN(n9471) );
  XNOR2_X1 U10684 ( .A(n9466), .B(n9465), .ZN(n9469) );
  AOI222_X1 U10685 ( .A1(n10266), .A2(n9469), .B1(n9468), .B2(n10264), .C1(
        n9467), .C2(n10263), .ZN(n9584) );
  NOR2_X1 U10686 ( .A1(n9584), .A2(n4483), .ZN(n9470) );
  AOI211_X1 U10687 ( .C1(n9582), .C2(n10282), .A(n9471), .B(n9470), .ZN(n9472)
         );
  OAI21_X1 U10688 ( .B1(n9585), .B2(n9481), .A(n9472), .ZN(P1_U3274) );
  NAND2_X1 U10689 ( .A1(n9474), .A2(n9473), .ZN(n9475) );
  XNOR2_X1 U10690 ( .A(n9475), .B(n9479), .ZN(n9476) );
  OAI222_X1 U10691 ( .A1(n10128), .A2(n9478), .B1(n10129), .B2(n10093), .C1(
        n9477), .C2(n9476), .ZN(n9588) );
  INV_X1 U10692 ( .A(n9588), .ZN(n9493) );
  AND2_X1 U10693 ( .A1(n9480), .A2(n9479), .ZN(n9586) );
  OR3_X1 U10694 ( .A1(n9587), .A2(n9586), .A3(n9481), .ZN(n9492) );
  AOI211_X1 U10695 ( .C1(n9483), .C2(n9504), .A(n10325), .B(n9482), .ZN(n9589)
         );
  NOR2_X1 U10696 ( .A1(n9485), .A2(n9484), .ZN(n9489) );
  OAI22_X1 U10697 ( .A1(n9508), .A2(n9487), .B1(n9486), .B2(n9505), .ZN(n9488)
         );
  AOI211_X1 U10698 ( .C1(n9589), .C2(n9490), .A(n9489), .B(n9488), .ZN(n9491)
         );
  OAI211_X1 U10699 ( .C1(n4483), .C2(n9493), .A(n9492), .B(n9491), .ZN(
        P1_U3275) );
  XNOR2_X1 U10700 ( .A(n9495), .B(n9494), .ZN(n9501) );
  OAI22_X1 U10701 ( .A1(n10109), .A2(n10129), .B1(n10128), .B2(n9496), .ZN(
        n9500) );
  XNOR2_X1 U10702 ( .A(n9498), .B(n9497), .ZN(n9597) );
  NOR2_X1 U10703 ( .A1(n9597), .A2(n10272), .ZN(n9499) );
  AOI211_X1 U10704 ( .C1(n10266), .C2(n9501), .A(n9500), .B(n9499), .ZN(n9596)
         );
  INV_X1 U10705 ( .A(n9597), .ZN(n9514) );
  NAND2_X1 U10706 ( .A1(n9502), .A2(n9510), .ZN(n9503) );
  NAND2_X1 U10707 ( .A1(n9504), .A2(n9503), .ZN(n9593) );
  OAI22_X1 U10708 ( .A1(n9508), .A2(n9507), .B1(n9506), .B2(n9505), .ZN(n9509)
         );
  AOI21_X1 U10709 ( .B1(n9510), .B2(n10276), .A(n9509), .ZN(n9511) );
  OAI21_X1 U10710 ( .B1(n9593), .B2(n9512), .A(n9511), .ZN(n9513) );
  AOI21_X1 U10711 ( .B1(n9514), .B2(n10283), .A(n9513), .ZN(n9515) );
  OAI21_X1 U10712 ( .B1(n9596), .B2(n4483), .A(n9515), .ZN(P1_U3276) );
  AOI21_X1 U10713 ( .B1(n9516), .B2(n10164), .A(n10145), .ZN(n9517) );
  OAI21_X1 U10714 ( .B1(n9518), .B2(n10325), .A(n9517), .ZN(n9599) );
  MUX2_X1 U10715 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9599), .S(n10341), .Z(
        P1_U3554) );
  INV_X1 U10716 ( .A(n10298), .ZN(n10320) );
  NAND2_X1 U10717 ( .A1(n9519), .A2(n10320), .ZN(n9524) );
  NOR2_X1 U10718 ( .A1(n9520), .A2(n10325), .ZN(n9522) );
  MUX2_X1 U10719 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9600), .S(n10341), .Z(
        P1_U3552) );
  NOR2_X1 U10720 ( .A1(n9526), .A2(n9525), .ZN(n9527) );
  OAI211_X1 U10721 ( .C1(n9529), .C2(n10298), .A(n9528), .B(n9527), .ZN(n9601)
         );
  MUX2_X1 U10722 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9601), .S(n10341), .Z(
        P1_U3551) );
  AOI21_X1 U10723 ( .B1(n10164), .B2(n9531), .A(n9530), .ZN(n9532) );
  OAI211_X1 U10724 ( .C1(n9534), .C2(n10298), .A(n9533), .B(n9532), .ZN(n9602)
         );
  MUX2_X1 U10725 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9602), .S(n10341), .Z(
        P1_U3550) );
  AOI21_X1 U10726 ( .B1(n10164), .B2(n9536), .A(n9535), .ZN(n9537) );
  OAI211_X1 U10727 ( .C1(n9539), .C2(n10298), .A(n9538), .B(n9537), .ZN(n9603)
         );
  MUX2_X1 U10728 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9603), .S(n10341), .Z(
        P1_U3549) );
  AOI22_X1 U10729 ( .A1(n9541), .A2(n10165), .B1(n10164), .B2(n9540), .ZN(
        n9542) );
  OAI211_X1 U10730 ( .C1(n9544), .C2(n10298), .A(n9543), .B(n9542), .ZN(n9604)
         );
  MUX2_X1 U10731 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9604), .S(n10341), .Z(
        P1_U3548) );
  AOI211_X1 U10732 ( .C1(n10164), .C2(n9547), .A(n9546), .B(n9545), .ZN(n9548)
         );
  OAI21_X1 U10733 ( .B1(n9549), .B2(n10298), .A(n9548), .ZN(n9605) );
  MUX2_X1 U10734 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9605), .S(n10341), .Z(
        P1_U3547) );
  AOI22_X1 U10735 ( .A1(n9551), .A2(n10165), .B1(n10164), .B2(n9550), .ZN(
        n9552) );
  OAI211_X1 U10736 ( .C1(n9554), .C2(n10298), .A(n9553), .B(n9552), .ZN(n9606)
         );
  MUX2_X1 U10737 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9606), .S(n10341), .Z(
        P1_U3546) );
  NAND2_X1 U10738 ( .A1(n9555), .A2(n10320), .ZN(n9560) );
  INV_X1 U10739 ( .A(n9556), .ZN(n9558) );
  NAND4_X1 U10740 ( .A1(n9560), .A2(n9559), .A3(n9558), .A4(n9557), .ZN(n9607)
         );
  MUX2_X1 U10741 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9607), .S(n10341), .Z(
        P1_U3545) );
  AOI211_X1 U10742 ( .C1(n10164), .C2(n9563), .A(n9562), .B(n9561), .ZN(n9564)
         );
  OAI21_X1 U10743 ( .B1(n9565), .B2(n10298), .A(n9564), .ZN(n9608) );
  MUX2_X1 U10744 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9608), .S(n10341), .Z(
        P1_U3544) );
  AOI22_X1 U10745 ( .A1(n9567), .A2(n10165), .B1(n10164), .B2(n9566), .ZN(
        n9568) );
  OAI211_X1 U10746 ( .C1(n9570), .C2(n10298), .A(n9569), .B(n9568), .ZN(n9609)
         );
  MUX2_X1 U10747 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9609), .S(n10341), .Z(
        P1_U3543) );
  AOI211_X1 U10748 ( .C1(n10164), .C2(n9573), .A(n9572), .B(n9571), .ZN(n9574)
         );
  OAI21_X1 U10749 ( .B1(n9575), .B2(n10298), .A(n9574), .ZN(n9610) );
  MUX2_X1 U10750 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9610), .S(n10341), .Z(
        P1_U3542) );
  AOI211_X1 U10751 ( .C1(n10164), .C2(n9578), .A(n9577), .B(n9576), .ZN(n9579)
         );
  OAI21_X1 U10752 ( .B1(n9580), .B2(n10298), .A(n9579), .ZN(n9611) );
  MUX2_X1 U10753 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9611), .S(n10341), .Z(
        P1_U3541) );
  AOI22_X1 U10754 ( .A1(n9582), .A2(n10165), .B1(n10164), .B2(n9581), .ZN(
        n9583) );
  OAI211_X1 U10755 ( .C1(n9585), .C2(n10298), .A(n9584), .B(n9583), .ZN(n9612)
         );
  MUX2_X1 U10756 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9612), .S(n10341), .Z(
        P1_U3540) );
  NOR3_X1 U10757 ( .A1(n9587), .A2(n9586), .A3(n10298), .ZN(n9591) );
  MUX2_X1 U10758 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9613), .S(n10341), .Z(
        P1_U3539) );
  OAI22_X1 U10759 ( .A1(n9593), .A2(n10325), .B1(n9592), .B2(n10323), .ZN(
        n9594) );
  INV_X1 U10760 ( .A(n9594), .ZN(n9595) );
  OAI211_X1 U10761 ( .C1(n9597), .C2(n10170), .A(n9596), .B(n9595), .ZN(n9614)
         );
  MUX2_X1 U10762 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9614), .S(n10341), .Z(
        P1_U3538) );
  MUX2_X1 U10763 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9598), .S(n10341), .Z(
        P1_U3523) );
  MUX2_X1 U10764 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9599), .S(n10333), .Z(
        P1_U3522) );
  MUX2_X1 U10765 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9600), .S(n10333), .Z(
        P1_U3520) );
  MUX2_X1 U10766 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9601), .S(n10333), .Z(
        P1_U3519) );
  MUX2_X1 U10767 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9602), .S(n10333), .Z(
        P1_U3518) );
  MUX2_X1 U10768 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9603), .S(n10333), .Z(
        P1_U3517) );
  MUX2_X1 U10769 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9604), .S(n10333), .Z(
        P1_U3516) );
  MUX2_X1 U10770 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9605), .S(n10333), .Z(
        P1_U3515) );
  MUX2_X1 U10771 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9606), .S(n10333), .Z(
        P1_U3514) );
  MUX2_X1 U10772 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9607), .S(n10333), .Z(
        P1_U3513) );
  MUX2_X1 U10773 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9608), .S(n10333), .Z(
        P1_U3512) );
  MUX2_X1 U10774 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9609), .S(n10333), .Z(
        P1_U3511) );
  MUX2_X1 U10775 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9610), .S(n10333), .Z(
        P1_U3510) );
  MUX2_X1 U10776 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9611), .S(n10333), .Z(
        P1_U3508) );
  MUX2_X1 U10777 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9612), .S(n10333), .Z(
        P1_U3505) );
  MUX2_X1 U10778 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9613), .S(n10333), .Z(
        P1_U3502) );
  MUX2_X1 U10779 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9614), .S(n10333), .Z(
        P1_U3499) );
  NOR4_X1 U10780 ( .A1(n9615), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5755), .A4(
        P1_U3084), .ZN(n9616) );
  AOI21_X1 U10781 ( .B1(n9617), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9616), .ZN(
        n9618) );
  OAI21_X1 U10782 ( .B1(n9619), .B2(n9624), .A(n9618), .ZN(P1_U3322) );
  INV_X1 U10783 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9621) );
  OAI222_X1 U10784 ( .A1(n9622), .A2(n9621), .B1(n9624), .B2(n9620), .C1(n5739), .C2(P1_U3084), .ZN(P1_U3323) );
  INV_X1 U10785 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9926) );
  OAI222_X1 U10786 ( .A1(n9626), .A2(n9926), .B1(P1_U3084), .B2(n9625), .C1(
        n9624), .C2(n9623), .ZN(P1_U3324) );
  MUX2_X1 U10787 ( .A(n9627), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10788 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10492) );
  NOR2_X1 U10789 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9628) );
  AOI21_X1 U10790 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9628), .ZN(n10459) );
  NOR2_X1 U10791 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9629) );
  AOI21_X1 U10792 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9629), .ZN(n10462) );
  NOR2_X1 U10793 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9630) );
  AOI21_X1 U10794 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9630), .ZN(n10465) );
  NOR2_X1 U10795 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9631) );
  AOI21_X1 U10796 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9631), .ZN(n10468) );
  NOR2_X1 U10797 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9632) );
  AOI21_X1 U10798 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9632), .ZN(n10471) );
  NOR2_X1 U10799 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9638) );
  XNOR2_X1 U10800 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10499) );
  NAND2_X1 U10801 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9636) );
  XOR2_X1 U10802 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10497) );
  NAND2_X1 U10803 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9634) );
  XOR2_X1 U10804 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10486) );
  AOI21_X1 U10805 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10453) );
  INV_X1 U10806 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10025) );
  NAND3_X1 U10807 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10455) );
  OAI21_X1 U10808 ( .B1(n10453), .B2(n10025), .A(n10455), .ZN(n10485) );
  NAND2_X1 U10809 ( .A1(n10486), .A2(n10485), .ZN(n9633) );
  NAND2_X1 U10810 ( .A1(n9634), .A2(n9633), .ZN(n10496) );
  NAND2_X1 U10811 ( .A1(n10497), .A2(n10496), .ZN(n9635) );
  NAND2_X1 U10812 ( .A1(n9636), .A2(n9635), .ZN(n10498) );
  NOR2_X1 U10813 ( .A1(n10499), .A2(n10498), .ZN(n9637) );
  NOR2_X1 U10814 ( .A1(n9638), .A2(n9637), .ZN(n9639) );
  NOR2_X1 U10815 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9639), .ZN(n10488) );
  AND2_X1 U10816 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9639), .ZN(n10487) );
  NOR2_X1 U10817 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10487), .ZN(n9640) );
  NOR2_X1 U10818 ( .A1(n10488), .A2(n9640), .ZN(n9641) );
  NAND2_X1 U10819 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n9641), .ZN(n9643) );
  XOR2_X1 U10820 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n9641), .Z(n10495) );
  NAND2_X1 U10821 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10495), .ZN(n9642) );
  NAND2_X1 U10822 ( .A1(n9643), .A2(n9642), .ZN(n9644) );
  NAND2_X1 U10823 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9644), .ZN(n9646) );
  XOR2_X1 U10824 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9644), .Z(n10484) );
  NAND2_X1 U10825 ( .A1(n10484), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9645) );
  NAND2_X1 U10826 ( .A1(n9646), .A2(n9645), .ZN(n9647) );
  NAND2_X1 U10827 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9647), .ZN(n9649) );
  XOR2_X1 U10828 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9647), .Z(n10494) );
  NAND2_X1 U10829 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10494), .ZN(n9648) );
  NAND2_X1 U10830 ( .A1(n9649), .A2(n9648), .ZN(n9650) );
  AND2_X1 U10831 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9650), .ZN(n9651) );
  XNOR2_X1 U10832 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9650), .ZN(n10483) );
  NAND2_X1 U10833 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9652) );
  OAI21_X1 U10834 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9652), .ZN(n10479) );
  NAND2_X1 U10835 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9653) );
  OAI21_X1 U10836 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9653), .ZN(n10476) );
  AOI21_X1 U10837 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10475), .ZN(n10474) );
  NOR2_X1 U10838 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9654) );
  AOI21_X1 U10839 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9654), .ZN(n10473) );
  NAND2_X1 U10840 ( .A1(n10474), .A2(n10473), .ZN(n10472) );
  OAI21_X1 U10841 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10472), .ZN(n10470) );
  NAND2_X1 U10842 ( .A1(n10471), .A2(n10470), .ZN(n10469) );
  OAI21_X1 U10843 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10469), .ZN(n10467) );
  NAND2_X1 U10844 ( .A1(n10468), .A2(n10467), .ZN(n10466) );
  OAI21_X1 U10845 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10466), .ZN(n10464) );
  NAND2_X1 U10846 ( .A1(n10465), .A2(n10464), .ZN(n10463) );
  OAI21_X1 U10847 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10463), .ZN(n10461) );
  NAND2_X1 U10848 ( .A1(n10462), .A2(n10461), .ZN(n10460) );
  OAI21_X1 U10849 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10460), .ZN(n10458) );
  NAND2_X1 U10850 ( .A1(n10459), .A2(n10458), .ZN(n10457) );
  OAI21_X1 U10851 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10457), .ZN(n10491) );
  NOR2_X1 U10852 ( .A1(n10492), .A2(n10491), .ZN(n9655) );
  NAND2_X1 U10853 ( .A1(n10492), .A2(n10491), .ZN(n10490) );
  OAI21_X1 U10854 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n9655), .A(n10490), .ZN(
        n10013) );
  INV_X1 U10855 ( .A(SI_0_), .ZN(n10011) );
  XNOR2_X1 U10856 ( .A(keyinput_g54), .B(n10359), .ZN(n9662) );
  AOI22_X1 U10857 ( .A1(SI_29_), .A2(keyinput_g3), .B1(SI_15_), .B2(
        keyinput_g17), .ZN(n9656) );
  OAI221_X1 U10858 ( .B1(SI_29_), .B2(keyinput_g3), .C1(SI_15_), .C2(
        keyinput_g17), .A(n9656), .ZN(n9661) );
  AOI22_X1 U10859 ( .A1(SI_9_), .A2(keyinput_g23), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_g71), .ZN(n9657) );
  OAI221_X1 U10860 ( .B1(SI_9_), .B2(keyinput_g23), .C1(
        P2_DATAO_REG_25__SCAN_IN), .C2(keyinput_g71), .A(n9657), .ZN(n9660) );
  AOI22_X1 U10861 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_g42), .B1(
        SI_14_), .B2(keyinput_g18), .ZN(n9658) );
  OAI221_X1 U10862 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .C1(
        SI_14_), .C2(keyinput_g18), .A(n9658), .ZN(n9659) );
  NOR4_X1 U10863 ( .A1(n9662), .A2(n9661), .A3(n9660), .A4(n9659), .ZN(n9690)
         );
  AOI22_X1 U10864 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .ZN(n9663) );
  OAI221_X1 U10865 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_g50), .A(n9663), .ZN(n9670) );
  AOI22_X1 U10866 ( .A1(SI_12_), .A2(keyinput_g20), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_g77), .ZN(n9664) );
  OAI221_X1 U10867 ( .B1(SI_12_), .B2(keyinput_g20), .C1(
        P2_DATAO_REG_19__SCAN_IN), .C2(keyinput_g77), .A(n9664), .ZN(n9669) );
  AOI22_X1 U10868 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(keyinput_g81), .B1(
        P1_D_REG_2__SCAN_IN), .B2(keyinput_g125), .ZN(n9665) );
  OAI221_X1 U10869 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_g81), .C1(
        P1_D_REG_2__SCAN_IN), .C2(keyinput_g125), .A(n9665), .ZN(n9668) );
  AOI22_X1 U10870 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_g93), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput_g101), .ZN(n9666) );
  OAI221_X1 U10871 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_g93), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput_g101), .A(n9666), .ZN(n9667) );
  NOR4_X1 U10872 ( .A1(n9670), .A2(n9669), .A3(n9668), .A4(n9667), .ZN(n9689)
         );
  AOI22_X1 U10873 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_g52), .B1(
        P2_REG3_REG_8__SCAN_IN), .B2(keyinput_g43), .ZN(n9671) );
  OAI221_X1 U10874 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_g52), .C1(
        P2_REG3_REG_8__SCAN_IN), .C2(keyinput_g43), .A(n9671), .ZN(n9678) );
  AOI22_X1 U10875 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput_g98), .ZN(n9672) );
  OAI221_X1 U10876 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput_g98), .A(n9672), .ZN(n9677) );
  AOI22_X1 U10877 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(keyinput_g68), .B1(
        SI_17_), .B2(keyinput_g15), .ZN(n9673) );
  OAI221_X1 U10878 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_g68), .C1(
        SI_17_), .C2(keyinput_g15), .A(n9673), .ZN(n9676) );
  AOI22_X1 U10879 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_g87), .B1(
        SI_27_), .B2(keyinput_g5), .ZN(n9674) );
  OAI221_X1 U10880 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_g87), .C1(
        SI_27_), .C2(keyinput_g5), .A(n9674), .ZN(n9675) );
  NOR4_X1 U10881 ( .A1(n9678), .A2(n9677), .A3(n9676), .A4(n9675), .ZN(n9688)
         );
  AOI22_X1 U10882 ( .A1(SI_3_), .A2(keyinput_g29), .B1(SI_10_), .B2(
        keyinput_g22), .ZN(n9679) );
  OAI221_X1 U10883 ( .B1(SI_3_), .B2(keyinput_g29), .C1(SI_10_), .C2(
        keyinput_g22), .A(n9679), .ZN(n9686) );
  AOI22_X1 U10884 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_g39), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_g78), .ZN(n9680) );
  OAI221_X1 U10885 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .C1(
        P2_DATAO_REG_18__SCAN_IN), .C2(keyinput_g78), .A(n9680), .ZN(n9685) );
  AOI22_X1 U10886 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n9681) );
  OAI221_X1 U10887 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n9681), .ZN(n9684) );
  AOI22_X1 U10888 ( .A1(P2_B_REG_SCAN_IN), .A2(keyinput_g64), .B1(
        P1_IR_REG_21__SCAN_IN), .B2(keyinput_g112), .ZN(n9682) );
  OAI221_X1 U10889 ( .B1(P2_B_REG_SCAN_IN), .B2(keyinput_g64), .C1(
        P1_IR_REG_21__SCAN_IN), .C2(keyinput_g112), .A(n9682), .ZN(n9683) );
  NOR4_X1 U10890 ( .A1(n9686), .A2(n9685), .A3(n9684), .A4(n9683), .ZN(n9687)
         );
  NAND4_X1 U10891 ( .A1(n9690), .A2(n9689), .A3(n9688), .A4(n9687), .ZN(n9831)
         );
  AOI22_X1 U10892 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(SI_4_), 
        .B2(keyinput_g28), .ZN(n9691) );
  OAI221_X1 U10893 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(SI_4_), .C2(keyinput_g28), .A(n9691), .ZN(n9698) );
  AOI22_X1 U10894 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_g84), .ZN(n9692) );
  OAI221_X1 U10895 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(
        P2_DATAO_REG_12__SCAN_IN), .C2(keyinput_g84), .A(n9692), .ZN(n9697) );
  AOI22_X1 U10896 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(keyinput_g82), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput_g110), .ZN(n9693) );
  OAI221_X1 U10897 ( .B1(P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_g82), .C1(
        P1_IR_REG_19__SCAN_IN), .C2(keyinput_g110), .A(n9693), .ZN(n9696) );
  AOI22_X1 U10898 ( .A1(SI_13_), .A2(keyinput_g19), .B1(P1_IR_REG_13__SCAN_IN), 
        .B2(keyinput_g104), .ZN(n9694) );
  OAI221_X1 U10899 ( .B1(SI_13_), .B2(keyinput_g19), .C1(P1_IR_REG_13__SCAN_IN), .C2(keyinput_g104), .A(n9694), .ZN(n9695) );
  NOR4_X1 U10900 ( .A1(n9698), .A2(n9697), .A3(n9696), .A4(n9695), .ZN(n9728)
         );
  AOI22_X1 U10901 ( .A1(SI_16_), .A2(keyinput_g16), .B1(P1_D_REG_0__SCAN_IN), 
        .B2(keyinput_g123), .ZN(n9699) );
  OAI221_X1 U10902 ( .B1(SI_16_), .B2(keyinput_g16), .C1(P1_D_REG_0__SCAN_IN), 
        .C2(keyinput_g123), .A(n9699), .ZN(n9706) );
  AOI22_X1 U10903 ( .A1(SI_1_), .A2(keyinput_g31), .B1(P1_IR_REG_6__SCAN_IN), 
        .B2(keyinput_g97), .ZN(n9700) );
  OAI221_X1 U10904 ( .B1(SI_1_), .B2(keyinput_g31), .C1(P1_IR_REG_6__SCAN_IN), 
        .C2(keyinput_g97), .A(n9700), .ZN(n9705) );
  AOI22_X1 U10905 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput_g79), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_g76), .ZN(n9701) );
  OAI221_X1 U10906 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .C1(
        P2_DATAO_REG_20__SCAN_IN), .C2(keyinput_g76), .A(n9701), .ZN(n9704) );
  AOI22_X1 U10907 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_g36), .B1(SI_8_), .B2(keyinput_g24), .ZN(n9702) );
  OAI221_X1 U10908 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .C1(
        SI_8_), .C2(keyinput_g24), .A(n9702), .ZN(n9703) );
  NOR4_X1 U10909 ( .A1(n9706), .A2(n9705), .A3(n9704), .A4(n9703), .ZN(n9727)
         );
  AOI22_X1 U10910 ( .A1(SI_6_), .A2(keyinput_g26), .B1(P1_D_REG_3__SCAN_IN), 
        .B2(keyinput_g126), .ZN(n9707) );
  OAI221_X1 U10911 ( .B1(SI_6_), .B2(keyinput_g26), .C1(P1_D_REG_3__SCAN_IN), 
        .C2(keyinput_g126), .A(n9707), .ZN(n9714) );
  AOI22_X1 U10912 ( .A1(SI_18_), .A2(keyinput_g14), .B1(P1_IR_REG_31__SCAN_IN), 
        .B2(keyinput_g122), .ZN(n9708) );
  OAI221_X1 U10913 ( .B1(SI_18_), .B2(keyinput_g14), .C1(P1_IR_REG_31__SCAN_IN), .C2(keyinput_g122), .A(n9708), .ZN(n9713) );
  AOI22_X1 U10914 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_g124), .B1(
        P1_IR_REG_22__SCAN_IN), .B2(keyinput_g113), .ZN(n9709) );
  OAI221_X1 U10915 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_g124), .C1(
        P1_IR_REG_22__SCAN_IN), .C2(keyinput_g113), .A(n9709), .ZN(n9712) );
  AOI22_X1 U10916 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(keyinput_g72), .B1(
        P1_IR_REG_26__SCAN_IN), .B2(keyinput_g117), .ZN(n9710) );
  OAI221_X1 U10917 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_g72), .C1(
        P1_IR_REG_26__SCAN_IN), .C2(keyinput_g117), .A(n9710), .ZN(n9711) );
  NOR4_X1 U10918 ( .A1(n9714), .A2(n9713), .A3(n9712), .A4(n9711), .ZN(n9726)
         );
  AOI22_X1 U10919 ( .A1(n5488), .A2(keyinput_g75), .B1(n5519), .B2(
        keyinput_g73), .ZN(n9715) );
  OAI221_X1 U10920 ( .B1(n5488), .B2(keyinput_g75), .C1(n5519), .C2(
        keyinput_g73), .A(n9715), .ZN(n9724) );
  AOI22_X1 U10921 ( .A1(SI_28_), .A2(keyinput_g4), .B1(n5750), .B2(
        keyinput_g109), .ZN(n9716) );
  OAI221_X1 U10922 ( .B1(SI_28_), .B2(keyinput_g4), .C1(n5750), .C2(
        keyinput_g109), .A(n9716), .ZN(n9723) );
  AOI22_X1 U10923 ( .A1(n9718), .A2(keyinput_g12), .B1(keyinput_g49), .B2(
        n9924), .ZN(n9717) );
  OAI221_X1 U10924 ( .B1(n9718), .B2(keyinput_g12), .C1(n9924), .C2(
        keyinput_g49), .A(n9717), .ZN(n9722) );
  XNOR2_X1 U10925 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_g34), .ZN(n9720) );
  XNOR2_X1 U10926 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_g33), .ZN(n9719) );
  NAND2_X1 U10927 ( .A1(n9720), .A2(n9719), .ZN(n9721) );
  NOR4_X1 U10928 ( .A1(n9724), .A2(n9723), .A3(n9722), .A4(n9721), .ZN(n9725)
         );
  NAND4_X1 U10929 ( .A1(n9728), .A2(n9727), .A3(n9726), .A4(n9725), .ZN(n9830)
         );
  INV_X1 U10930 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9952) );
  AOI22_X1 U10931 ( .A1(n9926), .A2(keyinput_g67), .B1(n9952), .B2(
        keyinput_g100), .ZN(n9729) );
  OAI221_X1 U10932 ( .B1(n9926), .B2(keyinput_g67), .C1(n9952), .C2(
        keyinput_g100), .A(n9729), .ZN(n9738) );
  AOI22_X1 U10933 ( .A1(n9929), .A2(keyinput_g74), .B1(n9731), .B2(keyinput_g6), .ZN(n9730) );
  OAI221_X1 U10934 ( .B1(n9929), .B2(keyinput_g74), .C1(n9731), .C2(
        keyinput_g6), .A(n9730), .ZN(n9737) );
  XOR2_X1 U10935 ( .A(n5275), .B(keyinput_g35), .Z(n9735) );
  XNOR2_X1 U10936 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_g120), .ZN(n9734)
         );
  XNOR2_X1 U10937 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_g88), .ZN(n9733)
         );
  XNOR2_X1 U10938 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_g115), .ZN(n9732)
         );
  NAND4_X1 U10939 ( .A1(n9735), .A2(n9734), .A3(n9733), .A4(n9732), .ZN(n9736)
         );
  NOR3_X1 U10940 ( .A1(n9738), .A2(n9737), .A3(n9736), .ZN(n9775) );
  INV_X1 U10941 ( .A(SI_7_), .ZN(n9927) );
  AOI22_X1 U10942 ( .A1(n9740), .A2(keyinput_g65), .B1(n9927), .B2(
        keyinput_g25), .ZN(n9739) );
  OAI221_X1 U10943 ( .B1(n9740), .B2(keyinput_g65), .C1(n9927), .C2(
        keyinput_g25), .A(n9739), .ZN(n9750) );
  AOI22_X1 U10944 ( .A1(n9742), .A2(keyinput_g13), .B1(n5729), .B2(
        keyinput_g96), .ZN(n9741) );
  OAI221_X1 U10945 ( .B1(n9742), .B2(keyinput_g13), .C1(n5729), .C2(
        keyinput_g96), .A(n9741), .ZN(n9749) );
  AOI22_X1 U10946 ( .A1(n4866), .A2(keyinput_g119), .B1(keyinput_g55), .B2(
        n9744), .ZN(n9743) );
  OAI221_X1 U10947 ( .B1(n4866), .B2(keyinput_g119), .C1(n9744), .C2(
        keyinput_g55), .A(n9743), .ZN(n9748) );
  XNOR2_X1 U10948 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_g105), .ZN(n9746)
         );
  XNOR2_X1 U10949 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_g66), .ZN(n9745)
         );
  NAND2_X1 U10950 ( .A1(n9746), .A2(n9745), .ZN(n9747) );
  NOR4_X1 U10951 ( .A1(n9750), .A2(n9749), .A3(n9748), .A4(n9747), .ZN(n9774)
         );
  AOI22_X1 U10952 ( .A1(n9752), .A2(keyinput_g51), .B1(n5735), .B2(
        keyinput_g121), .ZN(n9751) );
  OAI221_X1 U10953 ( .B1(n9752), .B2(keyinput_g51), .C1(n5735), .C2(
        keyinput_g121), .A(n9751), .ZN(n9761) );
  AOI22_X1 U10954 ( .A1(n4625), .A2(keyinput_g92), .B1(keyinput_g45), .B2(
        n9955), .ZN(n9753) );
  OAI221_X1 U10955 ( .B1(n4625), .B2(keyinput_g92), .C1(n9955), .C2(
        keyinput_g45), .A(n9753), .ZN(n9760) );
  AOI22_X1 U10956 ( .A1(n5558), .A2(keyinput_g47), .B1(keyinput_g37), .B2(
        n9755), .ZN(n9754) );
  OAI221_X1 U10957 ( .B1(n5558), .B2(keyinput_g47), .C1(n9755), .C2(
        keyinput_g37), .A(n9754), .ZN(n9759) );
  XOR2_X1 U10958 ( .A(n5185), .B(keyinput_g41), .Z(n9757) );
  XNOR2_X1 U10959 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_g118), .ZN(n9756)
         );
  NAND2_X1 U10960 ( .A1(n9757), .A2(n9756), .ZN(n9758) );
  NOR4_X1 U10961 ( .A1(n9761), .A2(n9760), .A3(n9759), .A4(n9758), .ZN(n9773)
         );
  INV_X1 U10962 ( .A(SI_11_), .ZN(n9975) );
  AOI22_X1 U10963 ( .A1(n9975), .A2(keyinput_g21), .B1(keyinput_g58), .B2(
        n5342), .ZN(n9762) );
  OAI221_X1 U10964 ( .B1(n9975), .B2(keyinput_g21), .C1(n5342), .C2(
        keyinput_g58), .A(n9762), .ZN(n9771) );
  AOI22_X1 U10965 ( .A1(n5531), .A2(keyinput_g38), .B1(n4886), .B2(
        keyinput_g103), .ZN(n9763) );
  OAI221_X1 U10966 ( .B1(n5531), .B2(keyinput_g38), .C1(n4886), .C2(
        keyinput_g103), .A(n9763), .ZN(n9770) );
  AOI22_X1 U10967 ( .A1(n9991), .A2(keyinput_g10), .B1(n9765), .B2(keyinput_g7), .ZN(n9764) );
  OAI221_X1 U10968 ( .B1(n9991), .B2(keyinput_g10), .C1(n9765), .C2(
        keyinput_g7), .A(n9764), .ZN(n9769) );
  XOR2_X1 U10969 ( .A(n5309), .B(keyinput_g53), .Z(n9767) );
  XNOR2_X1 U10970 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_g95), .ZN(n9766) );
  NAND2_X1 U10971 ( .A1(n9767), .A2(n9766), .ZN(n9768) );
  NOR4_X1 U10972 ( .A1(n9771), .A2(n9770), .A3(n9769), .A4(n9768), .ZN(n9772)
         );
  NAND4_X1 U10973 ( .A1(n9775), .A2(n9774), .A3(n9773), .A4(n9772), .ZN(n9829)
         );
  AOI22_X1 U10974 ( .A1(n6128), .A2(keyinput_g108), .B1(keyinput_g69), .B2(
        n9777), .ZN(n9776) );
  OAI221_X1 U10975 ( .B1(n6128), .B2(keyinput_g108), .C1(n9777), .C2(
        keyinput_g69), .A(n9776), .ZN(n9787) );
  AOI22_X1 U10976 ( .A1(n7282), .A2(keyinput_g56), .B1(n9779), .B2(
        keyinput_g62), .ZN(n9778) );
  OAI221_X1 U10977 ( .B1(n7282), .B2(keyinput_g56), .C1(n9779), .C2(
        keyinput_g62), .A(n9778), .ZN(n9786) );
  AOI22_X1 U10978 ( .A1(n9978), .A2(keyinput_g70), .B1(keyinput_g60), .B2(
        n9781), .ZN(n9780) );
  OAI221_X1 U10979 ( .B1(n9978), .B2(keyinput_g70), .C1(n9781), .C2(
        keyinput_g60), .A(n9780), .ZN(n9785) );
  XNOR2_X1 U10980 ( .A(SI_2_), .B(keyinput_g30), .ZN(n9783) );
  XNOR2_X1 U10981 ( .A(SI_31_), .B(keyinput_g1), .ZN(n9782) );
  NAND2_X1 U10982 ( .A1(n9783), .A2(n9782), .ZN(n9784) );
  NOR4_X1 U10983 ( .A1(n9787), .A2(n9786), .A3(n9785), .A4(n9784), .ZN(n9827)
         );
  AOI22_X1 U10984 ( .A1(n9789), .A2(keyinput_g46), .B1(n5728), .B2(
        keyinput_g94), .ZN(n9788) );
  OAI221_X1 U10985 ( .B1(n9789), .B2(keyinput_g46), .C1(n5728), .C2(
        keyinput_g94), .A(n9788), .ZN(n9799) );
  INV_X1 U10986 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9791) );
  AOI22_X1 U10987 ( .A1(n9792), .A2(keyinput_g83), .B1(n9791), .B2(
        keyinput_g127), .ZN(n9790) );
  OAI221_X1 U10988 ( .B1(n9792), .B2(keyinput_g83), .C1(n9791), .C2(
        keyinput_g127), .A(n9790), .ZN(n9798) );
  INV_X1 U10989 ( .A(SI_24_), .ZN(n9923) );
  XOR2_X1 U10990 ( .A(n9923), .B(keyinput_g8), .Z(n9796) );
  XNOR2_X1 U10991 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_g48), .ZN(n9795)
         );
  XNOR2_X1 U10992 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_g99), .ZN(n9794) );
  XNOR2_X1 U10993 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_g114), .ZN(n9793)
         );
  NAND4_X1 U10994 ( .A1(n9796), .A2(n9795), .A3(n9794), .A4(n9793), .ZN(n9797)
         );
  NOR3_X1 U10995 ( .A1(n9799), .A2(n9798), .A3(n9797), .ZN(n9826) );
  AOI22_X1 U10996 ( .A1(n9802), .A2(keyinput_g90), .B1(keyinput_g40), .B2(
        n9801), .ZN(n9800) );
  OAI221_X1 U10997 ( .B1(n9802), .B2(keyinput_g90), .C1(n9801), .C2(
        keyinput_g40), .A(n9800), .ZN(n9812) );
  AOI22_X1 U10998 ( .A1(n9805), .A2(keyinput_g85), .B1(n9804), .B2(
        keyinput_g80), .ZN(n9803) );
  OAI221_X1 U10999 ( .B1(n9805), .B2(keyinput_g85), .C1(n9804), .C2(
        keyinput_g80), .A(n9803), .ZN(n9811) );
  XNOR2_X1 U11000 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_g89), .ZN(n9809)
         );
  XNOR2_X1 U11001 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_g106), .ZN(n9808)
         );
  XNOR2_X1 U11002 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_g102), .ZN(n9807)
         );
  XNOR2_X1 U11003 ( .A(SI_5_), .B(keyinput_g27), .ZN(n9806) );
  NAND4_X1 U11004 ( .A1(n9809), .A2(n9808), .A3(n9807), .A4(n9806), .ZN(n9810)
         );
  NOR3_X1 U11005 ( .A1(n9812), .A2(n9811), .A3(n9810), .ZN(n9825) );
  INV_X1 U11006 ( .A(SI_21_), .ZN(n9953) );
  AOI22_X1 U11007 ( .A1(n9953), .A2(keyinput_g11), .B1(n5749), .B2(
        keyinput_g111), .ZN(n9813) );
  OAI221_X1 U11008 ( .B1(n9953), .B2(keyinput_g11), .C1(n5749), .C2(
        keyinput_g111), .A(n9813), .ZN(n9823) );
  INV_X1 U11009 ( .A(SI_30_), .ZN(n9815) );
  AOI22_X1 U11010 ( .A1(n9992), .A2(keyinput_g107), .B1(keyinput_g2), .B2(
        n9815), .ZN(n9814) );
  OAI221_X1 U11011 ( .B1(n9992), .B2(keyinput_g107), .C1(n9815), .C2(
        keyinput_g2), .A(n9814), .ZN(n9822) );
  AOI22_X1 U11012 ( .A1(n5759), .A2(keyinput_g116), .B1(keyinput_g9), .B2(
        n9817), .ZN(n9816) );
  OAI221_X1 U11013 ( .B1(n5759), .B2(keyinput_g116), .C1(n9817), .C2(
        keyinput_g9), .A(n9816), .ZN(n9821) );
  XNOR2_X1 U11014 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_g91), .ZN(n9819) );
  XNOR2_X1 U11015 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_g86), .ZN(n9818)
         );
  NAND2_X1 U11016 ( .A1(n9819), .A2(n9818), .ZN(n9820) );
  NOR4_X1 U11017 ( .A1(n9823), .A2(n9822), .A3(n9821), .A4(n9820), .ZN(n9824)
         );
  NAND4_X1 U11018 ( .A1(n9827), .A2(n9826), .A3(n9825), .A4(n9824), .ZN(n9828)
         );
  NOR4_X1 U11019 ( .A1(n9831), .A2(n9830), .A3(n9829), .A4(n9828), .ZN(n10010)
         );
  OAI22_X1 U11020 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput_f115), .B1(
        keyinput_f65), .B2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9832) );
  AOI221_X1 U11021 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(keyinput_f115), .C1(
        P2_DATAO_REG_31__SCAN_IN), .C2(keyinput_f65), .A(n9832), .ZN(n9839) );
  OAI22_X1 U11022 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_f96), .B1(
        keyinput_f87), .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9833) );
  AOI221_X1 U11023 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_f96), .C1(
        P2_DATAO_REG_9__SCAN_IN), .C2(keyinput_f87), .A(n9833), .ZN(n9838) );
  OAI22_X1 U11024 ( .A1(SI_19_), .A2(keyinput_f13), .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .ZN(n9834) );
  AOI221_X1 U11025 ( .B1(SI_19_), .B2(keyinput_f13), .C1(keyinput_f53), .C2(
        P2_REG3_REG_9__SCAN_IN), .A(n9834), .ZN(n9837) );
  OAI22_X1 U11026 ( .A1(SI_4_), .A2(keyinput_f28), .B1(keyinput_f1), .B2(
        SI_31_), .ZN(n9835) );
  AOI221_X1 U11027 ( .B1(SI_4_), .B2(keyinput_f28), .C1(SI_31_), .C2(
        keyinput_f1), .A(n9835), .ZN(n9836) );
  NAND4_X1 U11028 ( .A1(n9839), .A2(n9838), .A3(n9837), .A4(n9836), .ZN(n9867)
         );
  OAI22_X1 U11029 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_f99), .B1(
        keyinput_f80), .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n9840) );
  AOI221_X1 U11030 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput_f99), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput_f80), .A(n9840), .ZN(n9847) );
  OAI22_X1 U11031 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput_f127), .B1(
        keyinput_f121), .B2(P1_IR_REG_30__SCAN_IN), .ZN(n9841) );
  AOI221_X1 U11032 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput_f127), .C1(
        P1_IR_REG_30__SCAN_IN), .C2(keyinput_f121), .A(n9841), .ZN(n9846) );
  OAI22_X1 U11033 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput_f112), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .ZN(n9842) );
  AOI221_X1 U11034 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput_f112), .C1(
        keyinput_f57), .C2(P2_REG3_REG_22__SCAN_IN), .A(n9842), .ZN(n9845) );
  OAI22_X1 U11035 ( .A1(SI_27_), .A2(keyinput_f5), .B1(keyinput_f42), .B2(
        P2_REG3_REG_28__SCAN_IN), .ZN(n9843) );
  AOI221_X1 U11036 ( .B1(SI_27_), .B2(keyinput_f5), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n9843), .ZN(n9844) );
  NAND4_X1 U11037 ( .A1(n9847), .A2(n9846), .A3(n9845), .A4(n9844), .ZN(n9866)
         );
  OAI22_X1 U11038 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_f58), .B1(
        keyinput_f0), .B2(P2_WR_REG_SCAN_IN), .ZN(n9848) );
  AOI221_X1 U11039 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .C1(
        P2_WR_REG_SCAN_IN), .C2(keyinput_f0), .A(n9848), .ZN(n9855) );
  OAI22_X1 U11040 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_f38), .B1(
        keyinput_f61), .B2(P2_REG3_REG_6__SCAN_IN), .ZN(n9849) );
  AOI221_X1 U11041 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .C1(
        P2_REG3_REG_6__SCAN_IN), .C2(keyinput_f61), .A(n9849), .ZN(n9854) );
  OAI22_X1 U11042 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(
        P2_REG3_REG_7__SCAN_IN), .B2(keyinput_f35), .ZN(n9850) );
  AOI221_X1 U11043 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        keyinput_f35), .C2(P2_REG3_REG_7__SCAN_IN), .A(n9850), .ZN(n9853) );
  OAI22_X1 U11044 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_f124), .B1(SI_30_), 
        .B2(keyinput_f2), .ZN(n9851) );
  AOI221_X1 U11045 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_f124), .C1(
        keyinput_f2), .C2(SI_30_), .A(n9851), .ZN(n9852) );
  NAND4_X1 U11046 ( .A1(n9855), .A2(n9854), .A3(n9853), .A4(n9852), .ZN(n9865)
         );
  OAI22_X1 U11047 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput_f117), .B1(SI_2_), 
        .B2(keyinput_f30), .ZN(n9856) );
  AOI221_X1 U11048 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput_f117), .C1(
        keyinput_f30), .C2(SI_2_), .A(n9856), .ZN(n9863) );
  OAI22_X1 U11049 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput_f119), .B1(SI_23_), .B2(keyinput_f9), .ZN(n9857) );
  AOI221_X1 U11050 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput_f119), .C1(
        keyinput_f9), .C2(SI_23_), .A(n9857), .ZN(n9862) );
  OAI22_X1 U11051 ( .A1(SI_25_), .A2(keyinput_f7), .B1(SI_10_), .B2(
        keyinput_f22), .ZN(n9858) );
  AOI221_X1 U11052 ( .B1(SI_25_), .B2(keyinput_f7), .C1(keyinput_f22), .C2(
        SI_10_), .A(n9858), .ZN(n9861) );
  OAI22_X1 U11053 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput_f98), .B1(SI_3_), 
        .B2(keyinput_f29), .ZN(n9859) );
  AOI221_X1 U11054 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput_f98), .C1(
        keyinput_f29), .C2(SI_3_), .A(n9859), .ZN(n9860) );
  NAND4_X1 U11055 ( .A1(n9863), .A2(n9862), .A3(n9861), .A4(n9860), .ZN(n9864)
         );
  NOR4_X1 U11056 ( .A1(n9867), .A2(n9866), .A3(n9865), .A4(n9864), .ZN(n10006)
         );
  OAI22_X1 U11057 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput_f86), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_f89), .ZN(n9868) );
  AOI221_X1 U11058 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_f86), .C1(
        keyinput_f89), .C2(P2_DATAO_REG_7__SCAN_IN), .A(n9868), .ZN(n9875) );
  OAI22_X1 U11059 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(keyinput_f83), .B1(
        keyinput_f34), .B2(P2_STATE_REG_SCAN_IN), .ZN(n9869) );
  AOI221_X1 U11060 ( .B1(P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_f83), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_f34), .A(n9869), .ZN(n9874) );
  OAI22_X1 U11061 ( .A1(P1_D_REG_0__SCAN_IN), .A2(keyinput_f123), .B1(
        keyinput_f26), .B2(SI_6_), .ZN(n9870) );
  AOI221_X1 U11062 ( .B1(P1_D_REG_0__SCAN_IN), .B2(keyinput_f123), .C1(SI_6_), 
        .C2(keyinput_f26), .A(n9870), .ZN(n9873) );
  OAI22_X1 U11063 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput_f101), .B1(SI_20_), .B2(keyinput_f12), .ZN(n9871) );
  AOI221_X1 U11064 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput_f101), .C1(
        keyinput_f12), .C2(SI_20_), .A(n9871), .ZN(n9872) );
  NAND4_X1 U11065 ( .A1(n9875), .A2(n9874), .A3(n9873), .A4(n9872), .ZN(n10004) );
  OAI22_X1 U11066 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_f110), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_f84), .ZN(n9876) );
  AOI221_X1 U11067 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_f110), .C1(
        keyinput_f84), .C2(P2_DATAO_REG_12__SCAN_IN), .A(n9876), .ZN(n9901) );
  OAI22_X1 U11068 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput_f122), .B1(SI_29_), .B2(keyinput_f3), .ZN(n9877) );
  AOI221_X1 U11069 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput_f122), .C1(
        keyinput_f3), .C2(SI_29_), .A(n9877), .ZN(n9880) );
  OAI22_X1 U11070 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(keyinput_f90), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .ZN(n9878) );
  AOI221_X1 U11071 ( .B1(P2_DATAO_REG_6__SCAN_IN), .B2(keyinput_f90), .C1(
        keyinput_f51), .C2(P2_REG3_REG_24__SCAN_IN), .A(n9878), .ZN(n9879) );
  OAI211_X1 U11072 ( .C1(n10359), .C2(keyinput_f54), .A(n9880), .B(n9879), 
        .ZN(n9881) );
  AOI21_X1 U11073 ( .B1(n10359), .B2(keyinput_f54), .A(n9881), .ZN(n9900) );
  AOI22_X1 U11074 ( .A1(SI_9_), .A2(keyinput_f23), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_f72), .ZN(n9882) );
  OAI221_X1 U11075 ( .B1(SI_9_), .B2(keyinput_f23), .C1(
        P2_DATAO_REG_24__SCAN_IN), .C2(keyinput_f72), .A(n9882), .ZN(n9889) );
  AOI22_X1 U11076 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_f37), .B1(
        P1_D_REG_2__SCAN_IN), .B2(keyinput_f125), .ZN(n9883) );
  OAI221_X1 U11077 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .C1(
        P1_D_REG_2__SCAN_IN), .C2(keyinput_f125), .A(n9883), .ZN(n9888) );
  AOI22_X1 U11078 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(keyinput_f69), .B1(
        P1_IR_REG_20__SCAN_IN), .B2(keyinput_f111), .ZN(n9884) );
  OAI221_X1 U11079 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_f69), .C1(
        P1_IR_REG_20__SCAN_IN), .C2(keyinput_f111), .A(n9884), .ZN(n9887) );
  AOI22_X1 U11080 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_f52), .B1(
        P2_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .ZN(n9885) );
  OAI221_X1 U11081 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .C1(
        P2_REG3_REG_8__SCAN_IN), .C2(keyinput_f43), .A(n9885), .ZN(n9886) );
  NOR4_X1 U11082 ( .A1(n9889), .A2(n9888), .A3(n9887), .A4(n9886), .ZN(n9899)
         );
  AOI22_X1 U11083 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(keyinput_f81), .B1(
        SI_26_), .B2(keyinput_f6), .ZN(n9890) );
  OAI221_X1 U11084 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_f81), .C1(
        SI_26_), .C2(keyinput_f6), .A(n9890), .ZN(n9897) );
  AOI22_X1 U11085 ( .A1(SI_8_), .A2(keyinput_f24), .B1(SI_17_), .B2(
        keyinput_f15), .ZN(n9891) );
  OAI221_X1 U11086 ( .B1(SI_8_), .B2(keyinput_f24), .C1(SI_17_), .C2(
        keyinput_f15), .A(n9891), .ZN(n9896) );
  AOI22_X1 U11087 ( .A1(SI_1_), .A2(keyinput_f31), .B1(SI_5_), .B2(
        keyinput_f27), .ZN(n9892) );
  OAI221_X1 U11088 ( .B1(SI_1_), .B2(keyinput_f31), .C1(SI_5_), .C2(
        keyinput_f27), .A(n9892), .ZN(n9895) );
  AOI22_X1 U11089 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_f41), .B1(
        P1_IR_REG_27__SCAN_IN), .B2(keyinput_f118), .ZN(n9893) );
  OAI221_X1 U11090 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .C1(
        P1_IR_REG_27__SCAN_IN), .C2(keyinput_f118), .A(n9893), .ZN(n9894) );
  NOR4_X1 U11091 ( .A1(n9897), .A2(n9896), .A3(n9895), .A4(n9894), .ZN(n9898)
         );
  NAND4_X1 U11092 ( .A1(n9901), .A2(n9900), .A3(n9899), .A4(n9898), .ZN(n10003) );
  AOI22_X1 U11093 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_f85), .ZN(n9902) );
  OAI221_X1 U11094 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(
        P2_DATAO_REG_11__SCAN_IN), .C2(keyinput_f85), .A(n9902), .ZN(n9909) );
  AOI22_X1 U11095 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput_f126), .B1(
        P1_IR_REG_13__SCAN_IN), .B2(keyinput_f104), .ZN(n9903) );
  OAI221_X1 U11096 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput_f126), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput_f104), .A(n9903), .ZN(n9908) );
  AOI22_X1 U11097 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput_f66), .B1(
        SI_13_), .B2(keyinput_f19), .ZN(n9904) );
  OAI221_X1 U11098 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_f66), .C1(
        SI_13_), .C2(keyinput_f19), .A(n9904), .ZN(n9907) );
  AOI22_X1 U11099 ( .A1(SI_12_), .A2(keyinput_f20), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_f76), .ZN(n9905) );
  OAI221_X1 U11100 ( .B1(SI_12_), .B2(keyinput_f20), .C1(
        P2_DATAO_REG_20__SCAN_IN), .C2(keyinput_f76), .A(n9905), .ZN(n9906) );
  NOR4_X1 U11101 ( .A1(n9909), .A2(n9908), .A3(n9907), .A4(n9906), .ZN(n9948)
         );
  AOI22_X1 U11102 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(keyinput_f68), .B1(
        SI_15_), .B2(keyinput_f17), .ZN(n9910) );
  OAI221_X1 U11103 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_f68), .C1(
        SI_15_), .C2(keyinput_f17), .A(n9910), .ZN(n9918) );
  AOI22_X1 U11104 ( .A1(SI_14_), .A2(keyinput_f18), .B1(P1_IR_REG_25__SCAN_IN), 
        .B2(keyinput_f116), .ZN(n9911) );
  OAI221_X1 U11105 ( .B1(SI_14_), .B2(keyinput_f18), .C1(P1_IR_REG_25__SCAN_IN), .C2(keyinput_f116), .A(n9911), .ZN(n9917) );
  AOI22_X1 U11106 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_f59), .B1(
        P1_IR_REG_17__SCAN_IN), .B2(keyinput_f108), .ZN(n9912) );
  OAI221_X1 U11107 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_f59), .C1(
        P1_IR_REG_17__SCAN_IN), .C2(keyinput_f108), .A(n9912), .ZN(n9916) );
  AOI22_X1 U11108 ( .A1(n9914), .A2(keyinput_f82), .B1(keyinput_f44), .B2(
        n10024), .ZN(n9913) );
  OAI221_X1 U11109 ( .B1(n9914), .B2(keyinput_f82), .C1(n10024), .C2(
        keyinput_f44), .A(n9913), .ZN(n9915) );
  NOR4_X1 U11110 ( .A1(n9918), .A2(n9917), .A3(n9916), .A4(n9915), .ZN(n9947)
         );
  AOI22_X1 U11111 ( .A1(n9921), .A2(keyinput_f71), .B1(keyinput_f78), .B2(
        n9920), .ZN(n9919) );
  OAI221_X1 U11112 ( .B1(n9921), .B2(keyinput_f71), .C1(n9920), .C2(
        keyinput_f78), .A(n9919), .ZN(n9933) );
  AOI22_X1 U11113 ( .A1(n9924), .A2(keyinput_f49), .B1(n9923), .B2(keyinput_f8), .ZN(n9922) );
  OAI221_X1 U11114 ( .B1(n9924), .B2(keyinput_f49), .C1(n9923), .C2(
        keyinput_f8), .A(n9922), .ZN(n9932) );
  AOI22_X1 U11115 ( .A1(n9927), .A2(keyinput_f25), .B1(keyinput_f67), .B2(
        n9926), .ZN(n9925) );
  OAI221_X1 U11116 ( .B1(n9927), .B2(keyinput_f25), .C1(n9926), .C2(
        keyinput_f67), .A(n9925), .ZN(n9931) );
  AOI22_X1 U11117 ( .A1(n9929), .A2(keyinput_f74), .B1(keyinput_f63), .B2(
        n8340), .ZN(n9928) );
  OAI221_X1 U11118 ( .B1(n9929), .B2(keyinput_f74), .C1(n8340), .C2(
        keyinput_f63), .A(n9928), .ZN(n9930) );
  NOR4_X1 U11119 ( .A1(n9933), .A2(n9932), .A3(n9931), .A4(n9930), .ZN(n9946)
         );
  AOI22_X1 U11120 ( .A1(n9935), .A2(keyinput_f36), .B1(n4625), .B2(
        keyinput_f92), .ZN(n9934) );
  OAI221_X1 U11121 ( .B1(n9935), .B2(keyinput_f36), .C1(n4625), .C2(
        keyinput_f92), .A(n9934), .ZN(n9944) );
  AOI22_X1 U11122 ( .A1(n4886), .A2(keyinput_f103), .B1(keyinput_f79), .B2(
        n9937), .ZN(n9936) );
  OAI221_X1 U11123 ( .B1(n4886), .B2(keyinput_f103), .C1(n9937), .C2(
        keyinput_f79), .A(n9936), .ZN(n9943) );
  XNOR2_X1 U11124 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_f60), .ZN(n9941)
         );
  XNOR2_X1 U11125 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_f91), .ZN(n9940) );
  XNOR2_X1 U11126 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_f97), .ZN(n9939) );
  XNOR2_X1 U11127 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_f62), .ZN(n9938)
         );
  NAND4_X1 U11128 ( .A1(n9941), .A2(n9940), .A3(n9939), .A4(n9938), .ZN(n9942)
         );
  NOR3_X1 U11129 ( .A1(n9944), .A2(n9943), .A3(n9942), .ZN(n9945) );
  NAND4_X1 U11130 ( .A1(n9948), .A2(n9947), .A3(n9946), .A4(n9945), .ZN(n10002) );
  AOI22_X1 U11131 ( .A1(n9950), .A2(keyinput_f77), .B1(n5750), .B2(
        keyinput_f109), .ZN(n9949) );
  OAI221_X1 U11132 ( .B1(n9950), .B2(keyinput_f77), .C1(n5750), .C2(
        keyinput_f109), .A(n9949), .ZN(n9962) );
  AOI22_X1 U11133 ( .A1(n9953), .A2(keyinput_f11), .B1(n9952), .B2(
        keyinput_f100), .ZN(n9951) );
  OAI221_X1 U11134 ( .B1(n9953), .B2(keyinput_f11), .C1(n9952), .C2(
        keyinput_f100), .A(n9951), .ZN(n9961) );
  AOI22_X1 U11135 ( .A1(n9956), .A2(keyinput_f64), .B1(keyinput_f45), .B2(
        n9955), .ZN(n9954) );
  OAI221_X1 U11136 ( .B1(n9956), .B2(keyinput_f64), .C1(n9955), .C2(
        keyinput_f45), .A(n9954), .ZN(n9960) );
  XNOR2_X1 U11137 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_f114), .ZN(n9958)
         );
  XNOR2_X1 U11138 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_f55), .ZN(n9957)
         );
  NAND2_X1 U11139 ( .A1(n9958), .A2(n9957), .ZN(n9959) );
  NOR4_X1 U11140 ( .A1(n9962), .A2(n9961), .A3(n9960), .A4(n9959), .ZN(n10000)
         );
  XNOR2_X1 U11141 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_f106), .ZN(n9966)
         );
  XNOR2_X1 U11142 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_f46), .ZN(n9965)
         );
  XNOR2_X1 U11143 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_f95), .ZN(n9964) );
  XNOR2_X1 U11144 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_f48), .ZN(n9963)
         );
  NAND4_X1 U11145 ( .A1(n9966), .A2(n9965), .A3(n9964), .A4(n9963), .ZN(n9972)
         );
  XNOR2_X1 U11146 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_f120), .ZN(n9970)
         );
  XNOR2_X1 U11147 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_f33), .ZN(n9969) );
  XNOR2_X1 U11148 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_f102), .ZN(n9968)
         );
  XNOR2_X1 U11149 ( .A(SI_16_), .B(keyinput_f16), .ZN(n9967) );
  NAND4_X1 U11150 ( .A1(n9970), .A2(n9969), .A3(n9968), .A4(n9967), .ZN(n9971)
         );
  NOR2_X1 U11151 ( .A1(n9972), .A2(n9971), .ZN(n9999) );
  AOI22_X1 U11152 ( .A1(n5488), .A2(keyinput_f75), .B1(keyinput_f56), .B2(
        n7282), .ZN(n9973) );
  OAI221_X1 U11153 ( .B1(n5488), .B2(keyinput_f75), .C1(n7282), .C2(
        keyinput_f56), .A(n9973), .ZN(n9984) );
  AOI22_X1 U11154 ( .A1(n5519), .A2(keyinput_f73), .B1(keyinput_f21), .B2(
        n9975), .ZN(n9974) );
  OAI221_X1 U11155 ( .B1(n5519), .B2(keyinput_f73), .C1(n9975), .C2(
        keyinput_f21), .A(n9974), .ZN(n9983) );
  AOI22_X1 U11156 ( .A1(n9978), .A2(keyinput_f70), .B1(keyinput_f39), .B2(
        n9977), .ZN(n9976) );
  OAI221_X1 U11157 ( .B1(n9978), .B2(keyinput_f70), .C1(n9977), .C2(
        keyinput_f39), .A(n9976), .ZN(n9982) );
  XOR2_X1 U11158 ( .A(n5441), .B(keyinput_f50), .Z(n9980) );
  XNOR2_X1 U11159 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_f105), .ZN(n9979)
         );
  NAND2_X1 U11160 ( .A1(n9980), .A2(n9979), .ZN(n9981) );
  NOR4_X1 U11161 ( .A1(n9984), .A2(n9983), .A3(n9982), .A4(n9981), .ZN(n9998)
         );
  AOI22_X1 U11162 ( .A1(n5727), .A2(keyinput_f93), .B1(keyinput_f4), .B2(n5626), .ZN(n9985) );
  OAI221_X1 U11163 ( .B1(n5727), .B2(keyinput_f93), .C1(n5626), .C2(
        keyinput_f4), .A(n9985), .ZN(n9996) );
  INV_X1 U11164 ( .A(SI_18_), .ZN(n9988) );
  AOI22_X1 U11165 ( .A1(n9988), .A2(keyinput_f14), .B1(keyinput_f88), .B2(
        n9987), .ZN(n9986) );
  OAI221_X1 U11166 ( .B1(n9988), .B2(keyinput_f14), .C1(n9987), .C2(
        keyinput_f88), .A(n9986), .ZN(n9995) );
  AOI22_X1 U11167 ( .A1(n5767), .A2(keyinput_f113), .B1(keyinput_f94), .B2(
        n5728), .ZN(n9989) );
  OAI221_X1 U11168 ( .B1(n5767), .B2(keyinput_f113), .C1(n5728), .C2(
        keyinput_f94), .A(n9989), .ZN(n9994) );
  AOI22_X1 U11169 ( .A1(n9992), .A2(keyinput_f107), .B1(keyinput_f10), .B2(
        n9991), .ZN(n9990) );
  OAI221_X1 U11170 ( .B1(n9992), .B2(keyinput_f107), .C1(n9991), .C2(
        keyinput_f10), .A(n9990), .ZN(n9993) );
  NOR4_X1 U11171 ( .A1(n9996), .A2(n9995), .A3(n9994), .A4(n9993), .ZN(n9997)
         );
  NAND4_X1 U11172 ( .A1(n10000), .A2(n9999), .A3(n9998), .A4(n9997), .ZN(
        n10001) );
  NOR4_X1 U11173 ( .A1(n10004), .A2(n10003), .A3(n10002), .A4(n10001), .ZN(
        n10005) );
  AOI22_X1 U11174 ( .A1(n10006), .A2(n10005), .B1(keyinput_f32), .B2(SI_0_), 
        .ZN(n10007) );
  OAI21_X1 U11175 ( .B1(keyinput_f32), .B2(SI_0_), .A(n10007), .ZN(n10008) );
  OAI21_X1 U11176 ( .B1(n10011), .B2(keyinput_g32), .A(n10008), .ZN(n10009) );
  AOI211_X1 U11177 ( .C1(n10011), .C2(keyinput_g32), .A(n10010), .B(n10009), 
        .ZN(n10012) );
  XNOR2_X1 U11178 ( .A(n10013), .B(n10012), .ZN(n10017) );
  NOR2_X1 U11179 ( .A1(n10015), .A2(n10014), .ZN(n10016) );
  XOR2_X1 U11180 ( .A(n10017), .B(n10016), .Z(ADD_1071_U4) );
  NAND2_X1 U11181 ( .A1(n10355), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10018) );
  NAND2_X1 U11182 ( .A1(n10019), .A2(n10018), .ZN(n10022) );
  INV_X1 U11183 ( .A(n10020), .ZN(n10021) );
  NAND2_X1 U11184 ( .A1(n10022), .A2(n10021), .ZN(n10030) );
  NAND2_X1 U11185 ( .A1(n10042), .A2(n10023), .ZN(n10029) );
  OAI22_X1 U11186 ( .A1(n10026), .A2(n10025), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10024), .ZN(n10027) );
  INV_X1 U11187 ( .A(n10027), .ZN(n10028) );
  OAI211_X1 U11188 ( .C1(n10030), .C2(n10347), .A(n10029), .B(n10028), .ZN(
        n10031) );
  INV_X1 U11189 ( .A(n10031), .ZN(n10036) );
  NOR2_X1 U11190 ( .A1(n10353), .A2(n5203), .ZN(n10034) );
  OAI211_X1 U11191 ( .C1(n10034), .C2(n10033), .A(n10342), .B(n10032), .ZN(
        n10035) );
  NAND2_X1 U11192 ( .A1(n10036), .A2(n10035), .ZN(P2_U3246) );
  AOI22_X1 U11193 ( .A1(n10350), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10048) );
  AOI211_X1 U11194 ( .C1(n10039), .C2(n10038), .A(n10037), .B(n10347), .ZN(
        n10040) );
  AOI21_X1 U11195 ( .B1(n10042), .B2(n10041), .A(n10040), .ZN(n10047) );
  OAI211_X1 U11196 ( .C1(n10045), .C2(n10044), .A(n10342), .B(n10043), .ZN(
        n10046) );
  NAND3_X1 U11197 ( .A1(n10048), .A2(n10047), .A3(n10046), .ZN(P2_U3247) );
  NAND2_X1 U11198 ( .A1(n10050), .A2(n10049), .ZN(n10051) );
  AOI21_X1 U11199 ( .B1(n10052), .B2(n10330), .A(n10051), .ZN(n10053) );
  AND2_X1 U11200 ( .A1(n10054), .A2(n10053), .ZN(n10056) );
  INV_X1 U11201 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10055) );
  AOI22_X1 U11202 ( .A1(n10333), .A2(n10056), .B1(n10055), .B2(n10331), .ZN(
        P1_U3484) );
  AOI22_X1 U11203 ( .A1(n10341), .A2(n10056), .B1(n6885), .B2(n10339), .ZN(
        P1_U3533) );
  INV_X1 U11204 ( .A(n10057), .ZN(n10058) );
  OAI21_X1 U11205 ( .B1(n10092), .B2(n10059), .A(n10058), .ZN(n10063) );
  NOR2_X1 U11206 ( .A1(n10061), .A2(n10060), .ZN(n10062) );
  NOR2_X1 U11207 ( .A1(n10063), .A2(n10062), .ZN(n10070) );
  OAI21_X1 U11208 ( .B1(n10065), .B2(n4572), .A(n10064), .ZN(n10068) );
  NOR2_X1 U11209 ( .A1(n10066), .A2(n10323), .ZN(n10160) );
  AOI22_X1 U11210 ( .A1(n10068), .A2(n10101), .B1(n10067), .B2(n10160), .ZN(
        n10069) );
  OAI211_X1 U11211 ( .C1(n10106), .C2(n10071), .A(n10070), .B(n10069), .ZN(
        P1_U3222) );
  OAI21_X1 U11212 ( .B1(n10073), .B2(n10434), .A(n10072), .ZN(n10074) );
  AOI21_X1 U11213 ( .B1(n10075), .B2(n8951), .A(n10074), .ZN(n10085) );
  INV_X1 U11214 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10076) );
  AOI22_X1 U11215 ( .A1(n10452), .A2(n10085), .B1(n10076), .B2(n10450), .ZN(
        P2_U3550) );
  INV_X1 U11216 ( .A(n10077), .ZN(n10423) );
  INV_X1 U11217 ( .A(n10078), .ZN(n10084) );
  INV_X1 U11218 ( .A(n10079), .ZN(n10080) );
  OAI22_X1 U11219 ( .A1(n10081), .A2(n10436), .B1(n10080), .B2(n10434), .ZN(
        n10083) );
  AOI211_X1 U11220 ( .C1(n10423), .C2(n10084), .A(n10083), .B(n10082), .ZN(
        n10087) );
  AOI22_X1 U11221 ( .A1(n10452), .A2(n10087), .B1(n5377), .B2(n10450), .ZN(
        P2_U3533) );
  AOI22_X1 U11222 ( .A1(n10444), .A2(n10085), .B1(n5677), .B2(n10442), .ZN(
        P2_U3518) );
  INV_X1 U11223 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10086) );
  AOI22_X1 U11224 ( .A1(n10444), .A2(n10087), .B1(n10086), .B2(n10442), .ZN(
        P2_U3490) );
  NOR2_X1 U11225 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10088), .ZN(n10198) );
  AOI21_X1 U11226 ( .B1(n10090), .B2(n10089), .A(n10198), .ZN(n10091) );
  OAI21_X1 U11227 ( .B1(n10093), .B2(n10092), .A(n10091), .ZN(n10094) );
  AOI21_X1 U11228 ( .B1(n10096), .B2(n10095), .A(n10094), .ZN(n10104) );
  XNOR2_X1 U11229 ( .A(n10098), .B(n10097), .ZN(n10099) );
  XNOR2_X1 U11230 ( .A(n10100), .B(n10099), .ZN(n10102) );
  NAND2_X1 U11231 ( .A1(n10102), .A2(n10101), .ZN(n10103) );
  OAI211_X1 U11232 ( .C1(n10106), .C2(n10105), .A(n10104), .B(n10103), .ZN(
        P1_U3213) );
  OAI21_X1 U11233 ( .B1(n10113), .B2(n10108), .A(n10107), .ZN(n10116) );
  OAI22_X1 U11234 ( .A1(n10127), .A2(n10129), .B1(n10128), .B2(n10109), .ZN(
        n10115) );
  NAND2_X1 U11235 ( .A1(n10111), .A2(n10110), .ZN(n10112) );
  XOR2_X1 U11236 ( .A(n10113), .B(n10112), .Z(n10156) );
  NOR2_X1 U11237 ( .A1(n10156), .A2(n10272), .ZN(n10114) );
  AOI211_X1 U11238 ( .C1(n10266), .C2(n10116), .A(n10115), .B(n10114), .ZN(
        n10155) );
  INV_X1 U11239 ( .A(n10117), .ZN(n10118) );
  AOI222_X1 U11240 ( .A1(n10122), .A2(n10276), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n4483), .C1(n10275), .C2(n10118), .ZN(n10125) );
  INV_X1 U11241 ( .A(n10156), .ZN(n10123) );
  INV_X1 U11242 ( .A(n10119), .ZN(n10121) );
  AOI21_X1 U11243 ( .B1(n10122), .B2(n10121), .A(n10120), .ZN(n10153) );
  AOI22_X1 U11244 ( .A1(n10123), .A2(n10283), .B1(n10282), .B2(n10153), .ZN(
        n10124) );
  OAI211_X1 U11245 ( .C1(n4483), .C2(n10155), .A(n10125), .B(n10124), .ZN(
        P1_U3278) );
  XNOR2_X1 U11246 ( .A(n10126), .B(n4857), .ZN(n10135) );
  OAI22_X1 U11247 ( .A1(n10130), .A2(n10129), .B1(n10128), .B2(n10127), .ZN(
        n10134) );
  XNOR2_X1 U11248 ( .A(n10132), .B(n10131), .ZN(n10169) );
  NOR2_X1 U11249 ( .A1(n10169), .A2(n10272), .ZN(n10133) );
  AOI211_X1 U11250 ( .C1(n10135), .C2(n10266), .A(n10134), .B(n10133), .ZN(
        n10168) );
  INV_X1 U11251 ( .A(n10136), .ZN(n10137) );
  AOI222_X1 U11252 ( .A1(n10163), .A2(n10276), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n4483), .C1(n10137), .C2(n10275), .ZN(n10142) );
  INV_X1 U11253 ( .A(n10169), .ZN(n10140) );
  AOI21_X1 U11254 ( .B1(n10163), .B2(n10139), .A(n10138), .ZN(n10166) );
  AOI22_X1 U11255 ( .A1(n10140), .A2(n10283), .B1(n10282), .B2(n10166), .ZN(
        n10141) );
  OAI211_X1 U11256 ( .C1(n4483), .C2(n10168), .A(n10142), .B(n10141), .ZN(
        P1_U3280) );
  NOR2_X1 U11257 ( .A1(n10143), .A2(n10325), .ZN(n10144) );
  AOI22_X1 U11258 ( .A1(n10341), .A2(n10173), .B1(n8075), .B2(n10339), .ZN(
        P1_U3553) );
  OAI21_X1 U11259 ( .B1(n10148), .B2(n10323), .A(n10147), .ZN(n10149) );
  AOI211_X1 U11260 ( .C1(n10151), .C2(n10320), .A(n10150), .B(n10149), .ZN(
        n10175) );
  AOI22_X1 U11261 ( .A1(n10341), .A2(n10175), .B1(n9183), .B2(n10339), .ZN(
        P1_U3537) );
  AOI21_X1 U11262 ( .B1(n10153), .B2(n10165), .A(n10152), .ZN(n10154) );
  OAI211_X1 U11263 ( .C1(n10170), .C2(n10156), .A(n10155), .B(n10154), .ZN(
        n10157) );
  INV_X1 U11264 ( .A(n10157), .ZN(n10177) );
  AOI22_X1 U11265 ( .A1(n10341), .A2(n10177), .B1(n9182), .B2(n10339), .ZN(
        P1_U3536) );
  NOR2_X1 U11266 ( .A1(n10158), .A2(n10170), .ZN(n10161) );
  NOR4_X1 U11267 ( .A1(n10162), .A2(n10161), .A3(n10160), .A4(n10159), .ZN(
        n10179) );
  AOI22_X1 U11268 ( .A1(n10341), .A2(n10179), .B1(n6009), .B2(n10339), .ZN(
        P1_U3535) );
  AOI22_X1 U11269 ( .A1(n10166), .A2(n10165), .B1(n10164), .B2(n10163), .ZN(
        n10167) );
  OAI211_X1 U11270 ( .C1(n10170), .C2(n10169), .A(n10168), .B(n10167), .ZN(
        n10171) );
  INV_X1 U11271 ( .A(n10171), .ZN(n10181) );
  AOI22_X1 U11272 ( .A1(n10341), .A2(n10181), .B1(n6971), .B2(n10339), .ZN(
        P1_U3534) );
  INV_X1 U11273 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U11274 ( .A1(n10333), .A2(n10173), .B1(n10172), .B2(n10331), .ZN(
        P1_U3521) );
  INV_X1 U11275 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U11276 ( .A1(n10333), .A2(n10175), .B1(n10174), .B2(n10331), .ZN(
        P1_U3496) );
  INV_X1 U11277 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U11278 ( .A1(n10333), .A2(n10177), .B1(n10176), .B2(n10331), .ZN(
        P1_U3493) );
  INV_X1 U11279 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10178) );
  AOI22_X1 U11280 ( .A1(n10333), .A2(n10179), .B1(n10178), .B2(n10331), .ZN(
        P1_U3490) );
  INV_X1 U11281 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U11282 ( .A1(n10333), .A2(n10181), .B1(n10180), .B2(n10331), .ZN(
        P1_U3487) );
  XNOR2_X1 U11283 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U11284 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10194) );
  AOI211_X1 U11285 ( .C1(n10184), .C2(n10183), .A(n10182), .B(n10245), .ZN(
        n10185) );
  AOI211_X1 U11286 ( .C1(n10251), .C2(n10187), .A(n10186), .B(n10185), .ZN(
        n10193) );
  AOI21_X1 U11287 ( .B1(n10190), .B2(n10189), .A(n10188), .ZN(n10191) );
  OR2_X1 U11288 ( .A1(n10191), .A2(n10257), .ZN(n10192) );
  OAI211_X1 U11289 ( .C1(n10194), .C2(n10260), .A(n10193), .B(n10192), .ZN(
        P1_U3254) );
  INV_X1 U11290 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10206) );
  AOI211_X1 U11291 ( .C1(n10196), .C2(n7906), .A(n10195), .B(n10245), .ZN(
        n10197) );
  AOI211_X1 U11292 ( .C1(n10251), .C2(n10199), .A(n10198), .B(n10197), .ZN(
        n10205) );
  AOI21_X1 U11293 ( .B1(n10202), .B2(n10201), .A(n10200), .ZN(n10203) );
  OR2_X1 U11294 ( .A1(n10257), .A2(n10203), .ZN(n10204) );
  OAI211_X1 U11295 ( .C1(n10206), .C2(n10260), .A(n10205), .B(n10204), .ZN(
        P1_U3255) );
  INV_X1 U11296 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10217) );
  INV_X1 U11297 ( .A(n10207), .ZN(n10211) );
  AOI211_X1 U11298 ( .C1(n10209), .C2(n9507), .A(n10208), .B(n10245), .ZN(
        n10210) );
  AOI211_X1 U11299 ( .C1(n10212), .C2(n10251), .A(n10211), .B(n10210), .ZN(
        n10216) );
  OAI211_X1 U11300 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n10214), .A(n10238), 
        .B(n10213), .ZN(n10215) );
  OAI211_X1 U11301 ( .C1(n10217), .C2(n10260), .A(n10216), .B(n10215), .ZN(
        P1_U3256) );
  INV_X1 U11302 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10229) );
  INV_X1 U11303 ( .A(n10218), .ZN(n10222) );
  AOI211_X1 U11304 ( .C1(n4568), .C2(n10220), .A(n10219), .B(n10245), .ZN(
        n10221) );
  AOI211_X1 U11305 ( .C1(n10223), .C2(n10251), .A(n10222), .B(n10221), .ZN(
        n10228) );
  OAI211_X1 U11306 ( .C1(n10226), .C2(n10225), .A(n10238), .B(n10224), .ZN(
        n10227) );
  OAI211_X1 U11307 ( .C1(n10229), .C2(n10260), .A(n10228), .B(n10227), .ZN(
        P1_U3257) );
  INV_X1 U11308 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10243) );
  INV_X1 U11309 ( .A(n10230), .ZN(n10235) );
  AOI211_X1 U11310 ( .C1(n10233), .C2(n10232), .A(n10231), .B(n10245), .ZN(
        n10234) );
  AOI211_X1 U11311 ( .C1(n10236), .C2(n10251), .A(n10235), .B(n10234), .ZN(
        n10242) );
  OAI211_X1 U11312 ( .C1(n10240), .C2(n10239), .A(n10238), .B(n10237), .ZN(
        n10241) );
  OAI211_X1 U11313 ( .C1(n10243), .C2(n10260), .A(n10242), .B(n10241), .ZN(
        P1_U3258) );
  INV_X1 U11314 ( .A(n10244), .ZN(n10250) );
  AOI211_X1 U11315 ( .C1(n10248), .C2(n10247), .A(n10246), .B(n10245), .ZN(
        n10249) );
  AOI211_X1 U11316 ( .C1(n10252), .C2(n10251), .A(n10250), .B(n10249), .ZN(
        n10259) );
  AOI21_X1 U11317 ( .B1(n10255), .B2(n10254), .A(n10253), .ZN(n10256) );
  OR2_X1 U11318 ( .A1(n10257), .A2(n10256), .ZN(n10258) );
  OAI211_X1 U11319 ( .C1(n10492), .C2(n10260), .A(n10259), .B(n10258), .ZN(
        P1_U3259) );
  XOR2_X1 U11320 ( .A(n10268), .B(n10261), .Z(n10278) );
  AOI22_X1 U11321 ( .A1(n10265), .A2(n10264), .B1(n10263), .B2(n10262), .ZN(
        n10271) );
  OAI211_X1 U11322 ( .C1(n10269), .C2(n10268), .A(n10267), .B(n10266), .ZN(
        n10270) );
  OAI211_X1 U11323 ( .C1(n10278), .C2(n10272), .A(n10271), .B(n10270), .ZN(
        n10327) );
  INV_X1 U11324 ( .A(n10327), .ZN(n10286) );
  INV_X1 U11325 ( .A(n10273), .ZN(n10274) );
  AOI222_X1 U11326 ( .A1(n10277), .A2(n10276), .B1(P1_REG2_REG_9__SCAN_IN), 
        .B2(n4483), .C1(n10275), .C2(n10274), .ZN(n10285) );
  INV_X1 U11327 ( .A(n10278), .ZN(n10329) );
  OAI21_X1 U11328 ( .B1(n10280), .B2(n10324), .A(n10279), .ZN(n10326) );
  INV_X1 U11329 ( .A(n10326), .ZN(n10281) );
  AOI22_X1 U11330 ( .A1(n10329), .A2(n10283), .B1(n10282), .B2(n10281), .ZN(
        n10284) );
  OAI211_X1 U11331 ( .C1(n4483), .C2(n10286), .A(n10285), .B(n10284), .ZN(
        P1_U3282) );
  NAND2_X1 U11332 ( .A1(n10288), .A2(n10287), .ZN(n10289) );
  AND2_X1 U11333 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10289), .ZN(P1_U3292) );
  AND2_X1 U11334 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10289), .ZN(P1_U3293) );
  AND2_X1 U11335 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10289), .ZN(P1_U3294) );
  AND2_X1 U11336 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10289), .ZN(P1_U3295) );
  AND2_X1 U11337 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10289), .ZN(P1_U3296) );
  AND2_X1 U11338 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10289), .ZN(P1_U3297) );
  AND2_X1 U11339 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10289), .ZN(P1_U3298) );
  AND2_X1 U11340 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10289), .ZN(P1_U3299) );
  AND2_X1 U11341 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10289), .ZN(P1_U3300) );
  AND2_X1 U11342 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10289), .ZN(P1_U3301) );
  AND2_X1 U11343 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10289), .ZN(P1_U3302) );
  AND2_X1 U11344 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10289), .ZN(P1_U3303) );
  AND2_X1 U11345 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10289), .ZN(P1_U3304) );
  AND2_X1 U11346 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10289), .ZN(P1_U3305) );
  AND2_X1 U11347 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10289), .ZN(P1_U3306) );
  AND2_X1 U11348 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10289), .ZN(P1_U3307) );
  AND2_X1 U11349 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10289), .ZN(P1_U3308) );
  AND2_X1 U11350 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10289), .ZN(P1_U3309) );
  AND2_X1 U11351 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10289), .ZN(P1_U3310) );
  AND2_X1 U11352 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10289), .ZN(P1_U3311) );
  AND2_X1 U11353 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10289), .ZN(P1_U3312) );
  AND2_X1 U11354 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10289), .ZN(P1_U3313) );
  AND2_X1 U11355 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10289), .ZN(P1_U3314) );
  AND2_X1 U11356 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10289), .ZN(P1_U3315) );
  AND2_X1 U11357 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10289), .ZN(P1_U3316) );
  AND2_X1 U11358 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10289), .ZN(P1_U3317) );
  AND2_X1 U11359 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10289), .ZN(P1_U3318) );
  AND2_X1 U11360 ( .A1(n10289), .A2(P1_D_REG_4__SCAN_IN), .ZN(P1_U3319) );
  AND2_X1 U11361 ( .A1(n10289), .A2(P1_D_REG_3__SCAN_IN), .ZN(P1_U3320) );
  AND2_X1 U11362 ( .A1(n10289), .A2(P1_D_REG_2__SCAN_IN), .ZN(P1_U3321) );
  INV_X1 U11363 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U11364 ( .A1(n10333), .A2(n10291), .B1(n10290), .B2(n10331), .ZN(
        P1_U3457) );
  OAI22_X1 U11365 ( .A1(n10293), .A2(n10325), .B1(n10292), .B2(n10323), .ZN(
        n10295) );
  AOI211_X1 U11366 ( .C1(n10330), .C2(n10296), .A(n10295), .B(n10294), .ZN(
        n10334) );
  INV_X1 U11367 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U11368 ( .A1(n10333), .A2(n10334), .B1(n10297), .B2(n10331), .ZN(
        P1_U3463) );
  NOR2_X1 U11369 ( .A1(n10299), .A2(n10298), .ZN(n10303) );
  NOR4_X1 U11370 ( .A1(n10303), .A2(n10302), .A3(n10301), .A4(n10300), .ZN(
        n10335) );
  AOI22_X1 U11371 ( .A1(n10333), .A2(n10335), .B1(n5867), .B2(n10331), .ZN(
        P1_U3469) );
  OAI22_X1 U11372 ( .A1(n10305), .A2(n10325), .B1(n10304), .B2(n10323), .ZN(
        n10307) );
  AOI211_X1 U11373 ( .C1(n10330), .C2(n10308), .A(n10307), .B(n10306), .ZN(
        n10336) );
  INV_X1 U11374 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U11375 ( .A1(n10333), .A2(n10336), .B1(n10309), .B2(n10331), .ZN(
        P1_U3472) );
  OAI211_X1 U11376 ( .C1(n10312), .C2(n10323), .A(n10311), .B(n10310), .ZN(
        n10313) );
  AOI21_X1 U11377 ( .B1(n10320), .B2(n10314), .A(n10313), .ZN(n10337) );
  INV_X1 U11378 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10315) );
  AOI22_X1 U11379 ( .A1(n10333), .A2(n10337), .B1(n10315), .B2(n10331), .ZN(
        P1_U3475) );
  OAI22_X1 U11380 ( .A1(n10317), .A2(n10325), .B1(n10316), .B2(n10323), .ZN(
        n10318) );
  AOI211_X1 U11381 ( .C1(n10321), .C2(n10320), .A(n10319), .B(n10318), .ZN(
        n10338) );
  INV_X1 U11382 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10322) );
  AOI22_X1 U11383 ( .A1(n10333), .A2(n10338), .B1(n10322), .B2(n10331), .ZN(
        P1_U3478) );
  OAI22_X1 U11384 ( .A1(n10326), .A2(n10325), .B1(n10324), .B2(n10323), .ZN(
        n10328) );
  AOI211_X1 U11385 ( .C1(n10330), .C2(n10329), .A(n10328), .B(n10327), .ZN(
        n10340) );
  INV_X1 U11386 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U11387 ( .A1(n10333), .A2(n10340), .B1(n10332), .B2(n10331), .ZN(
        P1_U3481) );
  AOI22_X1 U11388 ( .A1(n10341), .A2(n10334), .B1(n6642), .B2(n10339), .ZN(
        P1_U3526) );
  AOI22_X1 U11389 ( .A1(n10341), .A2(n10335), .B1(n5866), .B2(n10339), .ZN(
        P1_U3528) );
  AOI22_X1 U11390 ( .A1(n10341), .A2(n10336), .B1(n6644), .B2(n10339), .ZN(
        P1_U3529) );
  AOI22_X1 U11391 ( .A1(n10341), .A2(n10337), .B1(n5910), .B2(n10339), .ZN(
        P1_U3530) );
  AOI22_X1 U11392 ( .A1(n10341), .A2(n10338), .B1(n5930), .B2(n10339), .ZN(
        P1_U3531) );
  AOI22_X1 U11393 ( .A1(n10341), .A2(n10340), .B1(n5953), .B2(n10339), .ZN(
        P1_U3532) );
  AOI22_X1 U11394 ( .A1(n10343), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10342), .ZN(n10354) );
  OR2_X1 U11395 ( .A1(n10344), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10345) );
  OAI211_X1 U11396 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n10347), .A(n10346), .B(
        n10345), .ZN(n10348) );
  INV_X1 U11397 ( .A(n10348), .ZN(n10352) );
  AOI22_X1 U11398 ( .A1(n10350), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10351) );
  OAI221_X1 U11399 ( .B1(n10355), .B2(n10354), .C1(n10353), .C2(n10352), .A(
        n10351), .ZN(P2_U3245) );
  AOI21_X1 U11400 ( .B1(n10357), .B2(n10409), .A(n10356), .ZN(n10411) );
  OAI22_X1 U11401 ( .A1(n7188), .A2(n10360), .B1(n10359), .B2(n10358), .ZN(
        n10365) );
  AOI21_X1 U11402 ( .B1(n10363), .B2(n10362), .A(n10361), .ZN(n10364) );
  AOI211_X1 U11403 ( .C1(n10366), .C2(n10409), .A(n10365), .B(n10364), .ZN(
        n10367) );
  OAI21_X1 U11404 ( .B1(n8877), .B2(n10411), .A(n10367), .ZN(P2_U3296) );
  NOR2_X1 U11405 ( .A1(n10369), .A2(n10368), .ZN(n10383) );
  INV_X1 U11406 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n10370) );
  NOR2_X1 U11407 ( .A1(n10405), .A2(n10370), .ZN(P2_U3297) );
  INV_X1 U11408 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n10371) );
  NOR2_X1 U11409 ( .A1(n10405), .A2(n10371), .ZN(P2_U3298) );
  INV_X1 U11410 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10372) );
  NOR2_X1 U11411 ( .A1(n10405), .A2(n10372), .ZN(P2_U3299) );
  INV_X1 U11412 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10373) );
  NOR2_X1 U11413 ( .A1(n10383), .A2(n10373), .ZN(P2_U3300) );
  INV_X1 U11414 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10374) );
  NOR2_X1 U11415 ( .A1(n10383), .A2(n10374), .ZN(P2_U3301) );
  INV_X1 U11416 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10375) );
  NOR2_X1 U11417 ( .A1(n10383), .A2(n10375), .ZN(P2_U3302) );
  INV_X1 U11418 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10376) );
  NOR2_X1 U11419 ( .A1(n10383), .A2(n10376), .ZN(P2_U3303) );
  INV_X1 U11420 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10377) );
  NOR2_X1 U11421 ( .A1(n10383), .A2(n10377), .ZN(P2_U3304) );
  INV_X1 U11422 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10378) );
  NOR2_X1 U11423 ( .A1(n10383), .A2(n10378), .ZN(P2_U3305) );
  INV_X1 U11424 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10379) );
  NOR2_X1 U11425 ( .A1(n10383), .A2(n10379), .ZN(P2_U3306) );
  INV_X1 U11426 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10380) );
  NOR2_X1 U11427 ( .A1(n10383), .A2(n10380), .ZN(P2_U3307) );
  INV_X1 U11428 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10381) );
  NOR2_X1 U11429 ( .A1(n10383), .A2(n10381), .ZN(P2_U3308) );
  INV_X1 U11430 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n10382) );
  NOR2_X1 U11431 ( .A1(n10383), .A2(n10382), .ZN(P2_U3309) );
  INV_X1 U11432 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10384) );
  NOR2_X1 U11433 ( .A1(n10405), .A2(n10384), .ZN(P2_U3310) );
  INV_X1 U11434 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10385) );
  NOR2_X1 U11435 ( .A1(n10405), .A2(n10385), .ZN(P2_U3311) );
  INV_X1 U11436 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10386) );
  NOR2_X1 U11437 ( .A1(n10405), .A2(n10386), .ZN(P2_U3312) );
  INV_X1 U11438 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10387) );
  NOR2_X1 U11439 ( .A1(n10405), .A2(n10387), .ZN(P2_U3313) );
  INV_X1 U11440 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10388) );
  NOR2_X1 U11441 ( .A1(n10405), .A2(n10388), .ZN(P2_U3314) );
  INV_X1 U11442 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10389) );
  NOR2_X1 U11443 ( .A1(n10405), .A2(n10389), .ZN(P2_U3315) );
  INV_X1 U11444 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10390) );
  NOR2_X1 U11445 ( .A1(n10405), .A2(n10390), .ZN(P2_U3316) );
  INV_X1 U11446 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10391) );
  NOR2_X1 U11447 ( .A1(n10405), .A2(n10391), .ZN(P2_U3317) );
  INV_X1 U11448 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10392) );
  NOR2_X1 U11449 ( .A1(n10405), .A2(n10392), .ZN(P2_U3318) );
  INV_X1 U11450 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10393) );
  NOR2_X1 U11451 ( .A1(n10405), .A2(n10393), .ZN(P2_U3319) );
  INV_X1 U11452 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10394) );
  NOR2_X1 U11453 ( .A1(n10405), .A2(n10394), .ZN(P2_U3320) );
  INV_X1 U11454 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10395) );
  NOR2_X1 U11455 ( .A1(n10405), .A2(n10395), .ZN(P2_U3321) );
  INV_X1 U11456 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10396) );
  NOR2_X1 U11457 ( .A1(n10405), .A2(n10396), .ZN(P2_U3322) );
  NOR2_X1 U11458 ( .A1(n10405), .A2(n10397), .ZN(P2_U3323) );
  NOR2_X1 U11459 ( .A1(n10405), .A2(n10398), .ZN(P2_U3324) );
  NOR2_X1 U11460 ( .A1(n10405), .A2(n10399), .ZN(P2_U3325) );
  NOR2_X1 U11461 ( .A1(n10405), .A2(n10400), .ZN(P2_U3326) );
  OAI22_X1 U11462 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n10405), .B1(n10404), .B2(
        n10401), .ZN(n10402) );
  INV_X1 U11463 ( .A(n10402), .ZN(P2_U3437) );
  OAI22_X1 U11464 ( .A1(P2_D_REG_1__SCAN_IN), .A2(n10405), .B1(n10404), .B2(
        n10403), .ZN(n10406) );
  INV_X1 U11465 ( .A(n10406), .ZN(P2_U3438) );
  AOI22_X1 U11466 ( .A1(n10409), .A2(n10440), .B1(n10408), .B2(n10407), .ZN(
        n10410) );
  AND2_X1 U11467 ( .A1(n10411), .A2(n10410), .ZN(n10445) );
  AOI22_X1 U11468 ( .A1(n10444), .A2(n10445), .B1(n5202), .B2(n10442), .ZN(
        P2_U3451) );
  OAI21_X1 U11469 ( .B1(n10413), .B2(n10434), .A(n10412), .ZN(n10414) );
  AOI21_X1 U11470 ( .B1(n10415), .B2(n10440), .A(n10414), .ZN(n10417) );
  AND2_X1 U11471 ( .A1(n10417), .A2(n10416), .ZN(n10446) );
  AOI22_X1 U11472 ( .A1(n10444), .A2(n10446), .B1(n5192), .B2(n10442), .ZN(
        P2_U3454) );
  OAI21_X1 U11473 ( .B1(n10419), .B2(n10434), .A(n10418), .ZN(n10421) );
  AOI211_X1 U11474 ( .C1(n10423), .C2(n10422), .A(n10421), .B(n10420), .ZN(
        n10447) );
  AOI22_X1 U11475 ( .A1(n10444), .A2(n10447), .B1(n5228), .B2(n10442), .ZN(
        P2_U3460) );
  OAI211_X1 U11476 ( .C1(n10426), .C2(n10434), .A(n10425), .B(n10424), .ZN(
        n10427) );
  AOI21_X1 U11477 ( .B1(n10440), .B2(n10428), .A(n10427), .ZN(n10448) );
  AOI22_X1 U11478 ( .A1(n10444), .A2(n10448), .B1(n5274), .B2(n10442), .ZN(
        P2_U3472) );
  OAI22_X1 U11479 ( .A1(n10430), .A2(n10436), .B1(n10429), .B2(n10434), .ZN(
        n10432) );
  AOI211_X1 U11480 ( .C1(n10440), .C2(n10433), .A(n10432), .B(n10431), .ZN(
        n10449) );
  AOI22_X1 U11481 ( .A1(n10444), .A2(n10449), .B1(n5312), .B2(n10442), .ZN(
        P2_U3478) );
  OAI22_X1 U11482 ( .A1(n10437), .A2(n10436), .B1(n10435), .B2(n10434), .ZN(
        n10439) );
  AOI211_X1 U11483 ( .C1(n10441), .C2(n10440), .A(n10439), .B(n10438), .ZN(
        n10451) );
  INV_X1 U11484 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U11485 ( .A1(n10444), .A2(n10451), .B1(n10443), .B2(n10442), .ZN(
        P2_U3484) );
  AOI22_X1 U11486 ( .A1(n10452), .A2(n10445), .B1(n5203), .B2(n10450), .ZN(
        P2_U3520) );
  AOI22_X1 U11487 ( .A1(n10452), .A2(n10446), .B1(n6800), .B2(n10450), .ZN(
        P2_U3521) );
  AOI22_X1 U11488 ( .A1(n10452), .A2(n10447), .B1(n6798), .B2(n10450), .ZN(
        P2_U3523) );
  AOI22_X1 U11489 ( .A1(n10452), .A2(n10448), .B1(n6857), .B2(n10450), .ZN(
        P2_U3527) );
  AOI22_X1 U11490 ( .A1(n10452), .A2(n10449), .B1(n7029), .B2(n10450), .ZN(
        P2_U3529) );
  AOI22_X1 U11491 ( .A1(n10452), .A2(n10451), .B1(n7097), .B2(n10450), .ZN(
        P2_U3531) );
  INV_X1 U11492 ( .A(n10453), .ZN(n10454) );
  NAND2_X1 U11493 ( .A1(n10455), .A2(n10454), .ZN(n10456) );
  XNOR2_X1 U11494 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10456), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11495 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11496 ( .B1(n10459), .B2(n10458), .A(n10457), .ZN(ADD_1071_U56) );
  OAI21_X1 U11497 ( .B1(n10462), .B2(n10461), .A(n10460), .ZN(ADD_1071_U57) );
  OAI21_X1 U11498 ( .B1(n10465), .B2(n10464), .A(n10463), .ZN(ADD_1071_U58) );
  OAI21_X1 U11499 ( .B1(n10468), .B2(n10467), .A(n10466), .ZN(ADD_1071_U59) );
  OAI21_X1 U11500 ( .B1(n10471), .B2(n10470), .A(n10469), .ZN(ADD_1071_U60) );
  OAI21_X1 U11501 ( .B1(n10474), .B2(n10473), .A(n10472), .ZN(ADD_1071_U61) );
  AOI21_X1 U11502 ( .B1(n10477), .B2(n10476), .A(n10475), .ZN(ADD_1071_U62) );
  AOI21_X1 U11503 ( .B1(n10480), .B2(n10479), .A(n10478), .ZN(ADD_1071_U63) );
  AOI21_X1 U11504 ( .B1(n10483), .B2(n10482), .A(n10481), .ZN(ADD_1071_U47) );
  XOR2_X1 U11505 ( .A(n10484), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11506 ( .A(n10486), .B(n10485), .Z(ADD_1071_U54) );
  NOR2_X1 U11507 ( .A1(n10488), .A2(n10487), .ZN(n10489) );
  XOR2_X1 U11508 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10489), .Z(ADD_1071_U51) );
  OAI21_X1 U11509 ( .B1(n10492), .B2(n10491), .A(n10490), .ZN(n10493) );
  XNOR2_X1 U11510 ( .A(n10493), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11511 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10494), .Z(ADD_1071_U48) );
  XOR2_X1 U11512 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10495), .Z(ADD_1071_U50) );
  XOR2_X1 U11513 ( .A(n10497), .B(n10496), .Z(ADD_1071_U53) );
  XNOR2_X1 U11514 ( .A(n10499), .B(n10498), .ZN(ADD_1071_U52) );
  INV_X2 U5026 ( .A(n6513), .ZN(n6488) );
  CLKBUF_X2 U5137 ( .A(n5888), .Z(n4485) );
endmodule

