

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, 
        HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3628, n3629, n3630, n3631, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659;

  NAND2_X1 U3662 ( .A1(n5005), .A2(n4891), .ZN(n5350) );
  CLKBUF_X2 U3663 ( .A(n3778), .Z(n3634) );
  CLKBUF_X2 U3664 ( .A(n3886), .Z(n4682) );
  CLKBUF_X2 U3665 ( .A(n3937), .Z(n5133) );
  CLKBUF_X2 U3666 ( .A(n3907), .Z(n3637) );
  CLKBUF_X2 U3667 ( .A(n3777), .Z(n4635) );
  AND2_X2 U3668 ( .A1(n4974), .A2(n5128), .ZN(n3850) );
  CLKBUF_X2 U3669 ( .A(n3980), .Z(n3938) );
  INV_X1 U3671 ( .A(n4189), .ZN(n5054) );
  CLKBUF_X1 U3674 ( .A(n7523), .Z(n3628) );
  AOI21_X1 U3675 ( .B1(n7529), .B2(STATE_REG_0__SCAN_IN), .A(n7174), .ZN(n7523) );
  AND2_X2 U3676 ( .A1(n5138), .A2(n5131), .ZN(n3902) );
  INV_X1 U3677 ( .A(n4827), .ZN(n4858) );
  NAND4_X1 U3678 ( .A1(n3712), .A2(n3711), .A3(n3710), .A4(n3709), .ZN(n3802)
         );
  INV_X1 U3679 ( .A(n4647), .ZN(n4701) );
  NOR2_X2 U3680 ( .A1(n6500), .A2(n6115), .ZN(n6114) );
  AND2_X1 U3681 ( .A1(n4113), .A2(n6681), .ZN(n3643) );
  INV_X1 U3682 ( .A(n7324), .ZN(n7372) );
  INV_X1 U3683 ( .A(n7422), .ZN(n7442) );
  NAND2_X1 U3684 ( .A1(n3641), .A2(n6511), .ZN(n6500) );
  NAND2_X1 U3685 ( .A1(n6644), .A2(n6761), .ZN(n6586) );
  INV_X1 U3687 ( .A(n7211), .ZN(n7276) );
  INV_X2 U3688 ( .A(n7425), .ZN(n7445) );
  AND2_X2 U3689 ( .A1(n5132), .A2(n4974), .ZN(n4673) );
  AND2_X1 U3691 ( .A1(n5128), .A2(n5163), .ZN(n3629) );
  AND2_X1 U3692 ( .A1(n5128), .A2(n5163), .ZN(n3630) );
  AND2_X1 U3693 ( .A1(n4978), .A2(n3676), .ZN(n3631) );
  INV_X1 U3694 ( .A(n4188), .ZN(n5169) );
  BUF_X2 U3695 ( .A(n6724), .Z(n6741) );
  AOI21_X2 U3696 ( .B1(n5271), .B2(n4127), .A(n3918), .ZN(n7128) );
  NOR2_X4 U3697 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5138) );
  NOR2_X1 U3698 ( .A1(n6540), .A2(n6542), .ZN(n6526) );
  CLKBUF_X1 U3699 ( .A(n6540), .Z(n6541) );
  CLKBUF_X1 U3700 ( .A(n6559), .Z(n6573) );
  INV_X2 U3701 ( .A(n6751), .ZN(n6769) );
  OAI211_X1 U3702 ( .C1(n4647), .C2(n4246), .A(n4245), .B(n4244), .ZN(n5038)
         );
  OR2_X1 U3703 ( .A1(n4890), .A2(n5144), .ZN(n5005) );
  NAND2_X1 U3704 ( .A1(n4734), .A2(n7499), .ZN(n4890) );
  XNOR2_X1 U3705 ( .A(n5155), .B(n5153), .ZN(n5096) );
  INV_X1 U3706 ( .A(n4167), .ZN(n4145) );
  INV_X2 U3707 ( .A(n3655), .ZN(n3633) );
  BUF_X1 U3708 ( .A(n3802), .Z(n4174) );
  BUF_X2 U3709 ( .A(n4673), .Z(n4553) );
  NAND2_X1 U3710 ( .A1(n3645), .A2(n4107), .ZN(n6718) );
  CLKBUF_X1 U3711 ( .A(n6526), .Z(n6527) );
  OAI211_X1 U3712 ( .C1(n6118), .C2(n6030), .A(n6029), .B(n6028), .ZN(n6031)
         );
  XNOR2_X1 U3713 ( .A(n4866), .B(n6030), .ZN(n6113) );
  CLKBUF_X1 U3714 ( .A(n6027), .Z(n6498) );
  AND2_X1 U3715 ( .A1(n5022), .A2(n5038), .ZN(n4247) );
  AOI21_X1 U3716 ( .B1(n5169), .B2(n4346), .A(n4196), .ZN(n5030) );
  OAI21_X1 U3717 ( .B1(n4218), .B2(n4726), .A(n4013), .ZN(n4014) );
  INV_X1 U3718 ( .A(n3961), .ZN(n7129) );
  OR2_X2 U3719 ( .A1(n4172), .A2(n4171), .ZN(n6097) );
  BUF_X1 U3720 ( .A(n4202), .Z(n7454) );
  CLKBUF_X1 U3721 ( .A(n3876), .Z(n3969) );
  NAND2_X1 U3722 ( .A1(n4725), .A2(n4743), .ZN(n6100) );
  NAND2_X1 U3723 ( .A1(n3656), .A2(n4764), .ZN(n6023) );
  INV_X2 U3724 ( .A(n3926), .ZN(n3837) );
  CLKBUF_X1 U3725 ( .A(n4173), .Z(n4877) );
  AND2_X4 U3726 ( .A1(n3926), .A2(n3653), .ZN(n4781) );
  AND2_X2 U3727 ( .A1(n5054), .A2(n4192), .ZN(n4868) );
  AND2_X1 U3728 ( .A1(n3735), .A2(n3734), .ZN(n3799) );
  BUF_X1 U3729 ( .A(n5251), .Z(n3650) );
  AND2_X2 U3730 ( .A1(n3635), .A2(n4743), .ZN(n3915) );
  INV_X2 U3731 ( .A(n3798), .ZN(n5225) );
  CLKBUF_X2 U3732 ( .A(n4636), .Z(n4681) );
  AND4_X1 U3733 ( .A1(n3761), .A2(n3760), .A3(n3759), .A4(n3758), .ZN(n3767)
         );
  BUF_X2 U3734 ( .A(n3783), .Z(n4675) );
  BUF_X2 U3735 ( .A(n4519), .Z(n4674) );
  CLKBUF_X2 U3736 ( .A(n3902), .Z(n4683) );
  NOR2_X4 U3737 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5163) );
  AND2_X1 U3738 ( .A1(n4116), .A2(n3666), .ZN(n4117) );
  OAI21_X1 U3739 ( .B1(n6769), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n6708), 
        .ZN(n6698) );
  OR2_X1 U3740 ( .A1(n6708), .A2(n6050), .ZN(n4116) );
  OR2_X1 U3741 ( .A1(n6742), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6731)
         );
  AND2_X1 U3742 ( .A1(n4112), .A2(n6689), .ZN(n6681) );
  NAND2_X1 U3743 ( .A1(n6718), .A2(n4108), .ZN(n4110) );
  CLKBUF_X1 U3744 ( .A(n6741), .Z(n6779) );
  AND2_X2 U3745 ( .A1(n6643), .A2(n6642), .ZN(n6644) );
  NOR2_X1 U3746 ( .A1(n6027), .A2(n6116), .ZN(n6026) );
  CLKBUF_X1 U3747 ( .A(n6522), .Z(n6555) );
  AND2_X1 U3748 ( .A1(n6865), .A2(n4904), .ZN(n6847) );
  INV_X1 U3749 ( .A(n6906), .ZN(n6864) );
  NOR2_X2 U3750 ( .A1(n6896), .A2(n6646), .ZN(n6877) );
  CLKBUF_X1 U3751 ( .A(n5021), .Z(n5077) );
  INV_X1 U3752 ( .A(n4079), .ZN(n4082) );
  AOI21_X1 U3753 ( .B1(n4252), .B2(n4346), .A(n4251), .ZN(n5087) );
  NAND2_X1 U3754 ( .A1(n4217), .A2(n5032), .ZN(n5031) );
  OAI21_X1 U3755 ( .B1(n5067), .B2(n5072), .A(n5068), .ZN(n3997) );
  NAND2_X1 U3756 ( .A1(n4068), .A2(n4127), .ZN(n4079) );
  INV_X1 U3757 ( .A(n5030), .ZN(n4217) );
  AND2_X1 U3758 ( .A1(n4227), .A2(n4226), .ZN(n5078) );
  CLKBUF_X1 U3759 ( .A(n4197), .Z(n5381) );
  BUF_X1 U3760 ( .A(n3990), .Z(n5100) );
  NAND2_X1 U3761 ( .A1(n4800), .A2(n4799), .ZN(n5859) );
  NOR2_X1 U3762 ( .A1(n4604), .A2(n6531), .ZN(n4625) );
  CLKBUF_X1 U3763 ( .A(n5102), .Z(n6066) );
  OR2_X1 U3764 ( .A1(n4890), .A2(n6095), .ZN(n7233) );
  INV_X1 U3765 ( .A(n5516), .ZN(n4800) );
  INV_X2 U3766 ( .A(n4926), .ZN(n5176) );
  NOR2_X2 U3767 ( .A1(n5123), .A2(n5264), .ZN(n5518) );
  CLKBUF_X1 U3768 ( .A(n5103), .Z(n5415) );
  NAND2_X1 U3769 ( .A1(n4788), .A2(n4787), .ZN(n5123) );
  INV_X1 U3770 ( .A(n5092), .ZN(n4788) );
  OR2_X1 U3771 ( .A1(n4496), .A2(n4495), .ZN(n4516) );
  CLKBUF_X1 U3772 ( .A(n3873), .Z(n3874) );
  NAND2_X1 U3773 ( .A1(n3864), .A2(n3862), .ZN(n3871) );
  NAND2_X1 U3774 ( .A1(n3832), .A2(n3831), .ZN(n3864) );
  AOI21_X1 U3775 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n3848), .A(n4161), 
        .ZN(n4170) );
  NOR2_X1 U3776 ( .A1(n4461), .A2(n6780), .ZN(n4478) );
  AND2_X1 U3777 ( .A1(n3836), .A2(n3835), .ZN(n4874) );
  NOR2_X1 U3778 ( .A1(n3846), .A2(n3845), .ZN(n3847) );
  AND3_X2 U3779 ( .A1(n3819), .A2(n3818), .A3(n4876), .ZN(n4729) );
  BUF_X4 U3780 ( .A(n4781), .Z(n3655) );
  INV_X1 U3781 ( .A(n4158), .ZN(n4168) );
  NAND2_X1 U3782 ( .A1(n3947), .A2(n3881), .ZN(n4167) );
  AND2_X1 U3783 ( .A1(n3837), .A2(n5251), .ZN(n4876) );
  INV_X1 U3784 ( .A(n3799), .ZN(n4867) );
  AND2_X1 U3785 ( .A1(n3799), .A2(n3738), .ZN(n4912) );
  OR2_X1 U3786 ( .A1(n3944), .A2(n3943), .ZN(n4084) );
  AND2_X1 U3787 ( .A1(n5225), .A2(n4174), .ZN(n4176) );
  AND2_X2 U3788 ( .A1(n4132), .A2(n3798), .ZN(n4157) );
  INV_X1 U3789 ( .A(n3653), .ZN(n3820) );
  AND3_X1 U3790 ( .A1(n3744), .A2(n3743), .A3(n3667), .ZN(n3660) );
  NOR2_X1 U3791 ( .A1(n4265), .A2(n5838), .ZN(n4319) );
  INV_X1 U3792 ( .A(n3653), .ZN(n3635) );
  AND4_X1 U3793 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), .ZN(n3769)
         );
  AND4_X1 U3794 ( .A1(n3717), .A2(n3716), .A3(n3715), .A4(n3714), .ZN(n3723)
         );
  AND4_X1 U3795 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3768)
         );
  AND4_X1 U3796 ( .A1(n3721), .A2(n3720), .A3(n3719), .A4(n3718), .ZN(n3722)
         );
  AND4_X1 U3797 ( .A1(n3782), .A2(n3781), .A3(n3780), .A4(n3779), .ZN(n3795)
         );
  AND4_X1 U3798 ( .A1(n3708), .A2(n3707), .A3(n3706), .A4(n3705), .ZN(n3709)
         );
  AND4_X1 U3799 ( .A1(n3776), .A2(n3775), .A3(n3774), .A4(n3773), .ZN(n3796)
         );
  AND4_X1 U3800 ( .A1(n3704), .A2(n3703), .A3(n3702), .A4(n3701), .ZN(n3710)
         );
  AND4_X1 U3801 ( .A1(n3765), .A2(n3764), .A3(n3763), .A4(n3762), .ZN(n3766)
         );
  AND4_X1 U3802 ( .A1(n3700), .A2(n3699), .A3(n3698), .A4(n3697), .ZN(n3711)
         );
  AND4_X1 U3803 ( .A1(n3696), .A2(n3695), .A3(n3694), .A4(n3693), .ZN(n3712)
         );
  AND4_X1 U3804 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(n3793)
         );
  AND4_X1 U3805 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(n3794)
         );
  BUF_X2 U3806 ( .A(n4433), .Z(n4636) );
  NAND2_X2 U3807 ( .A1(n7174), .A2(n7533), .ZN(n7071) );
  BUF_X2 U3808 ( .A(n3931), .Z(n4676) );
  BUF_X2 U3809 ( .A(n3788), .Z(n3636) );
  AND2_X2 U3810 ( .A1(n3670), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4978)
         );
  NOR3_X1 U3811 ( .A1(n6619), .A2(n4182), .A3(n6607), .ZN(n4221) );
  BUF_X2 U3812 ( .A(n3887), .Z(n3638) );
  AND2_X2 U3813 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5131) );
  INV_X1 U3814 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3670) );
  CLKBUF_X1 U3815 ( .A(n5067), .Z(n3639) );
  CLKBUF_X1 U3816 ( .A(n7136), .Z(n3640) );
  XNOR2_X1 U3817 ( .A(n4014), .B(n4765), .ZN(n7136) );
  NAND2_X1 U3818 ( .A1(n3965), .A2(n3964), .ZN(n5067) );
  AND2_X1 U3819 ( .A1(n6501), .A2(n4630), .ZN(n3641) );
  NOR2_X1 U3820 ( .A1(n6528), .A2(n6512), .ZN(n6499) );
  AND2_X1 U3821 ( .A1(n6526), .A2(n4607), .ZN(n6511) );
  AND2_X2 U3822 ( .A1(n3922), .A2(n3869), .ZN(n3896) );
  AND2_X2 U3823 ( .A1(n5128), .A2(n5131), .ZN(n3887) );
  NAND2_X1 U3824 ( .A1(n4037), .A2(n3991), .ZN(n4188) );
  AOI211_X1 U3825 ( .C1(n5169), .C2(n7520), .A(n5440), .B(n5171), .ZN(n5172)
         );
  NAND2_X1 U3826 ( .A1(n7137), .A2(n3640), .ZN(n3642) );
  INV_X1 U3827 ( .A(n4106), .ZN(n3644) );
  NOR2_X1 U3828 ( .A1(n6719), .A2(n3644), .ZN(n3645) );
  INV_X1 U3829 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3646) );
  CLKBUF_X1 U3830 ( .A(n5851), .Z(n3647) );
  INV_X1 U3831 ( .A(n3849), .ZN(n3648) );
  OR2_X1 U3832 ( .A1(n6727), .A2(n6751), .ZN(n3649) );
  NAND2_X1 U3833 ( .A1(n3649), .A2(n6874), .ZN(n6753) );
  AND2_X4 U3834 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5128) );
  AND2_X2 U3835 ( .A1(n5132), .A2(n5163), .ZN(n3777) );
  AND2_X2 U3836 ( .A1(n6061), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5132)
         );
  OAI211_X1 U3837 ( .C1(n3816), .C2(n3817), .A(n3838), .B(n3739), .ZN(n3771)
         );
  NAND2_X1 U3838 ( .A1(n3849), .A2(n3848), .ZN(n3919) );
  NAND4_X1 U3839 ( .A1(n3769), .A2(n3768), .A3(n3767), .A4(n3766), .ZN(n3654)
         );
  NAND2_X1 U3840 ( .A1(n4189), .A2(n3802), .ZN(n5063) );
  NAND4_X4 U3841 ( .A1(n3769), .A2(n3768), .A3(n3767), .A4(n3766), .ZN(n3653)
         );
  AND2_X1 U3842 ( .A1(n3926), .A2(n3653), .ZN(n3651) );
  AND2_X2 U3843 ( .A1(n5132), .A2(n5131), .ZN(n3778) );
  OR2_X1 U3844 ( .A1(n4010), .A2(n4039), .ZN(n4011) );
  AND2_X2 U3845 ( .A1(n3997), .A2(n3996), .ZN(n7137) );
  OR2_X2 U3846 ( .A1(n6898), .A2(n6899), .ZN(n6896) );
  AND2_X1 U3847 ( .A1(n4974), .A2(n5128), .ZN(n3652) );
  AND2_X1 U3848 ( .A1(n4974), .A2(n5128), .ZN(n3657) );
  NAND2_X4 U3849 ( .A1(n3660), .A2(n3749), .ZN(n3926) );
  AND4_X2 U3850 ( .A1(n3748), .A2(n3747), .A3(n3746), .A4(n3745), .ZN(n3749)
         );
  AOI21_X2 U3851 ( .B1(n5096), .B2(n3848), .A(n3988), .ZN(n3990) );
  INV_X1 U3852 ( .A(n4781), .ZN(n3656) );
  AND2_X1 U3853 ( .A1(n4743), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4132) );
  NAND2_X1 U3854 ( .A1(n5025), .A2(n5027), .ZN(n5026) );
  AND2_X1 U3855 ( .A1(n4977), .A2(n4875), .ZN(n5137) );
  INV_X1 U3856 ( .A(n3802), .ZN(n3738) );
  CLKBUF_X1 U3857 ( .A(n4192), .Z(n4193) );
  AOI21_X1 U3858 ( .B1(n4170), .B2(n4169), .A(n4168), .ZN(n4172) );
  NOR2_X1 U3859 ( .A1(n4170), .A2(n4717), .ZN(n4171) );
  INV_X1 U3860 ( .A(n4037), .ZN(n4040) );
  AND2_X1 U3861 ( .A1(n4052), .A2(n4051), .ZN(n4055) );
  AND2_X2 U3862 ( .A1(n3671), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3676)
         );
  AND2_X2 U3863 ( .A1(n4978), .A2(n5138), .ZN(n3783) );
  INV_X1 U3864 ( .A(n3987), .ZN(n3988) );
  NAND2_X1 U3865 ( .A1(n4874), .A2(n3847), .ZN(n3862) );
  NOR2_X1 U3866 ( .A1(n4743), .A2(n3654), .ZN(n5735) );
  NAND2_X1 U3867 ( .A1(n6559), .A2(n6560), .ZN(n6540) );
  INV_X1 U3868 ( .A(n5814), .ZN(n4390) );
  NOR2_X2 U3869 ( .A1(n7123), .A2(n4770), .ZN(n5025) );
  NOR2_X1 U3870 ( .A1(n4781), .A2(n4753), .ZN(n4854) );
  OR2_X1 U3871 ( .A1(n3827), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3828)
         );
  INV_X1 U3872 ( .A(n4725), .ZN(n4990) );
  AOI22_X1 U3873 ( .A1(n3652), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3777), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U3874 ( .A1(n4433), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3778), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U3875 ( .A1(n4519), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3886), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3674) );
  OR2_X1 U3876 ( .A1(n7190), .A2(n5712), .ZN(n7301) );
  NOR2_X1 U3877 ( .A1(n6097), .A2(n4921), .ZN(n5708) );
  OR2_X1 U3878 ( .A1(n6100), .A2(n7517), .ZN(n4921) );
  NAND2_X1 U3879 ( .A1(n4625), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4649)
         );
  OR2_X1 U3880 ( .A1(n6716), .A2(n4220), .ZN(n4585) );
  OAI21_X1 U3881 ( .B1(n4197), .B2(n4388), .A(n4403), .ZN(n4961) );
  NAND2_X1 U3882 ( .A1(n4113), .A2(n6681), .ZN(n4708) );
  NAND2_X1 U3883 ( .A1(n6698), .A2(n6835), .ZN(n6697) );
  NOR2_X2 U3884 ( .A1(n7112), .A2(n7111), .ZN(n7114) );
  AND2_X1 U3885 ( .A1(n6751), .A2(n7268), .ZN(n6003) );
  NOR2_X1 U3886 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5112), .ZN(n5413) );
  INV_X1 U3887 ( .A(n5413), .ZN(n5303) );
  INV_X1 U3888 ( .A(n4174), .ZN(n5901) );
  NAND2_X1 U3889 ( .A1(n7301), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U3890 ( .A1(n7126), .A2(n6086), .ZN(n6647) );
  AND2_X1 U3891 ( .A1(n4915), .A2(n7499), .ZN(n7126) );
  AND2_X1 U3892 ( .A1(n7491), .A2(n7490), .ZN(n7518) );
  OR2_X1 U3893 ( .A1(n3653), .A2(n4712), .ZN(n3815) );
  NAND2_X1 U3894 ( .A1(n3797), .A2(n3650), .ZN(n3833) );
  AND2_X1 U3895 ( .A1(n3841), .A2(n3635), .ZN(n3770) );
  INV_X1 U3896 ( .A(n4056), .ZN(n4054) );
  OR2_X1 U3897 ( .A1(n4025), .A2(n4024), .ZN(n4058) );
  OR2_X1 U3898 ( .A1(n4007), .A2(n4006), .ZN(n4029) );
  AOI22_X1 U3899 ( .A1(n3657), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3777), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3730) );
  NAND2_X1 U3900 ( .A1(n4673), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U3901 ( .A1(n3937), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3717) );
  NOR2_X1 U3902 ( .A1(n4392), .A2(n6018), .ZN(n4421) );
  AND2_X1 U3903 ( .A1(n4240), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4229)
         );
  XNOR2_X1 U3904 ( .A(n4028), .B(n4038), .ZN(n4239) );
  NOR2_X1 U3905 ( .A1(n6751), .A2(n4101), .ZN(n4103) );
  NAND2_X1 U3906 ( .A1(n5518), .A2(n5517), .ZN(n5516) );
  OR2_X1 U3907 ( .A1(n4050), .A2(n4049), .ZN(n4070) );
  NAND2_X1 U3908 ( .A1(n3866), .A2(n3661), .ZN(n3867) );
  NAND2_X1 U3909 ( .A1(n3650), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3881) );
  NOR2_X1 U3910 ( .A1(n4157), .A2(n4718), .ZN(n4159) );
  AND2_X1 U3911 ( .A1(n4874), .A2(n4873), .ZN(n4977) );
  NAND2_X1 U3912 ( .A1(n3875), .A2(n3874), .ZN(n3966) );
  NAND2_X1 U3913 ( .A1(n4444), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4461)
         );
  INV_X1 U3914 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6607) );
  NAND2_X1 U3915 ( .A1(n7114), .A2(n5990), .ZN(n6898) );
  AND2_X1 U3916 ( .A1(n4809), .A2(n4808), .ZN(n5723) );
  NAND2_X1 U3917 ( .A1(n5515), .A2(n4355), .ZN(n4356) );
  INV_X1 U3918 ( .A(n7024), .ZN(n4942) );
  INV_X1 U3919 ( .A(n5061), .ZN(n5052) );
  AND2_X1 U3920 ( .A1(n7188), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4700) );
  OR2_X1 U3921 ( .A1(n4629), .A2(n4628), .ZN(n6512) );
  INV_X1 U3922 ( .A(n6529), .ZN(n4607) );
  NAND2_X1 U3923 ( .A1(n4184), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4583)
         );
  INV_X1 U3924 ( .A(n6527), .ZN(n6543) );
  NAND2_X1 U3925 ( .A1(n4183), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4547)
         );
  OR2_X1 U3926 ( .A1(n4547), .A2(n4546), .ZN(n4552) );
  CLKBUF_X1 U3927 ( .A(n6571), .Z(n6572) );
  CLKBUF_X1 U3928 ( .A(n5986), .Z(n5987) );
  AND2_X1 U3929 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n4421), .ZN(n4444)
         );
  CLKBUF_X1 U3930 ( .A(n5983), .Z(n5984) );
  NAND2_X1 U3931 ( .A1(n4374), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4392)
         );
  CLKBUF_X1 U3932 ( .A(n5875), .Z(n5876) );
  AND2_X1 U3933 ( .A1(n4368), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4374)
         );
  CLKBUF_X1 U3934 ( .A(n5812), .Z(n5813) );
  CLKBUF_X1 U3935 ( .A(n5754), .Z(n5755) );
  NOR2_X1 U3936 ( .A1(n4347), .A2(n5729), .ZN(n4368) );
  NAND2_X1 U3937 ( .A1(n4271), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4347)
         );
  NOR2_X1 U3938 ( .A1(n4301), .A2(n5821), .ZN(n4286) );
  NAND2_X1 U3939 ( .A1(n4319), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4301)
         );
  INV_X1 U3940 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U3941 ( .A1(n4248), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4265)
         );
  AND2_X1 U3942 ( .A1(n4229), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4248)
         );
  NAND2_X1 U3943 ( .A1(n4238), .A2(n4237), .ZN(n5022) );
  AND2_X1 U3944 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n4221), .ZN(n4240)
         );
  OR2_X1 U3945 ( .A1(n6522), .A2(n6523), .ZN(n6525) );
  NOR2_X2 U3946 ( .A1(n6525), .A2(n6519), .ZN(n6518) );
  AND2_X1 U3947 ( .A1(n6577), .A2(n6561), .ZN(n6552) );
  NOR2_X2 U3948 ( .A1(n6593), .A2(n6575), .ZN(n6577) );
  AOI21_X1 U3949 ( .B1(n6751), .B2(n6726), .A(n6725), .ZN(n6763) );
  CLKBUF_X1 U3950 ( .A(n6786), .Z(n6787) );
  NAND2_X1 U3951 ( .A1(n4817), .A2(n4816), .ZN(n5881) );
  INV_X1 U3952 ( .A(n5817), .ZN(n4817) );
  AND2_X1 U3953 ( .A1(n5767), .A2(n5723), .ZN(n5758) );
  NOR2_X2 U3954 ( .A1(n5859), .A2(n5765), .ZN(n5767) );
  NAND2_X1 U3955 ( .A1(n4779), .A2(n4778), .ZN(n5092) );
  INV_X1 U3956 ( .A(n5026), .ZN(n4779) );
  NAND2_X1 U3957 ( .A1(n4967), .A2(n4966), .ZN(n4965) );
  NAND2_X1 U3958 ( .A1(n3821), .A2(n4868), .ZN(n4739) );
  NOR2_X1 U3959 ( .A1(n3838), .A2(n5901), .ZN(n7452) );
  CLKBUF_X1 U3960 ( .A(n5098), .Z(n5099) );
  NAND2_X1 U3961 ( .A1(n3968), .A2(n3967), .ZN(n5155) );
  INV_X1 U3962 ( .A(n3966), .ZN(n3968) );
  NAND2_X1 U3963 ( .A1(n3975), .A2(n3974), .ZN(n5153) );
  INV_X1 U3964 ( .A(n3817), .ZN(n3818) );
  AND3_X1 U3965 ( .A1(n4995), .A2(n4994), .A3(n4993), .ZN(n7472) );
  CLKBUF_X1 U3966 ( .A(n5096), .Z(n5097) );
  AND2_X1 U3967 ( .A1(n5440), .A2(n5663), .ZN(n7581) );
  INV_X1 U3968 ( .A(n5114), .ZN(n5629) );
  INV_X1 U3969 ( .A(n6935), .ZN(n5419) );
  INV_X1 U3970 ( .A(n4743), .ZN(n5251) );
  BUF_X1 U3971 ( .A(n3799), .Z(n5230) );
  AOI22_X1 U3972 ( .A1(n3907), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3887), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3679) );
  OR3_X1 U3973 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5112), .A3(n7508), .ZN(n5252) );
  AOI21_X1 U3974 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7576), .A(n5303), .ZN(
        n7587) );
  NAND2_X1 U3975 ( .A1(n5739), .A2(n5722), .ZN(n7421) );
  AND2_X1 U3976 ( .A1(n7301), .A2(n5730), .ZN(n7411) );
  INV_X1 U3977 ( .A(n7421), .ZN(n7441) );
  INV_X1 U3978 ( .A(n6647), .ZN(n7124) );
  AND2_X1 U3979 ( .A1(n6085), .A2(n4868), .ZN(n7550) );
  AND2_X1 U3980 ( .A1(n6085), .A2(n5902), .ZN(n7554) );
  INV_X1 U3981 ( .A(n6085), .ZN(n7553) );
  NAND2_X1 U3982 ( .A1(n5062), .A2(n5061), .ZN(n6085) );
  NAND2_X1 U3983 ( .A1(n5060), .A2(n7499), .ZN(n5062) );
  OR2_X1 U3984 ( .A1(n5059), .A2(n5058), .ZN(n5060) );
  OR2_X1 U3985 ( .A1(n7553), .A2(n5064), .ZN(n5848) );
  NOR2_X1 U3987 ( .A1(n4697), .A2(n6104), .ZN(n4185) );
  AND2_X1 U3988 ( .A1(n5040), .A2(n5039), .ZN(n7306) );
  AND2_X1 U3989 ( .A1(n7447), .A2(n4179), .ZN(n7158) );
  INV_X1 U3990 ( .A(n7169), .ZN(n7154) );
  NAND2_X1 U3991 ( .A1(n7483), .A2(n7499), .ZN(n7447) );
  OAI21_X1 U3992 ( .B1(n3643), .B2(n6751), .A(n4117), .ZN(n4119) );
  OAI21_X1 U3993 ( .B1(n4710), .B2(n6751), .A(n4709), .ZN(n4711) );
  NAND2_X1 U3994 ( .A1(n6700), .A2(n6699), .ZN(n6701) );
  NAND2_X1 U3995 ( .A1(n6698), .A2(n6751), .ZN(n6699) );
  NAND2_X1 U3996 ( .A1(n6697), .A2(n6769), .ZN(n6700) );
  NAND2_X1 U3997 ( .A1(n6753), .A2(n6728), .ZN(n6732) );
  CLKBUF_X1 U3998 ( .A(n6012), .Z(n6013) );
  CLKBUF_X1 U3999 ( .A(n6000), .Z(n6001) );
  CLKBUF_X1 U4000 ( .A(n5959), .Z(n5960) );
  NAND2_X1 U4001 ( .A1(n5857), .A2(n5888), .ZN(n7197) );
  INV_X1 U4002 ( .A(n6892), .ZN(n7278) );
  INV_X1 U4003 ( .A(n5415), .ZN(n7557) );
  INV_X1 U4004 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5411) );
  INV_X1 U4005 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7480) );
  AND2_X1 U4006 ( .A1(n5168), .A2(n5303), .ZN(n6992) );
  INV_X1 U4007 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n7455) );
  NOR2_X1 U4008 ( .A1(n7508), .A2(n6097), .ZN(n6059) );
  INV_X1 U4009 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n7465) );
  NOR2_X1 U4010 ( .A1(n5282), .A2(n5415), .ZN(n5911) );
  INV_X1 U4011 ( .A(n5538), .ZN(n5597) );
  INV_X1 U4012 ( .A(n5674), .ZN(n5699) );
  AND2_X1 U4013 ( .A1(n7581), .A2(n5415), .ZN(n7652) );
  AND2_X1 U4014 ( .A1(n5440), .A2(n5439), .ZN(n7644) );
  NOR2_X1 U4015 ( .A1(n5253), .A2(n5303), .ZN(n6936) );
  NOR2_X1 U4016 ( .A1(n5246), .A2(n5303), .ZN(n6941) );
  NOR2_X1 U4017 ( .A1(n5231), .A2(n5303), .ZN(n6946) );
  NOR2_X1 U4018 ( .A1(n5241), .A2(n5303), .ZN(n6951) );
  NOR2_X1 U4019 ( .A1(n6678), .A2(n5303), .ZN(n6956) );
  NOR2_X1 U4020 ( .A1(n6675), .A2(n5303), .ZN(n6966) );
  AND2_X1 U4021 ( .A1(n5383), .A2(n5415), .ZN(n5640) );
  AND2_X1 U4022 ( .A1(n5383), .A2(n7557), .ZN(n5639) );
  NOR2_X1 U4023 ( .A1(n6672), .A2(n5303), .ZN(n6973) );
  INV_X1 U4024 ( .A(n7597), .ZN(n5680) );
  INV_X1 U4025 ( .A(n6946), .ZN(n7610) );
  INV_X1 U4026 ( .A(n7605), .ZN(n5683) );
  INV_X1 U4027 ( .A(n6951), .ZN(n7618) );
  INV_X1 U4028 ( .A(n6956), .ZN(n7626) );
  INV_X1 U4029 ( .A(n7621), .ZN(n5692) );
  INV_X1 U4030 ( .A(n6961), .ZN(n7634) );
  INV_X1 U4031 ( .A(n7629), .ZN(n5689) );
  INV_X1 U4032 ( .A(n7637), .ZN(n5686) );
  INV_X1 U4033 ( .A(n6973), .ZN(n7658) );
  INV_X1 U4034 ( .A(n7650), .ZN(n5695) );
  NOR2_X1 U4035 ( .A1(n5252), .A2(n3837), .ZN(n7613) );
  NOR2_X1 U4036 ( .A1(n5252), .A2(n5901), .ZN(n7629) );
  AND2_X1 U4037 ( .A1(n4177), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7499) );
  AND2_X1 U4038 ( .A1(n7498), .A2(n7497), .ZN(n7506) );
  INV_X1 U4039 ( .A(n7506), .ZN(n7512) );
  INV_X1 U4040 ( .A(n4918), .ZN(n4919) );
  NAND2_X1 U4041 ( .A1(n6649), .A2(n4916), .ZN(n4920) );
  OAI22_X1 U4042 ( .A1(n6113), .A2(n6647), .B1(n4917), .B2(n7126), .ZN(n4918)
         );
  INV_X1 U4043 ( .A(n4388), .ZN(n4346) );
  AOI22_X1 U4044 ( .A1(n3816), .A2(n3915), .B1(n4176), .B2(n3651), .ZN(n3844)
         );
  AND2_X2 U4045 ( .A1(n3814), .A2(n4912), .ZN(n4725) );
  INV_X1 U4046 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3671) );
  INV_X1 U4047 ( .A(n4232), .ZN(n4647) );
  AND2_X1 U4048 ( .A1(n4039), .A2(n4038), .ZN(n3658) );
  NAND2_X1 U4049 ( .A1(n4176), .A2(n3653), .ZN(n3659) );
  OR2_X1 U4050 ( .A1(n3865), .A2(n3848), .ZN(n3661) );
  NAND2_X1 U4051 ( .A1(n4054), .A2(n4053), .ZN(n4068) );
  AND2_X1 U4052 ( .A1(n4464), .A2(n4463), .ZN(n3662) );
  AND2_X1 U4053 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3663) );
  INV_X1 U4054 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4118) );
  NOR2_X1 U4055 ( .A1(n4870), .A2(n4175), .ZN(n3664) );
  INV_X1 U4056 ( .A(n4220), .ZN(n5272) );
  NAND2_X1 U4057 ( .A1(n5350), .A2(n5349), .ZN(n3665) );
  NAND2_X1 U4058 ( .A1(n7126), .A2(n4193), .ZN(n6648) );
  INV_X1 U4059 ( .A(n6648), .ZN(n4916) );
  OR2_X1 U4060 ( .A1(n4890), .A2(n4742), .ZN(n7212) );
  OR2_X1 U4061 ( .A1(n6680), .A2(n4115), .ZN(n3666) );
  INV_X1 U4062 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4182) );
  NAND2_X1 U4063 ( .A1(n3880), .A2(n3879), .ZN(n3967) );
  AND3_X1 U4064 ( .A1(n3742), .A2(n3741), .A3(n3740), .ZN(n3667) );
  OR4_X1 U4065 ( .A1(n6801), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n6802), 
        .A4(n6050), .ZN(n3668) );
  NAND2_X1 U4066 ( .A1(n4999), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4998)
         );
  OR2_X1 U4067 ( .A1(n3986), .A2(n3985), .ZN(n3993) );
  OR2_X1 U4068 ( .A1(n3893), .A2(n3892), .ZN(n3901) );
  INV_X1 U4069 ( .A(n4055), .ZN(n4053) );
  NAND2_X1 U4070 ( .A1(n4040), .A2(n3658), .ZN(n4056) );
  OR2_X1 U4071 ( .A1(n3860), .A2(n3859), .ZN(n3925) );
  INV_X1 U4072 ( .A(n4130), .ZN(n4125) );
  AOI22_X1 U4073 ( .A1(n4673), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3631), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4074 ( .A1(n3783), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3902), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3678) );
  INV_X1 U4075 ( .A(n4552), .ZN(n4184) );
  INV_X1 U4076 ( .A(n4236), .ZN(n4237) );
  INV_X1 U4077 ( .A(n5094), .ZN(n4778) );
  NAND2_X1 U4078 ( .A1(n4056), .A2(n4055), .ZN(n4228) );
  NAND2_X1 U4079 ( .A1(n5225), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3947) );
  INV_X1 U4080 ( .A(n5124), .ZN(n4787) );
  INV_X1 U4081 ( .A(n6574), .ZN(n4551) );
  NAND2_X1 U4082 ( .A1(n4157), .A2(n4127), .ZN(n4158) );
  OAI22_X1 U4083 ( .A1(n4160), .A2(n4159), .B1(n4158), .B2(n4718), .ZN(n4161)
         );
  OR2_X1 U4084 ( .A1(n4649), .A2(n6503), .ZN(n4667) );
  INV_X1 U4085 ( .A(n4516), .ZN(n4183) );
  INV_X1 U4086 ( .A(n5754), .ZN(n4391) );
  INV_X1 U4087 ( .A(n5862), .ZN(n4799) );
  AND2_X1 U4088 ( .A1(n4786), .A2(n4785), .ZN(n5124) );
  XNOR2_X1 U4089 ( .A(n4068), .B(n4067), .ZN(n4252) );
  INV_X1 U4090 ( .A(n5057), .ZN(n3821) );
  AND4_X1 U4091 ( .A1(n3727), .A2(n3726), .A3(n3725), .A4(n3724), .ZN(n3735)
         );
  INV_X1 U4092 ( .A(n4966), .ZN(n4753) );
  INV_X1 U4093 ( .A(n6512), .ZN(n4630) );
  NAND2_X1 U4094 ( .A1(n4208), .A2(n4207), .ZN(n4968) );
  OR2_X1 U4095 ( .A1(n4667), .A2(n6119), .ZN(n4697) );
  OR2_X1 U4096 ( .A1(n4583), .A2(n6548), .ZN(n4604) );
  INV_X1 U4097 ( .A(n4645), .ZN(n4693) );
  AND2_X1 U4098 ( .A1(n7452), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4645) );
  AND4_X1 U4099 ( .A1(n4269), .A2(n4268), .A3(n4267), .A4(n4266), .ZN(n5121)
         );
  NAND2_X1 U4100 ( .A1(n4219), .A2(n4346), .ZN(n4227) );
  AND2_X1 U4101 ( .A1(n6751), .A2(n3663), .ZN(n6728) );
  INV_X1 U4102 ( .A(n5818), .ZN(n4816) );
  AND2_X1 U4103 ( .A1(n4806), .A2(n4805), .ZN(n5765) );
  AND2_X1 U4104 ( .A1(n3653), .A2(n4174), .ZN(n4127) );
  XNOR2_X1 U4105 ( .A(n3966), .B(n3967), .ZN(n5098) );
  NOR2_X1 U4106 ( .A1(n5169), .A2(n5271), .ZN(n5573) );
  INV_X1 U4107 ( .A(n6066), .ZN(n5663) );
  NOR2_X1 U4108 ( .A1(n5382), .A2(n5397), .ZN(n5462) );
  NOR2_X1 U4109 ( .A1(n6608), .A2(n7580), .ZN(n6927) );
  AOI21_X1 U4110 ( .B1(n7514), .B2(n5108), .A(n6059), .ZN(n5112) );
  OR2_X1 U4111 ( .A1(n4163), .A2(n4162), .ZN(n4718) );
  NAND2_X1 U4112 ( .A1(n4478), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4496)
         );
  AND2_X1 U4113 ( .A1(n4286), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4271)
         );
  INV_X1 U4114 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U4115 ( .A1(n5739), .A2(n5716), .ZN(n7324) );
  CLKBUF_X1 U4116 ( .A(n4753), .Z(n6022) );
  INV_X1 U4117 ( .A(n4910), .ZN(n4911) );
  INV_X1 U4118 ( .A(n6572), .ZN(n6589) );
  AND2_X1 U4119 ( .A1(n5515), .A2(n5514), .ZN(n5799) );
  INV_X1 U4120 ( .A(n7158), .ZN(n6791) );
  NAND2_X1 U4121 ( .A1(n3954), .A2(n3953), .ZN(n5103) );
  INV_X1 U4122 ( .A(n5911), .ZN(n5953) );
  AND2_X1 U4123 ( .A1(n5404), .A2(n5403), .ZN(n5537) );
  OR2_X1 U4124 ( .A1(n5381), .A2(n5101), .ZN(n5417) );
  INV_X1 U4125 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n7474) );
  INV_X1 U4126 ( .A(n5462), .ZN(n5509) );
  INV_X1 U4127 ( .A(n5639), .ZN(n5486) );
  AND2_X1 U4128 ( .A1(n7455), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4177) );
  INV_X1 U4129 ( .A(n6072), .ZN(n5739) );
  AND2_X1 U4130 ( .A1(n7301), .A2(STATE2_REG_3__SCAN_IN), .ZN(n7439) );
  CLKBUF_X1 U4131 ( .A(n5025), .Z(n5043) );
  INV_X1 U4132 ( .A(n7126), .ZN(n6636) );
  INV_X1 U4133 ( .A(n6669), .ZN(n7551) );
  AND2_X1 U4134 ( .A1(n4206), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4937) );
  AND2_X1 U4135 ( .A1(n6589), .A2(n6588), .ZN(n6758) );
  INV_X1 U4136 ( .A(n5987), .ZN(n6775) );
  AND2_X1 U4137 ( .A1(n5119), .A2(n5262), .ZN(n5515) );
  AND2_X1 U4138 ( .A1(n5091), .A2(n5024), .ZN(n7318) );
  INV_X1 U4139 ( .A(n7447), .ZN(n7166) );
  NOR2_X1 U4140 ( .A1(n6097), .A2(n4735), .ZN(n7483) );
  OAI21_X1 U4141 ( .B1(n6682), .B2(n6698), .A(n6681), .ZN(n6683) );
  NOR2_X1 U4142 ( .A1(n7261), .A2(n7197), .ZN(n7272) );
  XNOR2_X1 U4143 ( .A(n4087), .B(n4780), .ZN(n5347) );
  AND2_X1 U4144 ( .A1(n5169), .A2(n5381), .ZN(n5440) );
  AND2_X1 U4145 ( .A1(n5308), .A2(n7557), .ZN(n6974) );
  AND2_X1 U4146 ( .A1(n5283), .A2(n5415), .ZN(n6976) );
  AND2_X1 U4147 ( .A1(n5396), .A2(n5415), .ZN(n5698) );
  NOR2_X1 U4148 ( .A1(n5417), .A2(n5416), .ZN(n5658) );
  AND2_X1 U4149 ( .A1(n5565), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5304)
         );
  INV_X1 U4150 ( .A(n7563), .ZN(n7653) );
  AND2_X1 U4151 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5565) );
  INV_X1 U4152 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7576) );
  NOR2_X1 U4153 ( .A1(n5236), .A2(n5303), .ZN(n6961) );
  INV_X1 U4154 ( .A(n5369), .ZN(n5488) );
  NOR2_X1 U4155 ( .A1(n5252), .A2(n5230), .ZN(n7605) );
  NOR2_X1 U4156 ( .A1(n5252), .A2(n6086), .ZN(n7650) );
  INV_X1 U4157 ( .A(STATE_REG_2__SCAN_IN), .ZN(n7533) );
  OR2_X1 U4158 ( .A1(n5708), .A2(n5707), .ZN(n7190) );
  INV_X1 U4159 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n7520) );
  INV_X1 U4160 ( .A(n7439), .ZN(n7429) );
  NAND2_X1 U4161 ( .A1(n7301), .A2(n5713), .ZN(n7422) );
  INV_X1 U4162 ( .A(n7419), .ZN(n7435) );
  NAND2_X2 U4163 ( .A1(n6085), .A2(n5064), .ZN(n6669) );
  OR2_X1 U4164 ( .A1(n6097), .A2(n4941), .ZN(n7024) );
  NAND2_X1 U4165 ( .A1(n5708), .A2(n4922), .ZN(n5061) );
  OR2_X1 U4166 ( .A1(n7158), .A2(n5080), .ZN(n7169) );
  XNOR2_X1 U4167 ( .A(n4711), .B(n6050), .ZN(n6038) );
  OR2_X1 U4168 ( .A1(n7282), .A2(n4897), .ZN(n6906) );
  OR2_X1 U4169 ( .A1(n4890), .A2(n4738), .ZN(n6892) );
  INV_X1 U4170 ( .A(n7454), .ZN(n6045) );
  INV_X1 U4171 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n6061) );
  INV_X1 U4172 ( .A(n5111), .ZN(n5260) );
  INV_X1 U4173 ( .A(n6936), .ZN(n7594) );
  INV_X1 U4174 ( .A(n6941), .ZN(n7602) );
  INV_X1 U4175 ( .A(n6966), .ZN(n7642) );
  INV_X1 U4176 ( .A(n7582), .ZN(n5703) );
  INV_X1 U4177 ( .A(n7613), .ZN(n5677) );
  AND2_X1 U4178 ( .A1(n7587), .A2(n5307), .ZN(n5344) );
  INV_X1 U4179 ( .A(n7540), .ZN(n7174) );
  NAND2_X1 U4180 ( .A1(n4920), .A2(n4919), .ZN(U2829) );
  INV_X1 U4181 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4182 ( .A1(n4673), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3675) );
  AND2_X2 U4183 ( .A1(n4978), .A2(n5128), .ZN(n4519) );
  AND2_X4 U4184 ( .A1(n4974), .A2(n5138), .ZN(n3886) );
  AND2_X2 U4185 ( .A1(n4978), .A2(n5132), .ZN(n4433) );
  AND4_X2 U4186 ( .A1(n3675), .A2(n3674), .A3(n3673), .A4(n3672), .ZN(n3682)
         );
  AND2_X2 U4187 ( .A1(n4974), .A2(n3676), .ZN(n3931) );
  AND2_X2 U4188 ( .A1(n3676), .A2(n5163), .ZN(n3788) );
  AOI22_X1 U4189 ( .A1(n3931), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3788), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3680) );
  AND2_X2 U4190 ( .A1(n5138), .A2(n5163), .ZN(n3907) );
  AND2_X2 U4191 ( .A1(n3676), .A2(n5131), .ZN(n3937) );
  AOI22_X1 U4192 ( .A1(n3937), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3677) );
  AND4_X2 U4193 ( .A1(n3680), .A2(n3679), .A3(n3678), .A4(n3677), .ZN(n3681)
         );
  AND2_X4 U4194 ( .A1(n3682), .A2(n3681), .ZN(n4189) );
  AOI22_X1 U4195 ( .A1(n3657), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3777), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4196 ( .A1(n4519), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3886), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4197 ( .A1(n3931), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3783), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4198 ( .A1(n3788), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3683) );
  NAND4_X1 U4199 ( .A1(n3686), .A2(n3685), .A3(n3684), .A4(n3683), .ZN(n3692)
         );
  AOI22_X1 U4200 ( .A1(n4433), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3778), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4201 ( .A1(n3937), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3629), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4202 ( .A1(n3902), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3887), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3687) );
  NAND4_X1 U4203 ( .A1(n3690), .A2(n3688), .A3(n3689), .A4(n3687), .ZN(n3691)
         );
  OR2_X2 U4204 ( .A1(n3692), .A2(n3691), .ZN(n4192) );
  NAND2_X2 U4205 ( .A1(n4189), .A2(n4192), .ZN(n4173) );
  NAND2_X1 U4206 ( .A1(n3777), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3696) );
  NAND2_X1 U4207 ( .A1(n3657), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3695)
         );
  NAND2_X1 U4208 ( .A1(n4433), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3694)
         );
  NAND2_X1 U4209 ( .A1(n3886), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3693) );
  NAND2_X1 U4210 ( .A1(n4673), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3700) );
  NAND2_X1 U4211 ( .A1(n3931), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3699) );
  NAND2_X1 U4212 ( .A1(n3788), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3698) );
  NAND2_X1 U4213 ( .A1(n3887), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3697)
         );
  NAND2_X1 U4214 ( .A1(n3778), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3704)
         );
  NAND2_X1 U4215 ( .A1(n3772), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3703) );
  NAND2_X1 U4216 ( .A1(n3980), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3702)
         );
  NAND2_X1 U4217 ( .A1(n4519), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3701)
         );
  NAND2_X1 U4218 ( .A1(n3937), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3708) );
  NAND2_X1 U4219 ( .A1(n3783), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3707) );
  NAND2_X1 U4220 ( .A1(n3902), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3706) );
  NAND2_X1 U4221 ( .A1(n3907), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3705) );
  NAND2_X1 U4222 ( .A1(n4192), .A2(n3802), .ZN(n3713) );
  NAND2_X2 U4223 ( .A1(n4173), .A2(n3713), .ZN(n3813) );
  AOI22_X1 U4224 ( .A1(n3783), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3902), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4225 ( .A1(n3907), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3887), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4226 ( .A1(n3931), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3788), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4227 ( .A1(n3657), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3777), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4228 ( .A1(n4433), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3778), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4229 ( .A1(n4673), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4230 ( .A1(n4519), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3886), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3718) );
  NAND2_X2 U4231 ( .A1(n3723), .A2(n3722), .ZN(n3798) );
  NAND2_X2 U4232 ( .A1(n3813), .A2(n5225), .ZN(n3816) );
  AOI22_X1 U4233 ( .A1(n3783), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3902), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4234 ( .A1(n3931), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3788), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4235 ( .A1(n4433), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4236 ( .A1(n3907), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3887), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4237 ( .A1(n4673), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4519), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3728) );
  INV_X1 U4238 ( .A(n3728), .ZN(n3733) );
  AOI22_X1 U4239 ( .A1(n3778), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3886), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4240 ( .A1(n3937), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3729) );
  NAND3_X1 U4241 ( .A1(n3731), .A2(n3730), .A3(n3729), .ZN(n3732) );
  NOR2_X1 U4242 ( .A1(n3733), .A2(n3732), .ZN(n3734) );
  NAND2_X1 U4243 ( .A1(n4173), .A2(n4867), .ZN(n3817) );
  NAND2_X1 U4244 ( .A1(n3799), .A2(n3798), .ZN(n3736) );
  NOR2_X1 U4245 ( .A1(n4173), .A2(n3736), .ZN(n3737) );
  INV_X1 U4246 ( .A(n3737), .ZN(n3838) );
  NAND2_X1 U4247 ( .A1(n4912), .A2(n4868), .ZN(n3739) );
  AOI22_X1 U4248 ( .A1(n3931), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3783), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4249 ( .A1(n3907), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3887), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4250 ( .A1(n3937), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3902), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3741) );
  NAND2_X1 U4251 ( .A1(n3778), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3740)
         );
  AOI22_X1 U4252 ( .A1(n4636), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3886), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4253 ( .A1(n3657), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3777), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4254 ( .A1(n3788), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3629), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4255 ( .A1(n3631), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4519), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3745) );
  NAND2_X1 U4256 ( .A1(n5063), .A2(n3926), .ZN(n3841) );
  NAND2_X1 U4257 ( .A1(n4433), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3753)
         );
  NAND2_X1 U4258 ( .A1(n3657), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3752)
         );
  NAND2_X1 U4259 ( .A1(n4519), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3751)
         );
  NAND2_X1 U4260 ( .A1(n3778), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3750)
         );
  NAND2_X1 U4261 ( .A1(n4673), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3757) );
  NAND2_X1 U4262 ( .A1(n3931), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3756) );
  NAND2_X1 U4263 ( .A1(n3783), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3755) );
  NAND2_X1 U4264 ( .A1(n3902), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3754) );
  NAND2_X1 U4265 ( .A1(n3886), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3761) );
  NAND2_X1 U4266 ( .A1(n3631), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3760) );
  NAND2_X1 U4267 ( .A1(n3777), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3759) );
  NAND2_X1 U4268 ( .A1(n3630), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3758)
         );
  NAND2_X1 U4269 ( .A1(n3788), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3765) );
  NAND2_X1 U4270 ( .A1(n3937), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3764) );
  NAND2_X1 U4271 ( .A1(n3887), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3763)
         );
  NAND2_X1 U4272 ( .A1(n3907), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3762) );
  NAND2_X1 U4273 ( .A1(n3771), .A2(n3770), .ZN(n3797) );
  NAND2_X1 U4274 ( .A1(n4519), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3776)
         );
  NAND2_X1 U4275 ( .A1(n3772), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3775) );
  NAND2_X1 U4276 ( .A1(n4673), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3774) );
  NAND2_X1 U4277 ( .A1(n3886), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3773) );
  NAND2_X1 U4278 ( .A1(n3777), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3782) );
  NAND2_X1 U4279 ( .A1(n3652), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3781)
         );
  NAND2_X1 U4280 ( .A1(n4433), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3780)
         );
  NAND2_X1 U4281 ( .A1(n3778), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3779)
         );
  NAND2_X1 U4282 ( .A1(n3937), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3787) );
  NAND2_X1 U4283 ( .A1(n3783), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3786) );
  NAND2_X1 U4284 ( .A1(n3980), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3785)
         );
  NAND2_X1 U4285 ( .A1(n3902), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3784) );
  NAND2_X1 U4286 ( .A1(n3931), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3792) );
  NAND2_X1 U4287 ( .A1(n3788), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3791) );
  NAND2_X1 U4288 ( .A1(n3887), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3790)
         );
  NAND2_X1 U4289 ( .A1(n3907), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3789) );
  NAND4_X4 U4290 ( .A1(n3796), .A2(n3795), .A3(n3794), .A4(n3793), .ZN(n4743)
         );
  AND2_X1 U4291 ( .A1(n5230), .A2(n3926), .ZN(n3800) );
  OAI211_X1 U4292 ( .C1(n5063), .C2(n3798), .A(n3800), .B(n3813), .ZN(n4870)
         );
  INV_X1 U4293 ( .A(n4870), .ZN(n3804) );
  NAND2_X1 U4294 ( .A1(n7533), .A2(STATE_REG_1__SCAN_IN), .ZN(n7529) );
  INV_X1 U4295 ( .A(STATE_REG_1__SCAN_IN), .ZN(n7524) );
  NAND2_X1 U4296 ( .A1(n7524), .A2(STATE_REG_2__SCAN_IN), .ZN(n3801) );
  NAND2_X1 U4297 ( .A1(n7529), .A2(n3801), .ZN(n4712) );
  NAND2_X1 U4298 ( .A1(n3815), .A2(n5901), .ZN(n3803) );
  NAND4_X1 U4299 ( .A1(n3833), .A2(n3804), .A3(n3803), .A4(n3844), .ZN(n3805)
         );
  NAND2_X1 U4300 ( .A1(n3805), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3807) );
  NAND2_X1 U4301 ( .A1(n4157), .A2(n5063), .ZN(n3806) );
  NAND2_X1 U4302 ( .A1(n3807), .A2(n3806), .ZN(n3876) );
  NAND2_X1 U4303 ( .A1(n3876), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3825) );
  INV_X1 U4304 ( .A(n5565), .ZN(n3808) );
  NAND2_X1 U4305 ( .A1(n7474), .A2(n7576), .ZN(n6923) );
  NAND2_X1 U4306 ( .A1(n3808), .A2(n6923), .ZN(n5387) );
  NOR2_X1 U4307 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n7501) );
  NAND2_X1 U4308 ( .A1(n7501), .A2(n3848), .ZN(n4178) );
  OR2_X1 U4309 ( .A1(n5387), .A2(n4178), .ZN(n3811) );
  INV_X1 U4310 ( .A(n4177), .ZN(n3809) );
  NAND2_X1 U4311 ( .A1(n3809), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3810) );
  NAND2_X1 U4312 ( .A1(n3811), .A2(n3810), .ZN(n3827) );
  INV_X1 U4313 ( .A(n3827), .ZN(n3824) );
  NAND2_X1 U4314 ( .A1(n5063), .A2(n3798), .ZN(n3812) );
  NAND3_X1 U4315 ( .A1(n3813), .A2(n3926), .A3(n3812), .ZN(n3839) );
  INV_X1 U4316 ( .A(n3839), .ZN(n3814) );
  INV_X1 U4317 ( .A(n3815), .ZN(n3822) );
  INV_X1 U4318 ( .A(n3816), .ZN(n3819) );
  NAND2_X2 U4319 ( .A1(n4729), .A2(n3820), .ZN(n7460) );
  NAND3_X1 U4320 ( .A1(n4912), .A2(n5735), .A3(n3837), .ZN(n5057) );
  OAI211_X1 U4321 ( .C1(n6100), .C2(n3822), .A(n7460), .B(n4739), .ZN(n3823)
         );
  NAND2_X1 U4322 ( .A1(n3823), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3826) );
  NAND3_X1 U4323 ( .A1(n3825), .A2(n3824), .A3(n3826), .ZN(n3873) );
  INV_X1 U4324 ( .A(n3826), .ZN(n3829) );
  NAND2_X1 U4325 ( .A1(n3829), .A2(n3828), .ZN(n3830) );
  NAND2_X1 U4326 ( .A1(n3873), .A2(n3830), .ZN(n3870) );
  NAND2_X1 U4327 ( .A1(n3876), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3832) );
  MUX2_X1 U4328 ( .A(n4178), .B(n4177), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3831) );
  INV_X1 U4329 ( .A(n3833), .ZN(n3834) );
  NAND2_X1 U4330 ( .A1(n3834), .A2(n3659), .ZN(n3836) );
  NAND2_X1 U4331 ( .A1(n4867), .A2(n4743), .ZN(n3835) );
  NAND2_X1 U4332 ( .A1(n3839), .A2(n3654), .ZN(n3843) );
  NAND2_X1 U4333 ( .A1(n7501), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3840) );
  AOI21_X1 U4334 ( .B1(n3841), .B2(n3915), .A(n3840), .ZN(n3842) );
  OAI211_X1 U4335 ( .C1(n3926), .C2(n3838), .A(n3843), .B(n3842), .ZN(n3846)
         );
  INV_X1 U4336 ( .A(n3844), .ZN(n3845) );
  XNOR2_X1 U4337 ( .A(n3870), .B(n3871), .ZN(n4975) );
  INV_X1 U4338 ( .A(n4975), .ZN(n3849) );
  INV_X1 U4339 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4340 ( .A1(n3850), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4341 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n4553), .B1(n4674), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4342 ( .A1(n4676), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4675), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4343 ( .A1(n3936), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3902), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3851) );
  NAND4_X1 U4344 ( .A1(n3854), .A2(n3853), .A3(n3852), .A4(n3851), .ZN(n3860)
         );
  AOI22_X1 U4345 ( .A1(n4681), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4346 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n3636), .B1(n5133), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4347 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(n3886), .B1(n3938), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4348 ( .A1(n3637), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3855) );
  NAND4_X1 U4349 ( .A1(n3858), .A2(n3857), .A3(n3856), .A4(n3855), .ZN(n3859)
         );
  INV_X1 U4350 ( .A(n3925), .ZN(n3861) );
  OR2_X1 U4351 ( .A1(n3947), .A2(n3861), .ZN(n3868) );
  INV_X1 U4352 ( .A(n3862), .ZN(n3863) );
  XNOR2_X2 U4353 ( .A(n3864), .B(n3863), .ZN(n4202) );
  NAND2_X1 U4354 ( .A1(n4157), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3866) );
  NAND2_X1 U4355 ( .A1(n3650), .A2(n3925), .ZN(n3865) );
  AOI21_X2 U4356 ( .B1(n4202), .B2(n3848), .A(n3867), .ZN(n3920) );
  NAND2_X1 U4357 ( .A1(n3920), .A2(n3947), .ZN(n3869) );
  NAND3_X1 U4358 ( .A1(n3919), .A2(n3868), .A3(n3869), .ZN(n3922) );
  INV_X1 U4359 ( .A(n3870), .ZN(n3872) );
  NAND2_X1 U4360 ( .A1(n3872), .A2(n3871), .ZN(n3875) );
  NAND2_X1 U4361 ( .A1(n3969), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3880) );
  NOR2_X1 U4362 ( .A1(n5565), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3877)
         );
  NOR2_X1 U4363 ( .A1(n5304), .A2(n3877), .ZN(n5113) );
  INV_X1 U4364 ( .A(n4178), .ZN(n3973) );
  NOR2_X1 U4365 ( .A1(n4177), .A2(n5411), .ZN(n3878) );
  AOI21_X1 U4366 ( .B1(n5113), .B2(n3973), .A(n3878), .ZN(n3879) );
  NAND2_X1 U4367 ( .A1(n5098), .A2(n3848), .ZN(n3895) );
  AOI22_X1 U4368 ( .A1(n3634), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4369 ( .A1(n3936), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4674), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4370 ( .A1(n4676), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4675), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4371 ( .A1(n5133), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3882) );
  NAND4_X1 U4372 ( .A1(n3885), .A2(n3884), .A3(n3883), .A4(n3882), .ZN(n3893)
         );
  AOI22_X1 U4373 ( .A1(n4681), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3850), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4374 ( .A1(n4553), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4375 ( .A1(n3636), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4376 ( .A1(n3637), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3888) );
  NAND4_X1 U4377 ( .A1(n3891), .A2(n3890), .A3(n3889), .A4(n3888), .ZN(n3892)
         );
  AOI22_X1 U4378 ( .A1(n4167), .A2(n3901), .B1(n4157), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3894) );
  NAND2_X1 U4379 ( .A1(n3895), .A2(n3894), .ZN(n3897) );
  NAND2_X1 U4380 ( .A1(n3896), .A2(n3897), .ZN(n3989) );
  INV_X1 U4381 ( .A(n3896), .ZN(n3899) );
  INV_X1 U4382 ( .A(n3897), .ZN(n3898) );
  NAND2_X1 U4383 ( .A1(n3899), .A2(n3898), .ZN(n3900) );
  NAND2_X1 U4384 ( .A1(n3989), .A2(n3900), .ZN(n4197) );
  INV_X1 U4385 ( .A(n4197), .ZN(n5271) );
  INV_X1 U4386 ( .A(n3901), .ZN(n3914) );
  AOI22_X1 U4387 ( .A1(n3850), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4388 ( .A1(n4681), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4389 ( .A1(n4676), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4675), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4390 ( .A1(n4553), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3902), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3903) );
  NAND4_X1 U4391 ( .A1(n3906), .A2(n3905), .A3(n3904), .A4(n3903), .ZN(n3913)
         );
  AOI22_X1 U4392 ( .A1(n4674), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3886), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4393 ( .A1(n3636), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5133), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4394 ( .A1(n3631), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4395 ( .A1(n3637), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3908) );
  NAND4_X1 U4396 ( .A1(n3911), .A2(n3910), .A3(n3909), .A4(n3908), .ZN(n3912)
         );
  OR2_X1 U4397 ( .A1(n3913), .A2(n3912), .ZN(n3956) );
  NAND2_X1 U4398 ( .A1(n3925), .A2(n3956), .ZN(n3924) );
  NAND2_X1 U4399 ( .A1(n3924), .A2(n3914), .ZN(n3992) );
  OAI21_X1 U4400 ( .B1(n3914), .B2(n3924), .A(n3992), .ZN(n3916) );
  NAND2_X1 U4401 ( .A1(n3916), .A2(n3915), .ZN(n3917) );
  NAND2_X1 U4402 ( .A1(n3650), .A2(n3926), .ZN(n3955) );
  NAND2_X1 U4403 ( .A1(n3917), .A2(n3955), .ZN(n3918) );
  INV_X1 U4404 ( .A(n3919), .ZN(n3921) );
  NAND2_X1 U4405 ( .A1(n3921), .A2(n3920), .ZN(n3923) );
  NAND2_X1 U4406 ( .A1(n3923), .A2(n3922), .ZN(n5102) );
  NAND2_X1 U4407 ( .A1(n5102), .A2(n3653), .ZN(n3930) );
  OAI21_X1 U4408 ( .B1(n3956), .B2(n3925), .A(n3924), .ZN(n3927) );
  INV_X1 U4409 ( .A(n3915), .ZN(n4728) );
  OAI211_X1 U4410 ( .C1(n3927), .C2(n4728), .A(n4174), .B(n3926), .ZN(n3928)
         );
  INV_X1 U4411 ( .A(n3928), .ZN(n3929) );
  NAND2_X1 U4412 ( .A1(n3930), .A2(n3929), .ZN(n5010) );
  NAND2_X1 U4413 ( .A1(n4202), .A2(n3848), .ZN(n3954) );
  NAND2_X1 U4414 ( .A1(n4157), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3946) );
  AOI21_X1 U4415 ( .B1(n3650), .B2(n3956), .A(n3848), .ZN(n3945) );
  AOI22_X1 U4416 ( .A1(n3850), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4417 ( .A1(n3634), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3886), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4418 ( .A1(n4676), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3636), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4419 ( .A1(n3637), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3932) );
  NAND4_X1 U4420 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3944)
         );
  AOI22_X1 U4421 ( .A1(n4553), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4422 ( .A1(n4681), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4674), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4423 ( .A1(n5133), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4424 ( .A1(n4675), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3902), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3939) );
  NAND4_X1 U4425 ( .A1(n3942), .A2(n3941), .A3(n3940), .A4(n3939), .ZN(n3943)
         );
  NAND2_X1 U4426 ( .A1(n5225), .A2(n4084), .ZN(n4080) );
  NAND3_X1 U4427 ( .A1(n3946), .A2(n3945), .A3(n4080), .ZN(n3952) );
  INV_X1 U4428 ( .A(n3947), .ZN(n3950) );
  INV_X1 U4429 ( .A(n4084), .ZN(n3948) );
  XNOR2_X1 U4430 ( .A(n3948), .B(n3956), .ZN(n3949) );
  NAND2_X1 U4431 ( .A1(n3950), .A2(n3949), .ZN(n3951) );
  XNOR2_X1 U4432 ( .A(n3952), .B(n3951), .ZN(n3953) );
  INV_X1 U4433 ( .A(n4127), .ZN(n4726) );
  OAI21_X1 U4434 ( .B1(n4728), .B2(n3956), .A(n3955), .ZN(n3957) );
  INV_X1 U4435 ( .A(n3957), .ZN(n3958) );
  OAI21_X1 U4436 ( .B1(n5103), .B2(n4726), .A(n3958), .ZN(n4999) );
  INV_X1 U4437 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5014) );
  NOR2_X1 U4438 ( .A1(n4998), .A2(n5014), .ZN(n3960) );
  NAND2_X1 U4439 ( .A1(n4998), .A2(n5014), .ZN(n3959) );
  OAI21_X1 U4440 ( .B1(n5010), .B2(n3960), .A(n3959), .ZN(n3961) );
  NAND2_X1 U4441 ( .A1(n7129), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3962)
         );
  NAND2_X1 U4442 ( .A1(n7128), .A2(n3962), .ZN(n3965) );
  INV_X1 U4443 ( .A(n7129), .ZN(n3963) );
  INV_X1 U4444 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n7234) );
  NAND2_X1 U4445 ( .A1(n3963), .A2(n7234), .ZN(n3964) );
  INV_X1 U4446 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U4447 ( .A1(n3969), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3975) );
  NAND2_X1 U4448 ( .A1(n5304), .A2(n7480), .ZN(n5662) );
  INV_X1 U4449 ( .A(n5304), .ZN(n3970) );
  NAND2_X1 U4450 ( .A1(n3970), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3971) );
  NAND2_X1 U4451 ( .A1(n5662), .A2(n3971), .ZN(n5423) );
  NOR2_X1 U4452 ( .A1(n4177), .A2(n7480), .ZN(n3972) );
  AOI21_X1 U4453 ( .B1(n5423), .B2(n3973), .A(n3972), .ZN(n3974) );
  AOI22_X1 U4454 ( .A1(n3850), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4455 ( .A1(n4681), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4456 ( .A1(n4553), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3936), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4457 ( .A1(n4674), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3976) );
  NAND4_X1 U4458 ( .A1(n3979), .A2(n3978), .A3(n3977), .A4(n3976), .ZN(n3986)
         );
  AOI22_X1 U4459 ( .A1(n4676), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3636), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4460 ( .A1(n5133), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4461 ( .A1(n4675), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4462 ( .A1(n3637), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3981) );
  NAND4_X1 U4463 ( .A1(n3984), .A2(n3983), .A3(n3982), .A4(n3981), .ZN(n3985)
         );
  AOI22_X1 U4464 ( .A1(n4167), .A2(n3993), .B1(n4157), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3987) );
  NOR2_X2 U4465 ( .A1(n3989), .A2(n3990), .ZN(n4010) );
  INV_X1 U4466 ( .A(n4010), .ZN(n4037) );
  NAND2_X1 U4467 ( .A1(n5100), .A2(n3989), .ZN(n3991) );
  NAND2_X1 U4468 ( .A1(n3992), .A2(n3993), .ZN(n4031) );
  OAI211_X1 U4469 ( .C1(n3993), .C2(n3992), .A(n4031), .B(n3915), .ZN(n3994)
         );
  OAI21_X1 U4470 ( .B1(n4188), .B2(n4726), .A(n3994), .ZN(n3995) );
  INV_X1 U4471 ( .A(n3995), .ZN(n5068) );
  NAND2_X1 U4472 ( .A1(n5067), .A2(n5072), .ZN(n3996) );
  AOI22_X1 U4473 ( .A1(n3634), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4474 ( .A1(n4553), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4475 ( .A1(n4676), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5133), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4476 ( .A1(n3636), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3998) );
  NAND4_X1 U4477 ( .A1(n4001), .A2(n4000), .A3(n3999), .A4(n3998), .ZN(n4007)
         );
  AOI22_X1 U4478 ( .A1(n4681), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3850), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U4479 ( .A1(n3936), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4674), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4480 ( .A1(n4683), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4481 ( .A1(n4675), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4002) );
  NAND4_X1 U4482 ( .A1(n4005), .A2(n4004), .A3(n4003), .A4(n4002), .ZN(n4006)
         );
  NAND2_X1 U4483 ( .A1(n4167), .A2(n4029), .ZN(n4009) );
  NAND2_X1 U4484 ( .A1(n4157), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4008) );
  NAND2_X1 U4485 ( .A1(n4009), .A2(n4008), .ZN(n4039) );
  NAND2_X1 U4486 ( .A1(n4010), .A2(n4039), .ZN(n4028) );
  NAND2_X1 U4487 ( .A1(n4011), .A2(n4028), .ZN(n4218) );
  XNOR2_X1 U4488 ( .A(n4031), .B(n4029), .ZN(n4012) );
  NAND2_X1 U4489 ( .A1(n4012), .A2(n3915), .ZN(n4013) );
  INV_X1 U4490 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4765) );
  NAND2_X1 U4491 ( .A1(n7137), .A2(n7136), .ZN(n7135) );
  NAND2_X1 U4492 ( .A1(n4014), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4015)
         );
  NAND2_X1 U4493 ( .A1(n7135), .A2(n4015), .ZN(n7142) );
  AOI22_X1 U4494 ( .A1(n3850), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4495 ( .A1(n4681), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4496 ( .A1(n4553), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3936), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4497 ( .A1(n4674), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4016) );
  NAND4_X1 U4498 ( .A1(n4019), .A2(n4018), .A3(n4017), .A4(n4016), .ZN(n4025)
         );
  AOI22_X1 U4499 ( .A1(n4676), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3636), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4500 ( .A1(n5133), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4501 ( .A1(n4675), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4502 ( .A1(n3637), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4020) );
  NAND4_X1 U4503 ( .A1(n4023), .A2(n4022), .A3(n4021), .A4(n4020), .ZN(n4024)
         );
  NAND2_X1 U4504 ( .A1(n4167), .A2(n4058), .ZN(n4027) );
  NAND2_X1 U4505 ( .A1(n4157), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4026) );
  NAND2_X1 U4506 ( .A1(n4027), .A2(n4026), .ZN(n4038) );
  NAND2_X1 U4507 ( .A1(n4239), .A2(n4127), .ZN(n4034) );
  INV_X1 U4508 ( .A(n4029), .ZN(n4030) );
  OR2_X1 U4509 ( .A1(n4031), .A2(n4030), .ZN(n4057) );
  XNOR2_X1 U4510 ( .A(n4057), .B(n4058), .ZN(n4032) );
  NAND2_X1 U4511 ( .A1(n4032), .A2(n3915), .ZN(n4033) );
  NAND2_X1 U4512 ( .A1(n4034), .A2(n4033), .ZN(n4035) );
  INV_X1 U4513 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n7213) );
  XNOR2_X1 U4514 ( .A(n4035), .B(n7213), .ZN(n7144) );
  NAND2_X1 U4515 ( .A1(n7142), .A2(n7144), .ZN(n7143) );
  NAND2_X1 U4516 ( .A1(n4035), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4036)
         );
  NAND2_X1 U4517 ( .A1(n7143), .A2(n4036), .ZN(n7148) );
  AOI22_X1 U4518 ( .A1(n4553), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3936), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U4519 ( .A1(n4681), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4674), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U4520 ( .A1(n5133), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U4521 ( .A1(n3636), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4041) );
  NAND4_X1 U4522 ( .A1(n4044), .A2(n4043), .A3(n4042), .A4(n4041), .ZN(n4050)
         );
  AOI22_X1 U4523 ( .A1(n3850), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U4524 ( .A1(n3634), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U4525 ( .A1(n4675), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U4526 ( .A1(n4676), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4045) );
  NAND4_X1 U4527 ( .A1(n4048), .A2(n4047), .A3(n4046), .A4(n4045), .ZN(n4049)
         );
  NAND2_X1 U4528 ( .A1(n4167), .A2(n4070), .ZN(n4052) );
  NAND2_X1 U4529 ( .A1(n4157), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4051) );
  INV_X1 U4530 ( .A(n4228), .ZN(n4062) );
  INV_X1 U4531 ( .A(n4057), .ZN(n4059) );
  NAND2_X1 U4532 ( .A1(n4059), .A2(n4058), .ZN(n4069) );
  INV_X1 U4533 ( .A(n4070), .ZN(n4060) );
  XNOR2_X1 U4534 ( .A(n4069), .B(n4060), .ZN(n4061) );
  OAI22_X1 U4535 ( .A1(n4079), .A2(n4062), .B1(n4061), .B2(n4728), .ZN(n7150)
         );
  OAI21_X1 U4536 ( .B1(n7148), .B2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n7150), 
        .ZN(n4064) );
  NAND2_X1 U4537 ( .A1(n7148), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4063)
         );
  NAND2_X1 U4538 ( .A1(n4064), .A2(n4063), .ZN(n5360) );
  NAND2_X1 U4539 ( .A1(n4167), .A2(n4084), .ZN(n4066) );
  NAND2_X1 U4540 ( .A1(n4157), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4065) );
  NAND2_X1 U4541 ( .A1(n4066), .A2(n4065), .ZN(n4067) );
  NAND2_X1 U4542 ( .A1(n4252), .A2(n4127), .ZN(n4074) );
  INV_X1 U4543 ( .A(n4069), .ZN(n4071) );
  NAND2_X1 U4544 ( .A1(n4071), .A2(n4070), .ZN(n4083) );
  XNOR2_X1 U4545 ( .A(n4083), .B(n4084), .ZN(n4072) );
  NAND2_X1 U4546 ( .A1(n4072), .A2(n3915), .ZN(n4073) );
  NAND2_X1 U4547 ( .A1(n4074), .A2(n4073), .ZN(n4076) );
  INV_X1 U4548 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4075) );
  XNOR2_X1 U4549 ( .A(n4076), .B(n4075), .ZN(n5362) );
  NAND2_X1 U4550 ( .A1(n5360), .A2(n5362), .ZN(n4078) );
  NAND2_X1 U4551 ( .A1(n4076), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4077)
         );
  NAND2_X1 U4552 ( .A1(n4078), .A2(n4077), .ZN(n5345) );
  NOR2_X1 U4553 ( .A1(n4080), .A2(n3848), .ZN(n4081) );
  NAND2_X4 U4554 ( .A1(n4082), .A2(n4081), .ZN(n6751) );
  INV_X1 U4555 ( .A(n4083), .ZN(n4085) );
  NAND3_X1 U4556 ( .A1(n4085), .A2(n3915), .A3(n4084), .ZN(n4086) );
  NAND2_X1 U4557 ( .A1(n6751), .A2(n4086), .ZN(n4087) );
  INV_X1 U4558 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4780) );
  NAND2_X1 U4559 ( .A1(n5345), .A2(n5347), .ZN(n4089) );
  NAND2_X1 U4560 ( .A1(n4087), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4088)
         );
  NAND2_X1 U4561 ( .A1(n4089), .A2(n4088), .ZN(n5791) );
  XNOR2_X1 U4562 ( .A(n6751), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5793)
         );
  NAND2_X1 U4563 ( .A1(n5791), .A2(n5793), .ZN(n4091) );
  NAND2_X1 U4564 ( .A1(n6769), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4090)
         );
  NAND2_X1 U4565 ( .A1(n4091), .A2(n4090), .ZN(n5827) );
  INV_X1 U4566 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4790) );
  NAND2_X1 U4567 ( .A1(n6751), .A2(n4790), .ZN(n5829) );
  NAND2_X1 U4568 ( .A1(n5827), .A2(n5829), .ZN(n5851) );
  INV_X1 U4569 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n7198) );
  AND2_X1 U4570 ( .A1(n6751), .A2(n7198), .ZN(n5852) );
  INV_X1 U4571 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4801) );
  NAND2_X1 U4572 ( .A1(n6769), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U4573 ( .A1(n6769), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5850) );
  OAI211_X1 U4574 ( .C1(n6751), .C2(n4801), .A(n5884), .B(n5850), .ZN(n4092)
         );
  INV_X1 U4575 ( .A(n4092), .ZN(n4093) );
  OAI21_X1 U4576 ( .B1(n5851), .B2(n5852), .A(n4093), .ZN(n4095) );
  NAND2_X1 U4577 ( .A1(n6751), .A2(n4801), .ZN(n4094) );
  NAND2_X1 U4578 ( .A1(n4095), .A2(n4094), .ZN(n5959) );
  XNOR2_X1 U4579 ( .A(n6751), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5961)
         );
  NAND2_X1 U4580 ( .A1(n5959), .A2(n5961), .ZN(n4098) );
  INV_X1 U4581 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4096) );
  NAND2_X1 U4582 ( .A1(n6751), .A2(n4096), .ZN(n4097) );
  NAND2_X1 U4583 ( .A1(n4098), .A2(n4097), .ZN(n5967) );
  XNOR2_X1 U4584 ( .A(n6751), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5969)
         );
  NAND2_X1 U4585 ( .A1(n5967), .A2(n5969), .ZN(n4100) );
  INV_X1 U4586 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4810) );
  NAND2_X1 U4587 ( .A1(n6751), .A2(n4810), .ZN(n4099) );
  NAND2_X1 U4588 ( .A1(n4100), .A2(n4099), .ZN(n6000) );
  INV_X1 U4589 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n7268) );
  NAND2_X1 U4590 ( .A1(n6769), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6002) );
  OAI21_X2 U4591 ( .B1(n6000), .B2(n6003), .A(n6002), .ZN(n6012) );
  INV_X1 U4592 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4818) );
  NAND2_X1 U4593 ( .A1(n6751), .A2(n4818), .ZN(n6014) );
  NAND2_X1 U4594 ( .A1(n6012), .A2(n6014), .ZN(n6785) );
  NAND2_X1 U4595 ( .A1(n6769), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U4596 ( .A1(n6785), .A2(n6015), .ZN(n6786) );
  NOR2_X1 U4597 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4101) );
  NAND2_X1 U4598 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4897) );
  NAND2_X1 U4599 ( .A1(n6751), .A2(n4897), .ZN(n4102) );
  OAI21_X1 U4600 ( .B1(n6786), .B2(n4103), .A(n4102), .ZN(n6724) );
  NOR2_X1 U4601 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6889) );
  NOR2_X1 U4602 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6729) );
  INV_X1 U4603 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6860) );
  INV_X1 U4604 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6849) );
  NAND4_X1 U4605 ( .A1(n6889), .A2(n6729), .A3(n6860), .A4(n6849), .ZN(n4104)
         );
  NAND2_X1 U4606 ( .A1(n6769), .A2(n4104), .ZN(n4105) );
  NAND2_X1 U4607 ( .A1(n6724), .A2(n4105), .ZN(n4107) );
  AND2_X1 U4608 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6888) );
  AND2_X1 U4609 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4888) );
  AND2_X1 U4610 ( .A1(n6888), .A2(n4888), .ZN(n6857) );
  AND2_X1 U4611 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4901) );
  NAND2_X1 U4612 ( .A1(n6857), .A2(n4901), .ZN(n4883) );
  NAND2_X1 U4613 ( .A1(n6751), .A2(n4883), .ZN(n4106) );
  NAND2_X1 U4614 ( .A1(n4107), .A2(n4106), .ZN(n6720) );
  INV_X1 U4615 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6846) );
  XNOR2_X1 U4616 ( .A(n6751), .B(n6846), .ZN(n6719) );
  NAND2_X1 U4617 ( .A1(n6769), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4108) );
  NAND2_X1 U4618 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6682) );
  NAND2_X1 U4619 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4114) );
  NOR2_X1 U4620 ( .A1(n6682), .A2(n4114), .ZN(n4109) );
  NAND2_X1 U4621 ( .A1(n6708), .A2(n4109), .ZN(n4113) );
  OAI21_X1 U4622 ( .B1(n4110), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n6769), 
        .ZN(n4112) );
  INV_X1 U4623 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6835) );
  INV_X1 U4624 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6812) );
  NAND2_X1 U4625 ( .A1(n6835), .A2(n6812), .ZN(n4111) );
  NAND2_X1 U4626 ( .A1(n6769), .A2(n4111), .ZN(n6689) );
  INV_X1 U4627 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6050) );
  NOR2_X1 U4628 ( .A1(n6751), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6680)
         );
  NOR3_X1 U4629 ( .A1(n4114), .A2(n6682), .A3(n6050), .ZN(n4115) );
  XNOR2_X1 U4630 ( .A(n4119), .B(n4118), .ZN(n6053) );
  INV_X1 U4631 ( .A(n4157), .ZN(n4124) );
  XNOR2_X1 U4632 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4126) );
  NAND2_X1 U4633 ( .A1(n7576), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4130) );
  NAND2_X1 U4634 ( .A1(n4126), .A2(n4125), .ZN(n4121) );
  NAND2_X1 U4635 ( .A1(n7474), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4120) );
  NAND2_X1 U4636 ( .A1(n4121), .A2(n4120), .ZN(n4143) );
  XNOR2_X1 U4637 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4142) );
  NAND2_X1 U4638 ( .A1(n4143), .A2(n4142), .ZN(n4123) );
  NAND2_X1 U4639 ( .A1(n5411), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4122) );
  NAND2_X1 U4640 ( .A1(n4123), .A2(n4122), .ZN(n4154) );
  XNOR2_X1 U4641 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4153) );
  XNOR2_X1 U4642 ( .A(n4154), .B(n4153), .ZN(n4715) );
  NAND2_X1 U4643 ( .A1(n4124), .A2(n4715), .ZN(n4152) );
  XNOR2_X1 U4644 ( .A(n4126), .B(n4125), .ZN(n4713) );
  INV_X1 U4645 ( .A(n4713), .ZN(n4128) );
  AOI21_X1 U4646 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n4128), .A(n4168), .ZN(
        n4136) );
  INV_X1 U4647 ( .A(n4136), .ZN(n4141) );
  OAI21_X1 U4648 ( .B1(n4145), .B2(n3820), .A(n4174), .ZN(n4129) );
  AOI21_X1 U4649 ( .B1(n4157), .B2(n4713), .A(n4129), .ZN(n4137) );
  INV_X1 U4650 ( .A(n4137), .ZN(n4140) );
  OAI21_X1 U4651 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7576), .A(n4130), 
        .ZN(n4133) );
  INV_X1 U4652 ( .A(n4133), .ZN(n4131) );
  NAND2_X1 U4653 ( .A1(n4167), .A2(n4131), .ZN(n4138) );
  OAI21_X1 U4654 ( .B1(n4176), .B2(n4133), .A(n4132), .ZN(n4135) );
  NAND2_X1 U4655 ( .A1(n5901), .A2(n4743), .ZN(n4134) );
  NAND2_X1 U4656 ( .A1(n4134), .A2(n3820), .ZN(n4144) );
  AOI222_X1 U4657 ( .A1(n4138), .A2(n4158), .B1(n4137), .B2(n4136), .C1(n4135), 
        .C2(n4144), .ZN(n4139) );
  AOI21_X1 U4658 ( .B1(n4141), .B2(n4140), .A(n4139), .ZN(n4150) );
  XNOR2_X1 U4659 ( .A(n4143), .B(n4142), .ZN(n4714) );
  INV_X1 U4660 ( .A(n4144), .ZN(n4147) );
  NOR2_X1 U4661 ( .A1(n4145), .A2(n4714), .ZN(n4146) );
  AOI211_X1 U4662 ( .C1(n4157), .C2(n4714), .A(n4147), .B(n4146), .ZN(n4149)
         );
  NAND2_X1 U4663 ( .A1(n4167), .A2(n4147), .ZN(n4148) );
  OAI22_X1 U4664 ( .A1(n4150), .A2(n4149), .B1(n4714), .B2(n4148), .ZN(n4151)
         );
  AOI22_X1 U4665 ( .A1(n4152), .A2(n4151), .B1(n4168), .B2(n4715), .ZN(n4160)
         );
  NAND2_X1 U4666 ( .A1(n4154), .A2(n4153), .ZN(n4156) );
  NAND2_X1 U4667 ( .A1(n7480), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4155) );
  NAND2_X1 U4668 ( .A1(n4156), .A2(n4155), .ZN(n4163) );
  NAND2_X1 U4669 ( .A1(n7465), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4162) );
  NAND2_X1 U4670 ( .A1(n4163), .A2(n4162), .ZN(n4166) );
  INV_X1 U4671 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4164) );
  NAND2_X1 U4672 ( .A1(n4164), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4165) );
  NAND2_X1 U4673 ( .A1(n4166), .A2(n4165), .ZN(n4717) );
  NAND2_X1 U4674 ( .A1(n4167), .A2(n4717), .ZN(n4169) );
  INV_X1 U4675 ( .A(n4877), .ZN(n4205) );
  AOI21_X1 U4676 ( .B1(n4205), .B2(n4174), .A(n4743), .ZN(n4175) );
  NAND2_X1 U4677 ( .A1(n3664), .A2(n4176), .ZN(n4735) );
  NOR2_X1 U4678 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n7590) );
  INV_X1 U4679 ( .A(n7590), .ZN(n7580) );
  NAND2_X1 U4680 ( .A1(n7580), .A2(n4178), .ZN(n7191) );
  NAND2_X1 U4681 ( .A1(n7191), .A2(n3848), .ZN(n4179) );
  NAND2_X1 U4682 ( .A1(n3848), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4181) );
  NAND2_X1 U4683 ( .A1(n7520), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4180) );
  AND2_X1 U4684 ( .A1(n4181), .A2(n4180), .ZN(n5080) );
  INV_X1 U4685 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5729) );
  INV_X1 U4686 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6018) );
  INV_X1 U4687 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6780) );
  INV_X1 U4688 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4495) );
  INV_X1 U4689 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4546) );
  INV_X1 U4690 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6548) );
  INV_X1 U4691 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6531) );
  INV_X1 U4692 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6503) );
  INV_X1 U4693 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6119) );
  INV_X1 U4694 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6104) );
  XNOR2_X1 U4695 ( .A(n4185), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5719)
         );
  NAND2_X1 U4696 ( .A1(n7590), .A2(n7455), .ZN(n7178) );
  OR2_X2 U4697 ( .A1(n7178), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7211) );
  INV_X1 U4698 ( .A(REIP_REG_31__SCAN_IN), .ZN(n7070) );
  NOR2_X1 U4699 ( .A1(n7211), .A2(n7070), .ZN(n6046) );
  AOI21_X1 U4700 ( .B1(n7158), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n6046), 
        .ZN(n4186) );
  OAI21_X1 U4701 ( .B1(n7169), .B2(n5719), .A(n4186), .ZN(n4187) );
  INV_X1 U4702 ( .A(n4187), .ZN(n4707) );
  NAND2_X1 U4703 ( .A1(n4189), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4388) );
  NAND2_X1 U4704 ( .A1(n4868), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4224) );
  INV_X2 U4705 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n7188) );
  NAND2_X1 U4706 ( .A1(n7188), .A2(n7520), .ZN(n4220) );
  NAND2_X1 U4707 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4210) );
  INV_X1 U4708 ( .A(n4210), .ZN(n4191) );
  INV_X1 U4709 ( .A(n4221), .ZN(n4190) );
  OAI21_X1 U4710 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n4191), .A(n4190), 
        .ZN(n6606) );
  AOI22_X1 U4711 ( .A1(n5272), .A2(n6606), .B1(n4700), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4195) );
  NOR2_X2 U4712 ( .A1(n4193), .A2(n7188), .ZN(n4232) );
  NAND2_X1 U4713 ( .A1(n4232), .A2(EAX_REG_3__SCAN_IN), .ZN(n4194) );
  OAI211_X1 U4714 ( .C1(n4224), .C2(n3671), .A(n4195), .B(n4194), .ZN(n4196)
         );
  INV_X1 U4715 ( .A(n4700), .ZN(n4403) );
  NAND2_X1 U4716 ( .A1(n5102), .A2(n4346), .ZN(n4201) );
  INV_X1 U4717 ( .A(n4224), .ZN(n4209) );
  NAND2_X1 U4718 ( .A1(n4209), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4199) );
  AOI22_X1 U4719 ( .A1(n4701), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n7188), .ZN(n4198) );
  AND2_X1 U4720 ( .A1(n4199), .A2(n4198), .ZN(n4200) );
  NAND2_X1 U4721 ( .A1(n4201), .A2(n4200), .ZN(n4969) );
  INV_X1 U4722 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n7451) );
  NAND2_X1 U4723 ( .A1(n7454), .A2(n4346), .ZN(n4204) );
  AOI22_X1 U4724 ( .A1(n4701), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n7188), .ZN(n4203) );
  OAI211_X1 U4725 ( .C1(n4224), .C2(n7451), .A(n4204), .B(n4203), .ZN(n4936)
         );
  OR2_X1 U4726 ( .A1(n4936), .A2(n4220), .ZN(n4208) );
  NAND2_X1 U4727 ( .A1(n5103), .A2(n4205), .ZN(n4206) );
  NAND2_X1 U4728 ( .A1(n4936), .A2(n4937), .ZN(n4207) );
  NAND2_X1 U4729 ( .A1(n4969), .A2(n4968), .ZN(n4970) );
  NAND2_X1 U4730 ( .A1(n4209), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4214) );
  OAI21_X1 U4731 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n4210), .ZN(n7134) );
  NAND2_X1 U4732 ( .A1(n5272), .A2(n7134), .ZN(n4211) );
  OAI21_X1 U4733 ( .B1(n4182), .B2(n4403), .A(n4211), .ZN(n4212) );
  AOI21_X1 U4734 ( .B1(n4701), .B2(EAX_REG_2__SCAN_IN), .A(n4212), .ZN(n4213)
         );
  AND2_X1 U4735 ( .A1(n4214), .A2(n4213), .ZN(n4215) );
  NOR2_X1 U4736 ( .A1(n4970), .A2(n4215), .ZN(n4216) );
  NAND2_X1 U4737 ( .A1(n4970), .A2(n4215), .ZN(n4962) );
  OAI21_X1 U4738 ( .B1(n4961), .B2(n4216), .A(n4962), .ZN(n4960) );
  INV_X1 U4739 ( .A(n4960), .ZN(n5032) );
  INV_X1 U4740 ( .A(n4218), .ZN(n4219) );
  XNOR2_X1 U4741 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .B(n4221), .ZN(n7289) );
  OAI21_X1 U4742 ( .B1(n7520), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n7188), 
        .ZN(n4223) );
  NAND2_X1 U4743 ( .A1(n4701), .A2(EAX_REG_4__SCAN_IN), .ZN(n4222) );
  OAI211_X1 U4744 ( .C1(n4224), .C2(n7465), .A(n4223), .B(n4222), .ZN(n4225)
         );
  OAI21_X1 U4745 ( .B1(n4220), .B2(n7289), .A(n4225), .ZN(n4226) );
  NOR2_X2 U4746 ( .A1(n5031), .A2(n5078), .ZN(n5021) );
  NAND2_X1 U4747 ( .A1(n4228), .A2(n4346), .ZN(n4238) );
  INV_X1 U4748 ( .A(n4248), .ZN(n4231) );
  INV_X1 U4749 ( .A(n4229), .ZN(n4243) );
  INV_X1 U4750 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4233) );
  NAND2_X1 U4751 ( .A1(n4243), .A2(n4233), .ZN(n4230) );
  NAND2_X1 U4752 ( .A1(n4231), .A2(n4230), .ZN(n7321) );
  INV_X1 U4753 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4234) );
  OAI22_X1 U4754 ( .A1(n4647), .A2(n4234), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4233), .ZN(n4235) );
  MUX2_X1 U4755 ( .A(n7321), .B(n4235), .S(n4220), .Z(n4236) );
  INV_X1 U4756 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4246) );
  NAND2_X1 U4757 ( .A1(n4239), .A2(n4346), .ZN(n4245) );
  INV_X1 U4758 ( .A(n4240), .ZN(n4241) );
  INV_X1 U4759 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n7298) );
  NAND2_X1 U4760 ( .A1(n4241), .A2(n7298), .ZN(n4242) );
  NAND2_X1 U4761 ( .A1(n4243), .A2(n4242), .ZN(n7309) );
  AOI22_X1 U4762 ( .A1(n7309), .A2(n5272), .B1(n4700), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4244) );
  NAND2_X1 U4763 ( .A1(n5021), .A2(n4247), .ZN(n5020) );
  INV_X1 U4764 ( .A(n5020), .ZN(n4254) );
  INV_X1 U4765 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4250) );
  OAI21_X1 U4766 ( .B1(n4248), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n4265), 
        .ZN(n7326) );
  AOI22_X1 U4767 ( .A1(n7326), .A2(n5272), .B1(n4700), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4249) );
  OAI21_X1 U4768 ( .B1(n4647), .B2(n4250), .A(n4249), .ZN(n4251) );
  INV_X1 U4769 ( .A(n5087), .ZN(n4253) );
  NAND2_X1 U4770 ( .A1(n4254), .A2(n4253), .ZN(n5088) );
  AOI22_X1 U4771 ( .A1(n3634), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4258) );
  AOI22_X1 U4772 ( .A1(n4676), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3636), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4257) );
  AOI22_X1 U4773 ( .A1(n4675), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4256) );
  AOI22_X1 U4774 ( .A1(n3637), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4255) );
  NAND4_X1 U4775 ( .A1(n4258), .A2(n4257), .A3(n4256), .A4(n4255), .ZN(n4264)
         );
  AOI22_X1 U4776 ( .A1(n3850), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4262) );
  AOI22_X1 U4777 ( .A1(n4553), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3936), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4261) );
  AOI22_X1 U4778 ( .A1(n4681), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4674), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4260) );
  AOI22_X1 U4779 ( .A1(n5133), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4259) );
  NAND4_X1 U4780 ( .A1(n4262), .A2(n4261), .A3(n4260), .A4(n4259), .ZN(n4263)
         );
  OAI21_X1 U4781 ( .B1(n4264), .B2(n4263), .A(n4346), .ZN(n4269) );
  NAND2_X1 U4782 ( .A1(n4232), .A2(EAX_REG_8__SCAN_IN), .ZN(n4268) );
  XNOR2_X1 U4783 ( .A(n4265), .B(n5838), .ZN(n5841) );
  NAND2_X1 U4784 ( .A1(n5841), .A2(n5272), .ZN(n4267) );
  NAND2_X1 U4785 ( .A1(n4700), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4266)
         );
  NOR2_X2 U4786 ( .A1(n5088), .A2(n5121), .ZN(n5119) );
  INV_X1 U4787 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4270) );
  XNOR2_X1 U4788 ( .A(n4271), .B(n4270), .ZN(n7364) );
  INV_X1 U4789 ( .A(n7364), .ZN(n5896) );
  AOI22_X1 U4790 ( .A1(n4681), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4275) );
  AOI22_X1 U4791 ( .A1(n3936), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4519), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4274) );
  AOI22_X1 U4792 ( .A1(n4675), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3636), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4273) );
  AOI22_X1 U4793 ( .A1(n5133), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4272) );
  NAND4_X1 U4794 ( .A1(n4275), .A2(n4274), .A3(n4273), .A4(n4272), .ZN(n4281)
         );
  AOI22_X1 U4795 ( .A1(n3850), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4279) );
  AOI22_X1 U4796 ( .A1(n4553), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4278) );
  AOI22_X1 U4797 ( .A1(n4676), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U4798 ( .A1(n3637), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4276) );
  NAND4_X1 U4799 ( .A1(n4279), .A2(n4278), .A3(n4277), .A4(n4276), .ZN(n4280)
         );
  NOR2_X1 U4800 ( .A1(n4281), .A2(n4280), .ZN(n4284) );
  NAND2_X1 U4801 ( .A1(n4701), .A2(EAX_REG_12__SCAN_IN), .ZN(n4283) );
  NAND2_X1 U4802 ( .A1(n4700), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4282)
         );
  OAI211_X1 U4803 ( .C1(n4388), .C2(n4284), .A(n4283), .B(n4282), .ZN(n4285)
         );
  AOI21_X1 U4804 ( .B1(n5896), .B2(n5272), .A(n4285), .ZN(n5764) );
  INV_X1 U4805 ( .A(n5764), .ZN(n4300) );
  XOR2_X1 U4806 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n4286), .Z(n7350) );
  AOI22_X1 U4807 ( .A1(n3850), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4290) );
  AOI22_X1 U4808 ( .A1(n3936), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5133), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4289) );
  AOI22_X1 U4809 ( .A1(n4676), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4288) );
  AOI22_X1 U4810 ( .A1(n3636), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4287) );
  NAND4_X1 U4811 ( .A1(n4290), .A2(n4289), .A3(n4288), .A4(n4287), .ZN(n4296)
         );
  AOI22_X1 U4812 ( .A1(n4681), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4294) );
  AOI22_X1 U4813 ( .A1(n4674), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4293) );
  AOI22_X1 U4814 ( .A1(n4553), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4292) );
  AOI22_X1 U4815 ( .A1(n4675), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4291) );
  NAND4_X1 U4816 ( .A1(n4294), .A2(n4293), .A3(n4292), .A4(n4291), .ZN(n4295)
         );
  OR2_X1 U4817 ( .A1(n4296), .A2(n4295), .ZN(n4297) );
  AOI22_X1 U4818 ( .A1(n4346), .A2(n4297), .B1(n4700), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4299) );
  NAND2_X1 U4819 ( .A1(n4701), .A2(EAX_REG_11__SCAN_IN), .ZN(n4298) );
  OAI211_X1 U4820 ( .C1(n7350), .C2(n4220), .A(n4299), .B(n4298), .ZN(n5798)
         );
  AND2_X1 U4821 ( .A1(n4300), .A2(n5798), .ZN(n4318) );
  XNOR2_X1 U4822 ( .A(n4301), .B(n5821), .ZN(n5832) );
  NAND2_X1 U4823 ( .A1(n5832), .A2(n5272), .ZN(n4317) );
  AOI22_X1 U4824 ( .A1(n3850), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4305) );
  AOI22_X1 U4825 ( .A1(n4553), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4674), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4304) );
  AOI22_X1 U4826 ( .A1(n3936), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4303) );
  AOI22_X1 U4827 ( .A1(n3636), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4302) );
  NAND4_X1 U4828 ( .A1(n4305), .A2(n4304), .A3(n4303), .A4(n4302), .ZN(n4311)
         );
  AOI22_X1 U4829 ( .A1(n4681), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4309) );
  AOI22_X1 U4830 ( .A1(n4675), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5133), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4308) );
  AOI22_X1 U4831 ( .A1(n3634), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4307) );
  AOI22_X1 U4832 ( .A1(n4676), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4306) );
  NAND4_X1 U4833 ( .A1(n4309), .A2(n4308), .A3(n4307), .A4(n4306), .ZN(n4310)
         );
  NOR2_X1 U4834 ( .A1(n4311), .A2(n4310), .ZN(n4314) );
  NAND2_X1 U4835 ( .A1(n4232), .A2(EAX_REG_10__SCAN_IN), .ZN(n4313) );
  NAND2_X1 U4836 ( .A1(n4700), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4312)
         );
  OAI211_X1 U4837 ( .C1(n4388), .C2(n4314), .A(n4313), .B(n4312), .ZN(n4315)
         );
  INV_X1 U4838 ( .A(n4315), .ZN(n4316) );
  NAND2_X1 U4839 ( .A1(n4317), .A2(n4316), .ZN(n5514) );
  AND2_X1 U4840 ( .A1(n4318), .A2(n5514), .ZN(n4333) );
  XOR2_X1 U4841 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n4319), .Z(n7339) );
  AOI22_X1 U4842 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n4553), .B1(n3936), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4323) );
  AOI22_X1 U4843 ( .A1(n4674), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4322) );
  AOI22_X1 U4844 ( .A1(n4676), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4321) );
  AOI22_X1 U4845 ( .A1(n3636), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4320) );
  NAND4_X1 U4846 ( .A1(n4323), .A2(n4322), .A3(n4321), .A4(n4320), .ZN(n4329)
         );
  AOI22_X1 U4847 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n4635), .B1(n3850), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4327) );
  AOI22_X1 U4848 ( .A1(n4681), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4326) );
  AOI22_X1 U4849 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5133), .B1(n3938), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4325) );
  AOI22_X1 U4850 ( .A1(n4675), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4324) );
  NAND4_X1 U4851 ( .A1(n4327), .A2(n4326), .A3(n4325), .A4(n4324), .ZN(n4328)
         );
  OR2_X1 U4852 ( .A1(n4329), .A2(n4328), .ZN(n4330) );
  AOI22_X1 U4853 ( .A1(n4346), .A2(n4330), .B1(n4700), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4332) );
  NAND2_X1 U4854 ( .A1(n4232), .A2(EAX_REG_9__SCAN_IN), .ZN(n4331) );
  OAI211_X1 U4855 ( .C1(n7339), .C2(n4220), .A(n4332), .B(n4331), .ZN(n5262)
         );
  AND2_X1 U4856 ( .A1(n4333), .A2(n5262), .ZN(n4334) );
  NAND2_X1 U4857 ( .A1(n5119), .A2(n4334), .ZN(n5761) );
  AOI22_X1 U4858 ( .A1(n3850), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4338) );
  AOI22_X1 U4859 ( .A1(n4674), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4337) );
  AOI22_X1 U4860 ( .A1(n4675), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3636), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4336) );
  AOI22_X1 U4861 ( .A1(n4553), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4335) );
  NAND4_X1 U4862 ( .A1(n4338), .A2(n4337), .A3(n4336), .A4(n4335), .ZN(n4344)
         );
  AOI22_X1 U4863 ( .A1(n4681), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4342) );
  AOI22_X1 U4864 ( .A1(n3936), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5133), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4341) );
  AOI22_X1 U4865 ( .A1(n4676), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4340) );
  AOI22_X1 U4866 ( .A1(n3637), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4339) );
  NAND4_X1 U4867 ( .A1(n4342), .A2(n4341), .A3(n4340), .A4(n4339), .ZN(n4343)
         );
  OR2_X1 U4868 ( .A1(n4344), .A2(n4343), .ZN(n4345) );
  AND2_X1 U4869 ( .A1(n4346), .A2(n4345), .ZN(n4351) );
  XNOR2_X2 U4870 ( .A(n5761), .B(n4351), .ZN(n5704) );
  NAND2_X1 U4871 ( .A1(n4701), .A2(EAX_REG_13__SCAN_IN), .ZN(n4350) );
  INV_X1 U4872 ( .A(n4347), .ZN(n4348) );
  XNOR2_X1 U4873 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n4348), .ZN(n5962)
         );
  AOI22_X1 U4874 ( .A1(n5272), .A2(n5962), .B1(n4700), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4349) );
  NAND2_X1 U4875 ( .A1(n4350), .A2(n4349), .ZN(n5706) );
  NAND2_X1 U4876 ( .A1(n5704), .A2(n5706), .ZN(n4357) );
  INV_X1 U4877 ( .A(n4351), .ZN(n4352) );
  NOR2_X1 U4878 ( .A1(n5764), .A2(n4352), .ZN(n4353) );
  AND2_X1 U4879 ( .A1(n4353), .A2(n5798), .ZN(n4354) );
  AND2_X1 U4880 ( .A1(n4354), .A2(n5514), .ZN(n4355) );
  NAND2_X1 U4881 ( .A1(n4357), .A2(n4356), .ZN(n5753) );
  AOI22_X1 U4882 ( .A1(n3850), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4361) );
  AOI22_X1 U4883 ( .A1(n4674), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4360) );
  AOI22_X1 U4884 ( .A1(n4553), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4359) );
  AOI22_X1 U4885 ( .A1(n3636), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4358) );
  NAND4_X1 U4886 ( .A1(n4361), .A2(n4360), .A3(n4359), .A4(n4358), .ZN(n4367)
         );
  AOI22_X1 U4887 ( .A1(n4681), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4365) );
  AOI22_X1 U4888 ( .A1(n3936), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5133), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4364) );
  AOI22_X1 U4889 ( .A1(n4675), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4363) );
  AOI22_X1 U4890 ( .A1(n4676), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4362) );
  NAND4_X1 U4891 ( .A1(n4365), .A2(n4364), .A3(n4363), .A4(n4362), .ZN(n4366)
         );
  NOR2_X1 U4892 ( .A1(n4367), .A2(n4366), .ZN(n4373) );
  INV_X1 U4893 ( .A(n4368), .ZN(n4369) );
  XNOR2_X1 U4894 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4369), .ZN(n7377)
         );
  INV_X1 U4895 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5976) );
  OAI22_X1 U4896 ( .A1(n7377), .A2(n4220), .B1(n4403), .B2(n5976), .ZN(n4370)
         );
  INV_X1 U4897 ( .A(n4370), .ZN(n4372) );
  NAND2_X1 U4898 ( .A1(n4701), .A2(EAX_REG_14__SCAN_IN), .ZN(n4371) );
  OAI211_X1 U4899 ( .C1(n4388), .C2(n4373), .A(n4372), .B(n4371), .ZN(n5752)
         );
  NAND2_X1 U4900 ( .A1(n5753), .A2(n5752), .ZN(n5754) );
  XOR2_X1 U4901 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4374), .Z(n6008) );
  INV_X1 U4902 ( .A(n6008), .ZN(n5865) );
  AOI22_X1 U4903 ( .A1(n3850), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4378) );
  AOI22_X1 U4904 ( .A1(n4681), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4377) );
  AOI22_X1 U4905 ( .A1(n4676), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4675), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4376) );
  AOI22_X1 U4906 ( .A1(n4674), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4375) );
  NAND4_X1 U4907 ( .A1(n4378), .A2(n4377), .A3(n4376), .A4(n4375), .ZN(n4384)
         );
  AOI22_X1 U4908 ( .A1(n4553), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4382) );
  AOI22_X1 U4909 ( .A1(n3936), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5133), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4381) );
  AOI22_X1 U4910 ( .A1(n3636), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4380) );
  AOI22_X1 U4911 ( .A1(n3637), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4379) );
  NAND4_X1 U4912 ( .A1(n4382), .A2(n4381), .A3(n4380), .A4(n4379), .ZN(n4383)
         );
  NOR2_X1 U4913 ( .A1(n4384), .A2(n4383), .ZN(n4387) );
  NAND2_X1 U4914 ( .A1(n4701), .A2(EAX_REG_15__SCAN_IN), .ZN(n4386) );
  NAND2_X1 U4915 ( .A1(n4700), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4385)
         );
  OAI211_X1 U4916 ( .C1(n4388), .C2(n4387), .A(n4386), .B(n4385), .ZN(n4389)
         );
  AOI21_X1 U4917 ( .B1(n5865), .B2(n5272), .A(n4389), .ZN(n5814) );
  NAND2_X1 U4918 ( .A1(n4391), .A2(n4390), .ZN(n5812) );
  XNOR2_X1 U4919 ( .A(n4392), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n7388)
         );
  AOI22_X1 U4920 ( .A1(n4681), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4396) );
  AOI22_X1 U4921 ( .A1(n3936), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4674), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4395) );
  AOI22_X1 U4922 ( .A1(n5133), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4394) );
  AOI22_X1 U4923 ( .A1(n4675), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4393) );
  NAND4_X1 U4924 ( .A1(n4396), .A2(n4395), .A3(n4394), .A4(n4393), .ZN(n4402)
         );
  AOI22_X1 U4925 ( .A1(n3850), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4400) );
  AOI22_X1 U4926 ( .A1(n4553), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4399) );
  AOI22_X1 U4927 ( .A1(n4676), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4398) );
  AOI22_X1 U4928 ( .A1(n3636), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4397) );
  NAND4_X1 U4929 ( .A1(n4400), .A2(n4399), .A3(n4398), .A4(n4397), .ZN(n4401)
         );
  OR2_X1 U4930 ( .A1(n4402), .A2(n4401), .ZN(n4405) );
  INV_X1 U4931 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5223) );
  OAI22_X1 U4932 ( .A1(n4647), .A2(n5223), .B1(n4403), .B2(n6018), .ZN(n4404)
         );
  AOI21_X1 U4933 ( .B1(n4645), .B2(n4405), .A(n4404), .ZN(n4406) );
  OAI21_X1 U4934 ( .B1(n7388), .B2(n4220), .A(n4406), .ZN(n5878) );
  INV_X1 U4935 ( .A(n5878), .ZN(n4407) );
  NOR2_X2 U4936 ( .A1(n5812), .A2(n4407), .ZN(n5875) );
  AOI22_X1 U4937 ( .A1(n3850), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U4938 ( .A1(n4681), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4410) );
  AOI22_X1 U4939 ( .A1(n4674), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4409) );
  AOI22_X1 U4940 ( .A1(n3936), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4408) );
  NAND4_X1 U4941 ( .A1(n4411), .A2(n4410), .A3(n4409), .A4(n4408), .ZN(n4417)
         );
  AOI22_X1 U4942 ( .A1(n4676), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4675), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4415) );
  AOI22_X1 U4943 ( .A1(n4553), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4414) );
  AOI22_X1 U4944 ( .A1(n3636), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4413) );
  AOI22_X1 U4945 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n5133), .B1(n4683), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4412) );
  NAND4_X1 U4946 ( .A1(n4415), .A2(n4414), .A3(n4413), .A4(n4412), .ZN(n4416)
         );
  NOR2_X1 U4947 ( .A1(n4417), .A2(n4416), .ZN(n4418) );
  OR2_X1 U4948 ( .A1(n4693), .A2(n4418), .ZN(n4428) );
  OAI21_X1 U4949 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n7520), .A(n7188), 
        .ZN(n4419) );
  INV_X1 U4950 ( .A(n4419), .ZN(n4420) );
  AOI21_X1 U4951 ( .B1(n4232), .B2(EAX_REG_17__SCAN_IN), .A(n4420), .ZN(n4427)
         );
  INV_X1 U4952 ( .A(n4444), .ZN(n4425) );
  INV_X1 U4953 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4423) );
  INV_X1 U4954 ( .A(n4421), .ZN(n4422) );
  NAND2_X1 U4955 ( .A1(n4423), .A2(n4422), .ZN(n4424) );
  NAND2_X1 U4956 ( .A1(n4425), .A2(n4424), .ZN(n7401) );
  NOR2_X1 U4957 ( .A1(n7401), .A2(n4220), .ZN(n4426) );
  AOI21_X1 U4958 ( .B1(n4428), .B2(n4427), .A(n4426), .ZN(n7109) );
  NAND2_X1 U4959 ( .A1(n5875), .A2(n7109), .ZN(n5983) );
  AOI22_X1 U4960 ( .A1(n4674), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4432) );
  AOI22_X1 U4961 ( .A1(n3936), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4431) );
  AOI22_X1 U4962 ( .A1(n4553), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3636), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4430) );
  AOI22_X1 U4963 ( .A1(n4676), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4429) );
  NAND4_X1 U4964 ( .A1(n4432), .A2(n4431), .A3(n4430), .A4(n4429), .ZN(n4441)
         );
  AOI22_X1 U4965 ( .A1(n3850), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n5133), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4439) );
  NAND2_X1 U4966 ( .A1(n4433), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4435)
         );
  NAND2_X1 U4967 ( .A1(n3638), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4434) );
  AND3_X1 U4968 ( .A1(n4435), .A2(n4220), .A3(n4434), .ZN(n4438) );
  AOI22_X1 U4969 ( .A1(n4675), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4437) );
  AOI22_X1 U4970 ( .A1(n3637), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4436) );
  NAND4_X1 U4971 ( .A1(n4439), .A2(n4438), .A3(n4437), .A4(n4436), .ZN(n4440)
         );
  NAND2_X1 U4972 ( .A1(n4693), .A2(n4220), .ZN(n4511) );
  OAI21_X1 U4973 ( .B1(n4441), .B2(n4440), .A(n4511), .ZN(n4443) );
  AOI22_X1 U4974 ( .A1(n4701), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n7188), .ZN(n4442) );
  NAND2_X1 U4975 ( .A1(n4443), .A2(n4442), .ZN(n4446) );
  INV_X1 U4976 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6790) );
  XNOR2_X1 U4977 ( .A(n4444), .B(n6790), .ZN(n6793) );
  NAND2_X1 U4978 ( .A1(n6793), .A2(n5272), .ZN(n4445) );
  NAND2_X1 U4979 ( .A1(n4446), .A2(n4445), .ZN(n5985) );
  NOR2_X2 U4980 ( .A1(n5983), .A2(n5985), .ZN(n5986) );
  AOI22_X1 U4981 ( .A1(n3850), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4450) );
  AOI22_X1 U4982 ( .A1(n4681), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4449) );
  AOI22_X1 U4983 ( .A1(n3936), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5133), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4448) );
  AOI22_X1 U4984 ( .A1(n4676), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4447) );
  NAND4_X1 U4985 ( .A1(n4450), .A2(n4449), .A3(n4448), .A4(n4447), .ZN(n4456)
         );
  AOI22_X1 U4986 ( .A1(n4674), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4454) );
  AOI22_X1 U4987 ( .A1(n4553), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4453) );
  AOI22_X1 U4988 ( .A1(n3636), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4452) );
  AOI22_X1 U4989 ( .A1(n4675), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4451) );
  NAND4_X1 U4990 ( .A1(n4454), .A2(n4453), .A3(n4452), .A4(n4451), .ZN(n4455)
         );
  NOR2_X1 U4991 ( .A1(n4456), .A2(n4455), .ZN(n4460) );
  OAI21_X1 U4992 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n7520), .A(n7188), 
        .ZN(n4457) );
  INV_X1 U4993 ( .A(n4457), .ZN(n4458) );
  AOI21_X1 U4994 ( .B1(n4232), .B2(EAX_REG_19__SCAN_IN), .A(n4458), .ZN(n4459)
         );
  OAI21_X1 U4995 ( .B1(n4693), .B2(n4460), .A(n4459), .ZN(n4464) );
  AND2_X1 U4996 ( .A1(n4461), .A2(n6780), .ZN(n4462) );
  OR2_X1 U4997 ( .A1(n4462), .A2(n4478), .ZN(n7415) );
  INV_X1 U4998 ( .A(n7415), .ZN(n6782) );
  NAND2_X1 U4999 ( .A1(n6782), .A2(n5272), .ZN(n4463) );
  AND2_X2 U5000 ( .A1(n5986), .A2(n3662), .ZN(n6643) );
  AOI22_X1 U5001 ( .A1(n4681), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5133), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4470) );
  AOI22_X1 U5002 ( .A1(n4553), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4675), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4469) );
  NAND2_X1 U5003 ( .A1(n4635), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4466)
         );
  NAND2_X1 U5004 ( .A1(n3638), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4465) );
  AND3_X1 U5005 ( .A1(n4466), .A2(n4220), .A3(n4465), .ZN(n4468) );
  AOI22_X1 U5006 ( .A1(n3637), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4467) );
  NAND4_X1 U5007 ( .A1(n4470), .A2(n4469), .A3(n4468), .A4(n4467), .ZN(n4476)
         );
  AOI22_X1 U5008 ( .A1(n3850), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4674), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4474) );
  AOI22_X1 U5009 ( .A1(n3936), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3636), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4473) );
  AOI22_X1 U5010 ( .A1(n4676), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4472) );
  AOI22_X1 U5011 ( .A1(n4682), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4471) );
  NAND4_X1 U5012 ( .A1(n4474), .A2(n4473), .A3(n4472), .A4(n4471), .ZN(n4475)
         );
  OR2_X1 U5013 ( .A1(n4476), .A2(n4475), .ZN(n4477) );
  NAND2_X1 U5014 ( .A1(n4511), .A2(n4477), .ZN(n4481) );
  AOI22_X1 U5015 ( .A1(n4701), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n7188), .ZN(n4480) );
  INV_X1 U5016 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n7430) );
  XNOR2_X1 U5017 ( .A(n4478), .B(n7430), .ZN(n7426) );
  AND2_X1 U5018 ( .A1(n7426), .A2(n5272), .ZN(n4479) );
  AOI21_X1 U5019 ( .B1(n4481), .B2(n4480), .A(n4479), .ZN(n6642) );
  AOI22_X1 U5020 ( .A1(n4681), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4553), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4485) );
  AOI22_X1 U5021 ( .A1(n3850), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4484) );
  AOI22_X1 U5022 ( .A1(n4676), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4483) );
  AOI22_X1 U5023 ( .A1(n3636), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4482) );
  NAND4_X1 U5024 ( .A1(n4485), .A2(n4484), .A3(n4483), .A4(n4482), .ZN(n4491)
         );
  AOI22_X1 U5025 ( .A1(n3634), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4489) );
  AOI22_X1 U5026 ( .A1(n3936), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4674), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4488) );
  AOI22_X1 U5027 ( .A1(n5133), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4487) );
  AOI22_X1 U5028 ( .A1(n4675), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4486) );
  NAND4_X1 U5029 ( .A1(n4489), .A2(n4488), .A3(n4487), .A4(n4486), .ZN(n4490)
         );
  NOR2_X1 U5030 ( .A1(n4491), .A2(n4490), .ZN(n4492) );
  OR2_X1 U5031 ( .A1(n4693), .A2(n4492), .ZN(n4500) );
  NAND2_X1 U5032 ( .A1(n7188), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4493)
         );
  NAND2_X1 U5033 ( .A1(n4220), .A2(n4493), .ZN(n4494) );
  AOI21_X1 U5034 ( .B1(n4232), .B2(EAX_REG_21__SCAN_IN), .A(n4494), .ZN(n4499)
         );
  NAND2_X1 U5035 ( .A1(n4496), .A2(n4495), .ZN(n4497) );
  NAND2_X1 U5036 ( .A1(n4516), .A2(n4497), .ZN(n7446) );
  NOR2_X1 U5037 ( .A1(n7446), .A2(n4220), .ZN(n4498) );
  AOI21_X1 U5038 ( .B1(n4500), .B2(n4499), .A(n4498), .ZN(n6761) );
  AOI22_X1 U5039 ( .A1(n4681), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4504) );
  AOI22_X1 U5040 ( .A1(n4635), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4503) );
  AOI22_X1 U5041 ( .A1(n3936), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4502) );
  AOI22_X1 U5042 ( .A1(n5133), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4501) );
  NAND4_X1 U5043 ( .A1(n4504), .A2(n4503), .A3(n4502), .A4(n4501), .ZN(n4513)
         );
  AOI22_X1 U5044 ( .A1(n3850), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4510) );
  AOI22_X1 U5045 ( .A1(n3634), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4675), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4509) );
  AOI22_X1 U5046 ( .A1(n4676), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4674), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4508) );
  NAND2_X1 U5047 ( .A1(n4553), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4506)
         );
  NAND2_X1 U5048 ( .A1(n3636), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4505) );
  AND3_X1 U5049 ( .A1(n4506), .A2(n4505), .A3(n4220), .ZN(n4507) );
  NAND4_X1 U5050 ( .A1(n4510), .A2(n4509), .A3(n4508), .A4(n4507), .ZN(n4512)
         );
  OAI21_X1 U5051 ( .B1(n4513), .B2(n4512), .A(n4511), .ZN(n4515) );
  AOI22_X1 U5052 ( .A1(n4701), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n7188), .ZN(n4514) );
  NAND2_X1 U5053 ( .A1(n4515), .A2(n4514), .ZN(n4518) );
  XNOR2_X1 U5054 ( .A(n4516), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6757)
         );
  NAND2_X1 U5055 ( .A1(n6757), .A2(n5272), .ZN(n4517) );
  NAND2_X1 U5056 ( .A1(n4518), .A2(n4517), .ZN(n6587) );
  NOR2_X2 U5057 ( .A1(n6586), .A2(n6587), .ZN(n6571) );
  AOI22_X1 U5058 ( .A1(n3850), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4523) );
  AOI22_X1 U5059 ( .A1(n4636), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4522) );
  AOI22_X1 U5060 ( .A1(n4553), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3936), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4521) );
  AOI22_X1 U5061 ( .A1(n4674), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4520) );
  NAND4_X1 U5062 ( .A1(n4523), .A2(n4522), .A3(n4521), .A4(n4520), .ZN(n4529)
         );
  AOI22_X1 U5063 ( .A1(n4676), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3636), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4527) );
  AOI22_X1 U5064 ( .A1(n5133), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4526) );
  AOI22_X1 U5065 ( .A1(n4675), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4525) );
  AOI22_X1 U5066 ( .A1(n3637), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4524) );
  NAND4_X1 U5067 ( .A1(n4527), .A2(n4526), .A3(n4525), .A4(n4524), .ZN(n4528)
         );
  OR2_X1 U5068 ( .A1(n4529), .A2(n4528), .ZN(n4541) );
  AOI22_X1 U5069 ( .A1(n3850), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4533) );
  AOI22_X1 U5070 ( .A1(n4636), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4532) );
  AOI22_X1 U5071 ( .A1(n4553), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3936), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4531) );
  AOI22_X1 U5072 ( .A1(n4674), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4530) );
  NAND4_X1 U5073 ( .A1(n4533), .A2(n4532), .A3(n4531), .A4(n4530), .ZN(n4539)
         );
  AOI22_X1 U5074 ( .A1(n4676), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3636), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4537) );
  AOI22_X1 U5075 ( .A1(n5133), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4536) );
  AOI22_X1 U5076 ( .A1(n4675), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4535) );
  AOI22_X1 U5077 ( .A1(n3637), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4534) );
  NAND4_X1 U5078 ( .A1(n4537), .A2(n4536), .A3(n4535), .A4(n4534), .ZN(n4538)
         );
  OR2_X1 U5079 ( .A1(n4539), .A2(n4538), .ZN(n4540) );
  NAND2_X1 U5080 ( .A1(n4540), .A2(n4541), .ZN(n4577) );
  OAI21_X1 U5081 ( .B1(n4541), .B2(n4540), .A(n4577), .ZN(n4545) );
  NAND2_X1 U5082 ( .A1(n7188), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4542)
         );
  NAND2_X1 U5083 ( .A1(n4220), .A2(n4542), .ZN(n4543) );
  AOI21_X1 U5084 ( .B1(n4232), .B2(EAX_REG_23__SCAN_IN), .A(n4543), .ZN(n4544)
         );
  OAI21_X1 U5085 ( .B1(n4693), .B2(n4545), .A(n4544), .ZN(n4550) );
  NAND2_X1 U5086 ( .A1(n4547), .A2(n4546), .ZN(n4548) );
  AND2_X1 U5087 ( .A1(n4552), .A2(n4548), .ZN(n6745) );
  NAND2_X1 U5088 ( .A1(n6745), .A2(n5272), .ZN(n4549) );
  NAND2_X1 U5089 ( .A1(n4550), .A2(n4549), .ZN(n6574) );
  AND2_X2 U5090 ( .A1(n6571), .A2(n4551), .ZN(n6559) );
  XNOR2_X1 U5091 ( .A(n4552), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6736)
         );
  AOI22_X1 U5092 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n4682), .B1(n4635), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4557) );
  AOI22_X1 U5093 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4553), .B1(n4675), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4556) );
  AOI22_X1 U5094 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4676), .B1(n3636), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4555) );
  AOI22_X1 U5095 ( .A1(n3637), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4554) );
  NAND4_X1 U5096 ( .A1(n4557), .A2(n4556), .A3(n4555), .A4(n4554), .ZN(n4563)
         );
  AOI22_X1 U5097 ( .A1(n4636), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3850), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4561) );
  AOI22_X1 U5098 ( .A1(n4674), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4560) );
  AOI22_X1 U5099 ( .A1(n3936), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4559) );
  AOI22_X1 U5100 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n5133), .B1(n4683), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4558) );
  NAND4_X1 U5101 ( .A1(n4561), .A2(n4560), .A3(n4559), .A4(n4558), .ZN(n4562)
         );
  NOR2_X1 U5102 ( .A1(n4563), .A2(n4562), .ZN(n4578) );
  XNOR2_X1 U5103 ( .A(n4577), .B(n4578), .ZN(n4564) );
  OR2_X1 U5104 ( .A1(n4693), .A2(n4564), .ZN(n4566) );
  AOI22_X1 U5105 ( .A1(n4701), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n4700), .ZN(n4565) );
  OAI211_X1 U5106 ( .C1(n6736), .C2(n4220), .A(n4566), .B(n4565), .ZN(n6560)
         );
  AOI22_X1 U5107 ( .A1(n3850), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4570) );
  AOI22_X1 U5108 ( .A1(n4636), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4569) );
  AOI22_X1 U5109 ( .A1(n4553), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3936), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5110 ( .A1(n4674), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4567) );
  NAND4_X1 U5111 ( .A1(n4570), .A2(n4569), .A3(n4568), .A4(n4567), .ZN(n4576)
         );
  AOI22_X1 U5112 ( .A1(n4676), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3636), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4574) );
  AOI22_X1 U5113 ( .A1(n5133), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4573) );
  AOI22_X1 U5114 ( .A1(n4675), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4572) );
  AOI22_X1 U5115 ( .A1(n3637), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4571) );
  NAND4_X1 U5116 ( .A1(n4574), .A2(n4573), .A3(n4572), .A4(n4571), .ZN(n4575)
         );
  OR2_X1 U5117 ( .A1(n4576), .A2(n4575), .ZN(n4587) );
  NOR2_X1 U5118 ( .A1(n4578), .A2(n4577), .ZN(n4588) );
  XNOR2_X1 U5119 ( .A(n4587), .B(n4588), .ZN(n4582) );
  NAND2_X1 U5120 ( .A1(n7188), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4579)
         );
  NAND2_X1 U5121 ( .A1(n4220), .A2(n4579), .ZN(n4580) );
  AOI21_X1 U5122 ( .B1(n4232), .B2(EAX_REG_25__SCAN_IN), .A(n4580), .ZN(n4581)
         );
  OAI21_X1 U5123 ( .B1(n4693), .B2(n4582), .A(n4581), .ZN(n4586) );
  NAND2_X1 U5124 ( .A1(n4583), .A2(n6548), .ZN(n4584) );
  NAND2_X1 U5125 ( .A1(n4604), .A2(n4584), .ZN(n6716) );
  NAND2_X1 U5126 ( .A1(n4586), .A2(n4585), .ZN(n6542) );
  NAND2_X1 U5127 ( .A1(n4588), .A2(n4587), .ZN(n4608) );
  AOI22_X1 U5128 ( .A1(n3850), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4592) );
  AOI22_X1 U5129 ( .A1(n4553), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3936), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4591) );
  AOI22_X1 U5130 ( .A1(n4636), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4590) );
  AOI22_X1 U5131 ( .A1(n5133), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4589) );
  NAND4_X1 U5132 ( .A1(n4592), .A2(n4591), .A3(n4590), .A4(n4589), .ZN(n4598)
         );
  AOI22_X1 U5133 ( .A1(n4674), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4596) );
  AOI22_X1 U5134 ( .A1(n4676), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4675), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4595) );
  AOI22_X1 U5135 ( .A1(n4683), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4594) );
  AOI22_X1 U5136 ( .A1(n3636), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4593) );
  NAND4_X1 U5137 ( .A1(n4596), .A2(n4595), .A3(n4594), .A4(n4593), .ZN(n4597)
         );
  NOR2_X1 U5138 ( .A1(n4598), .A2(n4597), .ZN(n4609) );
  XOR2_X1 U5139 ( .A(n4608), .B(n4609), .Z(n4599) );
  NAND2_X1 U5140 ( .A1(n4599), .A2(n4645), .ZN(n4603) );
  NAND2_X1 U5141 ( .A1(n7188), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4600)
         );
  NAND2_X1 U5142 ( .A1(n4220), .A2(n4600), .ZN(n4601) );
  AOI21_X1 U5143 ( .B1(n4232), .B2(EAX_REG_26__SCAN_IN), .A(n4601), .ZN(n4602)
         );
  NAND2_X1 U5144 ( .A1(n4603), .A2(n4602), .ZN(n4606) );
  XNOR2_X1 U5145 ( .A(n4604), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6530)
         );
  NAND2_X1 U5146 ( .A1(n6530), .A2(n5272), .ZN(n4605) );
  NAND2_X1 U5147 ( .A1(n4606), .A2(n4605), .ZN(n6529) );
  NOR2_X1 U5148 ( .A1(n4609), .A2(n4608), .ZN(n4644) );
  AOI22_X1 U5149 ( .A1(n3850), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4613) );
  AOI22_X1 U5150 ( .A1(n4636), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4612) );
  AOI22_X1 U5151 ( .A1(n4553), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3936), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4611) );
  AOI22_X1 U5152 ( .A1(n4674), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4610) );
  NAND4_X1 U5153 ( .A1(n4613), .A2(n4612), .A3(n4611), .A4(n4610), .ZN(n4619)
         );
  AOI22_X1 U5154 ( .A1(n4676), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3636), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4617) );
  AOI22_X1 U5155 ( .A1(n5133), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4616) );
  AOI22_X1 U5156 ( .A1(n4675), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4615) );
  AOI22_X1 U5157 ( .A1(n3637), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4614) );
  NAND4_X1 U5158 ( .A1(n4617), .A2(n4616), .A3(n4615), .A4(n4614), .ZN(n4618)
         );
  OR2_X1 U5159 ( .A1(n4619), .A2(n4618), .ZN(n4643) );
  INV_X1 U5160 ( .A(n4643), .ZN(n4620) );
  XNOR2_X1 U5161 ( .A(n4644), .B(n4620), .ZN(n4624) );
  INV_X1 U5162 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4622) );
  NAND2_X1 U5163 ( .A1(n7188), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4621)
         );
  OAI211_X1 U5164 ( .C1(n4647), .C2(n4622), .A(n4220), .B(n4621), .ZN(n4623)
         );
  AOI21_X1 U5165 ( .B1(n4624), .B2(n4645), .A(n4623), .ZN(n4629) );
  INV_X1 U5166 ( .A(n4625), .ZN(n4626) );
  INV_X1 U5167 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6513) );
  NAND2_X1 U5168 ( .A1(n4626), .A2(n6513), .ZN(n4627) );
  NAND2_X1 U5169 ( .A1(n4649), .A2(n4627), .ZN(n6703) );
  NOR2_X1 U5170 ( .A1(n6703), .A2(n4220), .ZN(n4628) );
  AOI22_X1 U5171 ( .A1(n3634), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4634) );
  AOI22_X1 U5172 ( .A1(n4675), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3636), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4633) );
  AOI22_X1 U5173 ( .A1(n4674), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4632) );
  AOI22_X1 U5174 ( .A1(n3637), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4631) );
  NAND4_X1 U5175 ( .A1(n4634), .A2(n4633), .A3(n4632), .A4(n4631), .ZN(n4642)
         );
  AOI22_X1 U5176 ( .A1(n3850), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4640) );
  AOI22_X1 U5177 ( .A1(n4636), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4553), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4639) );
  AOI22_X1 U5178 ( .A1(n3936), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5133), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4638) );
  AOI22_X1 U5179 ( .A1(n4676), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4637) );
  NAND4_X1 U5180 ( .A1(n4640), .A2(n4639), .A3(n4638), .A4(n4637), .ZN(n4641)
         );
  NOR2_X1 U5181 ( .A1(n4642), .A2(n4641), .ZN(n4653) );
  NAND2_X1 U5182 ( .A1(n4644), .A2(n4643), .ZN(n4652) );
  XOR2_X1 U5183 ( .A(n4653), .B(n4652), .Z(n4646) );
  NAND2_X1 U5184 ( .A1(n4646), .A2(n4645), .ZN(n4651) );
  AOI21_X1 U5185 ( .B1(n6503), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4648) );
  AOI21_X1 U5186 ( .B1(n4232), .B2(EAX_REG_28__SCAN_IN), .A(n4648), .ZN(n4650)
         );
  XNOR2_X1 U5187 ( .A(n4649), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6502)
         );
  AOI22_X1 U5188 ( .A1(n4651), .A2(n4650), .B1(n5272), .B2(n6502), .ZN(n6501)
         );
  NOR2_X1 U5189 ( .A1(n4653), .A2(n4652), .ZN(n4672) );
  AOI22_X1 U5190 ( .A1(n4681), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4553), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4657) );
  AOI22_X1 U5191 ( .A1(n3936), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5133), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4656) );
  AOI22_X1 U5192 ( .A1(n4676), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3636), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4655) );
  AOI22_X1 U5193 ( .A1(n4675), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4683), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4654) );
  NAND4_X1 U5194 ( .A1(n4657), .A2(n4656), .A3(n4655), .A4(n4654), .ZN(n4663)
         );
  AOI22_X1 U5195 ( .A1(n3850), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4661) );
  AOI22_X1 U5196 ( .A1(n3634), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4682), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4660) );
  AOI22_X1 U5197 ( .A1(n4674), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4659) );
  AOI22_X1 U5198 ( .A1(n3637), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4658) );
  NAND4_X1 U5199 ( .A1(n4661), .A2(n4660), .A3(n4659), .A4(n4658), .ZN(n4662)
         );
  OR2_X1 U5200 ( .A1(n4663), .A2(n4662), .ZN(n4671) );
  XNOR2_X1 U5201 ( .A(n4672), .B(n4671), .ZN(n4664) );
  NOR2_X1 U5202 ( .A1(n4664), .A2(n4693), .ZN(n4670) );
  INV_X1 U5203 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4666) );
  NAND2_X1 U5204 ( .A1(n7188), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4665)
         );
  OAI211_X1 U5205 ( .C1(n4647), .C2(n4666), .A(n4220), .B(n4665), .ZN(n4669)
         );
  NAND2_X1 U5206 ( .A1(n4667), .A2(n6119), .ZN(n4668) );
  NAND2_X1 U5207 ( .A1(n4697), .A2(n4668), .ZN(n6686) );
  OAI22_X1 U5208 ( .A1(n4670), .A2(n4669), .B1(n6686), .B2(n4220), .ZN(n6115)
         );
  NAND2_X1 U5209 ( .A1(n4672), .A2(n4671), .ZN(n4690) );
  AOI22_X1 U5210 ( .A1(n3850), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4680) );
  AOI22_X1 U5211 ( .A1(n4674), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4553), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4679) );
  AOI22_X1 U5212 ( .A1(n3629), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3936), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4678) );
  AOI22_X1 U5213 ( .A1(n4676), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4675), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4677) );
  NAND4_X1 U5214 ( .A1(n4680), .A2(n4679), .A3(n4678), .A4(n4677), .ZN(n4689)
         );
  AOI22_X1 U5215 ( .A1(n4681), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4687) );
  AOI22_X1 U5216 ( .A1(n4682), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5133), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4686) );
  AOI22_X1 U5217 ( .A1(n4683), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3636), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4685) );
  AOI22_X1 U5218 ( .A1(n3638), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4684) );
  NAND4_X1 U5219 ( .A1(n4687), .A2(n4686), .A3(n4685), .A4(n4684), .ZN(n4688)
         );
  NOR2_X1 U5220 ( .A1(n4689), .A2(n4688), .ZN(n4691) );
  NAND2_X1 U5221 ( .A1(n4690), .A2(n4691), .ZN(n4695) );
  NOR2_X1 U5222 ( .A1(n4691), .A2(n4690), .ZN(n4692) );
  NOR2_X1 U5223 ( .A1(n4693), .A2(n4692), .ZN(n4694) );
  NAND2_X1 U5224 ( .A1(n4695), .A2(n4694), .ZN(n4699) );
  AOI21_X1 U5225 ( .B1(n6104), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4696) );
  AOI21_X1 U5226 ( .B1(n4232), .B2(EAX_REG_30__SCAN_IN), .A(n4696), .ZN(n4698)
         );
  XNOR2_X1 U5227 ( .A(n4697), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6033)
         );
  AOI22_X1 U5228 ( .A1(n4699), .A2(n4698), .B1(n5272), .B2(n6033), .ZN(n4910)
         );
  NAND2_X1 U5229 ( .A1(n6114), .A2(n4910), .ZN(n4704) );
  AOI22_X1 U5230 ( .A1(n4701), .A2(EAX_REG_31__SCAN_IN), .B1(n4700), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4702) );
  INV_X1 U5231 ( .A(n4702), .ZN(n4703) );
  XNOR2_X2 U5232 ( .A(n4704), .B(n4703), .ZN(n6087) );
  NOR2_X1 U5233 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7455), .ZN(n5709) );
  NAND2_X1 U5234 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n5709), .ZN(n7185) );
  INV_X1 U5235 ( .A(n7185), .ZN(n4705) );
  NAND2_X1 U5236 ( .A1(n7590), .A2(n4705), .ZN(n6797) );
  INV_X2 U5237 ( .A(n6797), .ZN(n7165) );
  NAND2_X1 U5238 ( .A1(n6087), .A2(n7165), .ZN(n4706) );
  OAI211_X1 U5239 ( .C1(n6053), .C2(n7447), .A(n4707), .B(n4706), .ZN(U2955)
         );
  INV_X1 U5240 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6802) );
  NOR2_X1 U5241 ( .A1(n4708), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4710)
         );
  NAND2_X1 U5242 ( .A1(n3643), .A2(n6751), .ZN(n4709) );
  INV_X1 U5243 ( .A(STATE_REG_0__SCAN_IN), .ZN(n7535) );
  NAND2_X1 U5244 ( .A1(n4712), .A2(n7535), .ZN(n7183) );
  INV_X1 U5245 ( .A(READY_N), .ZN(n7502) );
  NOR3_X1 U5246 ( .A1(n4715), .A2(n4714), .A3(n4713), .ZN(n4716) );
  OR2_X1 U5247 ( .A1(n4717), .A2(n4716), .ZN(n4719) );
  NAND2_X1 U5248 ( .A1(n4719), .A2(n4718), .ZN(n6098) );
  NAND2_X1 U5249 ( .A1(n7502), .A2(n6098), .ZN(n4983) );
  AOI21_X1 U5250 ( .B1(n3653), .B2(n7183), .A(n4983), .ZN(n4722) );
  NOR2_X1 U5251 ( .A1(n4868), .A2(n3650), .ZN(n4720) );
  NOR2_X1 U5252 ( .A1(n6097), .A2(n4720), .ZN(n4721) );
  MUX2_X1 U5253 ( .A(n4722), .B(n4721), .S(n5230), .Z(n4723) );
  INV_X1 U5254 ( .A(n4723), .ZN(n4733) );
  INV_X1 U5255 ( .A(n7183), .ZN(n4939) );
  OR2_X1 U5256 ( .A1(n3653), .A2(n4939), .ZN(n5715) );
  NAND2_X1 U5257 ( .A1(n5715), .A2(n7502), .ZN(n4724) );
  OR2_X1 U5258 ( .A1(n6097), .A2(n4724), .ZN(n4989) );
  NOR2_X1 U5259 ( .A1(n3838), .A2(n4726), .ZN(n4875) );
  NAND2_X1 U5260 ( .A1(n3816), .A2(n4743), .ZN(n4727) );
  MUX2_X1 U5261 ( .A(n4728), .B(n4727), .S(n5063), .Z(n4872) );
  AOI21_X1 U5262 ( .B1(n4872), .B2(n3664), .A(n4729), .ZN(n4986) );
  AOI21_X1 U5263 ( .B1(n6097), .B2(n4875), .A(n4986), .ZN(n4730) );
  OAI21_X1 U5264 ( .B1(n4989), .B2(n4990), .A(n4730), .ZN(n4731) );
  INV_X1 U5265 ( .A(n4731), .ZN(n4732) );
  NAND2_X1 U5266 ( .A1(n4733), .A2(n4732), .ZN(n4734) );
  NAND2_X1 U5267 ( .A1(n3664), .A2(n5735), .ZN(n5135) );
  NAND2_X1 U5268 ( .A1(n5135), .A2(n4735), .ZN(n6091) );
  AND2_X4 U5269 ( .A1(n3653), .A2(n4743), .ZN(n4966) );
  NAND2_X1 U5270 ( .A1(n4725), .A2(n4966), .ZN(n4736) );
  OAI211_X1 U5271 ( .C1(n5225), .C2(n4739), .A(n7460), .B(n4736), .ZN(n4737)
         );
  NOR2_X1 U5272 ( .A1(n6091), .A2(n4737), .ZN(n4738) );
  NAND2_X1 U5273 ( .A1(n4725), .A2(n3915), .ZN(n7496) );
  INV_X1 U5274 ( .A(n4739), .ZN(n4740) );
  NAND2_X1 U5275 ( .A1(n4740), .A2(n5225), .ZN(n4741) );
  AND2_X1 U5276 ( .A1(n7496), .A2(n4741), .ZN(n4742) );
  INV_X2 U5277 ( .A(n7212), .ZN(n7269) );
  NAND2_X1 U5278 ( .A1(n3837), .A2(n4743), .ZN(n4764) );
  OAI22_X1 U5279 ( .A1(n6023), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n6022), .ZN(n6024) );
  INV_X1 U5280 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4746) );
  NAND2_X1 U5281 ( .A1(n4966), .A2(n4746), .ZN(n4745) );
  NAND2_X1 U5282 ( .A1(n4764), .A2(n5014), .ZN(n4744) );
  NAND3_X1 U5283 ( .A1(n4745), .A2(n4744), .A3(n3656), .ZN(n4748) );
  NAND2_X1 U5284 ( .A1(n4781), .A2(n4746), .ZN(n4747) );
  NAND2_X1 U5285 ( .A1(n4748), .A2(n4747), .ZN(n4750) );
  NAND2_X1 U5286 ( .A1(n4764), .A2(EBX_REG_0__SCAN_IN), .ZN(n4749) );
  OAI21_X1 U5287 ( .B1(n4781), .B2(EBX_REG_0__SCAN_IN), .A(n4749), .ZN(n4935)
         );
  XNOR2_X1 U5288 ( .A(n4750), .B(n4935), .ZN(n4967) );
  INV_X1 U5289 ( .A(n4750), .ZN(n4751) );
  NAND2_X1 U5290 ( .A1(n4751), .A2(n4935), .ZN(n4752) );
  NAND2_X1 U5291 ( .A1(n4965), .A2(n4752), .ZN(n4963) );
  MUX2_X1 U5292 ( .A(n4854), .B(n3655), .S(EBX_REG_3__SCAN_IN), .Z(n4755) );
  NOR2_X1 U5293 ( .A1(n6023), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4754)
         );
  NOR2_X2 U5294 ( .A1(n4755), .A2(n4754), .ZN(n5033) );
  OAI21_X1 U5295 ( .B1(n3655), .B2(n7234), .A(n4858), .ZN(n4757) );
  INV_X1 U5296 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4758) );
  NAND2_X1 U5297 ( .A1(n4966), .A2(n4758), .ZN(n4756) );
  NAND2_X1 U5298 ( .A1(n4757), .A2(n4756), .ZN(n4760) );
  NAND2_X1 U5299 ( .A1(n3655), .A2(n4758), .ZN(n4759) );
  NAND2_X1 U5300 ( .A1(n4760), .A2(n4759), .ZN(n5034) );
  NAND2_X1 U5301 ( .A1(n5033), .A2(n5034), .ZN(n4761) );
  OR2_X2 U5302 ( .A1(n4963), .A2(n4761), .ZN(n7123) );
  INV_X1 U5303 ( .A(EBX_REG_5__SCAN_IN), .ZN(n5045) );
  MUX2_X1 U5304 ( .A(n3655), .B(n4854), .S(n5045), .Z(n4763) );
  NOR2_X1 U5305 ( .A1(n6023), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4762)
         );
  NOR2_X1 U5306 ( .A1(n4763), .A2(n4762), .ZN(n5041) );
  INV_X1 U5307 ( .A(n4764), .ZN(n4827) );
  NAND2_X1 U5308 ( .A1(n4858), .A2(n4765), .ZN(n4767) );
  INV_X1 U5309 ( .A(EBX_REG_4__SCAN_IN), .ZN(n7297) );
  NAND2_X1 U5310 ( .A1(n4966), .A2(n7297), .ZN(n4766) );
  NAND3_X1 U5311 ( .A1(n4767), .A2(n3633), .A3(n4766), .ZN(n4769) );
  NAND2_X1 U5312 ( .A1(n3655), .A2(n7297), .ZN(n4768) );
  NAND2_X1 U5313 ( .A1(n4769), .A2(n4768), .ZN(n7122) );
  NAND2_X1 U5314 ( .A1(n5041), .A2(n7122), .ZN(n4770) );
  INV_X1 U5315 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4771) );
  NAND2_X1 U5316 ( .A1(n4858), .A2(n4771), .ZN(n4773) );
  INV_X1 U5317 ( .A(EBX_REG_6__SCAN_IN), .ZN(n7312) );
  NAND2_X1 U5318 ( .A1(n4966), .A2(n7312), .ZN(n4772) );
  NAND3_X1 U5319 ( .A1(n4773), .A2(n3633), .A3(n4772), .ZN(n4775) );
  NAND2_X1 U5320 ( .A1(n3655), .A2(n7312), .ZN(n4774) );
  NAND2_X1 U5321 ( .A1(n4775), .A2(n4774), .ZN(n5027) );
  INV_X1 U5322 ( .A(n4854), .ZN(n4861) );
  MUX2_X1 U5323 ( .A(n4861), .B(n3633), .S(EBX_REG_7__SCAN_IN), .Z(n4777) );
  INV_X1 U5324 ( .A(n6023), .ZN(n4807) );
  NAND2_X1 U5325 ( .A1(n4807), .A2(n4075), .ZN(n4776) );
  NAND2_X1 U5326 ( .A1(n4777), .A2(n4776), .ZN(n5094) );
  NAND2_X1 U5327 ( .A1(n4858), .A2(n4780), .ZN(n4783) );
  INV_X1 U5328 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4784) );
  NAND2_X1 U5329 ( .A1(n4966), .A2(n4784), .ZN(n4782) );
  NAND3_X1 U5330 ( .A1(n4783), .A2(n3633), .A3(n4782), .ZN(n4786) );
  NAND2_X1 U5331 ( .A1(n3655), .A2(n4784), .ZN(n4785) );
  MUX2_X1 U5332 ( .A(n4861), .B(n3633), .S(EBX_REG_9__SCAN_IN), .Z(n4789) );
  OAI21_X1 U5333 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n6023), .A(n4789), 
        .ZN(n5264) );
  NAND2_X1 U5334 ( .A1(n4858), .A2(n4790), .ZN(n4792) );
  INV_X1 U5335 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4793) );
  NAND2_X1 U5336 ( .A1(n4966), .A2(n4793), .ZN(n4791) );
  NAND3_X1 U5337 ( .A1(n4792), .A2(n3633), .A3(n4791), .ZN(n4795) );
  NAND2_X1 U5338 ( .A1(n3655), .A2(n4793), .ZN(n4794) );
  NAND2_X1 U5339 ( .A1(n4795), .A2(n4794), .ZN(n5517) );
  INV_X1 U5340 ( .A(EBX_REG_11__SCAN_IN), .ZN(n7108) );
  NAND2_X1 U5341 ( .A1(n4854), .A2(n7108), .ZN(n4798) );
  NAND2_X1 U5342 ( .A1(n4966), .A2(n7108), .ZN(n4796) );
  OAI211_X1 U5343 ( .C1(n3655), .C2(n7198), .A(n4796), .B(n4858), .ZN(n4797)
         );
  NAND2_X1 U5344 ( .A1(n4798), .A2(n4797), .ZN(n5862) );
  NAND2_X1 U5345 ( .A1(n4858), .A2(n4801), .ZN(n4803) );
  INV_X1 U5346 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4804) );
  NAND2_X1 U5347 ( .A1(n4966), .A2(n4804), .ZN(n4802) );
  NAND3_X1 U5348 ( .A1(n4803), .A2(n3633), .A3(n4802), .ZN(n4806) );
  NAND2_X1 U5349 ( .A1(n3655), .A2(n4804), .ZN(n4805) );
  MUX2_X1 U5350 ( .A(n4861), .B(n3633), .S(EBX_REG_13__SCAN_IN), .Z(n4809) );
  NAND2_X1 U5351 ( .A1(n4807), .A2(n4096), .ZN(n4808) );
  NAND2_X1 U5352 ( .A1(n4858), .A2(n4810), .ZN(n4812) );
  INV_X1 U5353 ( .A(EBX_REG_14__SCAN_IN), .ZN(n7380) );
  NAND2_X1 U5354 ( .A1(n4966), .A2(n7380), .ZN(n4811) );
  NAND3_X1 U5355 ( .A1(n4812), .A2(n3633), .A3(n4811), .ZN(n4814) );
  NAND2_X1 U5356 ( .A1(n3655), .A2(n7380), .ZN(n4813) );
  NAND2_X1 U5357 ( .A1(n4814), .A2(n4813), .ZN(n5757) );
  NAND2_X1 U5358 ( .A1(n5758), .A2(n5757), .ZN(n5817) );
  MUX2_X1 U5359 ( .A(n4861), .B(n3633), .S(EBX_REG_15__SCAN_IN), .Z(n4815) );
  OAI21_X1 U5360 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n6023), .A(n4815), 
        .ZN(n5818) );
  NAND2_X1 U5361 ( .A1(n4858), .A2(n4818), .ZN(n4820) );
  INV_X1 U5362 ( .A(EBX_REG_16__SCAN_IN), .ZN(n7391) );
  NAND2_X1 U5363 ( .A1(n4966), .A2(n7391), .ZN(n4819) );
  NAND3_X1 U5364 ( .A1(n4820), .A2(n3633), .A3(n4819), .ZN(n4822) );
  NAND2_X1 U5365 ( .A1(n3655), .A2(n7391), .ZN(n4821) );
  AND2_X1 U5366 ( .A1(n4822), .A2(n4821), .ZN(n5882) );
  OR2_X2 U5367 ( .A1(n5881), .A2(n5882), .ZN(n7112) );
  INV_X1 U5368 ( .A(EBX_REG_17__SCAN_IN), .ZN(n7116) );
  NAND2_X1 U5369 ( .A1(n4854), .A2(n7116), .ZN(n4826) );
  INV_X1 U5370 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4824) );
  NAND2_X1 U5371 ( .A1(n4966), .A2(n7116), .ZN(n4823) );
  OAI211_X1 U5372 ( .C1(n3655), .C2(n4824), .A(n4823), .B(n4858), .ZN(n4825)
         );
  NAND2_X1 U5373 ( .A1(n4826), .A2(n4825), .ZN(n7111) );
  INV_X1 U5374 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6907) );
  NAND2_X1 U5375 ( .A1(n4858), .A2(n6907), .ZN(n4829) );
  INV_X1 U5376 ( .A(EBX_REG_18__SCAN_IN), .ZN(n4830) );
  NAND2_X1 U5377 ( .A1(n4966), .A2(n4830), .ZN(n4828) );
  NAND3_X1 U5378 ( .A1(n4829), .A2(n3633), .A3(n4828), .ZN(n4832) );
  NAND2_X1 U5379 ( .A1(n3655), .A2(n4830), .ZN(n4831) );
  NAND2_X1 U5380 ( .A1(n4832), .A2(n4831), .ZN(n5990) );
  INV_X1 U5381 ( .A(EBX_REG_19__SCAN_IN), .ZN(n7409) );
  NAND2_X1 U5382 ( .A1(n4854), .A2(n7409), .ZN(n4835) );
  INV_X1 U5383 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6767) );
  NAND2_X1 U5384 ( .A1(n4966), .A2(n7409), .ZN(n4833) );
  OAI211_X1 U5385 ( .C1(n3655), .C2(n6767), .A(n4833), .B(n4858), .ZN(n4834)
         );
  NAND2_X1 U5386 ( .A1(n4835), .A2(n4834), .ZN(n6899) );
  INV_X1 U5387 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6884) );
  OAI21_X1 U5388 ( .B1(n3655), .B2(n6884), .A(n4858), .ZN(n4838) );
  INV_X1 U5389 ( .A(EBX_REG_20__SCAN_IN), .ZN(n4836) );
  NAND2_X1 U5390 ( .A1(n4966), .A2(n4836), .ZN(n4837) );
  AOI22_X1 U5391 ( .A1(n4838), .A2(n4837), .B1(n3655), .B2(n4836), .ZN(n6646)
         );
  INV_X1 U5392 ( .A(EBX_REG_21__SCAN_IN), .ZN(n7436) );
  NAND2_X1 U5393 ( .A1(n4854), .A2(n7436), .ZN(n4841) );
  INV_X1 U5394 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6727) );
  NAND2_X1 U5395 ( .A1(n4966), .A2(n7436), .ZN(n4839) );
  OAI211_X1 U5396 ( .C1(n3655), .C2(n6727), .A(n4839), .B(n4858), .ZN(n4840)
         );
  AND2_X1 U5397 ( .A1(n4841), .A2(n4840), .ZN(n6876) );
  NAND2_X1 U5398 ( .A1(n6877), .A2(n6876), .ZN(n6590) );
  INV_X1 U5399 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6867) );
  NAND2_X1 U5400 ( .A1(n4858), .A2(n6867), .ZN(n4843) );
  INV_X1 U5401 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U5402 ( .A1(n4966), .A2(n6641), .ZN(n4842) );
  NAND3_X1 U5403 ( .A1(n4843), .A2(n3633), .A3(n4842), .ZN(n4845) );
  NAND2_X1 U5404 ( .A1(n3655), .A2(n6641), .ZN(n4844) );
  AND2_X1 U5405 ( .A1(n4845), .A2(n4844), .ZN(n6591) );
  INV_X1 U5407 ( .A(EBX_REG_23__SCAN_IN), .ZN(n4846) );
  NAND2_X1 U5408 ( .A1(n4854), .A2(n4846), .ZN(n4849) );
  NAND2_X1 U5409 ( .A1(n4966), .A2(n4846), .ZN(n4847) );
  OAI211_X1 U5410 ( .C1(n3655), .C2(n6860), .A(n4847), .B(n4858), .ZN(n4848)
         );
  NAND2_X1 U5411 ( .A1(n4849), .A2(n4848), .ZN(n6575) );
  OAI21_X1 U5412 ( .B1(n3655), .B2(n6849), .A(n4858), .ZN(n4851) );
  INV_X1 U5413 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U5414 ( .A1(n4966), .A2(n6567), .ZN(n4850) );
  NAND2_X1 U5415 ( .A1(n4851), .A2(n4850), .ZN(n4853) );
  NAND2_X1 U5416 ( .A1(n3655), .A2(n6567), .ZN(n4852) );
  NAND2_X1 U5417 ( .A1(n4853), .A2(n4852), .ZN(n6561) );
  INV_X1 U5418 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6634) );
  NAND2_X1 U5419 ( .A1(n4854), .A2(n6634), .ZN(n4857) );
  NAND2_X1 U5420 ( .A1(n4966), .A2(n6634), .ZN(n4855) );
  OAI211_X1 U5421 ( .C1(n3655), .C2(n6846), .A(n4855), .B(n4858), .ZN(n4856)
         );
  AND2_X1 U5422 ( .A1(n4857), .A2(n4856), .ZN(n6553) );
  NAND2_X1 U5423 ( .A1(n6552), .A2(n6553), .ZN(n6522) );
  OAI21_X1 U5424 ( .B1(n3655), .B2(n6835), .A(n4858), .ZN(n4860) );
  INV_X1 U5425 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U5426 ( .A1(n4966), .A2(n6633), .ZN(n4859) );
  AOI22_X1 U5427 ( .A1(n4860), .A2(n4859), .B1(n3655), .B2(n6633), .ZN(n6523)
         );
  MUX2_X1 U5428 ( .A(n4861), .B(n3633), .S(EBX_REG_27__SCAN_IN), .Z(n4862) );
  OAI21_X1 U5429 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n6023), .A(n4862), 
        .ZN(n6519) );
  INV_X1 U5430 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6811) );
  NAND2_X1 U5431 ( .A1(n4858), .A2(n6811), .ZN(n4863) );
  OAI211_X1 U5432 ( .C1(EBX_REG_28__SCAN_IN), .C2(n6022), .A(n4863), .B(n3633), 
        .ZN(n4865) );
  INV_X1 U5433 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6631) );
  NAND2_X1 U5434 ( .A1(n3655), .A2(n6631), .ZN(n4864) );
  NAND2_X1 U5435 ( .A1(n4865), .A2(n4864), .ZN(n6496) );
  NAND2_X1 U5436 ( .A1(n6518), .A2(n6496), .ZN(n6027) );
  MUX2_X1 U5437 ( .A(n6024), .B(n3633), .S(n6027), .Z(n4866) );
  OAI22_X1 U5438 ( .A1(n6023), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n6022), .ZN(n6030) );
  INV_X1 U5439 ( .A(n6113), .ZN(n4886) );
  INV_X1 U5440 ( .A(REIP_REG_30__SCAN_IN), .ZN(n7068) );
  NOR2_X1 U5441 ( .A1(n7211), .A2(n7068), .ZN(n6034) );
  NAND3_X1 U5442 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n5971) );
  NOR2_X1 U5443 ( .A1(n4810), .A2(n5971), .ZN(n4893) );
  INV_X1 U5444 ( .A(n4893), .ZN(n7261) );
  NOR2_X1 U5445 ( .A1(n4780), .A2(n4075), .ZN(n7245) );
  NAND3_X1 U5446 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n7245), .ZN(n4881) );
  NAND2_X1 U5447 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n7219) );
  NOR3_X1 U5448 ( .A1(n4771), .A2(n7213), .A3(n7219), .ZN(n4880) );
  INV_X1 U5449 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5002) );
  OAI21_X1 U5450 ( .B1(n5014), .B2(n5002), .A(n7234), .ZN(n7232) );
  NAND2_X1 U5451 ( .A1(n4880), .A2(n7232), .ZN(n5352) );
  NOR2_X1 U5452 ( .A1(n4881), .A2(n5352), .ZN(n5857) );
  NAND2_X1 U5453 ( .A1(n3650), .A2(n3654), .ZN(n5738) );
  OR2_X1 U5454 ( .A1(n5738), .A2(n4867), .ZN(n4984) );
  OAI21_X1 U5455 ( .B1(n5230), .B2(n4868), .A(n4984), .ZN(n4869) );
  AOI21_X1 U5456 ( .B1(n4870), .B2(n6023), .A(n4869), .ZN(n4871) );
  AND2_X1 U5457 ( .A1(n4872), .A2(n4871), .ZN(n4873) );
  INV_X1 U5458 ( .A(n5137), .ZN(n6095) );
  NAND2_X1 U5459 ( .A1(n4729), .A2(n3654), .ZN(n5144) );
  INV_X1 U5460 ( .A(n4890), .ZN(n4879) );
  NAND2_X1 U5461 ( .A1(n7452), .A2(n4876), .ZN(n5145) );
  OAI211_X1 U5462 ( .C1(n5057), .C2(n4877), .A(n4977), .B(n5145), .ZN(n4878)
         );
  NAND2_X1 U5463 ( .A1(n4879), .A2(n4878), .ZN(n4891) );
  NAND2_X1 U5464 ( .A1(n5002), .A2(n5005), .ZN(n5012) );
  NAND2_X1 U5465 ( .A1(n5350), .A2(n5012), .ZN(n5071) );
  INV_X1 U5466 ( .A(n5071), .ZN(n7235) );
  NAND2_X1 U5467 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5070) );
  INV_X1 U5468 ( .A(n4880), .ZN(n5348) );
  OR2_X1 U5469 ( .A1(n5070), .A2(n5348), .ZN(n5349) );
  NOR2_X1 U5470 ( .A1(n4881), .A2(n5349), .ZN(n4889) );
  NAND2_X1 U5471 ( .A1(n7235), .A2(n4889), .ZN(n6910) );
  NAND2_X1 U5472 ( .A1(n7233), .A2(n6910), .ZN(n5888) );
  AND2_X1 U5473 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4882) );
  NAND2_X1 U5474 ( .A1(n7272), .A2(n4882), .ZN(n7282) );
  INV_X1 U5475 ( .A(n4883), .ZN(n4884) );
  NAND2_X1 U5476 ( .A1(n6864), .A2(n4884), .ZN(n6831) );
  NAND2_X1 U5477 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6832) );
  NOR2_X1 U5478 ( .A1(n6831), .A2(n6832), .ZN(n6809) );
  INV_X1 U5479 ( .A(n6682), .ZN(n6810) );
  NAND2_X1 U5480 ( .A1(n6809), .A2(n6810), .ZN(n6801) );
  NOR3_X1 U5481 ( .A1(n6801), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n6802), 
        .ZN(n4885) );
  AOI211_X1 U5482 ( .C1(n7269), .C2(n4886), .A(n6034), .B(n4885), .ZN(n4908)
         );
  NAND2_X1 U5483 ( .A1(n4891), .A2(n7233), .ZN(n5001) );
  INV_X1 U5484 ( .A(n5001), .ZN(n4887) );
  NAND2_X1 U5485 ( .A1(n4887), .A2(n5005), .ZN(n7260) );
  INV_X1 U5486 ( .A(n7260), .ZN(n7246) );
  INV_X1 U5487 ( .A(n6888), .ZN(n6726) );
  NOR2_X1 U5488 ( .A1(n6906), .A2(n6726), .ZN(n6873) );
  INV_X1 U5489 ( .A(n4888), .ZN(n4900) );
  INV_X1 U5490 ( .A(n4889), .ZN(n4892) );
  NAND2_X1 U5491 ( .A1(n7211), .A2(n4890), .ZN(n5016) );
  OAI21_X1 U5492 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n4891), .A(n5016), 
        .ZN(n5351) );
  AOI21_X1 U5493 ( .B1(n5350), .B2(n4892), .A(n5351), .ZN(n5856) );
  INV_X1 U5494 ( .A(n7233), .ZN(n5353) );
  NAND3_X1 U5495 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n4893), .ZN(n4895) );
  NAND2_X1 U5496 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5857), .ZN(n4894) );
  AOI222_X1 U5497 ( .A1(n5353), .A2(n4895), .B1(n5353), .B2(n4894), .C1(n4895), 
        .C2(n5350), .ZN(n4896) );
  NAND2_X1 U5498 ( .A1(n5856), .A2(n4896), .ZN(n7277) );
  AND2_X1 U5499 ( .A1(n7260), .A2(n4897), .ZN(n4898) );
  NOR2_X1 U5500 ( .A1(n7277), .A2(n4898), .ZN(n6895) );
  NAND2_X1 U5501 ( .A1(n7260), .A2(n6726), .ZN(n4899) );
  NAND2_X1 U5502 ( .A1(n6895), .A2(n4899), .ZN(n6880) );
  AOI21_X1 U5503 ( .B1(n6873), .B2(n4900), .A(n6880), .ZN(n6865) );
  NAND2_X1 U5504 ( .A1(n5071), .A2(n7233), .ZN(n4903) );
  INV_X1 U5505 ( .A(n4901), .ZN(n4902) );
  NAND2_X1 U5506 ( .A1(n4903), .A2(n4902), .ZN(n4904) );
  NAND2_X1 U5507 ( .A1(n6847), .A2(n7246), .ZN(n6049) );
  INV_X1 U5508 ( .A(n6832), .ZN(n4905) );
  NAND2_X1 U5509 ( .A1(n6847), .A2(n4905), .ZN(n4906) );
  NAND2_X1 U5510 ( .A1(n6049), .A2(n4906), .ZN(n6816) );
  OAI211_X1 U5511 ( .C1(n6810), .C2(n7246), .A(n6816), .B(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6799) );
  NAND3_X1 U5512 ( .A1(n6799), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n6049), .ZN(n4907) );
  AND2_X1 U5513 ( .A1(n4908), .A2(n4907), .ZN(n4909) );
  OAI21_X1 U5514 ( .B1(n6038), .B2(n6892), .A(n4909), .ZN(U2988) );
  XNOR2_X1 U5515 ( .A(n6114), .B(n4911), .ZN(n6649) );
  NAND2_X1 U5516 ( .A1(n6097), .A2(n5137), .ZN(n4988) );
  NOR2_X1 U5517 ( .A1(n3798), .A2(n4193), .ZN(n5055) );
  AND2_X1 U5518 ( .A1(n3837), .A2(n5054), .ZN(n4913) );
  NAND4_X1 U5519 ( .A1(n5055), .A2(n4913), .A3(n4912), .A4(n4966), .ZN(n4914)
         );
  NAND2_X1 U5520 ( .A1(n4988), .A2(n4914), .ZN(n4915) );
  INV_X1 U5521 ( .A(n4193), .ZN(n6086) );
  INV_X1 U5522 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4917) );
  AND3_X1 U5523 ( .A1(n4729), .A2(n7499), .A3(n6098), .ZN(n5707) );
  INV_X1 U5524 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7542) );
  INV_X1 U5525 ( .A(n7499), .ZN(n7517) );
  INV_X1 U5526 ( .A(n5708), .ZN(n4923) );
  OAI211_X1 U5527 ( .C1(n5707), .C2(n7542), .A(n4923), .B(n7178), .ZN(U2788)
         );
  INV_X1 U5528 ( .A(DATAI_15_), .ZN(n5849) );
  AND2_X1 U5529 ( .A1(n3654), .A2(n7502), .ZN(n4922) );
  INV_X1 U5530 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4925) );
  AOI21_X1 U5531 ( .B1(n3653), .B2(READY_N), .A(n4923), .ZN(n4926) );
  INV_X1 U5532 ( .A(EAX_REG_15__SCAN_IN), .ZN(n4924) );
  NAND2_X1 U5533 ( .A1(n5708), .A2(n3820), .ZN(n5224) );
  OAI222_X1 U5534 ( .A1(n5849), .A2(n5061), .B1(n4925), .B2(n4926), .C1(n4924), 
        .C2(n5224), .ZN(U2954) );
  INV_X2 U5535 ( .A(n5224), .ZN(n5201) );
  AOI22_X1 U5536 ( .A1(n5176), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n5201), .ZN(n4927) );
  NAND2_X1 U5537 ( .A1(n5052), .A2(DATAI_1_), .ZN(n5218) );
  NAND2_X1 U5538 ( .A1(n4927), .A2(n5218), .ZN(U2940) );
  AOI22_X1 U5539 ( .A1(n5176), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n5201), .ZN(n4928) );
  NAND2_X1 U5540 ( .A1(n5052), .A2(DATAI_3_), .ZN(n5179) );
  NAND2_X1 U5541 ( .A1(n4928), .A2(n5179), .ZN(U2942) );
  AOI22_X1 U5542 ( .A1(n5176), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n5201), .ZN(n4929) );
  NAND2_X1 U5543 ( .A1(n5052), .A2(DATAI_4_), .ZN(n5181) );
  NAND2_X1 U5544 ( .A1(n4929), .A2(n5181), .ZN(U2943) );
  AOI22_X1 U5545 ( .A1(n5176), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n5201), .ZN(n4930) );
  NAND2_X1 U5546 ( .A1(n5052), .A2(DATAI_14_), .ZN(n5183) );
  NAND2_X1 U5547 ( .A1(n4930), .A2(n5183), .ZN(U2938) );
  AOI22_X1 U5548 ( .A1(n5176), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n5201), .ZN(n4931) );
  NAND2_X1 U5549 ( .A1(n5052), .A2(DATAI_5_), .ZN(n5195) );
  NAND2_X1 U5550 ( .A1(n4931), .A2(n5195), .ZN(U2944) );
  AOI22_X1 U5551 ( .A1(n5176), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n5201), .ZN(n4932) );
  NAND2_X1 U5552 ( .A1(n5052), .A2(DATAI_2_), .ZN(n5177) );
  NAND2_X1 U5553 ( .A1(n4932), .A2(n5177), .ZN(U2941) );
  AOI22_X1 U5554 ( .A1(n5176), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n5201), .ZN(n4933) );
  NAND2_X1 U5555 ( .A1(n5052), .A2(DATAI_6_), .ZN(n5185) );
  NAND2_X1 U5556 ( .A1(n4933), .A2(n5185), .ZN(U2945) );
  AOI22_X1 U5557 ( .A1(n5176), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n5201), .ZN(n4934) );
  NAND2_X1 U5558 ( .A1(n5052), .A2(DATAI_0_), .ZN(n5221) );
  NAND2_X1 U5559 ( .A1(n4934), .A2(n5221), .ZN(U2939) );
  OAI21_X1 U5560 ( .B1(n6023), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4935), 
        .ZN(n5806) );
  XNOR2_X1 U5561 ( .A(n4937), .B(n4936), .ZN(n5811) );
  INV_X1 U5562 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4938) );
  OAI222_X1 U5563 ( .A1(n5806), .A2(n6647), .B1(n6648), .B2(n5811), .C1(n4938), 
        .C2(n7126), .ZN(U2859) );
  INV_X1 U5564 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4944) );
  NAND2_X1 U5565 ( .A1(n7496), .A2(n5144), .ZN(n4940) );
  NAND3_X1 U5566 ( .A1(n4940), .A2(n4939), .A3(n7499), .ZN(n4941) );
  NAND2_X1 U5567 ( .A1(n4942), .A2(n4743), .ZN(n5217) );
  AND2_X1 U5568 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5709), .ZN(n7192) );
  NOR2_X4 U5569 ( .A1(n7492), .A2(n4942), .ZN(n7003) );
  AOI22_X1 U5570 ( .A1(n7492), .A2(UWORD_REG_9__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4943) );
  OAI21_X1 U5571 ( .B1(n4944), .B2(n5217), .A(n4943), .ZN(U2898) );
  INV_X1 U5572 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4946) );
  AOI22_X1 U5573 ( .A1(n7492), .A2(UWORD_REG_5__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4945) );
  OAI21_X1 U5574 ( .B1(n4946), .B2(n5217), .A(n4945), .ZN(U2902) );
  INV_X1 U5575 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4948) );
  AOI22_X1 U5576 ( .A1(n7492), .A2(UWORD_REG_7__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4947) );
  OAI21_X1 U5577 ( .B1(n4948), .B2(n5217), .A(n4947), .ZN(U2900) );
  INV_X1 U5578 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4950) );
  AOI22_X1 U5579 ( .A1(n7492), .A2(UWORD_REG_12__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4949) );
  OAI21_X1 U5580 ( .B1(n4950), .B2(n5217), .A(n4949), .ZN(U2895) );
  INV_X1 U5581 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4952) );
  AOI22_X1 U5582 ( .A1(n7492), .A2(UWORD_REG_8__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4951) );
  OAI21_X1 U5583 ( .B1(n4952), .B2(n5217), .A(n4951), .ZN(U2899) );
  INV_X1 U5584 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4954) );
  AOI22_X1 U5585 ( .A1(n7492), .A2(UWORD_REG_10__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4953) );
  OAI21_X1 U5586 ( .B1(n4954), .B2(n5217), .A(n4953), .ZN(U2897) );
  INV_X1 U5587 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4956) );
  AOI22_X1 U5588 ( .A1(n7492), .A2(UWORD_REG_4__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4955) );
  OAI21_X1 U5589 ( .B1(n4956), .B2(n5217), .A(n4955), .ZN(U2903) );
  AOI22_X1 U5590 ( .A1(n7492), .A2(UWORD_REG_11__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4957) );
  OAI21_X1 U5591 ( .B1(n4622), .B2(n5217), .A(n4957), .ZN(U2896) );
  INV_X1 U5592 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4959) );
  AOI22_X1 U5593 ( .A1(n7492), .A2(UWORD_REG_6__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4958) );
  OAI21_X1 U5594 ( .B1(n4959), .B2(n5217), .A(n4958), .ZN(U2901) );
  OAI21_X1 U5595 ( .B1(n4962), .B2(n4961), .A(n4960), .ZN(n7127) );
  XNOR2_X1 U5596 ( .A(n4963), .B(n5034), .ZN(n7227) );
  AOI22_X1 U5597 ( .A1(n7124), .A2(n7227), .B1(EBX_REG_2__SCAN_IN), .B2(n6636), 
        .ZN(n4964) );
  OAI21_X1 U5598 ( .B1(n6648), .B2(n7127), .A(n4964), .ZN(U2857) );
  OAI21_X1 U5599 ( .B1(n4967), .B2(n4966), .A(n4965), .ZN(n6625) );
  INV_X1 U5600 ( .A(n6625), .ZN(n4973) );
  OR2_X1 U5601 ( .A1(n4969), .A2(n4968), .ZN(n4971) );
  AND2_X1 U5602 ( .A1(n4971), .A2(n4970), .ZN(n6620) );
  AOI22_X1 U5603 ( .A1(n4916), .A2(n6620), .B1(EBX_REG_1__SCAN_IN), .B2(n6636), 
        .ZN(n4972) );
  OAI21_X1 U5604 ( .B1(n4973), .B2(n6647), .A(n4972), .ZN(U2858) );
  INV_X1 U5605 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n7508) );
  INV_X1 U5606 ( .A(n6059), .ZN(n7513) );
  INV_X1 U5607 ( .A(n4974), .ZN(n4982) );
  AOI22_X1 U5608 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4118), .B2(n5014), .ZN(n6055)
         );
  NOR2_X1 U5609 ( .A1(n7455), .A2(n5002), .ZN(n6054) );
  INV_X1 U5610 ( .A(n6054), .ZN(n4981) );
  INV_X1 U5611 ( .A(n7501), .ZN(n7459) );
  INV_X1 U5612 ( .A(n3648), .ZN(n5273) );
  AND3_X1 U5613 ( .A1(n7460), .A2(n4990), .A3(n5057), .ZN(n4976) );
  NAND2_X1 U5614 ( .A1(n4977), .A2(n4976), .ZN(n7453) );
  OAI21_X1 U5615 ( .B1(n4978), .B2(n4974), .A(n7452), .ZN(n4979) );
  OAI21_X1 U5616 ( .B1(n5144), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n4979), 
        .ZN(n4980) );
  AOI21_X1 U5617 ( .B1(n5273), .B2(n7453), .A(n4980), .ZN(n7471) );
  OAI222_X1 U5618 ( .A1(n7513), .A2(n4982), .B1(n6055), .B2(n4981), .C1(n7459), 
        .C2(n7471), .ZN(n4996) );
  OAI22_X1 U5619 ( .A1(n6097), .A2(n5135), .B1(n4983), .B2(n7460), .ZN(n5059)
         );
  INV_X1 U5620 ( .A(n5059), .ZN(n4995) );
  INV_X1 U5621 ( .A(n4984), .ZN(n4985) );
  NOR2_X1 U5622 ( .A1(n4986), .A2(n4985), .ZN(n4987) );
  AND2_X1 U5623 ( .A1(n4988), .A2(n4987), .ZN(n4994) );
  INV_X1 U5624 ( .A(n4989), .ZN(n4992) );
  AOI22_X1 U5625 ( .A1(n6100), .A2(n7183), .B1(n5144), .B2(n4990), .ZN(n4991)
         );
  NAND2_X1 U5626 ( .A1(n4992), .A2(n4991), .ZN(n4993) );
  NOR2_X1 U5627 ( .A1(n7188), .A2(n7455), .ZN(n6039) );
  NAND2_X1 U5628 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6039), .ZN(n7507) );
  INV_X1 U5629 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7448) );
  OAI22_X1 U5630 ( .A1(n7472), .A2(n7517), .B1(n7507), .B2(n7448), .ZN(n7463)
         );
  AOI21_X1 U5631 ( .B1(n3848), .B2(STATE2_REG_3__SCAN_IN), .A(n7463), .ZN(
        n6920) );
  INV_X1 U5632 ( .A(n6920), .ZN(n7466) );
  OAI21_X1 U5633 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7513), .A(n7466), 
        .ZN(n7456) );
  AOI22_X1 U5634 ( .A1(n4996), .A2(n7466), .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n7456), .ZN(n4997) );
  INV_X1 U5635 ( .A(n4997), .ZN(U3460) );
  OAI21_X1 U5636 ( .B1(n4999), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4998), 
        .ZN(n5086) );
  INV_X1 U5637 ( .A(n5806), .ZN(n5004) );
  INV_X1 U5638 ( .A(REIP_REG_0__SCAN_IN), .ZN(n5000) );
  NOR2_X1 U5639 ( .A1(n7211), .A2(n5000), .ZN(n5082) );
  NAND2_X1 U5640 ( .A1(n5002), .A2(n5001), .ZN(n5015) );
  INV_X1 U5641 ( .A(n5015), .ZN(n5003) );
  AOI211_X1 U5642 ( .C1(n7269), .C2(n5004), .A(n5082), .B(n5003), .ZN(n5009)
         );
  INV_X1 U5643 ( .A(n5005), .ZN(n5007) );
  INV_X1 U5644 ( .A(n5016), .ZN(n5006) );
  OAI21_X1 U5645 ( .B1(n5007), .B2(n5006), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5008) );
  OAI211_X1 U5646 ( .C1(n6892), .C2(n5086), .A(n5009), .B(n5008), .ZN(U3018)
         );
  XNOR2_X1 U5647 ( .A(n4998), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5011)
         );
  XNOR2_X1 U5648 ( .A(n5010), .B(n5011), .ZN(n5783) );
  NAND3_X1 U5649 ( .A1(n7260), .A2(n5012), .A3(n5014), .ZN(n5019) );
  INV_X1 U5650 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5013) );
  NOR2_X1 U5651 ( .A1(n7211), .A2(n5013), .ZN(n5777) );
  AOI21_X1 U5652 ( .B1(n5016), .B2(n5015), .A(n5014), .ZN(n5017) );
  AOI211_X1 U5653 ( .C1(n7269), .C2(n6625), .A(n5777), .B(n5017), .ZN(n5018)
         );
  OAI211_X1 U5654 ( .C1(n5783), .C2(n6892), .A(n5019), .B(n5018), .ZN(U3017)
         );
  CLKBUF_X1 U5655 ( .A(n5020), .Z(n5091) );
  NAND2_X1 U5656 ( .A1(n5077), .A2(n5038), .ZN(n5040) );
  INV_X1 U5657 ( .A(n5022), .ZN(n5023) );
  NAND2_X1 U5658 ( .A1(n5040), .A2(n5023), .ZN(n5024) );
  INV_X1 U5659 ( .A(n7318), .ZN(n5066) );
  CLKBUF_X1 U5660 ( .A(n5026), .Z(n5093) );
  OAI21_X1 U5661 ( .B1(n5043), .B2(n5027), .A(n5093), .ZN(n7314) );
  INV_X1 U5662 ( .A(n7314), .ZN(n5028) );
  AOI22_X1 U5663 ( .A1(n7124), .A2(n5028), .B1(EBX_REG_6__SCAN_IN), .B2(n6636), 
        .ZN(n5029) );
  OAI21_X1 U5664 ( .B1(n5066), .B2(n6648), .A(n5029), .ZN(U2853) );
  OAI21_X1 U5665 ( .B1(n4217), .B2(n5032), .A(n5031), .ZN(n6617) );
  INV_X1 U5666 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6609) );
  INV_X1 U5667 ( .A(n4963), .ZN(n5035) );
  AOI21_X1 U5668 ( .B1(n5035), .B2(n5034), .A(n5033), .ZN(n5036) );
  INV_X1 U5669 ( .A(n7123), .ZN(n5042) );
  NOR2_X1 U5670 ( .A1(n5036), .A2(n5042), .ZN(n6612) );
  INV_X1 U5671 ( .A(n6612), .ZN(n5037) );
  OAI222_X1 U5672 ( .A1(n6617), .A2(n6648), .B1(n6609), .B2(n7126), .C1(n5037), 
        .C2(n6647), .ZN(U2856) );
  OR2_X1 U5673 ( .A1(n5077), .A2(n5038), .ZN(n5039) );
  INV_X1 U5674 ( .A(n7306), .ZN(n5065) );
  AOI21_X1 U5675 ( .B1(n5042), .B2(n7122), .A(n5041), .ZN(n5044) );
  OR2_X1 U5676 ( .A1(n5044), .A2(n5043), .ZN(n7299) );
  OAI222_X1 U5677 ( .A1(n5065), .A2(n6648), .B1(n5045), .B2(n7126), .C1(n6647), 
        .C2(n7299), .ZN(U2854) );
  AOI22_X1 U5678 ( .A1(n5176), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n5201), .ZN(n5046) );
  NAND2_X1 U5679 ( .A1(n5052), .A2(DATAI_12_), .ZN(n5199) );
  NAND2_X1 U5680 ( .A1(n5046), .A2(n5199), .ZN(U2936) );
  AOI22_X1 U5681 ( .A1(n5176), .A2(UWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_27__SCAN_IN), .B2(n5201), .ZN(n5047) );
  NAND2_X1 U5682 ( .A1(n5052), .A2(DATAI_11_), .ZN(n5197) );
  NAND2_X1 U5683 ( .A1(n5047), .A2(n5197), .ZN(U2935) );
  AOI22_X1 U5684 ( .A1(n5176), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n5201), .ZN(n5048) );
  NAND2_X1 U5685 ( .A1(n5052), .A2(DATAI_7_), .ZN(n5187) );
  NAND2_X1 U5686 ( .A1(n5048), .A2(n5187), .ZN(U2946) );
  AOI22_X1 U5687 ( .A1(n5176), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n5201), .ZN(n5049) );
  NAND2_X1 U5688 ( .A1(n5052), .A2(DATAI_10_), .ZN(n5193) );
  NAND2_X1 U5689 ( .A1(n5049), .A2(n5193), .ZN(U2949) );
  AOI22_X1 U5690 ( .A1(n5176), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n5201), .ZN(n5050) );
  NAND2_X1 U5691 ( .A1(n5052), .A2(DATAI_13_), .ZN(n5202) );
  NAND2_X1 U5692 ( .A1(n5050), .A2(n5202), .ZN(U2937) );
  AOI22_X1 U5693 ( .A1(n5176), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n5201), .ZN(n5051) );
  NAND2_X1 U5694 ( .A1(n5052), .A2(DATAI_8_), .ZN(n5189) );
  NAND2_X1 U5695 ( .A1(n5051), .A2(n5189), .ZN(U2947) );
  AOI22_X1 U5696 ( .A1(n5176), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n5201), .ZN(n5053) );
  NAND2_X1 U5697 ( .A1(n5052), .A2(DATAI_9_), .ZN(n5191) );
  NAND2_X1 U5698 ( .A1(n5053), .A2(n5191), .ZN(U2948) );
  NAND2_X1 U5699 ( .A1(n5055), .A2(n5054), .ZN(n5056) );
  NOR2_X1 U5700 ( .A1(n5057), .A2(n5056), .ZN(n5058) );
  NAND2_X1 U5701 ( .A1(n5063), .A2(n4193), .ZN(n5064) );
  INV_X1 U5702 ( .A(DATAI_2_), .ZN(n5231) );
  INV_X1 U5703 ( .A(EAX_REG_2__SCAN_IN), .ZN(n7000) );
  OAI222_X1 U5704 ( .A1(n5848), .A2(n5231), .B1(n6085), .B2(n7000), .C1(n6669), 
        .C2(n7127), .ZN(U2889) );
  INV_X1 U5705 ( .A(DATAI_3_), .ZN(n5241) );
  INV_X1 U5706 ( .A(EAX_REG_3__SCAN_IN), .ZN(n7002) );
  OAI222_X1 U5707 ( .A1(n5241), .A2(n5848), .B1(n6085), .B2(n7002), .C1(n6669), 
        .C2(n6617), .ZN(U2888) );
  INV_X1 U5708 ( .A(DATAI_0_), .ZN(n5253) );
  INV_X1 U5709 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6996) );
  OAI222_X1 U5710 ( .A1(n5848), .A2(n5253), .B1(n6085), .B2(n6996), .C1(n6669), 
        .C2(n5811), .ZN(U2891) );
  INV_X1 U5711 ( .A(DATAI_1_), .ZN(n5246) );
  INV_X1 U5712 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6998) );
  INV_X1 U5713 ( .A(n6620), .ZN(n5780) );
  OAI222_X1 U5714 ( .A1(n5246), .A2(n5848), .B1(n6085), .B2(n6998), .C1(n6669), 
        .C2(n5780), .ZN(U2890) );
  INV_X1 U5715 ( .A(DATAI_5_), .ZN(n5236) );
  OAI222_X1 U5716 ( .A1(n5236), .A2(n5848), .B1(n6085), .B2(n4246), .C1(n6669), 
        .C2(n5065), .ZN(U2886) );
  INV_X1 U5717 ( .A(DATAI_6_), .ZN(n6675) );
  OAI222_X1 U5718 ( .A1(n5848), .A2(n6675), .B1(n6085), .B2(n4234), .C1(n6669), 
        .C2(n5066), .ZN(U2885) );
  XNOR2_X1 U5719 ( .A(n5068), .B(n5072), .ZN(n5069) );
  XNOR2_X1 U5720 ( .A(n3639), .B(n5069), .ZN(n5751) );
  AOI21_X1 U5721 ( .B1(n5350), .B2(n5070), .A(n5351), .ZN(n7228) );
  OAI21_X1 U5722 ( .B1(n7232), .B2(n7233), .A(n7228), .ZN(n7208) );
  OAI21_X1 U5723 ( .B1(n5071), .B2(n5070), .A(n7233), .ZN(n7210) );
  NAND2_X1 U5724 ( .A1(n7232), .A2(n7210), .ZN(n7218) );
  INV_X1 U5725 ( .A(n7218), .ZN(n5073) );
  AOI22_X1 U5726 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n7208), .B1(n5073), 
        .B2(n5072), .ZN(n5076) );
  INV_X1 U5727 ( .A(REIP_REG_3__SCAN_IN), .ZN(n5074) );
  NOR2_X1 U5728 ( .A1(n7211), .A2(n5074), .ZN(n5746) );
  AOI21_X1 U5729 ( .B1(n7269), .B2(n6612), .A(n5746), .ZN(n5075) );
  OAI211_X1 U5730 ( .C1(n5751), .C2(n6892), .A(n5076), .B(n5075), .ZN(U3015)
         );
  AOI21_X1 U5731 ( .B1(n5078), .B2(n5031), .A(n5077), .ZN(n7139) );
  INV_X1 U5732 ( .A(n7139), .ZN(n7291) );
  INV_X1 U5733 ( .A(EAX_REG_4__SCAN_IN), .ZN(n7005) );
  INV_X1 U5734 ( .A(DATAI_4_), .ZN(n6678) );
  OAI222_X1 U5735 ( .A1(n7291), .A2(n6669), .B1(n6085), .B2(n7005), .C1(n5848), 
        .C2(n6678), .ZN(U2887) );
  INV_X1 U5736 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n5079) );
  AOI21_X1 U5737 ( .B1(n6791), .B2(n5080), .A(n5079), .ZN(n5081) );
  INV_X1 U5738 ( .A(n5081), .ZN(n5085) );
  INV_X1 U5739 ( .A(n5811), .ZN(n5083) );
  AOI21_X1 U5740 ( .B1(n5083), .B2(n7165), .A(n5082), .ZN(n5084) );
  OAI211_X1 U5741 ( .C1(n5086), .C2(n7447), .A(n5085), .B(n5084), .ZN(U2986)
         );
  CLKBUF_X1 U5742 ( .A(n5088), .Z(n5089) );
  INV_X1 U5743 ( .A(n5089), .ZN(n5090) );
  AOI21_X1 U5744 ( .B1(n5087), .B2(n5091), .A(n5090), .ZN(n7328) );
  INV_X1 U5745 ( .A(n7328), .ZN(n5261) );
  AOI21_X1 U5746 ( .B1(n5094), .B2(n5093), .A(n4788), .ZN(n7322) );
  AOI22_X1 U5747 ( .A1(n7124), .A2(n7322), .B1(EBX_REG_7__SCAN_IN), .B2(n6636), 
        .ZN(n5095) );
  OAI21_X1 U5748 ( .B1(n5261), .B2(n6648), .A(n5095), .ZN(U2852) );
  NAND3_X1 U5749 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n7480), .ZN(n5632) );
  NOR2_X1 U5750 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5632), .ZN(n5257)
         );
  INV_X1 U5751 ( .A(n5097), .ZN(n6608) );
  INV_X1 U5752 ( .A(n6927), .ZN(n5107) );
  NAND2_X1 U5753 ( .A1(n5099), .A2(n5273), .ZN(n5114) );
  NOR2_X1 U5754 ( .A1(n5629), .A2(n7580), .ZN(n5371) );
  INV_X1 U5755 ( .A(n5371), .ZN(n5106) );
  INV_X1 U5756 ( .A(n5100), .ZN(n5101) );
  NAND2_X1 U5757 ( .A1(n6066), .A2(n5415), .ZN(n5574) );
  NOR2_X2 U5758 ( .A1(n5417), .A2(n5574), .ZN(n5659) );
  INV_X1 U5759 ( .A(n5659), .ZN(n5104) );
  NOR2_X1 U5760 ( .A1(n5417), .A2(n6066), .ZN(n5396) );
  NAND2_X1 U5761 ( .A1(n5396), .A2(n7557), .ZN(n5674) );
  AOI21_X1 U5762 ( .B1(n5104), .B2(n5674), .A(n7520), .ZN(n5105) );
  AOI21_X1 U5763 ( .B1(n5107), .B2(n5106), .A(n5105), .ZN(n5109) );
  NAND2_X1 U5764 ( .A1(n7188), .A2(n7455), .ZN(n7514) );
  INV_X1 U5765 ( .A(n6039), .ZN(n5108) );
  OR2_X1 U5766 ( .A1(n5113), .A2(n7188), .ZN(n6931) );
  NAND2_X1 U5767 ( .A1(n5413), .A2(n6931), .ZN(n5395) );
  NOR2_X1 U5768 ( .A1(n5109), .A2(n5395), .ZN(n5110) );
  OR2_X1 U5769 ( .A1(n5387), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5912)
         );
  NAND2_X1 U5770 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5912), .ZN(n5908) );
  OAI211_X1 U5771 ( .C1(n5257), .C2(n7508), .A(n5110), .B(n5908), .ZN(n5111)
         );
  INV_X1 U5772 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5118) );
  AND2_X1 U5773 ( .A1(n7165), .A2(DATAI_31_), .ZN(n7651) );
  INV_X1 U5774 ( .A(n7651), .ZN(n5940) );
  AND2_X1 U5775 ( .A1(n7165), .A2(DATAI_23_), .ZN(n7654) );
  INV_X1 U5776 ( .A(DATAI_7_), .ZN(n6672) );
  OR2_X1 U5777 ( .A1(n5097), .A2(n7580), .ZN(n6935) );
  NAND2_X1 U5778 ( .A1(n5113), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5412) );
  OAI22_X1 U5779 ( .A1(n6935), .A2(n5114), .B1(n5912), .B2(n5412), .ZN(n5254)
         );
  AOI22_X1 U5780 ( .A1(n5659), .A2(n7654), .B1(n6973), .B2(n5254), .ZN(n5115)
         );
  OAI21_X1 U5781 ( .B1(n5940), .B2(n5674), .A(n5115), .ZN(n5116) );
  AOI21_X1 U5782 ( .B1(n7650), .B2(n5257), .A(n5116), .ZN(n5117) );
  OAI21_X1 U5783 ( .B1(n5260), .B2(n5118), .A(n5117), .ZN(U3075) );
  CLKBUF_X1 U5784 ( .A(n5119), .Z(n5120) );
  AND2_X1 U5785 ( .A1(n5089), .A2(n5121), .ZN(n5122) );
  NOR2_X1 U5786 ( .A1(n5120), .A2(n5122), .ZN(n5787) );
  INV_X1 U5787 ( .A(n5787), .ZN(n5847) );
  CLKBUF_X1 U5788 ( .A(n5123), .Z(n5265) );
  NAND2_X1 U5789 ( .A1(n5092), .A2(n5124), .ZN(n5125) );
  NAND2_X1 U5790 ( .A1(n5265), .A2(n5125), .ZN(n5842) );
  INV_X1 U5791 ( .A(n5842), .ZN(n5126) );
  AOI22_X1 U5792 ( .A1(n7124), .A2(n5126), .B1(EBX_REG_8__SCAN_IN), .B2(n6636), 
        .ZN(n5127) );
  OAI21_X1 U5793 ( .B1(n5847), .B2(n6648), .A(n5127), .ZN(U2851) );
  NAND2_X1 U5794 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n7448), .ZN(n5162) );
  INV_X1 U5795 ( .A(n5128), .ZN(n5161) );
  NAND2_X1 U5796 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5130) );
  INV_X1 U5797 ( .A(n5130), .ZN(n5129) );
  MUX2_X1 U5798 ( .A(n5130), .B(n5129), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n5134) );
  CLKBUF_X1 U5799 ( .A(n5131), .Z(n5143) );
  INV_X1 U5800 ( .A(n5143), .ZN(n6060) );
  AOI211_X1 U5801 ( .C1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n6060), .A(n5132), .B(n5133), .ZN(n6918) );
  OAI22_X1 U5802 ( .A1(n5144), .A2(n5134), .B1(n5145), .B2(n6918), .ZN(n5141)
         );
  INV_X1 U5803 ( .A(n5135), .ZN(n5136) );
  NOR2_X1 U5804 ( .A1(n5137), .A2(n5136), .ZN(n5151) );
  MUX2_X1 U5805 ( .A(n5138), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5143), 
        .Z(n5139) );
  NOR3_X1 U5806 ( .A1(n5151), .A2(n5128), .A3(n5139), .ZN(n5140) );
  AOI211_X1 U5807 ( .C1(n5097), .C2(n7453), .A(n5141), .B(n5140), .ZN(n6919)
         );
  NAND2_X1 U5808 ( .A1(n7472), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5142) );
  OAI21_X1 U5809 ( .B1(n7472), .B2(n6919), .A(n5142), .ZN(n7479) );
  XNOR2_X1 U5810 ( .A(n5143), .B(n3646), .ZN(n5150) );
  NAND2_X1 U5811 ( .A1(n5099), .A2(n7453), .ZN(n5149) );
  INV_X1 U5812 ( .A(n5144), .ZN(n7450) );
  XNOR2_X1 U5813 ( .A(n3646), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5147)
         );
  INV_X1 U5814 ( .A(n5145), .ZN(n5146) );
  AOI22_X1 U5815 ( .A1(n7450), .A2(n5147), .B1(n5146), .B2(n5150), .ZN(n5148)
         );
  OAI211_X1 U5816 ( .C1(n5151), .C2(n5150), .A(n5149), .B(n5148), .ZN(n6058)
         );
  MUX2_X1 U5817 ( .A(n6058), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(n7472), 
        .Z(n7467) );
  NAND3_X1 U5818 ( .A1(n7455), .A2(n7479), .A3(n7467), .ZN(n5160) );
  NAND2_X1 U5819 ( .A1(n7472), .A2(n7455), .ZN(n5152) );
  NAND2_X1 U5820 ( .A1(n5152), .A2(n5162), .ZN(n5159) );
  INV_X1 U5821 ( .A(n5153), .ZN(n5154) );
  OR2_X1 U5822 ( .A1(n5155), .A2(n5154), .ZN(n5156) );
  XNOR2_X1 U5823 ( .A(n5156), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n7461)
         );
  NOR2_X1 U5824 ( .A1(n7460), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5157) );
  AND2_X1 U5825 ( .A1(n7461), .A2(n5157), .ZN(n5158) );
  AOI21_X1 U5826 ( .B1(n5159), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n5158), 
        .ZN(n5164) );
  OAI211_X1 U5827 ( .C1(n5162), .C2(n5161), .A(n5160), .B(n5164), .ZN(n7489)
         );
  NAND2_X1 U5828 ( .A1(n5164), .A2(n5163), .ZN(n5165) );
  NAND2_X1 U5829 ( .A1(n7489), .A2(n5165), .ZN(n6040) );
  NAND2_X1 U5830 ( .A1(n6040), .A2(n7448), .ZN(n5167) );
  INV_X1 U5831 ( .A(n7507), .ZN(n5166) );
  NAND2_X1 U5832 ( .A1(n5167), .A2(n5166), .ZN(n5168) );
  INV_X1 U5833 ( .A(n6992), .ZN(n5173) );
  OAI21_X1 U5834 ( .B1(n7455), .B2(STATE2_REG_3__SCAN_IN), .A(n5173), .ZN(
        n6069) );
  NOR2_X1 U5835 ( .A1(n6992), .A2(n7580), .ZN(n6065) );
  INV_X1 U5836 ( .A(n6065), .ZN(n5174) );
  INV_X1 U5837 ( .A(n5417), .ZN(n5664) );
  NAND2_X1 U5838 ( .A1(n6066), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6064) );
  INV_X1 U5839 ( .A(n6064), .ZN(n5566) );
  NAND2_X1 U5840 ( .A1(n5664), .A2(n5566), .ZN(n5626) );
  OR2_X1 U5841 ( .A1(n5100), .A2(n6066), .ZN(n5170) );
  NOR2_X1 U5842 ( .A1(n5381), .A2(n5170), .ZN(n5383) );
  NAND2_X1 U5843 ( .A1(n5383), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5608) );
  NAND2_X1 U5844 ( .A1(n5626), .A2(n5608), .ZN(n5171) );
  OAI222_X1 U5845 ( .A1(n5173), .A2(n7480), .B1(n6069), .B2(n6608), .C1(n5174), 
        .C2(n5172), .ZN(U3462) );
  XNOR2_X1 U5846 ( .A(n5381), .B(n6064), .ZN(n5175) );
  INV_X1 U5847 ( .A(n5099), .ZN(n5741) );
  OAI222_X1 U5848 ( .A1(n5175), .A2(n5174), .B1(n6069), .B2(n5741), .C1(n5411), 
        .C2(n5173), .ZN(U3463) );
  AOI22_X1 U5849 ( .A1(n5176), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n5201), .ZN(n5178) );
  NAND2_X1 U5850 ( .A1(n5178), .A2(n5177), .ZN(U2926) );
  AOI22_X1 U5851 ( .A1(n5176), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n5201), .ZN(n5180) );
  NAND2_X1 U5852 ( .A1(n5180), .A2(n5179), .ZN(U2927) );
  AOI22_X1 U5853 ( .A1(n5176), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n5201), .ZN(n5182) );
  NAND2_X1 U5854 ( .A1(n5182), .A2(n5181), .ZN(U2928) );
  AOI22_X1 U5855 ( .A1(n5176), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n5201), .ZN(n5184) );
  NAND2_X1 U5856 ( .A1(n5184), .A2(n5183), .ZN(U2953) );
  AOI22_X1 U5857 ( .A1(n5176), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n5201), .ZN(n5186) );
  NAND2_X1 U5858 ( .A1(n5186), .A2(n5185), .ZN(U2930) );
  AOI22_X1 U5859 ( .A1(n5176), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n5201), .ZN(n5188) );
  NAND2_X1 U5860 ( .A1(n5188), .A2(n5187), .ZN(U2931) );
  AOI22_X1 U5861 ( .A1(n5176), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n5201), .ZN(n5190) );
  NAND2_X1 U5862 ( .A1(n5190), .A2(n5189), .ZN(U2932) );
  AOI22_X1 U5863 ( .A1(n5176), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n5201), .ZN(n5192) );
  NAND2_X1 U5864 ( .A1(n5192), .A2(n5191), .ZN(U2933) );
  AOI22_X1 U5865 ( .A1(n5176), .A2(UWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_26__SCAN_IN), .B2(n5201), .ZN(n5194) );
  NAND2_X1 U5866 ( .A1(n5194), .A2(n5193), .ZN(U2934) );
  AOI22_X1 U5867 ( .A1(n5176), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n5201), .ZN(n5196) );
  NAND2_X1 U5868 ( .A1(n5196), .A2(n5195), .ZN(U2929) );
  AOI22_X1 U5869 ( .A1(n5176), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n5201), .ZN(n5198) );
  NAND2_X1 U5870 ( .A1(n5198), .A2(n5197), .ZN(U2950) );
  AOI22_X1 U5871 ( .A1(n5176), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n5201), .ZN(n5200) );
  NAND2_X1 U5872 ( .A1(n5200), .A2(n5199), .ZN(U2951) );
  AOI22_X1 U5873 ( .A1(n5176), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n5201), .ZN(n5203) );
  NAND2_X1 U5874 ( .A1(n5203), .A2(n5202), .ZN(U2952) );
  INV_X1 U5875 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5207) );
  NOR2_X1 U5876 ( .A1(n5252), .A2(n4189), .ZN(n7637) );
  AND2_X1 U5877 ( .A1(n7165), .A2(DATAI_30_), .ZN(n7639) );
  INV_X1 U5878 ( .A(n7639), .ZN(n5920) );
  AND2_X1 U5879 ( .A1(n7165), .A2(DATAI_22_), .ZN(n7638) );
  AOI22_X1 U5880 ( .A1(n5659), .A2(n7638), .B1(n6966), .B2(n5254), .ZN(n5204)
         );
  OAI21_X1 U5881 ( .B1(n5920), .B2(n5674), .A(n5204), .ZN(n5205) );
  AOI21_X1 U5882 ( .B1(n7637), .B2(n5257), .A(n5205), .ZN(n5206) );
  OAI21_X1 U5883 ( .B1(n5260), .B2(n5207), .A(n5206), .ZN(U3074) );
  INV_X1 U5884 ( .A(EAX_REG_30__SCAN_IN), .ZN(n5209) );
  AOI22_X1 U5885 ( .A1(n7492), .A2(UWORD_REG_14__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5208) );
  OAI21_X1 U5886 ( .B1(n5209), .B2(n5217), .A(n5208), .ZN(U2893) );
  INV_X1 U5887 ( .A(EAX_REG_17__SCAN_IN), .ZN(n5220) );
  AOI22_X1 U5888 ( .A1(n7492), .A2(UWORD_REG_1__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5210) );
  OAI21_X1 U5889 ( .B1(n5220), .B2(n5217), .A(n5210), .ZN(U2906) );
  INV_X1 U5890 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5212) );
  AOI22_X1 U5891 ( .A1(n7492), .A2(UWORD_REG_2__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5211) );
  OAI21_X1 U5892 ( .B1(n5212), .B2(n5217), .A(n5211), .ZN(U2905) );
  INV_X1 U5893 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5214) );
  AOI22_X1 U5894 ( .A1(n7492), .A2(UWORD_REG_3__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5213) );
  OAI21_X1 U5895 ( .B1(n5214), .B2(n5217), .A(n5213), .ZN(U2904) );
  AOI22_X1 U5896 ( .A1(n7492), .A2(UWORD_REG_13__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n5215) );
  OAI21_X1 U5897 ( .B1(n4666), .B2(n5217), .A(n5215), .ZN(U2894) );
  AOI22_X1 U5898 ( .A1(n7492), .A2(UWORD_REG_0__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5216) );
  OAI21_X1 U5899 ( .B1(n5223), .B2(n5217), .A(n5216), .ZN(U2907) );
  NAND2_X1 U5900 ( .A1(n5176), .A2(UWORD_REG_1__SCAN_IN), .ZN(n5219) );
  OAI211_X1 U5901 ( .C1(n5224), .C2(n5220), .A(n5219), .B(n5218), .ZN(U2925)
         );
  NAND2_X1 U5902 ( .A1(n5176), .A2(UWORD_REG_0__SCAN_IN), .ZN(n5222) );
  OAI211_X1 U5903 ( .C1(n5224), .C2(n5223), .A(n5222), .B(n5221), .ZN(U2924)
         );
  INV_X1 U5904 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5229) );
  NOR2_X1 U5905 ( .A1(n5252), .A2(n5225), .ZN(n7621) );
  AND2_X1 U5906 ( .A1(n7165), .A2(DATAI_28_), .ZN(n7623) );
  INV_X1 U5907 ( .A(n7623), .ZN(n5925) );
  AND2_X1 U5908 ( .A1(n7165), .A2(DATAI_20_), .ZN(n7622) );
  AOI22_X1 U5909 ( .A1(n5659), .A2(n7622), .B1(n6956), .B2(n5254), .ZN(n5226)
         );
  OAI21_X1 U5910 ( .B1(n5925), .B2(n5674), .A(n5226), .ZN(n5227) );
  AOI21_X1 U5911 ( .B1(n7621), .B2(n5257), .A(n5227), .ZN(n5228) );
  OAI21_X1 U5912 ( .B1(n5260), .B2(n5229), .A(n5228), .ZN(U3072) );
  INV_X1 U5913 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5235) );
  AND2_X1 U5914 ( .A1(n7165), .A2(DATAI_26_), .ZN(n7607) );
  INV_X1 U5915 ( .A(n7607), .ZN(n5935) );
  AND2_X1 U5916 ( .A1(n7165), .A2(DATAI_18_), .ZN(n7606) );
  AOI22_X1 U5917 ( .A1(n5659), .A2(n7606), .B1(n6946), .B2(n5254), .ZN(n5232)
         );
  OAI21_X1 U5918 ( .B1(n5935), .B2(n5674), .A(n5232), .ZN(n5233) );
  AOI21_X1 U5919 ( .B1(n7605), .B2(n5257), .A(n5233), .ZN(n5234) );
  OAI21_X1 U5920 ( .B1(n5260), .B2(n5235), .A(n5234), .ZN(U3070) );
  INV_X1 U5921 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5240) );
  AND2_X1 U5922 ( .A1(n7165), .A2(DATAI_29_), .ZN(n7631) );
  INV_X1 U5923 ( .A(n7631), .ZN(n5915) );
  AND2_X1 U5924 ( .A1(n7165), .A2(DATAI_21_), .ZN(n7630) );
  AOI22_X1 U5925 ( .A1(n5659), .A2(n7630), .B1(n6961), .B2(n5254), .ZN(n5237)
         );
  OAI21_X1 U5926 ( .B1(n5915), .B2(n5674), .A(n5237), .ZN(n5238) );
  AOI21_X1 U5927 ( .B1(n7629), .B2(n5257), .A(n5238), .ZN(n5239) );
  OAI21_X1 U5928 ( .B1(n5260), .B2(n5240), .A(n5239), .ZN(U3073) );
  INV_X1 U5929 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5245) );
  AND2_X1 U5930 ( .A1(n7165), .A2(DATAI_27_), .ZN(n7614) );
  INV_X1 U5931 ( .A(n7614), .ZN(n5930) );
  AND2_X1 U5932 ( .A1(n7165), .A2(DATAI_19_), .ZN(n7615) );
  AOI22_X1 U5933 ( .A1(n5659), .A2(n7615), .B1(n6951), .B2(n5254), .ZN(n5242)
         );
  OAI21_X1 U5934 ( .B1(n5930), .B2(n5674), .A(n5242), .ZN(n5243) );
  AOI21_X1 U5935 ( .B1(n7613), .B2(n5257), .A(n5243), .ZN(n5244) );
  OAI21_X1 U5936 ( .B1(n5260), .B2(n5245), .A(n5244), .ZN(U3071) );
  INV_X1 U5937 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5250) );
  NOR2_X1 U5938 ( .A1(n5252), .A2(n3820), .ZN(n7597) );
  AND2_X1 U5939 ( .A1(n7165), .A2(DATAI_25_), .ZN(n7598) );
  INV_X1 U5940 ( .A(n7598), .ZN(n5952) );
  AND2_X1 U5941 ( .A1(n7165), .A2(DATAI_17_), .ZN(n7599) );
  AOI22_X1 U5942 ( .A1(n5659), .A2(n7599), .B1(n6941), .B2(n5254), .ZN(n5247)
         );
  OAI21_X1 U5943 ( .B1(n5952), .B2(n5674), .A(n5247), .ZN(n5248) );
  AOI21_X1 U5944 ( .B1(n7597), .B2(n5257), .A(n5248), .ZN(n5249) );
  OAI21_X1 U5945 ( .B1(n5260), .B2(n5250), .A(n5249), .ZN(U3069) );
  INV_X1 U5946 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5259) );
  NOR2_X1 U5947 ( .A1(n5252), .A2(n3650), .ZN(n7582) );
  AND2_X1 U5948 ( .A1(n7165), .A2(DATAI_24_), .ZN(n7583) );
  INV_X1 U5949 ( .A(n7583), .ZN(n5945) );
  AND2_X1 U5950 ( .A1(n7165), .A2(DATAI_16_), .ZN(n7591) );
  AOI22_X1 U5951 ( .A1(n5659), .A2(n7591), .B1(n6936), .B2(n5254), .ZN(n5255)
         );
  OAI21_X1 U5952 ( .B1(n5945), .B2(n5674), .A(n5255), .ZN(n5256) );
  AOI21_X1 U5953 ( .B1(n7582), .B2(n5257), .A(n5256), .ZN(n5258) );
  OAI21_X1 U5954 ( .B1(n5260), .B2(n5259), .A(n5258), .ZN(U3068) );
  OAI222_X1 U5955 ( .A1(n5848), .A2(n6672), .B1(n6085), .B2(n4250), .C1(n6669), 
        .C2(n5261), .ZN(U2884) );
  NOR2_X1 U5956 ( .A1(n5120), .A2(n5262), .ZN(n5263) );
  OR2_X1 U5957 ( .A1(n5515), .A2(n5263), .ZN(n7338) );
  INV_X1 U5958 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5268) );
  INV_X1 U5959 ( .A(n5518), .ZN(n5267) );
  NAND2_X1 U5960 ( .A1(n5265), .A2(n5264), .ZN(n5266) );
  NAND2_X1 U5961 ( .A1(n5267), .A2(n5266), .ZN(n7251) );
  OAI222_X1 U5962 ( .A1(n7338), .A2(n6648), .B1(n5268), .B2(n7126), .C1(n6647), 
        .C2(n7251), .ZN(U2850) );
  INV_X1 U5963 ( .A(DATAI_8_), .ZN(n5269) );
  INV_X1 U5964 ( .A(EAX_REG_8__SCAN_IN), .ZN(n7010) );
  OAI222_X1 U5965 ( .A1(n5848), .A2(n5269), .B1(n6085), .B2(n7010), .C1(n6669), 
        .C2(n5847), .ZN(U2883) );
  NAND2_X1 U5966 ( .A1(n7480), .A2(n5411), .ZN(n6922) );
  INV_X1 U5967 ( .A(n6922), .ZN(n5567) );
  NAND2_X1 U5968 ( .A1(n5567), .A2(n7474), .ZN(n5270) );
  NOR2_X1 U5969 ( .A1(n7576), .A2(n5270), .ZN(n5278) );
  INV_X1 U5970 ( .A(n5278), .ZN(n5302) );
  NAND2_X1 U5971 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5270), .ZN(n5279) );
  NAND2_X1 U5972 ( .A1(n5573), .A2(n5663), .ZN(n5282) );
  AOI21_X1 U5973 ( .B1(n5282), .B2(n7188), .A(n5272), .ZN(n5274) );
  OR2_X1 U5974 ( .A1(n5097), .A2(n6045), .ZN(n5627) );
  OR2_X1 U5975 ( .A1(n5099), .A2(n5273), .ZN(n6934) );
  NOR2_X1 U5976 ( .A1(n5627), .A2(n6934), .ZN(n5277) );
  NOR2_X1 U5977 ( .A1(n5274), .A2(n5277), .ZN(n5275) );
  OAI21_X1 U5978 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5275), .A(n5302), .ZN(
        n5276) );
  NAND3_X1 U5979 ( .A1(n5413), .A2(n5279), .A3(n5276), .ZN(n5299) );
  OAI21_X1 U5980 ( .B1(n5278), .B2(n5277), .A(n7508), .ZN(n5281) );
  INV_X1 U5981 ( .A(n5279), .ZN(n5280) );
  AOI21_X1 U5982 ( .B1(n7188), .B2(n5281), .A(n5280), .ZN(n5298) );
  AOI22_X1 U5983 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5299), .B1(n6946), 
        .B2(n5298), .ZN(n5285) );
  INV_X1 U5984 ( .A(n5282), .ZN(n5283) );
  AOI22_X1 U5985 ( .A1(n5911), .A2(n7606), .B1(n6976), .B2(n7607), .ZN(n5284)
         );
  OAI211_X1 U5986 ( .C1(n5302), .C2(n5683), .A(n5285), .B(n5284), .ZN(U3030)
         );
  AOI22_X1 U5987 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5299), .B1(n6956), 
        .B2(n5298), .ZN(n5287) );
  AOI22_X1 U5988 ( .A1(n5911), .A2(n7622), .B1(n6976), .B2(n7623), .ZN(n5286)
         );
  OAI211_X1 U5989 ( .C1(n5302), .C2(n5692), .A(n5287), .B(n5286), .ZN(U3032)
         );
  AOI22_X1 U5990 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5299), .B1(n6961), 
        .B2(n5298), .ZN(n5289) );
  AOI22_X1 U5991 ( .A1(n5911), .A2(n7630), .B1(n6976), .B2(n7631), .ZN(n5288)
         );
  OAI211_X1 U5992 ( .C1(n5302), .C2(n5689), .A(n5289), .B(n5288), .ZN(U3033)
         );
  AOI22_X1 U5993 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5299), .B1(n6973), 
        .B2(n5298), .ZN(n5291) );
  AOI22_X1 U5994 ( .A1(n5911), .A2(n7654), .B1(n6976), .B2(n7651), .ZN(n5290)
         );
  OAI211_X1 U5995 ( .C1(n5302), .C2(n5695), .A(n5291), .B(n5290), .ZN(U3035)
         );
  AOI22_X1 U5996 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5299), .B1(n6936), 
        .B2(n5298), .ZN(n5293) );
  AOI22_X1 U5997 ( .A1(n5911), .A2(n7591), .B1(n6976), .B2(n7583), .ZN(n5292)
         );
  OAI211_X1 U5998 ( .C1(n5302), .C2(n5703), .A(n5293), .B(n5292), .ZN(U3028)
         );
  AOI22_X1 U5999 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5299), .B1(n6951), 
        .B2(n5298), .ZN(n5295) );
  AOI22_X1 U6000 ( .A1(n5911), .A2(n7615), .B1(n6976), .B2(n7614), .ZN(n5294)
         );
  OAI211_X1 U6001 ( .C1(n5302), .C2(n5677), .A(n5295), .B(n5294), .ZN(U3031)
         );
  AOI22_X1 U6002 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5299), .B1(n6966), 
        .B2(n5298), .ZN(n5297) );
  AOI22_X1 U6003 ( .A1(n5911), .A2(n7638), .B1(n6976), .B2(n7639), .ZN(n5296)
         );
  OAI211_X1 U6004 ( .C1(n5302), .C2(n5686), .A(n5297), .B(n5296), .ZN(U3034)
         );
  AOI22_X1 U6005 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5299), .B1(n6941), 
        .B2(n5298), .ZN(n5301) );
  AOI22_X1 U6006 ( .A1(n5911), .A2(n7599), .B1(n6976), .B2(n7598), .ZN(n5300)
         );
  OAI211_X1 U6007 ( .C1(n5302), .C2(n5680), .A(n5301), .B(n5300), .ZN(U3029)
         );
  AND2_X1 U6008 ( .A1(n5097), .A2(n7454), .ZN(n7574) );
  AND2_X1 U6009 ( .A1(n5304), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5341)
         );
  AOI21_X1 U6010 ( .B1(n7574), .B2(n5629), .A(n5341), .ZN(n5309) );
  OR2_X1 U6011 ( .A1(n5663), .A2(n5100), .ZN(n5305) );
  NOR2_X1 U6012 ( .A1(n5381), .A2(n5305), .ZN(n5308) );
  NAND2_X1 U6013 ( .A1(n7590), .A2(n7520), .ZN(n7579) );
  OAI21_X1 U6014 ( .B1(n5308), .B2(n6797), .A(n7579), .ZN(n5306) );
  NAND3_X1 U6015 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5368) );
  AOI22_X1 U6016 ( .A1(n5309), .A2(n5306), .B1(n7580), .B2(n5368), .ZN(n5307)
         );
  INV_X1 U6017 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U6018 ( .A1(n5308), .A2(n5415), .ZN(n5369) );
  OAI22_X1 U6019 ( .A1(n5309), .A2(n7580), .B1(n5368), .B2(n7188), .ZN(n5338)
         );
  AOI22_X1 U6020 ( .A1(n6974), .A2(n7630), .B1(n6961), .B2(n5338), .ZN(n5310)
         );
  OAI21_X1 U6021 ( .B1(n5915), .B2(n5369), .A(n5310), .ZN(n5311) );
  AOI21_X1 U6022 ( .B1(n7629), .B2(n5341), .A(n5311), .ZN(n5312) );
  OAI21_X1 U6023 ( .B1(n5344), .B2(n5313), .A(n5312), .ZN(U3145) );
  INV_X1 U6024 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n5317) );
  AOI22_X1 U6025 ( .A1(n6974), .A2(n7591), .B1(n6936), .B2(n5338), .ZN(n5314)
         );
  OAI21_X1 U6026 ( .B1(n5945), .B2(n5369), .A(n5314), .ZN(n5315) );
  AOI21_X1 U6027 ( .B1(n7582), .B2(n5341), .A(n5315), .ZN(n5316) );
  OAI21_X1 U6028 ( .B1(n5344), .B2(n5317), .A(n5316), .ZN(U3140) );
  INV_X1 U6029 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5321) );
  AOI22_X1 U6030 ( .A1(n6974), .A2(n7606), .B1(n6946), .B2(n5338), .ZN(n5318)
         );
  OAI21_X1 U6031 ( .B1(n5935), .B2(n5369), .A(n5318), .ZN(n5319) );
  AOI21_X1 U6032 ( .B1(n7605), .B2(n5341), .A(n5319), .ZN(n5320) );
  OAI21_X1 U6033 ( .B1(n5344), .B2(n5321), .A(n5320), .ZN(U3142) );
  INV_X1 U6034 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5325) );
  AOI22_X1 U6035 ( .A1(n6974), .A2(n7638), .B1(n6966), .B2(n5338), .ZN(n5322)
         );
  OAI21_X1 U6036 ( .B1(n5920), .B2(n5369), .A(n5322), .ZN(n5323) );
  AOI21_X1 U6037 ( .B1(n7637), .B2(n5341), .A(n5323), .ZN(n5324) );
  OAI21_X1 U6038 ( .B1(n5344), .B2(n5325), .A(n5324), .ZN(U3146) );
  INV_X1 U6039 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5329) );
  AOI22_X1 U6040 ( .A1(n6974), .A2(n7622), .B1(n6956), .B2(n5338), .ZN(n5326)
         );
  OAI21_X1 U6041 ( .B1(n5925), .B2(n5369), .A(n5326), .ZN(n5327) );
  AOI21_X1 U6042 ( .B1(n7621), .B2(n5341), .A(n5327), .ZN(n5328) );
  OAI21_X1 U6043 ( .B1(n5344), .B2(n5329), .A(n5328), .ZN(U3144) );
  INV_X1 U6044 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5333) );
  AOI22_X1 U6045 ( .A1(n6974), .A2(n7599), .B1(n6941), .B2(n5338), .ZN(n5330)
         );
  OAI21_X1 U6046 ( .B1(n5952), .B2(n5369), .A(n5330), .ZN(n5331) );
  AOI21_X1 U6047 ( .B1(n7597), .B2(n5341), .A(n5331), .ZN(n5332) );
  OAI21_X1 U6048 ( .B1(n5344), .B2(n5333), .A(n5332), .ZN(U3141) );
  INV_X1 U6049 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5337) );
  AOI22_X1 U6050 ( .A1(n6974), .A2(n7615), .B1(n6951), .B2(n5338), .ZN(n5334)
         );
  OAI21_X1 U6051 ( .B1(n5930), .B2(n5369), .A(n5334), .ZN(n5335) );
  AOI21_X1 U6052 ( .B1(n7613), .B2(n5341), .A(n5335), .ZN(n5336) );
  OAI21_X1 U6053 ( .B1(n5344), .B2(n5337), .A(n5336), .ZN(U3143) );
  INV_X1 U6054 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5343) );
  AOI22_X1 U6055 ( .A1(n6974), .A2(n7654), .B1(n6973), .B2(n5338), .ZN(n5339)
         );
  OAI21_X1 U6056 ( .B1(n5940), .B2(n5369), .A(n5339), .ZN(n5340) );
  AOI21_X1 U6057 ( .B1(n7650), .B2(n5341), .A(n5340), .ZN(n5342) );
  OAI21_X1 U6058 ( .B1(n5344), .B2(n5343), .A(n5342), .ZN(U3147) );
  CLKBUF_X1 U6059 ( .A(n5345), .Z(n5346) );
  XNOR2_X1 U6060 ( .A(n5346), .B(n5347), .ZN(n5789) );
  NOR2_X1 U6061 ( .A1(n5348), .A2(n7218), .ZN(n7240) );
  AOI21_X1 U6062 ( .B1(n4780), .B2(n4075), .A(n7245), .ZN(n5357) );
  AOI21_X1 U6063 ( .B1(n5353), .B2(n5352), .A(n5351), .ZN(n5354) );
  NAND2_X1 U6064 ( .A1(n3665), .A2(n5354), .ZN(n5364) );
  INV_X1 U6065 ( .A(n5364), .ZN(n7244) );
  NOR2_X1 U6066 ( .A1(n7244), .A2(n4780), .ZN(n5356) );
  NAND2_X1 U6067 ( .A1(n7276), .A2(REIP_REG_8__SCAN_IN), .ZN(n5785) );
  OAI21_X1 U6068 ( .B1(n7212), .B2(n5842), .A(n5785), .ZN(n5355) );
  AOI211_X1 U6069 ( .C1(n7240), .C2(n5357), .A(n5356), .B(n5355), .ZN(n5358)
         );
  OAI21_X1 U6070 ( .B1(n5789), .B2(n6892), .A(n5358), .ZN(U3010) );
  INV_X1 U6071 ( .A(DATAI_9_), .ZN(n5359) );
  INV_X1 U6072 ( .A(EAX_REG_9__SCAN_IN), .ZN(n7012) );
  OAI222_X1 U6073 ( .A1(n5848), .A2(n5359), .B1(n6085), .B2(n7012), .C1(n6669), 
        .C2(n7338), .ZN(U2882) );
  CLKBUF_X1 U6074 ( .A(n5360), .Z(n5361) );
  XNOR2_X1 U6075 ( .A(n5361), .B(n5362), .ZN(n5775) );
  INV_X1 U6076 ( .A(REIP_REG_7__SCAN_IN), .ZN(n5363) );
  NOR2_X1 U6077 ( .A1(n7211), .A2(n5363), .ZN(n5771) );
  AOI22_X1 U6078 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n5364), .B1(n7240), 
        .B2(n4075), .ZN(n5365) );
  INV_X1 U6079 ( .A(n5365), .ZN(n5366) );
  AOI211_X1 U6080 ( .C1(n7269), .C2(n7322), .A(n5771), .B(n5366), .ZN(n5367)
         );
  OAI21_X1 U6081 ( .B1(n5775), .B2(n6892), .A(n5367), .ZN(U3011) );
  OR2_X1 U6082 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5368), .ZN(n5491)
         );
  NOR2_X1 U6083 ( .A1(n5387), .A2(n7480), .ZN(n7560) );
  NOR2_X1 U6084 ( .A1(n7560), .A2(n7188), .ZN(n7566) );
  AOI211_X1 U6085 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5491), .A(n7566), .B(
        n5395), .ZN(n5373) );
  OAI21_X1 U6086 ( .B1(n5488), .B2(n5639), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5370) );
  OAI21_X1 U6087 ( .B1(n5419), .B2(n5371), .A(n5370), .ZN(n5372) );
  NAND2_X1 U6088 ( .A1(n5373), .A2(n5372), .ZN(n5484) );
  NAND2_X1 U6089 ( .A1(n5484), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5376)
         );
  INV_X1 U6090 ( .A(n5412), .ZN(n5402) );
  AOI22_X1 U6091 ( .A1(n6927), .A2(n5629), .B1(n5402), .B2(n7560), .ZN(n5485)
         );
  OAI22_X1 U6092 ( .A1(n5486), .A2(n5940), .B1(n5485), .B2(n7658), .ZN(n5374)
         );
  AOI21_X1 U6093 ( .B1(n7654), .B2(n5488), .A(n5374), .ZN(n5375) );
  OAI211_X1 U6094 ( .C1(n5491), .C2(n5695), .A(n5376), .B(n5375), .ZN(U3139)
         );
  NAND2_X1 U6095 ( .A1(n5484), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5379)
         );
  OAI22_X1 U6096 ( .A1(n5486), .A2(n5920), .B1(n5485), .B2(n7642), .ZN(n5377)
         );
  AOI21_X1 U6097 ( .B1(n7638), .B2(n5488), .A(n5377), .ZN(n5378) );
  OAI211_X1 U6098 ( .C1(n5491), .C2(n5686), .A(n5379), .B(n5378), .ZN(U3138)
         );
  NOR3_X1 U6099 ( .A1(n5411), .A2(n7480), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5607) );
  NAND2_X1 U6100 ( .A1(n7576), .A2(n5607), .ZN(n5513) );
  AOI21_X1 U6101 ( .B1(n5387), .B2(n5423), .A(n7188), .ZN(n5414) );
  AOI211_X1 U6102 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5513), .A(n5414), .B(
        n5395), .ZN(n5386) );
  AND2_X1 U6103 ( .A1(n5099), .A2(n3648), .ZN(n5667) );
  NOR2_X1 U6104 ( .A1(n5667), .A2(n7580), .ZN(n5399) );
  INV_X1 U6105 ( .A(n5169), .ZN(n5382) );
  NAND2_X1 U6106 ( .A1(n6066), .A2(n7557), .ZN(n5416) );
  INV_X1 U6107 ( .A(n5416), .ZN(n5380) );
  NAND2_X1 U6108 ( .A1(n5381), .A2(n5380), .ZN(n5397) );
  OAI21_X1 U6109 ( .B1(n5462), .B2(n5640), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5384) );
  OAI21_X1 U6110 ( .B1(n5419), .B2(n5399), .A(n5384), .ZN(n5385) );
  NAND2_X1 U6111 ( .A1(n5386), .A2(n5385), .ZN(n5507) );
  NAND2_X1 U6112 ( .A1(n5507), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5391)
         );
  INV_X1 U6113 ( .A(n5387), .ZN(n5422) );
  NOR2_X1 U6114 ( .A1(n5412), .A2(n5422), .ZN(n5388) );
  AOI22_X1 U6115 ( .A1(n6927), .A2(n5667), .B1(n5388), .B2(n5423), .ZN(n5508)
         );
  OAI22_X1 U6116 ( .A1(n5509), .A2(n5920), .B1(n5508), .B2(n7642), .ZN(n5389)
         );
  AOI21_X1 U6117 ( .B1(n7638), .B2(n5640), .A(n5389), .ZN(n5390) );
  OAI211_X1 U6118 ( .C1(n5513), .C2(n5686), .A(n5391), .B(n5390), .ZN(U3122)
         );
  NAND2_X1 U6119 ( .A1(n5507), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5394)
         );
  OAI22_X1 U6120 ( .A1(n5509), .A2(n5940), .B1(n5508), .B2(n7658), .ZN(n5392)
         );
  AOI21_X1 U6121 ( .B1(n7654), .B2(n5640), .A(n5392), .ZN(n5393) );
  OAI211_X1 U6122 ( .C1(n5513), .C2(n5695), .A(n5394), .B(n5393), .ZN(U3123)
         );
  NAND3_X1 U6123 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7480), .A3(n7474), .ZN(n5671) );
  OR2_X1 U6124 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5671), .ZN(n5542)
         );
  NOR2_X1 U6125 ( .A1(n5423), .A2(n5422), .ZN(n6932) );
  NOR2_X1 U6126 ( .A1(n6932), .A2(n7188), .ZN(n6924) );
  AOI211_X1 U6127 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5542), .A(n6924), .B(
        n5395), .ZN(n5401) );
  OR2_X1 U6128 ( .A1(n5169), .A2(n5397), .ZN(n5538) );
  OAI21_X1 U6129 ( .B1(n5698), .B2(n5597), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5398) );
  OAI21_X1 U6130 ( .B1(n6927), .B2(n5399), .A(n5398), .ZN(n5400) );
  NAND2_X1 U6131 ( .A1(n5401), .A2(n5400), .ZN(n5536) );
  NAND2_X1 U6132 ( .A1(n5536), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U6133 ( .A1(n5419), .A2(n5667), .ZN(n5404) );
  NAND2_X1 U6134 ( .A1(n6932), .A2(n5402), .ZN(n5403) );
  OAI22_X1 U6135 ( .A1(n5538), .A2(n5920), .B1(n5537), .B2(n7642), .ZN(n5405)
         );
  AOI21_X1 U6136 ( .B1(n7638), .B2(n5698), .A(n5405), .ZN(n5406) );
  OAI211_X1 U6137 ( .C1(n5542), .C2(n5686), .A(n5407), .B(n5406), .ZN(U3058)
         );
  NAND2_X1 U6138 ( .A1(n5536), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5410) );
  OAI22_X1 U6139 ( .A1(n5538), .A2(n5940), .B1(n5537), .B2(n7658), .ZN(n5408)
         );
  AOI21_X1 U6140 ( .B1(n7654), .B2(n5698), .A(n5408), .ZN(n5409) );
  OAI211_X1 U6141 ( .C1(n5542), .C2(n5695), .A(n5410), .B(n5409), .ZN(U3059)
         );
  NAND2_X1 U6142 ( .A1(n5411), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7575) );
  OR2_X1 U6143 ( .A1(n6923), .A2(n7575), .ZN(n5564) );
  NAND2_X1 U6144 ( .A1(n5413), .A2(n5412), .ZN(n7565) );
  AOI211_X1 U6145 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5564), .A(n5414), .B(
        n7565), .ZN(n5421) );
  INV_X1 U6146 ( .A(n6934), .ZN(n7573) );
  NOR2_X1 U6147 ( .A1(n7573), .A2(n7580), .ZN(n6928) );
  OAI21_X1 U6148 ( .B1(n7652), .B2(n5658), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5418) );
  OAI21_X1 U6149 ( .B1(n5419), .B2(n6928), .A(n5418), .ZN(n5420) );
  NAND2_X1 U6150 ( .A1(n5421), .A2(n5420), .ZN(n5558) );
  NAND2_X1 U6151 ( .A1(n5558), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5427) );
  INV_X1 U6152 ( .A(n5658), .ZN(n5560) );
  NOR2_X1 U6153 ( .A1(n6931), .A2(n5422), .ZN(n5424) );
  AOI22_X1 U6154 ( .A1(n6927), .A2(n7573), .B1(n5424), .B2(n5423), .ZN(n5559)
         );
  OAI22_X1 U6155 ( .A1(n5560), .A2(n5920), .B1(n5559), .B2(n7642), .ZN(n5425)
         );
  AOI21_X1 U6156 ( .B1(n7652), .B2(n7638), .A(n5425), .ZN(n5426) );
  OAI211_X1 U6157 ( .C1(n5564), .C2(n5686), .A(n5427), .B(n5426), .ZN(U3090)
         );
  NAND2_X1 U6158 ( .A1(n5558), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5430) );
  OAI22_X1 U6159 ( .A1(n5560), .A2(n5940), .B1(n5559), .B2(n7658), .ZN(n5428)
         );
  AOI21_X1 U6160 ( .B1(n7652), .B2(n7654), .A(n5428), .ZN(n5429) );
  OAI211_X1 U6161 ( .C1(n5564), .C2(n5695), .A(n5430), .B(n5429), .ZN(U3091)
         );
  INV_X1 U6162 ( .A(n7575), .ZN(n5431) );
  NAND2_X1 U6163 ( .A1(n5565), .A2(n5431), .ZN(n5468) );
  OR2_X1 U6164 ( .A1(n7474), .A2(n7575), .ZN(n7564) );
  INV_X1 U6165 ( .A(n7564), .ZN(n5436) );
  AOI21_X1 U6166 ( .B1(n5440), .B2(n5566), .A(n7580), .ZN(n5438) );
  OR2_X1 U6167 ( .A1(n5099), .A2(n3648), .ZN(n5913) );
  INV_X1 U6168 ( .A(n5913), .ZN(n5432) );
  AND2_X1 U6169 ( .A1(n5432), .A2(n5097), .ZN(n7570) );
  NAND2_X1 U6170 ( .A1(n7570), .A2(n7454), .ZN(n5433) );
  NAND2_X1 U6171 ( .A1(n5433), .A2(n5468), .ZN(n5437) );
  INV_X1 U6172 ( .A(n5437), .ZN(n5434) );
  NAND2_X1 U6173 ( .A1(n5438), .A2(n5434), .ZN(n5435) );
  OAI211_X1 U6174 ( .C1(n7590), .C2(n5436), .A(n5435), .B(n7587), .ZN(n5466)
         );
  AOI22_X1 U6175 ( .A1(n5438), .A2(n5437), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5436), .ZN(n5464) );
  INV_X1 U6176 ( .A(n5574), .ZN(n5439) );
  AOI22_X1 U6177 ( .A1(n7651), .A2(n7644), .B1(n5462), .B2(n7654), .ZN(n5441)
         );
  OAI21_X1 U6178 ( .B1(n5464), .B2(n7658), .A(n5441), .ZN(n5442) );
  AOI21_X1 U6179 ( .B1(INSTQUEUE_REG_11__7__SCAN_IN), .B2(n5466), .A(n5442), 
        .ZN(n5443) );
  OAI21_X1 U6180 ( .B1(n5695), .B2(n5468), .A(n5443), .ZN(U3115) );
  AOI22_X1 U6181 ( .A1(n7598), .A2(n7644), .B1(n5462), .B2(n7599), .ZN(n5444)
         );
  OAI21_X1 U6182 ( .B1(n5464), .B2(n7602), .A(n5444), .ZN(n5445) );
  AOI21_X1 U6183 ( .B1(INSTQUEUE_REG_11__1__SCAN_IN), .B2(n5466), .A(n5445), 
        .ZN(n5446) );
  OAI21_X1 U6184 ( .B1(n5680), .B2(n5468), .A(n5446), .ZN(U3109) );
  AOI22_X1 U6185 ( .A1(n7583), .A2(n7644), .B1(n5462), .B2(n7591), .ZN(n5447)
         );
  OAI21_X1 U6186 ( .B1(n5464), .B2(n7594), .A(n5447), .ZN(n5448) );
  AOI21_X1 U6187 ( .B1(INSTQUEUE_REG_11__0__SCAN_IN), .B2(n5466), .A(n5448), 
        .ZN(n5449) );
  OAI21_X1 U6188 ( .B1(n5703), .B2(n5468), .A(n5449), .ZN(U3108) );
  AOI22_X1 U6189 ( .A1(n7614), .A2(n7644), .B1(n5462), .B2(n7615), .ZN(n5450)
         );
  OAI21_X1 U6190 ( .B1(n5464), .B2(n7618), .A(n5450), .ZN(n5451) );
  AOI21_X1 U6191 ( .B1(INSTQUEUE_REG_11__3__SCAN_IN), .B2(n5466), .A(n5451), 
        .ZN(n5452) );
  OAI21_X1 U6192 ( .B1(n5677), .B2(n5468), .A(n5452), .ZN(U3111) );
  AOI22_X1 U6193 ( .A1(n7631), .A2(n7644), .B1(n5462), .B2(n7630), .ZN(n5453)
         );
  OAI21_X1 U6194 ( .B1(n5464), .B2(n7634), .A(n5453), .ZN(n5454) );
  AOI21_X1 U6195 ( .B1(INSTQUEUE_REG_11__5__SCAN_IN), .B2(n5466), .A(n5454), 
        .ZN(n5455) );
  OAI21_X1 U6196 ( .B1(n5689), .B2(n5468), .A(n5455), .ZN(U3113) );
  AOI22_X1 U6197 ( .A1(n7639), .A2(n7644), .B1(n5462), .B2(n7638), .ZN(n5456)
         );
  OAI21_X1 U6198 ( .B1(n5464), .B2(n7642), .A(n5456), .ZN(n5457) );
  AOI21_X1 U6199 ( .B1(INSTQUEUE_REG_11__6__SCAN_IN), .B2(n5466), .A(n5457), 
        .ZN(n5458) );
  OAI21_X1 U6200 ( .B1(n5686), .B2(n5468), .A(n5458), .ZN(U3114) );
  AOI22_X1 U6201 ( .A1(n7607), .A2(n7644), .B1(n5462), .B2(n7606), .ZN(n5459)
         );
  OAI21_X1 U6202 ( .B1(n5464), .B2(n7610), .A(n5459), .ZN(n5460) );
  AOI21_X1 U6203 ( .B1(INSTQUEUE_REG_11__2__SCAN_IN), .B2(n5466), .A(n5460), 
        .ZN(n5461) );
  OAI21_X1 U6204 ( .B1(n5683), .B2(n5468), .A(n5461), .ZN(U3110) );
  AOI22_X1 U6205 ( .A1(n7623), .A2(n7644), .B1(n5462), .B2(n7622), .ZN(n5463)
         );
  OAI21_X1 U6206 ( .B1(n5464), .B2(n7626), .A(n5463), .ZN(n5465) );
  AOI21_X1 U6207 ( .B1(INSTQUEUE_REG_11__4__SCAN_IN), .B2(n5466), .A(n5465), 
        .ZN(n5467) );
  OAI21_X1 U6208 ( .B1(n5692), .B2(n5468), .A(n5467), .ZN(U3112) );
  NAND2_X1 U6209 ( .A1(n5484), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5471)
         );
  OAI22_X1 U6210 ( .A1(n5486), .A2(n5925), .B1(n5485), .B2(n7626), .ZN(n5469)
         );
  AOI21_X1 U6211 ( .B1(n7622), .B2(n5488), .A(n5469), .ZN(n5470) );
  OAI211_X1 U6212 ( .C1(n5491), .C2(n5692), .A(n5471), .B(n5470), .ZN(U3136)
         );
  NAND2_X1 U6213 ( .A1(n5484), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5474)
         );
  OAI22_X1 U6214 ( .A1(n5486), .A2(n5945), .B1(n5485), .B2(n7594), .ZN(n5472)
         );
  AOI21_X1 U6215 ( .B1(n7591), .B2(n5488), .A(n5472), .ZN(n5473) );
  OAI211_X1 U6216 ( .C1(n5703), .C2(n5491), .A(n5474), .B(n5473), .ZN(U3132)
         );
  NAND2_X1 U6217 ( .A1(n5484), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5477)
         );
  OAI22_X1 U6218 ( .A1(n5486), .A2(n5930), .B1(n5485), .B2(n7618), .ZN(n5475)
         );
  AOI21_X1 U6219 ( .B1(n7615), .B2(n5488), .A(n5475), .ZN(n5476) );
  OAI211_X1 U6220 ( .C1(n5491), .C2(n5677), .A(n5477), .B(n5476), .ZN(U3135)
         );
  NAND2_X1 U6221 ( .A1(n5484), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5480)
         );
  OAI22_X1 U6222 ( .A1(n5486), .A2(n5952), .B1(n5485), .B2(n7602), .ZN(n5478)
         );
  AOI21_X1 U6223 ( .B1(n7599), .B2(n5488), .A(n5478), .ZN(n5479) );
  OAI211_X1 U6224 ( .C1(n5491), .C2(n5680), .A(n5480), .B(n5479), .ZN(U3133)
         );
  NAND2_X1 U6225 ( .A1(n5484), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5483)
         );
  OAI22_X1 U6226 ( .A1(n5486), .A2(n5935), .B1(n5485), .B2(n7610), .ZN(n5481)
         );
  AOI21_X1 U6227 ( .B1(n7606), .B2(n5488), .A(n5481), .ZN(n5482) );
  OAI211_X1 U6228 ( .C1(n5491), .C2(n5683), .A(n5483), .B(n5482), .ZN(U3134)
         );
  NAND2_X1 U6229 ( .A1(n5484), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5490)
         );
  OAI22_X1 U6230 ( .A1(n5486), .A2(n5915), .B1(n5485), .B2(n7634), .ZN(n5487)
         );
  AOI21_X1 U6231 ( .B1(n7630), .B2(n5488), .A(n5487), .ZN(n5489) );
  OAI211_X1 U6232 ( .C1(n5491), .C2(n5689), .A(n5490), .B(n5489), .ZN(U3137)
         );
  NAND2_X1 U6233 ( .A1(n5507), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5494)
         );
  OAI22_X1 U6234 ( .A1(n5509), .A2(n5925), .B1(n5508), .B2(n7626), .ZN(n5492)
         );
  AOI21_X1 U6235 ( .B1(n7622), .B2(n5640), .A(n5492), .ZN(n5493) );
  OAI211_X1 U6236 ( .C1(n5513), .C2(n5692), .A(n5494), .B(n5493), .ZN(U3120)
         );
  NAND2_X1 U6237 ( .A1(n5507), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5497)
         );
  OAI22_X1 U6238 ( .A1(n5509), .A2(n5945), .B1(n5508), .B2(n7594), .ZN(n5495)
         );
  AOI21_X1 U6239 ( .B1(n7591), .B2(n5640), .A(n5495), .ZN(n5496) );
  OAI211_X1 U6240 ( .C1(n5703), .C2(n5513), .A(n5497), .B(n5496), .ZN(U3116)
         );
  NAND2_X1 U6241 ( .A1(n5507), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5500)
         );
  OAI22_X1 U6242 ( .A1(n5509), .A2(n5935), .B1(n5508), .B2(n7610), .ZN(n5498)
         );
  AOI21_X1 U6243 ( .B1(n7606), .B2(n5640), .A(n5498), .ZN(n5499) );
  OAI211_X1 U6244 ( .C1(n5513), .C2(n5683), .A(n5500), .B(n5499), .ZN(U3118)
         );
  NAND2_X1 U6245 ( .A1(n5507), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5503)
         );
  OAI22_X1 U6246 ( .A1(n5509), .A2(n5915), .B1(n5508), .B2(n7634), .ZN(n5501)
         );
  AOI21_X1 U6247 ( .B1(n7630), .B2(n5640), .A(n5501), .ZN(n5502) );
  OAI211_X1 U6248 ( .C1(n5513), .C2(n5689), .A(n5503), .B(n5502), .ZN(U3121)
         );
  NAND2_X1 U6249 ( .A1(n5507), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5506)
         );
  OAI22_X1 U6250 ( .A1(n5509), .A2(n5952), .B1(n5508), .B2(n7602), .ZN(n5504)
         );
  AOI21_X1 U6251 ( .B1(n7599), .B2(n5640), .A(n5504), .ZN(n5505) );
  OAI211_X1 U6252 ( .C1(n5513), .C2(n5680), .A(n5506), .B(n5505), .ZN(U3117)
         );
  NAND2_X1 U6253 ( .A1(n5507), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5512)
         );
  OAI22_X1 U6254 ( .A1(n5509), .A2(n5930), .B1(n5508), .B2(n7618), .ZN(n5510)
         );
  AOI21_X1 U6255 ( .B1(n7615), .B2(n5640), .A(n5510), .ZN(n5511) );
  OAI211_X1 U6256 ( .C1(n5513), .C2(n5677), .A(n5512), .B(n5511), .ZN(U3119)
         );
  INV_X1 U6257 ( .A(n5799), .ZN(n5801) );
  OAI21_X1 U6258 ( .B1(n5515), .B2(n5514), .A(n5801), .ZN(n5836) );
  CLKBUF_X1 U6259 ( .A(n5516), .Z(n5861) );
  OAI21_X1 U6260 ( .B1(n5518), .B2(n5517), .A(n5861), .ZN(n5519) );
  INV_X1 U6261 ( .A(n5519), .ZN(n7243) );
  AOI22_X1 U6262 ( .A1(n7124), .A2(n7243), .B1(EBX_REG_10__SCAN_IN), .B2(n6636), .ZN(n5520) );
  OAI21_X1 U6263 ( .B1(n5836), .B2(n6648), .A(n5520), .ZN(U2849) );
  NAND2_X1 U6264 ( .A1(n5536), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5523) );
  OAI22_X1 U6265 ( .A1(n5538), .A2(n5925), .B1(n5537), .B2(n7626), .ZN(n5521)
         );
  AOI21_X1 U6266 ( .B1(n7622), .B2(n5698), .A(n5521), .ZN(n5522) );
  OAI211_X1 U6267 ( .C1(n5542), .C2(n5692), .A(n5523), .B(n5522), .ZN(U3056)
         );
  NAND2_X1 U6268 ( .A1(n5536), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5526) );
  OAI22_X1 U6269 ( .A1(n5538), .A2(n5945), .B1(n5537), .B2(n7594), .ZN(n5524)
         );
  AOI21_X1 U6270 ( .B1(n7591), .B2(n5698), .A(n5524), .ZN(n5525) );
  OAI211_X1 U6271 ( .C1(n5703), .C2(n5542), .A(n5526), .B(n5525), .ZN(U3052)
         );
  NAND2_X1 U6272 ( .A1(n5536), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5529) );
  OAI22_X1 U6273 ( .A1(n5538), .A2(n5935), .B1(n5537), .B2(n7610), .ZN(n5527)
         );
  AOI21_X1 U6274 ( .B1(n7606), .B2(n5698), .A(n5527), .ZN(n5528) );
  OAI211_X1 U6275 ( .C1(n5542), .C2(n5683), .A(n5529), .B(n5528), .ZN(U3054)
         );
  NAND2_X1 U6276 ( .A1(n5536), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5532) );
  OAI22_X1 U6277 ( .A1(n5538), .A2(n5930), .B1(n5537), .B2(n7618), .ZN(n5530)
         );
  AOI21_X1 U6278 ( .B1(n7615), .B2(n5698), .A(n5530), .ZN(n5531) );
  OAI211_X1 U6279 ( .C1(n5542), .C2(n5677), .A(n5532), .B(n5531), .ZN(U3055)
         );
  NAND2_X1 U6280 ( .A1(n5536), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5535) );
  OAI22_X1 U6281 ( .A1(n5538), .A2(n5952), .B1(n5537), .B2(n7602), .ZN(n5533)
         );
  AOI21_X1 U6282 ( .B1(n7599), .B2(n5698), .A(n5533), .ZN(n5534) );
  OAI211_X1 U6283 ( .C1(n5542), .C2(n5680), .A(n5535), .B(n5534), .ZN(U3053)
         );
  NAND2_X1 U6284 ( .A1(n5536), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5541) );
  OAI22_X1 U6285 ( .A1(n5538), .A2(n5915), .B1(n5537), .B2(n7634), .ZN(n5539)
         );
  AOI21_X1 U6286 ( .B1(n7630), .B2(n5698), .A(n5539), .ZN(n5540) );
  OAI211_X1 U6287 ( .C1(n5542), .C2(n5689), .A(n5541), .B(n5540), .ZN(U3057)
         );
  NAND2_X1 U6288 ( .A1(n5558), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5545) );
  OAI22_X1 U6289 ( .A1(n5560), .A2(n5925), .B1(n5559), .B2(n7626), .ZN(n5543)
         );
  AOI21_X1 U6290 ( .B1(n7652), .B2(n7622), .A(n5543), .ZN(n5544) );
  OAI211_X1 U6291 ( .C1(n5564), .C2(n5692), .A(n5545), .B(n5544), .ZN(U3088)
         );
  NAND2_X1 U6292 ( .A1(n5558), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5548) );
  OAI22_X1 U6293 ( .A1(n5560), .A2(n5945), .B1(n5559), .B2(n7594), .ZN(n5546)
         );
  AOI21_X1 U6294 ( .B1(n7652), .B2(n7591), .A(n5546), .ZN(n5547) );
  OAI211_X1 U6295 ( .C1(n5703), .C2(n5564), .A(n5548), .B(n5547), .ZN(U3084)
         );
  NAND2_X1 U6296 ( .A1(n5558), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5551) );
  OAI22_X1 U6297 ( .A1(n5560), .A2(n5935), .B1(n5559), .B2(n7610), .ZN(n5549)
         );
  AOI21_X1 U6298 ( .B1(n7652), .B2(n7606), .A(n5549), .ZN(n5550) );
  OAI211_X1 U6299 ( .C1(n5564), .C2(n5683), .A(n5551), .B(n5550), .ZN(U3086)
         );
  NAND2_X1 U6300 ( .A1(n5558), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5554) );
  OAI22_X1 U6301 ( .A1(n5560), .A2(n5930), .B1(n5559), .B2(n7618), .ZN(n5552)
         );
  AOI21_X1 U6302 ( .B1(n7652), .B2(n7615), .A(n5552), .ZN(n5553) );
  OAI211_X1 U6303 ( .C1(n5564), .C2(n5677), .A(n5554), .B(n5553), .ZN(U3087)
         );
  NAND2_X1 U6304 ( .A1(n5558), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5557) );
  OAI22_X1 U6305 ( .A1(n5560), .A2(n5952), .B1(n5559), .B2(n7602), .ZN(n5555)
         );
  AOI21_X1 U6306 ( .B1(n7652), .B2(n7599), .A(n5555), .ZN(n5556) );
  OAI211_X1 U6307 ( .C1(n5564), .C2(n5680), .A(n5557), .B(n5556), .ZN(U3085)
         );
  NAND2_X1 U6308 ( .A1(n5558), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5563) );
  OAI22_X1 U6309 ( .A1(n5560), .A2(n5915), .B1(n5559), .B2(n7634), .ZN(n5561)
         );
  AOI21_X1 U6310 ( .B1(n7652), .B2(n7630), .A(n5561), .ZN(n5562) );
  OAI211_X1 U6311 ( .C1(n5564), .C2(n5689), .A(n5563), .B(n5562), .ZN(U3089)
         );
  NAND2_X1 U6312 ( .A1(n5565), .A2(n5567), .ZN(n5603) );
  AOI21_X1 U6313 ( .B1(n5573), .B2(n5566), .A(n7580), .ZN(n5572) );
  INV_X1 U6314 ( .A(n5572), .ZN(n5569) );
  OAI21_X1 U6315 ( .B1(n5627), .B2(n5913), .A(n5603), .ZN(n5571) );
  NAND2_X1 U6316 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n5567), .ZN(n5906) );
  NAND2_X1 U6317 ( .A1(n5906), .A2(n7580), .ZN(n5568) );
  OAI211_X1 U6318 ( .C1(n5569), .C2(n5571), .A(n7587), .B(n5568), .ZN(n5601)
         );
  INV_X1 U6319 ( .A(n5906), .ZN(n5570) );
  AOI22_X1 U6320 ( .A1(n5572), .A2(n5571), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5570), .ZN(n5599) );
  INV_X1 U6321 ( .A(n5573), .ZN(n5575) );
  NOR2_X2 U6322 ( .A1(n5575), .A2(n5574), .ZN(n5950) );
  AOI22_X1 U6323 ( .A1(n5950), .A2(n7583), .B1(n7591), .B2(n5597), .ZN(n5576)
         );
  OAI21_X1 U6324 ( .B1(n5599), .B2(n7594), .A(n5576), .ZN(n5577) );
  AOI21_X1 U6325 ( .B1(INSTQUEUE_REG_3__0__SCAN_IN), .B2(n5601), .A(n5577), 
        .ZN(n5578) );
  OAI21_X1 U6326 ( .B1(n5703), .B2(n5603), .A(n5578), .ZN(U3044) );
  AOI22_X1 U6327 ( .A1(n5950), .A2(n7623), .B1(n7622), .B2(n5597), .ZN(n5579)
         );
  OAI21_X1 U6328 ( .B1(n5599), .B2(n7626), .A(n5579), .ZN(n5580) );
  AOI21_X1 U6329 ( .B1(INSTQUEUE_REG_3__4__SCAN_IN), .B2(n5601), .A(n5580), 
        .ZN(n5581) );
  OAI21_X1 U6330 ( .B1(n5692), .B2(n5603), .A(n5581), .ZN(U3048) );
  AOI22_X1 U6331 ( .A1(n5950), .A2(n7598), .B1(n7599), .B2(n5597), .ZN(n5582)
         );
  OAI21_X1 U6332 ( .B1(n5599), .B2(n7602), .A(n5582), .ZN(n5583) );
  AOI21_X1 U6333 ( .B1(INSTQUEUE_REG_3__1__SCAN_IN), .B2(n5601), .A(n5583), 
        .ZN(n5584) );
  OAI21_X1 U6334 ( .B1(n5680), .B2(n5603), .A(n5584), .ZN(U3045) );
  AOI22_X1 U6335 ( .A1(n5950), .A2(n7651), .B1(n7654), .B2(n5597), .ZN(n5585)
         );
  OAI21_X1 U6336 ( .B1(n5599), .B2(n7658), .A(n5585), .ZN(n5586) );
  AOI21_X1 U6337 ( .B1(INSTQUEUE_REG_3__7__SCAN_IN), .B2(n5601), .A(n5586), 
        .ZN(n5587) );
  OAI21_X1 U6338 ( .B1(n5695), .B2(n5603), .A(n5587), .ZN(U3051) );
  AOI22_X1 U6339 ( .A1(n5950), .A2(n7631), .B1(n7630), .B2(n5597), .ZN(n5588)
         );
  OAI21_X1 U6340 ( .B1(n5599), .B2(n7634), .A(n5588), .ZN(n5589) );
  AOI21_X1 U6341 ( .B1(INSTQUEUE_REG_3__5__SCAN_IN), .B2(n5601), .A(n5589), 
        .ZN(n5590) );
  OAI21_X1 U6342 ( .B1(n5689), .B2(n5603), .A(n5590), .ZN(U3049) );
  AOI22_X1 U6343 ( .A1(n5950), .A2(n7639), .B1(n7638), .B2(n5597), .ZN(n5591)
         );
  OAI21_X1 U6344 ( .B1(n5599), .B2(n7642), .A(n5591), .ZN(n5592) );
  AOI21_X1 U6345 ( .B1(INSTQUEUE_REG_3__6__SCAN_IN), .B2(n5601), .A(n5592), 
        .ZN(n5593) );
  OAI21_X1 U6346 ( .B1(n5686), .B2(n5603), .A(n5593), .ZN(U3050) );
  AOI22_X1 U6347 ( .A1(n5950), .A2(n7614), .B1(n7615), .B2(n5597), .ZN(n5594)
         );
  OAI21_X1 U6348 ( .B1(n5599), .B2(n7618), .A(n5594), .ZN(n5595) );
  AOI21_X1 U6349 ( .B1(INSTQUEUE_REG_3__3__SCAN_IN), .B2(n5601), .A(n5595), 
        .ZN(n5596) );
  OAI21_X1 U6350 ( .B1(n5677), .B2(n5603), .A(n5596), .ZN(U3047) );
  AOI22_X1 U6351 ( .A1(n5950), .A2(n7607), .B1(n7606), .B2(n5597), .ZN(n5598)
         );
  OAI21_X1 U6352 ( .B1(n5599), .B2(n7610), .A(n5598), .ZN(n5600) );
  AOI21_X1 U6353 ( .B1(INSTQUEUE_REG_3__2__SCAN_IN), .B2(n5601), .A(n5600), 
        .ZN(n5602) );
  OAI21_X1 U6354 ( .B1(n5683), .B2(n5603), .A(n5602), .ZN(U3046) );
  INV_X1 U6355 ( .A(DATAI_10_), .ZN(n5604) );
  INV_X1 U6356 ( .A(EAX_REG_10__SCAN_IN), .ZN(n7014) );
  OAI222_X1 U6357 ( .A1(n5848), .A2(n5604), .B1(n6085), .B2(n7014), .C1(n6669), 
        .C2(n5836), .ZN(U2881) );
  INV_X1 U6358 ( .A(n5607), .ZN(n5609) );
  NOR2_X1 U6359 ( .A1(n7576), .A2(n5609), .ZN(n5605) );
  INV_X1 U6360 ( .A(n5605), .ZN(n5643) );
  AOI21_X1 U6361 ( .B1(n7574), .B2(n5667), .A(n5605), .ZN(n5611) );
  NAND3_X1 U6362 ( .A1(n7590), .A2(n5611), .A3(n5608), .ZN(n5606) );
  OAI211_X1 U6363 ( .C1(n7590), .C2(n5607), .A(n7587), .B(n5606), .ZN(n5638)
         );
  NAND2_X1 U6364 ( .A1(n7590), .A2(n5608), .ZN(n5610) );
  OAI22_X1 U6365 ( .A1(n5611), .A2(n5610), .B1(n7188), .B2(n5609), .ZN(n5637)
         );
  AOI22_X1 U6366 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n5638), .B1(n6946), 
        .B2(n5637), .ZN(n5613) );
  AOI22_X1 U6367 ( .A1(n7607), .A2(n5640), .B1(n5639), .B2(n7606), .ZN(n5612)
         );
  OAI211_X1 U6368 ( .C1(n5683), .C2(n5643), .A(n5613), .B(n5612), .ZN(U3126)
         );
  AOI22_X1 U6369 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n5638), .B1(n6973), 
        .B2(n5637), .ZN(n5615) );
  AOI22_X1 U6370 ( .A1(n7651), .A2(n5640), .B1(n5639), .B2(n7654), .ZN(n5614)
         );
  OAI211_X1 U6371 ( .C1(n5695), .C2(n5643), .A(n5615), .B(n5614), .ZN(U3131)
         );
  AOI22_X1 U6372 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n5638), .B1(n6966), 
        .B2(n5637), .ZN(n5617) );
  AOI22_X1 U6373 ( .A1(n7639), .A2(n5640), .B1(n5639), .B2(n7638), .ZN(n5616)
         );
  OAI211_X1 U6374 ( .C1(n5686), .C2(n5643), .A(n5617), .B(n5616), .ZN(U3130)
         );
  AOI22_X1 U6375 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n5638), .B1(n6961), 
        .B2(n5637), .ZN(n5619) );
  AOI22_X1 U6376 ( .A1(n7631), .A2(n5640), .B1(n5639), .B2(n7630), .ZN(n5618)
         );
  OAI211_X1 U6377 ( .C1(n5689), .C2(n5643), .A(n5619), .B(n5618), .ZN(U3129)
         );
  AOI22_X1 U6378 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5638), .B1(n6936), 
        .B2(n5637), .ZN(n5621) );
  AOI22_X1 U6379 ( .A1(n7583), .A2(n5640), .B1(n5639), .B2(n7591), .ZN(n5620)
         );
  OAI211_X1 U6380 ( .C1(n5703), .C2(n5643), .A(n5621), .B(n5620), .ZN(U3124)
         );
  AOI22_X1 U6381 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5638), .B1(n6956), 
        .B2(n5637), .ZN(n5623) );
  AOI22_X1 U6382 ( .A1(n7623), .A2(n5640), .B1(n5639), .B2(n7622), .ZN(n5622)
         );
  OAI211_X1 U6383 ( .C1(n5692), .C2(n5643), .A(n5623), .B(n5622), .ZN(U3128)
         );
  AOI22_X1 U6384 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n5638), .B1(n6951), 
        .B2(n5637), .ZN(n5625) );
  AOI22_X1 U6385 ( .A1(n7614), .A2(n5640), .B1(n5639), .B2(n7615), .ZN(n5624)
         );
  OAI211_X1 U6386 ( .C1(n5677), .C2(n5643), .A(n5625), .B(n5624), .ZN(U3127)
         );
  NAND2_X1 U6387 ( .A1(n7590), .A2(n5626), .ZN(n5633) );
  INV_X1 U6388 ( .A(n5627), .ZN(n5668) );
  INV_X1 U6389 ( .A(n5662), .ZN(n5628) );
  AOI21_X1 U6390 ( .B1(n5668), .B2(n5629), .A(n5628), .ZN(n5634) );
  INV_X1 U6391 ( .A(n5634), .ZN(n5631) );
  NAND2_X1 U6392 ( .A1(n7580), .A2(n5632), .ZN(n5630) );
  OAI211_X1 U6393 ( .C1(n5633), .C2(n5631), .A(n7587), .B(n5630), .ZN(n5657)
         );
  OAI22_X1 U6394 ( .A1(n5634), .A2(n5633), .B1(n7188), .B2(n5632), .ZN(n5656)
         );
  AOI22_X1 U6395 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n5657), .B1(n6966), 
        .B2(n5656), .ZN(n5636) );
  AOI22_X1 U6396 ( .A1(n7639), .A2(n5659), .B1(n5658), .B2(n7638), .ZN(n5635)
         );
  OAI211_X1 U6397 ( .C1(n5662), .C2(n5686), .A(n5636), .B(n5635), .ZN(U3082)
         );
  AOI22_X1 U6398 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n5638), .B1(n6941), 
        .B2(n5637), .ZN(n5642) );
  AOI22_X1 U6399 ( .A1(n7598), .A2(n5640), .B1(n5639), .B2(n7599), .ZN(n5641)
         );
  OAI211_X1 U6400 ( .C1(n5680), .C2(n5643), .A(n5642), .B(n5641), .ZN(U3125)
         );
  AOI22_X1 U6401 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n5657), .B1(n6961), 
        .B2(n5656), .ZN(n5645) );
  AOI22_X1 U6402 ( .A1(n7631), .A2(n5659), .B1(n5658), .B2(n7630), .ZN(n5644)
         );
  OAI211_X1 U6403 ( .C1(n5662), .C2(n5689), .A(n5645), .B(n5644), .ZN(U3081)
         );
  AOI22_X1 U6404 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n5657), .B1(n6956), 
        .B2(n5656), .ZN(n5647) );
  AOI22_X1 U6405 ( .A1(n7623), .A2(n5659), .B1(n5658), .B2(n7622), .ZN(n5646)
         );
  OAI211_X1 U6406 ( .C1(n5662), .C2(n5692), .A(n5647), .B(n5646), .ZN(U3080)
         );
  AOI22_X1 U6407 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n5657), .B1(n6951), 
        .B2(n5656), .ZN(n5649) );
  AOI22_X1 U6408 ( .A1(n7614), .A2(n5659), .B1(n5658), .B2(n7615), .ZN(n5648)
         );
  OAI211_X1 U6409 ( .C1(n5662), .C2(n5677), .A(n5649), .B(n5648), .ZN(U3079)
         );
  AOI22_X1 U6410 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n5657), .B1(n6946), 
        .B2(n5656), .ZN(n5651) );
  AOI22_X1 U6411 ( .A1(n7607), .A2(n5659), .B1(n5658), .B2(n7606), .ZN(n5650)
         );
  OAI211_X1 U6412 ( .C1(n5662), .C2(n5683), .A(n5651), .B(n5650), .ZN(U3078)
         );
  AOI22_X1 U6413 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n5657), .B1(n6941), 
        .B2(n5656), .ZN(n5653) );
  AOI22_X1 U6414 ( .A1(n7598), .A2(n5659), .B1(n5658), .B2(n7599), .ZN(n5652)
         );
  OAI211_X1 U6415 ( .C1(n5662), .C2(n5680), .A(n5653), .B(n5652), .ZN(U3077)
         );
  AOI22_X1 U6416 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n5657), .B1(n6973), 
        .B2(n5656), .ZN(n5655) );
  AOI22_X1 U6417 ( .A1(n7651), .A2(n5659), .B1(n5658), .B2(n7654), .ZN(n5654)
         );
  OAI211_X1 U6418 ( .C1(n5662), .C2(n5695), .A(n5655), .B(n5654), .ZN(U3083)
         );
  AOI22_X1 U6419 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n5657), .B1(n6936), 
        .B2(n5656), .ZN(n5661) );
  AOI22_X1 U6420 ( .A1(n7583), .A2(n5659), .B1(n5658), .B2(n7591), .ZN(n5660)
         );
  OAI211_X1 U6421 ( .C1(n5662), .C2(n5703), .A(n5661), .B(n5660), .ZN(U3076)
         );
  NOR2_X1 U6422 ( .A1(n7576), .A2(n5671), .ZN(n5666) );
  INV_X1 U6423 ( .A(n5666), .ZN(n5702) );
  NAND3_X1 U6424 ( .A1(n5664), .A2(n5663), .A3(STATEBS16_REG_SCAN_IN), .ZN(
        n5665) );
  NAND2_X1 U6425 ( .A1(n5665), .A2(n7590), .ZN(n5672) );
  AOI21_X1 U6426 ( .B1(n5668), .B2(n5667), .A(n5666), .ZN(n5673) );
  INV_X1 U6427 ( .A(n5673), .ZN(n5670) );
  NAND2_X1 U6428 ( .A1(n7580), .A2(n5671), .ZN(n5669) );
  OAI211_X1 U6429 ( .C1(n5672), .C2(n5670), .A(n7587), .B(n5669), .ZN(n5697)
         );
  OAI22_X1 U6430 ( .A1(n5673), .A2(n5672), .B1(n7188), .B2(n5671), .ZN(n5696)
         );
  AOI22_X1 U6431 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n5697), .B1(n6951), 
        .B2(n5696), .ZN(n5676) );
  AOI22_X1 U6432 ( .A1(n5699), .A2(n7615), .B1(n5698), .B2(n7614), .ZN(n5675)
         );
  OAI211_X1 U6433 ( .C1(n5677), .C2(n5702), .A(n5676), .B(n5675), .ZN(U3063)
         );
  AOI22_X1 U6434 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n5697), .B1(n6941), 
        .B2(n5696), .ZN(n5679) );
  AOI22_X1 U6435 ( .A1(n5699), .A2(n7599), .B1(n5698), .B2(n7598), .ZN(n5678)
         );
  OAI211_X1 U6436 ( .C1(n5680), .C2(n5702), .A(n5679), .B(n5678), .ZN(U3061)
         );
  AOI22_X1 U6437 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n5697), .B1(n6946), 
        .B2(n5696), .ZN(n5682) );
  AOI22_X1 U6438 ( .A1(n5699), .A2(n7606), .B1(n5698), .B2(n7607), .ZN(n5681)
         );
  OAI211_X1 U6439 ( .C1(n5683), .C2(n5702), .A(n5682), .B(n5681), .ZN(U3062)
         );
  AOI22_X1 U6440 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n5697), .B1(n6966), 
        .B2(n5696), .ZN(n5685) );
  AOI22_X1 U6441 ( .A1(n5699), .A2(n7638), .B1(n5698), .B2(n7639), .ZN(n5684)
         );
  OAI211_X1 U6442 ( .C1(n5686), .C2(n5702), .A(n5685), .B(n5684), .ZN(U3066)
         );
  AOI22_X1 U6443 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n5697), .B1(n6961), 
        .B2(n5696), .ZN(n5688) );
  AOI22_X1 U6444 ( .A1(n5699), .A2(n7630), .B1(n5698), .B2(n7631), .ZN(n5687)
         );
  OAI211_X1 U6445 ( .C1(n5689), .C2(n5702), .A(n5688), .B(n5687), .ZN(U3065)
         );
  AOI22_X1 U6446 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5697), .B1(n6956), 
        .B2(n5696), .ZN(n5691) );
  AOI22_X1 U6447 ( .A1(n5699), .A2(n7622), .B1(n5698), .B2(n7623), .ZN(n5690)
         );
  OAI211_X1 U6448 ( .C1(n5692), .C2(n5702), .A(n5691), .B(n5690), .ZN(U3064)
         );
  AOI22_X1 U6449 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n5697), .B1(n6973), 
        .B2(n5696), .ZN(n5694) );
  AOI22_X1 U6450 ( .A1(n5699), .A2(n7654), .B1(n5698), .B2(n7651), .ZN(n5693)
         );
  OAI211_X1 U6451 ( .C1(n5695), .C2(n5702), .A(n5694), .B(n5693), .ZN(U3067)
         );
  AOI22_X1 U6452 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n5697), .B1(n6936), 
        .B2(n5696), .ZN(n5701) );
  AOI22_X1 U6453 ( .A1(n5699), .A2(n7591), .B1(n5698), .B2(n7583), .ZN(n5700)
         );
  OAI211_X1 U6454 ( .C1(n5703), .C2(n5702), .A(n5701), .B(n5700), .ZN(U3060)
         );
  CLKBUF_X1 U6455 ( .A(n5704), .Z(n5705) );
  XNOR2_X1 U6456 ( .A(n5705), .B(n5706), .ZN(n5966) );
  NOR3_X1 U6457 ( .A1(n3848), .A2(n7508), .A3(n7514), .ZN(n7509) );
  INV_X1 U6458 ( .A(n7509), .ZN(n5711) );
  INV_X1 U6459 ( .A(n5709), .ZN(n5710) );
  OR2_X1 U6460 ( .A1(n4220), .A2(n5710), .ZN(n7504) );
  NAND3_X1 U6461 ( .A1(n7211), .A2(n5711), .A3(n7504), .ZN(n5712) );
  NOR2_X1 U6462 ( .A1(n5719), .A2(n7455), .ZN(n5713) );
  NAND3_X1 U6463 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_11__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U6464 ( .A1(n7520), .A2(n7502), .ZN(n5725) );
  INV_X1 U6465 ( .A(n5725), .ZN(n5714) );
  AND3_X1 U6466 ( .A1(n5715), .A2(n4743), .A3(n5714), .ZN(n5716) );
  NAND2_X1 U6467 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n6613) );
  NOR2_X1 U6468 ( .A1(n6613), .A2(n5074), .ZN(n7286) );
  NAND2_X1 U6469 ( .A1(n7286), .A2(REIP_REG_4__SCAN_IN), .ZN(n7303) );
  INV_X1 U6470 ( .A(REIP_REG_5__SCAN_IN), .ZN(n7302) );
  NOR2_X1 U6471 ( .A1(n7303), .A2(n7302), .ZN(n7310) );
  NAND2_X1 U6472 ( .A1(n7310), .A2(REIP_REG_6__SCAN_IN), .ZN(n7323) );
  OR2_X1 U6473 ( .A1(n7323), .A2(n5363), .ZN(n5839) );
  INV_X1 U6474 ( .A(REIP_REG_8__SCAN_IN), .ZN(n7033) );
  NOR2_X1 U6475 ( .A1(n5839), .A2(n7033), .ZN(n5717) );
  NAND2_X1 U6476 ( .A1(n7372), .A2(n5717), .ZN(n7348) );
  NOR2_X1 U6477 ( .A1(n5867), .A2(n7348), .ZN(n5718) );
  INV_X1 U6478 ( .A(REIP_REG_12__SCAN_IN), .ZN(n7366) );
  NAND2_X1 U6479 ( .A1(n5718), .A2(n7366), .ZN(n7361) );
  INV_X1 U6480 ( .A(n5717), .ZN(n5868) );
  NAND2_X1 U6481 ( .A1(n7372), .A2(n5868), .ZN(n5840) );
  NAND2_X1 U6482 ( .A1(n5840), .A2(n7301), .ZN(n7337) );
  AOI21_X1 U6483 ( .B1(n7372), .B2(n5867), .A(n7337), .ZN(n7367) );
  NAND3_X1 U6484 ( .A1(n7361), .A2(n7367), .A3(REIP_REG_13__SCAN_IN), .ZN(
        n7374) );
  OAI221_X1 U6485 ( .B1(REIP_REG_13__SCAN_IN), .B2(REIP_REG_12__SCAN_IN), .C1(
        REIP_REG_13__SCAN_IN), .C2(n5718), .A(n7374), .ZN(n5734) );
  AND2_X1 U6486 ( .A1(n5719), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5720) );
  AND2_X2 U6487 ( .A1(n7301), .A2(n5720), .ZN(n7425) );
  INV_X1 U6488 ( .A(n5962), .ZN(n5732) );
  NAND2_X1 U6489 ( .A1(EBX_REG_31__SCAN_IN), .A2(n5725), .ZN(n5721) );
  NOR2_X1 U6490 ( .A1(n6022), .A2(n5721), .ZN(n5722) );
  NOR2_X1 U6491 ( .A1(n5767), .A2(n5723), .ZN(n5724) );
  OR2_X1 U6492 ( .A1(n5758), .A2(n5724), .ZN(n5770) );
  INV_X1 U6493 ( .A(n5770), .ZN(n7196) );
  OR2_X1 U6494 ( .A1(n7183), .A2(n5725), .ZN(n7495) );
  NAND2_X1 U6495 ( .A1(n3915), .A2(n7495), .ZN(n6070) );
  INV_X1 U6496 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6071) );
  NAND3_X1 U6497 ( .A1(n4743), .A2(n5725), .A3(n6071), .ZN(n5726) );
  AND2_X1 U6498 ( .A1(n6070), .A2(n5726), .ZN(n5727) );
  NOR2_X2 U6499 ( .A1(n6072), .A2(n5727), .ZN(n7419) );
  AOI22_X1 U6500 ( .A1(n7441), .A2(n7196), .B1(n7419), .B2(EBX_REG_13__SCAN_IN), .ZN(n5728) );
  OAI21_X1 U6501 ( .B1(n5729), .B2(n7429), .A(n5728), .ZN(n5731) );
  INV_X1 U6502 ( .A(n7178), .ZN(n5730) );
  AOI211_X1 U6503 ( .C1(n7425), .C2(n5732), .A(n5731), .B(n7411), .ZN(n5733)
         );
  OAI211_X1 U6504 ( .C1(n5966), .C2(n7422), .A(n5734), .B(n5733), .ZN(U2814)
         );
  INV_X1 U6505 ( .A(n5735), .ZN(n6096) );
  OAI21_X1 U6506 ( .B1(n6072), .B2(n6096), .A(n7422), .ZN(n7305) );
  INV_X1 U6507 ( .A(n7305), .ZN(n7290) );
  INV_X1 U6508 ( .A(REIP_REG_2__SCAN_IN), .ZN(n7026) );
  INV_X1 U6509 ( .A(n7134), .ZN(n5736) );
  NAND2_X1 U6510 ( .A1(n7425), .A2(n5736), .ZN(n5737) );
  OAI21_X1 U6511 ( .B1(n7026), .B2(n7301), .A(n5737), .ZN(n5743) );
  INV_X1 U6512 ( .A(n5738), .ZN(n6103) );
  NAND2_X1 U6513 ( .A1(n5739), .A2(n6103), .ZN(n6618) );
  XNOR2_X1 U6514 ( .A(REIP_REG_2__SCAN_IN), .B(REIP_REG_1__SCAN_IN), .ZN(n5740) );
  OAI22_X1 U6515 ( .A1(n5741), .A2(n6618), .B1(n7324), .B2(n5740), .ZN(n5742)
         );
  AOI211_X1 U6516 ( .C1(n7439), .C2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n5743), 
        .B(n5742), .ZN(n5745) );
  AOI22_X1 U6517 ( .A1(n7441), .A2(n7227), .B1(n7419), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n5744) );
  OAI211_X1 U6518 ( .C1(n7290), .C2(n7127), .A(n5745), .B(n5744), .ZN(U2825)
         );
  INV_X1 U6519 ( .A(n6617), .ZN(n5749) );
  AOI21_X1 U6520 ( .B1(n7158), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5746), 
        .ZN(n5747) );
  OAI21_X1 U6521 ( .B1(n7169), .B2(n6606), .A(n5747), .ZN(n5748) );
  AOI21_X1 U6522 ( .B1(n5749), .B2(n7165), .A(n5748), .ZN(n5750) );
  OAI21_X1 U6523 ( .B1(n5751), .B2(n7447), .A(n5750), .ZN(U2983) );
  OR2_X1 U6524 ( .A1(n5753), .A2(n5752), .ZN(n5756) );
  NAND2_X1 U6525 ( .A1(n5756), .A2(n5755), .ZN(n7375) );
  OR2_X1 U6526 ( .A1(n5758), .A2(n5757), .ZN(n5759) );
  AND2_X1 U6527 ( .A1(n5817), .A2(n5759), .ZN(n7368) );
  AOI22_X1 U6528 ( .A1(n7124), .A2(n7368), .B1(EBX_REG_14__SCAN_IN), .B2(n6636), .ZN(n5760) );
  OAI21_X1 U6529 ( .B1(n7375), .B2(n6648), .A(n5760), .ZN(U2845) );
  NAND2_X1 U6530 ( .A1(n5799), .A2(n5798), .ZN(n5763) );
  INV_X1 U6531 ( .A(n5761), .ZN(n5762) );
  AOI21_X1 U6532 ( .B1(n5764), .B2(n5763), .A(n5762), .ZN(n5898) );
  INV_X1 U6533 ( .A(n5898), .ZN(n7362) );
  AND2_X1 U6534 ( .A1(n5859), .A2(n5765), .ZN(n5766) );
  NOR2_X1 U6535 ( .A1(n5767), .A2(n5766), .ZN(n7355) );
  AOI22_X1 U6536 ( .A1(n7124), .A2(n7355), .B1(EBX_REG_12__SCAN_IN), .B2(n6636), .ZN(n5768) );
  OAI21_X1 U6537 ( .B1(n7362), .B2(n6648), .A(n5768), .ZN(U2847) );
  INV_X1 U6538 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5769) );
  OAI222_X1 U6539 ( .A1(n5770), .A2(n6647), .B1(n5769), .B2(n7126), .C1(n6648), 
        .C2(n5966), .ZN(U2846) );
  AOI21_X1 U6540 ( .B1(n7158), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5771), 
        .ZN(n5772) );
  OAI21_X1 U6541 ( .B1(n7169), .B2(n7326), .A(n5772), .ZN(n5773) );
  AOI21_X1 U6542 ( .B1(n7328), .B2(n7165), .A(n5773), .ZN(n5774) );
  OAI21_X1 U6543 ( .B1(n5775), .B2(n7447), .A(n5774), .ZN(U2979) );
  INV_X1 U6544 ( .A(DATAI_13_), .ZN(n5776) );
  INV_X1 U6545 ( .A(EAX_REG_13__SCAN_IN), .ZN(n7020) );
  OAI222_X1 U6546 ( .A1(n5848), .A2(n5776), .B1(n6669), .B2(n5966), .C1(n7020), 
        .C2(n6085), .ZN(U2878) );
  INV_X1 U6547 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U6548 ( .A1(n7158), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5779)
         );
  INV_X1 U6549 ( .A(n5777), .ZN(n5778) );
  OAI211_X1 U6550 ( .C1(n5780), .C2(n6797), .A(n5779), .B(n5778), .ZN(n5781)
         );
  AOI21_X1 U6551 ( .B1(n7154), .B2(n6619), .A(n5781), .ZN(n5782) );
  OAI21_X1 U6552 ( .B1(n5783), .B2(n7447), .A(n5782), .ZN(U2985) );
  NAND2_X1 U6553 ( .A1(n7158), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5784)
         );
  OAI211_X1 U6554 ( .C1(n7169), .C2(n5841), .A(n5785), .B(n5784), .ZN(n5786)
         );
  AOI21_X1 U6555 ( .B1(n5787), .B2(n7165), .A(n5786), .ZN(n5788) );
  OAI21_X1 U6556 ( .B1(n5789), .B2(n7447), .A(n5788), .ZN(U2978) );
  INV_X1 U6557 ( .A(DATAI_14_), .ZN(n5790) );
  INV_X1 U6558 ( .A(EAX_REG_14__SCAN_IN), .ZN(n7022) );
  OAI222_X1 U6559 ( .A1(n5848), .A2(n5790), .B1(n6085), .B2(n7022), .C1(n6669), 
        .C2(n7375), .ZN(U2877) );
  CLKBUF_X1 U6560 ( .A(n5791), .Z(n5792) );
  XOR2_X1 U6561 ( .A(n5792), .B(n5793), .Z(n7255) );
  NAND2_X1 U6562 ( .A1(n7255), .A2(n7166), .ZN(n5797) );
  INV_X1 U6563 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U6564 ( .A1(n7276), .A2(REIP_REG_9__SCAN_IN), .ZN(n7252) );
  OAI21_X1 U6565 ( .B1(n6791), .B2(n5794), .A(n7252), .ZN(n5795) );
  AOI21_X1 U6566 ( .B1(n7154), .B2(n7339), .A(n5795), .ZN(n5796) );
  OAI211_X1 U6567 ( .C1(n6797), .C2(n7338), .A(n5797), .B(n5796), .ZN(U2977)
         );
  INV_X1 U6568 ( .A(DATAI_11_), .ZN(n5804) );
  INV_X1 U6569 ( .A(EAX_REG_11__SCAN_IN), .ZN(n7016) );
  INV_X1 U6570 ( .A(n5798), .ZN(n5802) );
  AND2_X1 U6571 ( .A1(n5799), .A2(n5798), .ZN(n5800) );
  AOI21_X1 U6572 ( .B1(n5802), .B2(n5801), .A(n5800), .ZN(n7351) );
  INV_X1 U6573 ( .A(n7351), .ZN(n5803) );
  OAI222_X1 U6574 ( .A1(n5848), .A2(n5804), .B1(n6085), .B2(n7016), .C1(n6669), 
        .C2(n5803), .ZN(U2880) );
  INV_X1 U6575 ( .A(DATAI_12_), .ZN(n5805) );
  INV_X1 U6576 ( .A(EAX_REG_12__SCAN_IN), .ZN(n7018) );
  OAI222_X1 U6577 ( .A1(n5848), .A2(n5805), .B1(n6085), .B2(n7018), .C1(n6669), 
        .C2(n7362), .ZN(U2879) );
  AND2_X1 U6578 ( .A1(n7324), .A2(n7301), .ZN(n6075) );
  INV_X1 U6579 ( .A(n6075), .ZN(n6598) );
  OAI22_X1 U6580 ( .A1(n7435), .A2(n4938), .B1(n5806), .B2(n7421), .ZN(n5807)
         );
  AOI21_X1 U6581 ( .B1(REIP_REG_0__SCAN_IN), .B2(n6598), .A(n5807), .ZN(n5810)
         );
  INV_X1 U6582 ( .A(n6618), .ZN(n7283) );
  NAND2_X1 U6583 ( .A1(n7429), .A2(n7445), .ZN(n5808) );
  AOI22_X1 U6584 ( .A1(n7283), .A2(n7454), .B1(n5808), .B2(
        PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n5809) );
  OAI211_X1 U6585 ( .C1(n7290), .C2(n5811), .A(n5810), .B(n5809), .ZN(U2827)
         );
  NAND2_X1 U6586 ( .A1(n5755), .A2(n5814), .ZN(n5815) );
  NAND2_X1 U6587 ( .A1(n5813), .A2(n5815), .ZN(n6011) );
  INV_X1 U6588 ( .A(n5881), .ZN(n5816) );
  AOI21_X1 U6589 ( .B1(n5818), .B2(n5817), .A(n5816), .ZN(n7264) );
  AOI22_X1 U6590 ( .A1(n7264), .A2(n7124), .B1(EBX_REG_15__SCAN_IN), .B2(n6636), .ZN(n5819) );
  OAI21_X1 U6591 ( .B1(n6011), .B2(n6648), .A(n5819), .ZN(U2844) );
  INV_X1 U6592 ( .A(REIP_REG_9__SCAN_IN), .ZN(n7035) );
  NOR3_X1 U6593 ( .A1(REIP_REG_10__SCAN_IN), .A2(n7035), .A3(n7348), .ZN(n5825) );
  AOI22_X1 U6594 ( .A1(n7441), .A2(n7243), .B1(n7419), .B2(EBX_REG_10__SCAN_IN), .ZN(n5820) );
  INV_X1 U6595 ( .A(n7411), .ZN(n7315) );
  OAI211_X1 U6596 ( .C1(n7429), .C2(n5821), .A(n5820), .B(n7315), .ZN(n5824)
         );
  NOR2_X1 U6597 ( .A1(n7348), .A2(REIP_REG_9__SCAN_IN), .ZN(n7335) );
  OAI21_X1 U6598 ( .B1(n7335), .B2(n7337), .A(REIP_REG_10__SCAN_IN), .ZN(n5822) );
  OAI21_X1 U6599 ( .B1(n7445), .B2(n5832), .A(n5822), .ZN(n5823) );
  NOR3_X1 U6600 ( .A1(n5825), .A2(n5824), .A3(n5823), .ZN(n5826) );
  OAI21_X1 U6601 ( .B1(n5836), .B2(n7422), .A(n5826), .ZN(U2817) );
  CLKBUF_X1 U6602 ( .A(n5827), .Z(n5828) );
  NAND2_X1 U6603 ( .A1(n5850), .A2(n5829), .ZN(n5830) );
  XNOR2_X1 U6604 ( .A(n5828), .B(n5830), .ZN(n7247) );
  NAND2_X1 U6605 ( .A1(n7247), .A2(n7166), .ZN(n5835) );
  INV_X1 U6606 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5831) );
  NOR2_X1 U6607 ( .A1(n7211), .A2(n5831), .ZN(n7242) );
  NOR2_X1 U6608 ( .A1(n7169), .A2(n5832), .ZN(n5833) );
  AOI211_X1 U6609 ( .C1(n7158), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n7242), 
        .B(n5833), .ZN(n5834) );
  OAI211_X1 U6610 ( .C1(n6797), .C2(n5836), .A(n5835), .B(n5834), .ZN(U2976)
         );
  AOI22_X1 U6611 ( .A1(EBX_REG_8__SCAN_IN), .A2(n7419), .B1(
        REIP_REG_8__SCAN_IN), .B2(n7337), .ZN(n5837) );
  OAI211_X1 U6612 ( .C1(n7429), .C2(n5838), .A(n5837), .B(n7315), .ZN(n5845)
         );
  NOR2_X1 U6613 ( .A1(n5840), .A2(n5839), .ZN(n5844) );
  OAI22_X1 U6614 ( .A1(n7421), .A2(n5842), .B1(n7445), .B2(n5841), .ZN(n5843)
         );
  NOR3_X1 U6615 ( .A1(n5845), .A2(n5844), .A3(n5843), .ZN(n5846) );
  OAI21_X1 U6616 ( .B1(n7422), .B2(n5847), .A(n5846), .ZN(U2819) );
  OAI222_X1 U6617 ( .A1(n5849), .A2(n5848), .B1(n6085), .B2(n4924), .C1(n6669), 
        .C2(n6011), .ZN(U2876) );
  NAND2_X1 U6618 ( .A1(n3647), .A2(n5850), .ZN(n5855) );
  INV_X1 U6619 ( .A(n5884), .ZN(n5853) );
  NOR2_X1 U6620 ( .A1(n5853), .A2(n5852), .ZN(n5854) );
  NAND2_X1 U6621 ( .A1(n5855), .A2(n5854), .ZN(n5885) );
  OAI21_X1 U6622 ( .B1(n5855), .B2(n5854), .A(n5885), .ZN(n7157) );
  OAI21_X1 U6623 ( .B1(n5857), .B2(n7233), .A(n5856), .ZN(n7259) );
  INV_X1 U6624 ( .A(n7197), .ZN(n5858) );
  AOI22_X1 U6625 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n7259), .B1(n5858), .B2(n7198), .ZN(n5864) );
  INV_X1 U6626 ( .A(n5859), .ZN(n5860) );
  AOI21_X1 U6627 ( .B1(n5862), .B2(n5861), .A(n5860), .ZN(n7345) );
  AOI22_X1 U6628 ( .A1(n7269), .A2(n7345), .B1(n7276), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n5863) );
  OAI211_X1 U6629 ( .C1(n7157), .C2(n6892), .A(n5864), .B(n5863), .ZN(U3007)
         );
  INV_X1 U6630 ( .A(n7264), .ZN(n5866) );
  OAI22_X1 U6631 ( .A1(n5866), .A2(n7421), .B1(n7445), .B2(n5865), .ZN(n5873)
         );
  NOR2_X1 U6632 ( .A1(n5868), .A2(n5867), .ZN(n5869) );
  NAND4_X1 U6633 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .A3(
        REIP_REG_14__SCAN_IN), .A4(n5869), .ZN(n7371) );
  INV_X1 U6634 ( .A(n7371), .ZN(n5870) );
  NAND2_X1 U6635 ( .A1(n7372), .A2(n5870), .ZN(n7393) );
  INV_X1 U6636 ( .A(REIP_REG_15__SCAN_IN), .ZN(n7044) );
  INV_X1 U6637 ( .A(n7301), .ZN(n6626) );
  OAI21_X1 U6638 ( .B1(n6626), .B2(n7371), .A(n6598), .ZN(n7382) );
  AOI21_X1 U6639 ( .B1(n7439), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n7411), 
        .ZN(n5871) );
  OAI221_X1 U6640 ( .B1(REIP_REG_15__SCAN_IN), .B2(n7393), .C1(n7044), .C2(
        n7382), .A(n5871), .ZN(n5872) );
  AOI211_X1 U6641 ( .C1(EBX_REG_15__SCAN_IN), .C2(n7419), .A(n5873), .B(n5872), 
        .ZN(n5874) );
  OAI21_X1 U6642 ( .B1(n6011), .B2(n7422), .A(n5874), .ZN(U2812) );
  INV_X1 U6643 ( .A(n5813), .ZN(n5879) );
  INV_X1 U6644 ( .A(n5876), .ZN(n5877) );
  OAI21_X1 U6645 ( .B1(n5879), .B2(n5878), .A(n5877), .ZN(n7386) );
  INV_X1 U6646 ( .A(n7112), .ZN(n5880) );
  AOI21_X1 U6647 ( .B1(n5882), .B2(n5881), .A(n5880), .ZN(n7384) );
  AOI22_X1 U6648 ( .A1(n7384), .A2(n7124), .B1(EBX_REG_16__SCAN_IN), .B2(n6636), .ZN(n5883) );
  OAI21_X1 U6649 ( .B1(n7386), .B2(n6648), .A(n5883), .ZN(U2843) );
  NAND2_X1 U6650 ( .A1(n5885), .A2(n5884), .ZN(n5887) );
  XNOR2_X1 U6651 ( .A(n6751), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5886)
         );
  XNOR2_X1 U6652 ( .A(n5887), .B(n5886), .ZN(n5900) );
  NOR2_X1 U6653 ( .A1(n7211), .A2(n7366), .ZN(n5894) );
  NOR2_X1 U6654 ( .A1(n7198), .A2(n7197), .ZN(n5891) );
  AOI21_X1 U6655 ( .B1(n7198), .B2(n5888), .A(n7259), .ZN(n5889) );
  INV_X1 U6656 ( .A(n5889), .ZN(n5890) );
  MUX2_X1 U6657 ( .A(n5891), .B(n5890), .S(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .Z(n5892) );
  AOI211_X1 U6658 ( .C1(n7269), .C2(n7355), .A(n5894), .B(n5892), .ZN(n5893)
         );
  OAI21_X1 U6659 ( .B1(n5900), .B2(n6892), .A(n5893), .ZN(U3006) );
  AOI21_X1 U6660 ( .B1(n7158), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5894), 
        .ZN(n5895) );
  OAI21_X1 U6661 ( .B1(n7169), .B2(n5896), .A(n5895), .ZN(n5897) );
  AOI21_X1 U6662 ( .B1(n5898), .B2(n7165), .A(n5897), .ZN(n5899) );
  OAI21_X1 U6663 ( .B1(n5900), .B2(n7447), .A(n5899), .ZN(U2974) );
  AOI22_X1 U6664 ( .A1(n7550), .A2(DATAI_16_), .B1(n7553), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5904) );
  AND2_X1 U6665 ( .A1(n5901), .A2(n4193), .ZN(n5902) );
  NAND2_X1 U6666 ( .A1(n7554), .A2(DATAI_0_), .ZN(n5903) );
  OAI211_X1 U6667 ( .C1(n7386), .C2(n6669), .A(n5904), .B(n5903), .ZN(U2875)
         );
  OAI21_X1 U6668 ( .B1(n5911), .B2(n5950), .A(n7579), .ZN(n5905) );
  OAI21_X1 U6669 ( .B1(n5097), .B2(n5913), .A(n5905), .ZN(n5907) );
  NOR2_X1 U6670 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5906), .ZN(n5955)
         );
  AOI21_X1 U6671 ( .B1(n5907), .B2(n7508), .A(n5955), .ZN(n5910) );
  INV_X1 U6672 ( .A(n5908), .ZN(n5909) );
  NOR3_X2 U6673 ( .A1(n5910), .A2(n7565), .A3(n5909), .ZN(n5958) );
  INV_X1 U6674 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5918) );
  OAI22_X1 U6675 ( .A1(n6935), .A2(n5913), .B1(n5912), .B2(n6931), .ZN(n5949)
         );
  AOI22_X1 U6676 ( .A1(n5950), .A2(n7630), .B1(n6961), .B2(n5949), .ZN(n5914)
         );
  OAI21_X1 U6677 ( .B1(n5953), .B2(n5915), .A(n5914), .ZN(n5916) );
  AOI21_X1 U6678 ( .B1(n7629), .B2(n5955), .A(n5916), .ZN(n5917) );
  OAI21_X1 U6679 ( .B1(n5958), .B2(n5918), .A(n5917), .ZN(U3041) );
  INV_X1 U6680 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5923) );
  AOI22_X1 U6681 ( .A1(n5950), .A2(n7638), .B1(n6966), .B2(n5949), .ZN(n5919)
         );
  OAI21_X1 U6682 ( .B1(n5953), .B2(n5920), .A(n5919), .ZN(n5921) );
  AOI21_X1 U6683 ( .B1(n7637), .B2(n5955), .A(n5921), .ZN(n5922) );
  OAI21_X1 U6684 ( .B1(n5958), .B2(n5923), .A(n5922), .ZN(U3042) );
  INV_X1 U6685 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5928) );
  AOI22_X1 U6686 ( .A1(n5950), .A2(n7622), .B1(n6956), .B2(n5949), .ZN(n5924)
         );
  OAI21_X1 U6687 ( .B1(n5953), .B2(n5925), .A(n5924), .ZN(n5926) );
  AOI21_X1 U6688 ( .B1(n7621), .B2(n5955), .A(n5926), .ZN(n5927) );
  OAI21_X1 U6689 ( .B1(n5958), .B2(n5928), .A(n5927), .ZN(U3040) );
  INV_X1 U6690 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5933) );
  AOI22_X1 U6691 ( .A1(n5950), .A2(n7615), .B1(n6951), .B2(n5949), .ZN(n5929)
         );
  OAI21_X1 U6692 ( .B1(n5953), .B2(n5930), .A(n5929), .ZN(n5931) );
  AOI21_X1 U6693 ( .B1(n7613), .B2(n5955), .A(n5931), .ZN(n5932) );
  OAI21_X1 U6694 ( .B1(n5958), .B2(n5933), .A(n5932), .ZN(U3039) );
  INV_X1 U6695 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5938) );
  AOI22_X1 U6696 ( .A1(n5950), .A2(n7606), .B1(n6946), .B2(n5949), .ZN(n5934)
         );
  OAI21_X1 U6697 ( .B1(n5953), .B2(n5935), .A(n5934), .ZN(n5936) );
  AOI21_X1 U6698 ( .B1(n7605), .B2(n5955), .A(n5936), .ZN(n5937) );
  OAI21_X1 U6699 ( .B1(n5958), .B2(n5938), .A(n5937), .ZN(U3038) );
  INV_X1 U6700 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5943) );
  AOI22_X1 U6701 ( .A1(n5950), .A2(n7654), .B1(n6973), .B2(n5949), .ZN(n5939)
         );
  OAI21_X1 U6702 ( .B1(n5953), .B2(n5940), .A(n5939), .ZN(n5941) );
  AOI21_X1 U6703 ( .B1(n7650), .B2(n5955), .A(n5941), .ZN(n5942) );
  OAI21_X1 U6704 ( .B1(n5958), .B2(n5943), .A(n5942), .ZN(U3043) );
  INV_X1 U6705 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5948) );
  AOI22_X1 U6706 ( .A1(n5950), .A2(n7591), .B1(n6936), .B2(n5949), .ZN(n5944)
         );
  OAI21_X1 U6707 ( .B1(n5953), .B2(n5945), .A(n5944), .ZN(n5946) );
  AOI21_X1 U6708 ( .B1(n7582), .B2(n5955), .A(n5946), .ZN(n5947) );
  OAI21_X1 U6709 ( .B1(n5958), .B2(n5948), .A(n5947), .ZN(U3036) );
  INV_X1 U6710 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5957) );
  AOI22_X1 U6711 ( .A1(n5950), .A2(n7599), .B1(n6941), .B2(n5949), .ZN(n5951)
         );
  OAI21_X1 U6712 ( .B1(n5953), .B2(n5952), .A(n5951), .ZN(n5954) );
  AOI21_X1 U6713 ( .B1(n7597), .B2(n5955), .A(n5954), .ZN(n5956) );
  OAI21_X1 U6714 ( .B1(n5958), .B2(n5957), .A(n5956), .ZN(U3037) );
  XNOR2_X1 U6715 ( .A(n5960), .B(n5961), .ZN(n7200) );
  NAND2_X1 U6716 ( .A1(n7200), .A2(n7166), .ZN(n5965) );
  AND2_X1 U6717 ( .A1(n7276), .A2(REIP_REG_13__SCAN_IN), .ZN(n7195) );
  NOR2_X1 U6718 ( .A1(n7169), .A2(n5962), .ZN(n5963) );
  AOI211_X1 U6719 ( .C1(n7158), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n7195), 
        .B(n5963), .ZN(n5964) );
  OAI211_X1 U6720 ( .C1(n5966), .C2(n6797), .A(n5965), .B(n5964), .ZN(U2973)
         );
  CLKBUF_X1 U6721 ( .A(n5967), .Z(n5968) );
  XOR2_X1 U6722 ( .A(n5968), .B(n5969), .Z(n5982) );
  INV_X1 U6723 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5970) );
  NOR2_X1 U6724 ( .A1(n7211), .A2(n5970), .ZN(n5978) );
  NOR2_X1 U6725 ( .A1(n5971), .A2(n7197), .ZN(n5973) );
  AOI21_X1 U6726 ( .B1(n5971), .B2(n7260), .A(n7259), .ZN(n7203) );
  INV_X1 U6727 ( .A(n7203), .ZN(n5972) );
  MUX2_X1 U6728 ( .A(n5973), .B(n5972), .S(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .Z(n5974) );
  AOI211_X1 U6729 ( .C1(n7269), .C2(n7368), .A(n5978), .B(n5974), .ZN(n5975)
         );
  OAI21_X1 U6730 ( .B1(n5982), .B2(n6892), .A(n5975), .ZN(U3004) );
  NOR2_X1 U6731 ( .A1(n6791), .A2(n5976), .ZN(n5977) );
  AOI211_X1 U6732 ( .C1(n7154), .C2(n7377), .A(n5978), .B(n5977), .ZN(n5981)
         );
  INV_X1 U6733 ( .A(n7375), .ZN(n5979) );
  NAND2_X1 U6734 ( .A1(n5979), .A2(n7165), .ZN(n5980) );
  OAI211_X1 U6735 ( .C1(n5982), .C2(n7447), .A(n5981), .B(n5980), .ZN(U2972)
         );
  INV_X1 U6736 ( .A(n5984), .ZN(n5989) );
  INV_X1 U6737 ( .A(n5985), .ZN(n5988) );
  OAI21_X1 U6738 ( .B1(n5989), .B2(n5988), .A(n6775), .ZN(n6796) );
  NAND2_X1 U6739 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n7394) );
  INV_X1 U6740 ( .A(REIP_REG_17__SCAN_IN), .ZN(n7392) );
  NOR3_X1 U6741 ( .A1(n7371), .A2(n7394), .A3(n7392), .ZN(n6073) );
  OAI21_X1 U6742 ( .B1(n7324), .B2(n6073), .A(n7301), .ZN(n7402) );
  NAND2_X1 U6743 ( .A1(n7402), .A2(REIP_REG_18__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U6744 ( .A1(n7372), .A2(n6073), .ZN(n7404) );
  NOR2_X1 U6745 ( .A1(REIP_REG_18__SCAN_IN), .A2(n7404), .ZN(n7403) );
  NOR2_X1 U6746 ( .A1(n7411), .A2(n7403), .ZN(n5994) );
  AOI22_X1 U6747 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n7439), .B1(n7425), 
        .B2(n6793), .ZN(n5993) );
  OR2_X1 U6748 ( .A1(n7114), .A2(n5990), .ZN(n5991) );
  AND2_X1 U6749 ( .A1(n5991), .A2(n6898), .ZN(n6909) );
  AOI22_X1 U6750 ( .A1(n6909), .A2(n7441), .B1(n7419), .B2(EBX_REG_18__SCAN_IN), .ZN(n5992) );
  AND4_X1 U6751 ( .A1(n5995), .A2(n5994), .A3(n5993), .A4(n5992), .ZN(n5996)
         );
  OAI21_X1 U6752 ( .B1(n6796), .B2(n7422), .A(n5996), .ZN(U2809) );
  AOI22_X1 U6753 ( .A1(n6909), .A2(n7124), .B1(EBX_REG_18__SCAN_IN), .B2(n6636), .ZN(n5997) );
  OAI21_X1 U6754 ( .B1(n6796), .B2(n6648), .A(n5997), .ZN(U2841) );
  AOI22_X1 U6755 ( .A1(n7550), .A2(DATAI_18_), .B1(n7553), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U6756 ( .A1(n7554), .A2(DATAI_2_), .ZN(n5998) );
  OAI211_X1 U6757 ( .C1(n6796), .C2(n6669), .A(n5999), .B(n5998), .ZN(U2873)
         );
  INV_X1 U6758 ( .A(n6002), .ZN(n6004) );
  NOR2_X1 U6759 ( .A1(n6004), .A2(n6003), .ZN(n6005) );
  XNOR2_X1 U6760 ( .A(n6001), .B(n6005), .ZN(n7265) );
  NAND2_X1 U6761 ( .A1(n7265), .A2(n7166), .ZN(n6010) );
  INV_X1 U6762 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U6763 ( .A1(n7276), .A2(REIP_REG_15__SCAN_IN), .ZN(n7262) );
  OAI21_X1 U6764 ( .B1(n6791), .B2(n6006), .A(n7262), .ZN(n6007) );
  AOI21_X1 U6765 ( .B1(n7154), .B2(n6008), .A(n6007), .ZN(n6009) );
  OAI211_X1 U6766 ( .C1(n6797), .C2(n6011), .A(n6010), .B(n6009), .ZN(U2971)
         );
  NAND2_X1 U6767 ( .A1(n6015), .A2(n6014), .ZN(n6016) );
  XNOR2_X1 U6768 ( .A(n6013), .B(n6016), .ZN(n7270) );
  NAND2_X1 U6769 ( .A1(n7270), .A2(n7166), .ZN(n6021) );
  INV_X1 U6770 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6017) );
  OAI22_X1 U6771 ( .A1(n6791), .A2(n6018), .B1(n7211), .B2(n6017), .ZN(n6019)
         );
  AOI21_X1 U6772 ( .B1(n7154), .B2(n7388), .A(n6019), .ZN(n6020) );
  OAI211_X1 U6773 ( .C1(n6797), .C2(n7386), .A(n6021), .B(n6020), .ZN(U2970)
         );
  AOI22_X1 U6774 ( .A1(n6023), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6022), .ZN(n6032) );
  NAND2_X1 U6775 ( .A1(n6024), .A2(n3633), .ZN(n6025) );
  NAND2_X1 U6776 ( .A1(n3655), .A2(EBX_REG_29__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U6777 ( .A1(n6025), .A2(n6029), .ZN(n6116) );
  INV_X1 U6778 ( .A(n6026), .ZN(n6118) );
  NAND2_X1 U6779 ( .A1(n6498), .A2(n3655), .ZN(n6028) );
  XOR2_X1 U6780 ( .A(n6032), .B(n6031), .Z(n6084) );
  OAI22_X1 U6781 ( .A1(n6084), .A2(n6647), .B1(n7126), .B2(n6071), .ZN(U2828)
         );
  INV_X1 U6782 ( .A(n6033), .ZN(n6105) );
  AOI21_X1 U6783 ( .B1(n7158), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n6034), 
        .ZN(n6035) );
  OAI21_X1 U6784 ( .B1(n7169), .B2(n6105), .A(n6035), .ZN(n6036) );
  AOI21_X1 U6785 ( .B1(n6649), .B2(n7165), .A(n6036), .ZN(n6037) );
  OAI21_X1 U6786 ( .B1(n6038), .B2(n7447), .A(n6037), .ZN(U2956) );
  AND2_X1 U6787 ( .A1(n6040), .A2(n6039), .ZN(n7511) );
  INV_X1 U6788 ( .A(n7511), .ZN(n6042) );
  NAND2_X1 U6789 ( .A1(n6992), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6041) );
  OAI21_X1 U6790 ( .B1(n6992), .B2(n6042), .A(n6041), .ZN(n6043) );
  AOI21_X1 U6791 ( .B1(n6065), .B2(n7557), .A(n6043), .ZN(n6044) );
  OAI21_X1 U6792 ( .B1(n6045), .B2(n6069), .A(n6044), .ZN(U3465) );
  INV_X1 U6793 ( .A(n6046), .ZN(n6047) );
  OAI211_X1 U6794 ( .C1(n6084), .C2(n7212), .A(n6047), .B(n3668), .ZN(n6048)
         );
  INV_X1 U6795 ( .A(n6048), .ZN(n6052) );
  OAI211_X1 U6796 ( .C1(n6799), .C2(n6050), .A(INSTADDRPOINTER_REG_31__SCAN_IN), .B(n6049), .ZN(n6051) );
  OAI211_X1 U6797 ( .C1(n6053), .C2(n6892), .A(n6052), .B(n6051), .ZN(U2987)
         );
  AND2_X1 U6798 ( .A1(n6055), .A2(n6054), .ZN(n6057) );
  NOR3_X1 U6799 ( .A1(n6060), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n7513), 
        .ZN(n6056) );
  AOI211_X1 U6800 ( .C1(n6058), .C2(n7501), .A(n6057), .B(n6056), .ZN(n6063)
         );
  AOI21_X1 U6801 ( .B1(n6060), .B2(n6059), .A(n6920), .ZN(n6062) );
  OAI22_X1 U6802 ( .A1(n6063), .A2(n6920), .B1(n6062), .B2(n3646), .ZN(U3459)
         );
  OAI211_X1 U6803 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6066), .A(n6065), .B(
        n6064), .ZN(n6068) );
  NAND2_X1 U6804 ( .A1(n6992), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6067) );
  OAI211_X1 U6805 ( .C1(n6069), .C2(n3648), .A(n6068), .B(n6067), .ZN(U3464)
         );
  NAND2_X1 U6806 ( .A1(n6087), .A2(n7442), .ZN(n6083) );
  NOR3_X1 U6807 ( .A1(n6072), .A2(n6071), .A3(n6070), .ZN(n6081) );
  INV_X1 U6808 ( .A(REIP_REG_27__SCAN_IN), .ZN(n7061) );
  NAND3_X1 U6809 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .A3(
        REIP_REG_22__SCAN_IN), .ZN(n6579) );
  NAND3_X1 U6810 ( .A1(n6073), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n6578) );
  NOR2_X1 U6811 ( .A1(n6579), .A2(n6578), .ZN(n6074) );
  AND2_X1 U6812 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6074), .ZN(n6563) );
  NAND2_X1 U6813 ( .A1(n6563), .A2(REIP_REG_24__SCAN_IN), .ZN(n6546) );
  INV_X1 U6814 ( .A(REIP_REG_25__SCAN_IN), .ZN(n7058) );
  NOR2_X1 U6815 ( .A1(n6546), .A2(n7058), .ZN(n6533) );
  AND2_X1 U6816 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6533), .ZN(n6076) );
  INV_X1 U6817 ( .A(n6076), .ZN(n6514) );
  NOR3_X1 U6818 ( .A1(n7324), .A2(n7061), .A3(n6514), .ZN(n6504) );
  NAND3_X1 U6819 ( .A1(n6504), .A2(REIP_REG_29__SCAN_IN), .A3(
        REIP_REG_28__SCAN_IN), .ZN(n6108) );
  NOR2_X1 U6820 ( .A1(n6108), .A2(n7068), .ZN(n6079) );
  NAND2_X1 U6821 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_28__SCAN_IN), .ZN(
        n6077) );
  AOI21_X1 U6822 ( .B1(n6076), .B2(n7301), .A(n6075), .ZN(n6532) );
  AOI21_X1 U6823 ( .B1(n6598), .B2(n6077), .A(n6532), .ZN(n6505) );
  INV_X1 U6824 ( .A(REIP_REG_29__SCAN_IN), .ZN(n7066) );
  OAI21_X1 U6825 ( .B1(n7068), .B2(n7066), .A(n7372), .ZN(n6078) );
  NAND2_X1 U6826 ( .A1(n6505), .A2(n6078), .ZN(n6106) );
  MUX2_X1 U6827 ( .A(n6079), .B(n6106), .S(REIP_REG_31__SCAN_IN), .Z(n6080) );
  AOI211_X1 U6828 ( .C1(PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n7439), .A(n6081), 
        .B(n6080), .ZN(n6082) );
  OAI211_X1 U6829 ( .C1(n6084), .C2(n7421), .A(n6083), .B(n6082), .ZN(U2796)
         );
  NAND3_X1 U6830 ( .A1(n6087), .A2(n6086), .A3(n6085), .ZN(n6089) );
  AOI22_X1 U6831 ( .A1(n7550), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n7553), .ZN(n6088) );
  NAND2_X1 U6832 ( .A1(n6089), .A2(n6088), .ZN(U2860) );
  INV_X1 U6833 ( .A(n6098), .ZN(n6090) );
  NAND2_X1 U6834 ( .A1(n4729), .A2(n6090), .ZN(n6094) );
  INV_X1 U6835 ( .A(n6100), .ZN(n6092) );
  OAI21_X1 U6836 ( .B1(n6092), .B2(n6091), .A(n6097), .ZN(n6093) );
  OAI211_X1 U6837 ( .C1(n6097), .C2(n6095), .A(n6094), .B(n6093), .ZN(n7482)
         );
  NAND2_X1 U6838 ( .A1(n6097), .A2(n6096), .ZN(n6102) );
  NAND2_X1 U6839 ( .A1(n4729), .A2(n6098), .ZN(n6099) );
  NAND2_X1 U6840 ( .A1(n6100), .A2(n6099), .ZN(n6101) );
  NAND2_X1 U6841 ( .A1(n6102), .A2(n6101), .ZN(n7170) );
  OR2_X1 U6842 ( .A1(n3915), .A2(n6103), .ZN(n7175) );
  AOI21_X1 U6843 ( .B1(n7175), .B2(n7183), .A(READY_N), .ZN(n7186) );
  OR2_X1 U6844 ( .A1(n7170), .A2(n7186), .ZN(n7487) );
  AND2_X1 U6845 ( .A1(n7487), .A2(n7499), .ZN(n7449) );
  MUX2_X1 U6846 ( .A(MORE_REG_SCAN_IN), .B(n7482), .S(n7449), .Z(U3471) );
  NAND2_X1 U6847 ( .A1(n6649), .A2(n7442), .ZN(n6112) );
  OAI22_X1 U6848 ( .A1(n6105), .A2(n7445), .B1(n7429), .B2(n6104), .ZN(n6110)
         );
  INV_X1 U6849 ( .A(n6106), .ZN(n6107) );
  AOI21_X1 U6850 ( .B1(n7068), .B2(n6108), .A(n6107), .ZN(n6109) );
  AOI211_X1 U6851 ( .C1(EBX_REG_30__SCAN_IN), .C2(n7419), .A(n6110), .B(n6109), 
        .ZN(n6111) );
  OAI211_X1 U6852 ( .C1(n7421), .C2(n6113), .A(n6112), .B(n6111), .ZN(U2797)
         );
  AOI21_X1 U6853 ( .B1(n6115), .B2(n6500), .A(n6114), .ZN(n6629) );
  NAND2_X1 U6854 ( .A1(n6498), .A2(n6116), .ZN(n6117) );
  NAND2_X1 U6855 ( .A1(n6118), .A2(n6117), .ZN(n6798) );
  OAI22_X1 U6856 ( .A1(n6119), .A2(n7429), .B1(n7445), .B2(n6686), .ZN(n6120)
         );
  AOI21_X1 U6857 ( .B1(EBX_REG_29__SCAN_IN), .B2(n7419), .A(n6120), .ZN(n6123)
         );
  NAND2_X1 U6858 ( .A1(n6504), .A2(REIP_REG_28__SCAN_IN), .ZN(n6121) );
  MUX2_X1 U6859 ( .A(n6121), .B(n6505), .S(REIP_REG_29__SCAN_IN), .Z(n6122) );
  OAI211_X1 U6860 ( .C1(n6798), .C2(n7421), .A(n6123), .B(n6122), .ZN(n6124)
         );
  AOI21_X1 U6861 ( .B1(n6629), .B2(n7442), .A(n6124), .ZN(n6495) );
  XOR2_X1 U6862 ( .A(DATAI_31_), .B(keyinput_0), .Z(n6127) );
  XOR2_X1 U6863 ( .A(DATAI_30_), .B(keyinput_1), .Z(n6126) );
  XOR2_X1 U6864 ( .A(keyinput_2), .B(DATAI_29_), .Z(n6125) );
  AOI21_X1 U6865 ( .B1(n6127), .B2(n6126), .A(n6125), .ZN(n6130) );
  XNOR2_X1 U6866 ( .A(keyinput_3), .B(DATAI_28_), .ZN(n6129) );
  XNOR2_X1 U6867 ( .A(keyinput_4), .B(DATAI_27_), .ZN(n6128) );
  NOR3_X1 U6868 ( .A1(n6130), .A2(n6129), .A3(n6128), .ZN(n6133) );
  XOR2_X1 U6869 ( .A(keyinput_5), .B(DATAI_26_), .Z(n6132) );
  XNOR2_X1 U6870 ( .A(keyinput_6), .B(DATAI_25_), .ZN(n6131) );
  OAI21_X1 U6871 ( .B1(n6133), .B2(n6132), .A(n6131), .ZN(n6136) );
  XOR2_X1 U6872 ( .A(keyinput_7), .B(DATAI_24_), .Z(n6135) );
  XNOR2_X1 U6873 ( .A(keyinput_8), .B(DATAI_23_), .ZN(n6134) );
  NAND3_X1 U6874 ( .A1(n6136), .A2(n6135), .A3(n6134), .ZN(n6140) );
  XNOR2_X1 U6875 ( .A(keyinput_9), .B(DATAI_22_), .ZN(n6139) );
  XOR2_X1 U6876 ( .A(keyinput_10), .B(DATAI_21_), .Z(n6138) );
  XNOR2_X1 U6877 ( .A(keyinput_11), .B(DATAI_20_), .ZN(n6137) );
  AOI211_X1 U6878 ( .C1(n6140), .C2(n6139), .A(n6138), .B(n6137), .ZN(n6144)
         );
  XOR2_X1 U6879 ( .A(keyinput_12), .B(DATAI_19_), .Z(n6143) );
  XOR2_X1 U6880 ( .A(keyinput_14), .B(DATAI_17_), .Z(n6142) );
  XNOR2_X1 U6881 ( .A(keyinput_13), .B(DATAI_18_), .ZN(n6141) );
  OAI211_X1 U6882 ( .C1(n6144), .C2(n6143), .A(n6142), .B(n6141), .ZN(n6147)
         );
  XOR2_X1 U6883 ( .A(keyinput_15), .B(DATAI_16_), .Z(n6146) );
  XNOR2_X1 U6884 ( .A(keyinput_16), .B(DATAI_15_), .ZN(n6145) );
  AOI21_X1 U6885 ( .B1(n6147), .B2(n6146), .A(n6145), .ZN(n6150) );
  XOR2_X1 U6886 ( .A(DATAI_14_), .B(keyinput_17), .Z(n6149) );
  XOR2_X1 U6887 ( .A(keyinput_18), .B(DATAI_13_), .Z(n6148) );
  OAI21_X1 U6888 ( .B1(n6150), .B2(n6149), .A(n6148), .ZN(n6153) );
  XOR2_X1 U6889 ( .A(keyinput_19), .B(DATAI_12_), .Z(n6152) );
  XNOR2_X1 U6890 ( .A(keyinput_20), .B(DATAI_11_), .ZN(n6151) );
  NAND3_X1 U6891 ( .A1(n6153), .A2(n6152), .A3(n6151), .ZN(n6156) );
  XNOR2_X1 U6892 ( .A(keyinput_21), .B(DATAI_10_), .ZN(n6155) );
  XOR2_X1 U6893 ( .A(keyinput_22), .B(DATAI_9_), .Z(n6154) );
  AOI21_X1 U6894 ( .B1(n6156), .B2(n6155), .A(n6154), .ZN(n6159) );
  XOR2_X1 U6895 ( .A(keyinput_24), .B(DATAI_7_), .Z(n6158) );
  XNOR2_X1 U6896 ( .A(keyinput_23), .B(DATAI_8_), .ZN(n6157) );
  NOR3_X1 U6897 ( .A1(n6159), .A2(n6158), .A3(n6157), .ZN(n6162) );
  XOR2_X1 U6898 ( .A(keyinput_25), .B(DATAI_6_), .Z(n6161) );
  XOR2_X1 U6899 ( .A(keyinput_26), .B(DATAI_5_), .Z(n6160) );
  NOR3_X1 U6900 ( .A1(n6162), .A2(n6161), .A3(n6160), .ZN(n6168) );
  XNOR2_X1 U6901 ( .A(keyinput_27), .B(DATAI_4_), .ZN(n6167) );
  XOR2_X1 U6902 ( .A(keyinput_30), .B(DATAI_1_), .Z(n6165) );
  XNOR2_X1 U6903 ( .A(keyinput_28), .B(DATAI_3_), .ZN(n6164) );
  XNOR2_X1 U6904 ( .A(keyinput_29), .B(DATAI_2_), .ZN(n6163) );
  NOR3_X1 U6905 ( .A1(n6165), .A2(n6164), .A3(n6163), .ZN(n6166) );
  OAI21_X1 U6906 ( .B1(n6168), .B2(n6167), .A(n6166), .ZN(n6171) );
  XNOR2_X1 U6907 ( .A(keyinput_31), .B(DATAI_0_), .ZN(n6170) );
  XOR2_X1 U6908 ( .A(keyinput_32), .B(MEMORYFETCH_REG_SCAN_IN), .Z(n6169) );
  AOI21_X1 U6909 ( .B1(n6171), .B2(n6170), .A(n6169), .ZN(n6174) );
  XOR2_X1 U6910 ( .A(keyinput_33), .B(NA_N), .Z(n6173) );
  XNOR2_X1 U6911 ( .A(keyinput_34), .B(BS16_N), .ZN(n6172) );
  NOR3_X1 U6912 ( .A1(n6174), .A2(n6173), .A3(n6172), .ZN(n6177) );
  XNOR2_X1 U6913 ( .A(READY_N), .B(keyinput_35), .ZN(n6176) );
  XNOR2_X1 U6914 ( .A(keyinput_36), .B(HOLD), .ZN(n6175) );
  OAI21_X1 U6915 ( .B1(n6177), .B2(n6176), .A(n6175), .ZN(n6185) );
  INV_X1 U6916 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6994) );
  XNOR2_X1 U6917 ( .A(n6994), .B(keyinput_38), .ZN(n6181) );
  INV_X1 U6918 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n7179) );
  OAI22_X1 U6919 ( .A1(n7179), .A2(keyinput_37), .B1(CODEFETCH_REG_SCAN_IN), 
        .B2(keyinput_39), .ZN(n6178) );
  AOI21_X1 U6920 ( .B1(n7179), .B2(keyinput_37), .A(n6178), .ZN(n6179) );
  INV_X1 U6921 ( .A(n6179), .ZN(n6180) );
  AOI211_X1 U6922 ( .C1(CODEFETCH_REG_SCAN_IN), .C2(keyinput_39), .A(n6181), 
        .B(n6180), .ZN(n6184) );
  INV_X1 U6923 ( .A(D_C_N_REG_SCAN_IN), .ZN(n7172) );
  XNOR2_X1 U6924 ( .A(n7172), .B(keyinput_41), .ZN(n6183) );
  XNOR2_X1 U6925 ( .A(keyinput_40), .B(M_IO_N_REG_SCAN_IN), .ZN(n6182) );
  AOI211_X1 U6926 ( .C1(n6185), .C2(n6184), .A(n6183), .B(n6182), .ZN(n6189)
         );
  XNOR2_X1 U6927 ( .A(keyinput_42), .B(REQUESTPENDING_REG_SCAN_IN), .ZN(n6188)
         );
  XNOR2_X1 U6928 ( .A(n7520), .B(keyinput_43), .ZN(n6187) );
  XNOR2_X1 U6929 ( .A(keyinput_44), .B(MORE_REG_SCAN_IN), .ZN(n6186) );
  OAI211_X1 U6930 ( .C1(n6189), .C2(n6188), .A(n6187), .B(n6186), .ZN(n6192)
         );
  XOR2_X1 U6931 ( .A(keyinput_46), .B(W_R_N_REG_SCAN_IN), .Z(n6191) );
  XNOR2_X1 U6932 ( .A(keyinput_45), .B(FLUSH_REG_SCAN_IN), .ZN(n6190) );
  NAND3_X1 U6933 ( .A1(n6192), .A2(n6191), .A3(n6190), .ZN(n6203) );
  XOR2_X1 U6934 ( .A(keyinput_48), .B(BYTEENABLE_REG_1__SCAN_IN), .Z(n6196) );
  XNOR2_X1 U6935 ( .A(keyinput_47), .B(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6195)
         );
  XNOR2_X1 U6936 ( .A(keyinput_49), .B(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6194)
         );
  XNOR2_X1 U6937 ( .A(keyinput_50), .B(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6193)
         );
  NOR4_X1 U6938 ( .A1(n6196), .A2(n6195), .A3(n6194), .A4(n6193), .ZN(n6202)
         );
  XOR2_X1 U6939 ( .A(REIP_REG_31__SCAN_IN), .B(keyinput_51), .Z(n6200) );
  XOR2_X1 U6940 ( .A(REIP_REG_29__SCAN_IN), .B(keyinput_53), .Z(n6199) );
  XNOR2_X1 U6941 ( .A(REIP_REG_28__SCAN_IN), .B(keyinput_54), .ZN(n6198) );
  XNOR2_X1 U6942 ( .A(REIP_REG_30__SCAN_IN), .B(keyinput_52), .ZN(n6197) );
  NAND4_X1 U6943 ( .A1(n6200), .A2(n6199), .A3(n6198), .A4(n6197), .ZN(n6201)
         );
  AOI21_X1 U6944 ( .B1(n6203), .B2(n6202), .A(n6201), .ZN(n6216) );
  XNOR2_X1 U6945 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_60), .ZN(n6205) );
  XNOR2_X1 U6946 ( .A(keyinput_59), .B(REIP_REG_23__SCAN_IN), .ZN(n6204) );
  NOR2_X1 U6947 ( .A1(n6205), .A2(n6204), .ZN(n6212) );
  XNOR2_X1 U6948 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_58), .ZN(n6207) );
  XNOR2_X1 U6949 ( .A(REIP_REG_26__SCAN_IN), .B(keyinput_56), .ZN(n6206) );
  NOR2_X1 U6950 ( .A1(n6207), .A2(n6206), .ZN(n6211) );
  INV_X1 U6951 ( .A(keyinput_55), .ZN(n6208) );
  XNOR2_X1 U6952 ( .A(n6208), .B(REIP_REG_27__SCAN_IN), .ZN(n6210) );
  XNOR2_X1 U6953 ( .A(keyinput_57), .B(REIP_REG_25__SCAN_IN), .ZN(n6209) );
  NAND4_X1 U6954 ( .A1(n6212), .A2(n6211), .A3(n6210), .A4(n6209), .ZN(n6215)
         );
  XOR2_X1 U6955 ( .A(keyinput_61), .B(REIP_REG_21__SCAN_IN), .Z(n6214) );
  XNOR2_X1 U6956 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_62), .ZN(n6213) );
  OAI211_X1 U6957 ( .C1(n6216), .C2(n6215), .A(n6214), .B(n6213), .ZN(n6220)
         );
  XOR2_X1 U6958 ( .A(keyinput_63), .B(REIP_REG_19__SCAN_IN), .Z(n6219) );
  XOR2_X1 U6959 ( .A(keyinput_65), .B(REIP_REG_17__SCAN_IN), .Z(n6218) );
  XOR2_X1 U6960 ( .A(keyinput_64), .B(REIP_REG_18__SCAN_IN), .Z(n6217) );
  AOI211_X1 U6961 ( .C1(n6220), .C2(n6219), .A(n6218), .B(n6217), .ZN(n6224)
         );
  XOR2_X1 U6962 ( .A(keyinput_67), .B(BE_N_REG_3__SCAN_IN), .Z(n6223) );
  XNOR2_X1 U6963 ( .A(keyinput_68), .B(BE_N_REG_2__SCAN_IN), .ZN(n6222) );
  XNOR2_X1 U6964 ( .A(keyinput_66), .B(REIP_REG_16__SCAN_IN), .ZN(n6221) );
  NOR4_X1 U6965 ( .A1(n6224), .A2(n6223), .A3(n6222), .A4(n6221), .ZN(n6226)
         );
  XOR2_X1 U6966 ( .A(keyinput_69), .B(BE_N_REG_1__SCAN_IN), .Z(n6225) );
  NOR2_X1 U6967 ( .A1(n6226), .A2(n6225), .ZN(n6234) );
  XNOR2_X1 U6968 ( .A(keyinput_71), .B(ADDRESS_REG_29__SCAN_IN), .ZN(n6230) );
  XNOR2_X1 U6969 ( .A(keyinput_70), .B(BE_N_REG_0__SCAN_IN), .ZN(n6229) );
  XNOR2_X1 U6970 ( .A(keyinput_72), .B(ADDRESS_REG_28__SCAN_IN), .ZN(n6228) );
  XNOR2_X1 U6971 ( .A(keyinput_73), .B(ADDRESS_REG_27__SCAN_IN), .ZN(n6227) );
  NAND4_X1 U6972 ( .A1(n6230), .A2(n6229), .A3(n6228), .A4(n6227), .ZN(n6233)
         );
  INV_X1 U6973 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n7060) );
  XNOR2_X1 U6974 ( .A(n7060), .B(keyinput_74), .ZN(n6232) );
  XNOR2_X1 U6975 ( .A(keyinput_75), .B(ADDRESS_REG_25__SCAN_IN), .ZN(n6231) );
  OAI211_X1 U6976 ( .C1(n6234), .C2(n6233), .A(n6232), .B(n6231), .ZN(n6237)
         );
  INV_X1 U6977 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n7057) );
  XNOR2_X1 U6978 ( .A(n7057), .B(keyinput_76), .ZN(n6236) );
  XNOR2_X1 U6979 ( .A(keyinput_77), .B(ADDRESS_REG_23__SCAN_IN), .ZN(n6235) );
  AOI21_X1 U6980 ( .B1(n6237), .B2(n6236), .A(n6235), .ZN(n6241) );
  INV_X1 U6981 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n7054) );
  XNOR2_X1 U6982 ( .A(n7054), .B(keyinput_78), .ZN(n6240) );
  XNOR2_X1 U6983 ( .A(keyinput_79), .B(ADDRESS_REG_21__SCAN_IN), .ZN(n6239) );
  XNOR2_X1 U6984 ( .A(keyinput_80), .B(ADDRESS_REG_20__SCAN_IN), .ZN(n6238) );
  OAI211_X1 U6985 ( .C1(n6241), .C2(n6240), .A(n6239), .B(n6238), .ZN(n6245)
         );
  INV_X1 U6986 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n7049) );
  XNOR2_X1 U6987 ( .A(n7049), .B(keyinput_82), .ZN(n6244) );
  INV_X1 U6988 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n7050) );
  XNOR2_X1 U6989 ( .A(n7050), .B(keyinput_81), .ZN(n6243) );
  XNOR2_X1 U6990 ( .A(keyinput_83), .B(ADDRESS_REG_17__SCAN_IN), .ZN(n6242) );
  NAND4_X1 U6991 ( .A1(n6245), .A2(n6244), .A3(n6243), .A4(n6242), .ZN(n6249)
         );
  XNOR2_X1 U6992 ( .A(keyinput_84), .B(ADDRESS_REG_16__SCAN_IN), .ZN(n6248) );
  INV_X1 U6993 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n7043) );
  XNOR2_X1 U6994 ( .A(n7043), .B(keyinput_86), .ZN(n6247) );
  XNOR2_X1 U6995 ( .A(keyinput_85), .B(ADDRESS_REG_15__SCAN_IN), .ZN(n6246) );
  AOI211_X1 U6996 ( .C1(n6249), .C2(n6248), .A(n6247), .B(n6246), .ZN(n6252)
         );
  INV_X1 U6997 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n7041) );
  XNOR2_X1 U6998 ( .A(n7041), .B(keyinput_88), .ZN(n6251) );
  XNOR2_X1 U6999 ( .A(keyinput_87), .B(ADDRESS_REG_13__SCAN_IN), .ZN(n6250) );
  NOR3_X1 U7000 ( .A1(n6252), .A2(n6251), .A3(n6250), .ZN(n6259) );
  INV_X1 U7001 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n7039) );
  XNOR2_X1 U7002 ( .A(n7039), .B(keyinput_89), .ZN(n6255) );
  XNOR2_X1 U7003 ( .A(keyinput_90), .B(ADDRESS_REG_10__SCAN_IN), .ZN(n6254) );
  XNOR2_X1 U7004 ( .A(keyinput_91), .B(ADDRESS_REG_9__SCAN_IN), .ZN(n6253) );
  NAND3_X1 U7005 ( .A1(n6255), .A2(n6254), .A3(n6253), .ZN(n6258) );
  XNOR2_X1 U7006 ( .A(keyinput_93), .B(ADDRESS_REG_7__SCAN_IN), .ZN(n6257) );
  XNOR2_X1 U7007 ( .A(keyinput_92), .B(ADDRESS_REG_8__SCAN_IN), .ZN(n6256) );
  OAI211_X1 U7008 ( .C1(n6259), .C2(n6258), .A(n6257), .B(n6256), .ZN(n6262)
         );
  XOR2_X1 U7009 ( .A(keyinput_94), .B(ADDRESS_REG_6__SCAN_IN), .Z(n6261) );
  XOR2_X1 U7010 ( .A(keyinput_95), .B(ADDRESS_REG_5__SCAN_IN), .Z(n6260) );
  NAND3_X1 U7011 ( .A1(n6262), .A2(n6261), .A3(n6260), .ZN(n6265) );
  XNOR2_X1 U7012 ( .A(keyinput_96), .B(ADDRESS_REG_4__SCAN_IN), .ZN(n6264) );
  INV_X1 U7013 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n7029) );
  XNOR2_X1 U7014 ( .A(n7029), .B(keyinput_97), .ZN(n6263) );
  AOI21_X1 U7015 ( .B1(n6265), .B2(n6264), .A(n6263), .ZN(n6268) );
  XNOR2_X1 U7016 ( .A(keyinput_99), .B(ADDRESS_REG_1__SCAN_IN), .ZN(n6267) );
  XNOR2_X1 U7017 ( .A(keyinput_98), .B(ADDRESS_REG_2__SCAN_IN), .ZN(n6266) );
  NOR3_X1 U7018 ( .A1(n6268), .A2(n6267), .A3(n6266), .ZN(n6271) );
  INV_X1 U7019 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n7025) );
  XNOR2_X1 U7020 ( .A(n7025), .B(keyinput_100), .ZN(n6270) );
  XNOR2_X1 U7021 ( .A(STATE_REG_2__SCAN_IN), .B(keyinput_101), .ZN(n6269) );
  NOR3_X1 U7022 ( .A1(n6271), .A2(n6270), .A3(n6269), .ZN(n6274) );
  XNOR2_X1 U7023 ( .A(STATE_REG_1__SCAN_IN), .B(keyinput_102), .ZN(n6273) );
  XNOR2_X1 U7024 ( .A(n7535), .B(keyinput_103), .ZN(n6272) );
  OAI21_X1 U7025 ( .B1(n6274), .B2(n6273), .A(n6272), .ZN(n6277) );
  XOR2_X1 U7026 ( .A(keyinput_104), .B(DATAWIDTH_REG_0__SCAN_IN), .Z(n6276) );
  XOR2_X1 U7027 ( .A(keyinput_105), .B(DATAWIDTH_REG_1__SCAN_IN), .Z(n6275) );
  AOI21_X1 U7028 ( .B1(n6277), .B2(n6276), .A(n6275), .ZN(n6280) );
  XOR2_X1 U7029 ( .A(keyinput_106), .B(DATAWIDTH_REG_2__SCAN_IN), .Z(n6279) );
  XNOR2_X1 U7030 ( .A(keyinput_107), .B(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6278)
         );
  NOR3_X1 U7031 ( .A1(n6280), .A2(n6279), .A3(n6278), .ZN(n6286) );
  XNOR2_X1 U7032 ( .A(keyinput_108), .B(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6285)
         );
  XOR2_X1 U7033 ( .A(keyinput_111), .B(DATAWIDTH_REG_7__SCAN_IN), .Z(n6283) );
  INV_X1 U7034 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6984) );
  XNOR2_X1 U7035 ( .A(n6984), .B(keyinput_110), .ZN(n6282) );
  INV_X1 U7036 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6983) );
  XNOR2_X1 U7037 ( .A(n6983), .B(keyinput_109), .ZN(n6281) );
  NOR3_X1 U7038 ( .A1(n6283), .A2(n6282), .A3(n6281), .ZN(n6284) );
  OAI21_X1 U7039 ( .B1(n6286), .B2(n6285), .A(n6284), .ZN(n6289) );
  XOR2_X1 U7040 ( .A(keyinput_112), .B(DATAWIDTH_REG_8__SCAN_IN), .Z(n6288) );
  XNOR2_X1 U7041 ( .A(keyinput_113), .B(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6287)
         );
  NAND3_X1 U7042 ( .A1(n6289), .A2(n6288), .A3(n6287), .ZN(n6297) );
  XOR2_X1 U7043 ( .A(keyinput_116), .B(DATAWIDTH_REG_12__SCAN_IN), .Z(n6293)
         );
  XOR2_X1 U7044 ( .A(keyinput_117), .B(DATAWIDTH_REG_13__SCAN_IN), .Z(n6292)
         );
  INV_X1 U7045 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6986) );
  XNOR2_X1 U7046 ( .A(n6986), .B(keyinput_114), .ZN(n6291) );
  XNOR2_X1 U7047 ( .A(keyinput_115), .B(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6290)
         );
  NOR4_X1 U7048 ( .A1(n6293), .A2(n6292), .A3(n6291), .A4(n6290), .ZN(n6296)
         );
  XOR2_X1 U7049 ( .A(keyinput_119), .B(DATAWIDTH_REG_15__SCAN_IN), .Z(n6295)
         );
  INV_X1 U7050 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6987) );
  XNOR2_X1 U7051 ( .A(n6987), .B(keyinput_118), .ZN(n6294) );
  AOI211_X1 U7052 ( .C1(n6297), .C2(n6296), .A(n6295), .B(n6294), .ZN(n6301)
         );
  XOR2_X1 U7053 ( .A(keyinput_121), .B(DATAWIDTH_REG_17__SCAN_IN), .Z(n6300)
         );
  XNOR2_X1 U7054 ( .A(keyinput_122), .B(DATAWIDTH_REG_18__SCAN_IN), .ZN(n6299)
         );
  XNOR2_X1 U7055 ( .A(keyinput_120), .B(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6298)
         );
  NOR4_X1 U7056 ( .A1(n6301), .A2(n6300), .A3(n6299), .A4(n6298), .ZN(n6304)
         );
  XOR2_X1 U7057 ( .A(keyinput_123), .B(DATAWIDTH_REG_19__SCAN_IN), .Z(n6303)
         );
  XNOR2_X1 U7058 ( .A(keyinput_124), .B(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6302)
         );
  OAI21_X1 U7059 ( .B1(n6304), .B2(n6303), .A(n6302), .ZN(n6308) );
  INV_X1 U7060 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6990) );
  XNOR2_X1 U7061 ( .A(n6990), .B(keyinput_126), .ZN(n6307) );
  XNOR2_X1 U7062 ( .A(keyinput_127), .B(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6306)
         );
  XNOR2_X1 U7063 ( .A(DATAWIDTH_REG_21__SCAN_IN), .B(keyinput_125), .ZN(n6305)
         );
  NAND4_X1 U7064 ( .A1(n6308), .A2(n6307), .A3(n6306), .A4(n6305), .ZN(n6493)
         );
  XNOR2_X1 U7065 ( .A(DATAI_30_), .B(keyinput_129), .ZN(n6311) );
  XNOR2_X1 U7066 ( .A(DATAI_31_), .B(keyinput_128), .ZN(n6310) );
  XOR2_X1 U7067 ( .A(DATAI_29_), .B(keyinput_130), .Z(n6309) );
  OAI21_X1 U7068 ( .B1(n6311), .B2(n6310), .A(n6309), .ZN(n6314) );
  XOR2_X1 U7069 ( .A(DATAI_27_), .B(keyinput_132), .Z(n6313) );
  XNOR2_X1 U7070 ( .A(DATAI_28_), .B(keyinput_131), .ZN(n6312) );
  NAND3_X1 U7071 ( .A1(n6314), .A2(n6313), .A3(n6312), .ZN(n6317) );
  XNOR2_X1 U7072 ( .A(DATAI_26_), .B(keyinput_133), .ZN(n6316) );
  XOR2_X1 U7073 ( .A(DATAI_25_), .B(keyinput_134), .Z(n6315) );
  AOI21_X1 U7074 ( .B1(n6317), .B2(n6316), .A(n6315), .ZN(n6320) );
  XOR2_X1 U7075 ( .A(DATAI_24_), .B(keyinput_135), .Z(n6319) );
  XOR2_X1 U7076 ( .A(DATAI_23_), .B(keyinput_136), .Z(n6318) );
  NOR3_X1 U7077 ( .A1(n6320), .A2(n6319), .A3(n6318), .ZN(n6324) );
  XOR2_X1 U7078 ( .A(DATAI_22_), .B(keyinput_137), .Z(n6323) );
  XNOR2_X1 U7079 ( .A(DATAI_20_), .B(keyinput_139), .ZN(n6322) );
  XNOR2_X1 U7080 ( .A(DATAI_21_), .B(keyinput_138), .ZN(n6321) );
  OAI211_X1 U7081 ( .C1(n6324), .C2(n6323), .A(n6322), .B(n6321), .ZN(n6328)
         );
  XNOR2_X1 U7082 ( .A(DATAI_19_), .B(keyinput_140), .ZN(n6327) );
  XOR2_X1 U7083 ( .A(DATAI_17_), .B(keyinput_142), .Z(n6326) );
  XNOR2_X1 U7084 ( .A(DATAI_18_), .B(keyinput_141), .ZN(n6325) );
  AOI211_X1 U7085 ( .C1(n6328), .C2(n6327), .A(n6326), .B(n6325), .ZN(n6331)
         );
  XOR2_X1 U7086 ( .A(DATAI_16_), .B(keyinput_143), .Z(n6330) );
  XOR2_X1 U7087 ( .A(DATAI_15_), .B(keyinput_144), .Z(n6329) );
  OAI21_X1 U7088 ( .B1(n6331), .B2(n6330), .A(n6329), .ZN(n6334) );
  XNOR2_X1 U7089 ( .A(DATAI_14_), .B(keyinput_145), .ZN(n6333) );
  XOR2_X1 U7090 ( .A(DATAI_13_), .B(keyinput_146), .Z(n6332) );
  AOI21_X1 U7091 ( .B1(n6334), .B2(n6333), .A(n6332), .ZN(n6337) );
  XOR2_X1 U7092 ( .A(DATAI_12_), .B(keyinput_147), .Z(n6336) );
  XOR2_X1 U7093 ( .A(DATAI_11_), .B(keyinput_148), .Z(n6335) );
  NOR3_X1 U7094 ( .A1(n6337), .A2(n6336), .A3(n6335), .ZN(n6340) );
  XOR2_X1 U7095 ( .A(DATAI_10_), .B(keyinput_149), .Z(n6339) );
  XNOR2_X1 U7096 ( .A(DATAI_9_), .B(keyinput_150), .ZN(n6338) );
  OAI21_X1 U7097 ( .B1(n6340), .B2(n6339), .A(n6338), .ZN(n6343) );
  XNOR2_X1 U7098 ( .A(DATAI_8_), .B(keyinput_151), .ZN(n6342) );
  XNOR2_X1 U7099 ( .A(DATAI_7_), .B(keyinput_152), .ZN(n6341) );
  NAND3_X1 U7100 ( .A1(n6343), .A2(n6342), .A3(n6341), .ZN(n6346) );
  XOR2_X1 U7101 ( .A(DATAI_6_), .B(keyinput_153), .Z(n6345) );
  XNOR2_X1 U7102 ( .A(DATAI_5_), .B(keyinput_154), .ZN(n6344) );
  NAND3_X1 U7103 ( .A1(n6346), .A2(n6345), .A3(n6344), .ZN(n6352) );
  XNOR2_X1 U7104 ( .A(DATAI_4_), .B(keyinput_155), .ZN(n6351) );
  XNOR2_X1 U7105 ( .A(DATAI_1_), .B(keyinput_158), .ZN(n6349) );
  XNOR2_X1 U7106 ( .A(DATAI_2_), .B(keyinput_157), .ZN(n6348) );
  XNOR2_X1 U7107 ( .A(DATAI_3_), .B(keyinput_156), .ZN(n6347) );
  NAND3_X1 U7108 ( .A1(n6349), .A2(n6348), .A3(n6347), .ZN(n6350) );
  AOI21_X1 U7109 ( .B1(n6352), .B2(n6351), .A(n6350), .ZN(n6355) );
  XNOR2_X1 U7110 ( .A(DATAI_0_), .B(keyinput_159), .ZN(n6354) );
  XNOR2_X1 U7111 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(keyinput_160), .ZN(n6353)
         );
  OAI21_X1 U7112 ( .B1(n6355), .B2(n6354), .A(n6353), .ZN(n6358) );
  XOR2_X1 U7113 ( .A(NA_N), .B(keyinput_161), .Z(n6357) );
  XNOR2_X1 U7114 ( .A(BS16_N), .B(keyinput_162), .ZN(n6356) );
  NAND3_X1 U7115 ( .A1(n6358), .A2(n6357), .A3(n6356), .ZN(n6361) );
  XNOR2_X1 U7116 ( .A(n7502), .B(keyinput_163), .ZN(n6360) );
  XOR2_X1 U7117 ( .A(HOLD), .B(keyinput_164), .Z(n6359) );
  AOI21_X1 U7118 ( .B1(n6361), .B2(n6360), .A(n6359), .ZN(n6365) );
  XNOR2_X1 U7119 ( .A(n6994), .B(keyinput_166), .ZN(n6364) );
  XNOR2_X1 U7120 ( .A(READREQUEST_REG_SCAN_IN), .B(keyinput_165), .ZN(n6363)
         );
  XNOR2_X1 U7121 ( .A(CODEFETCH_REG_SCAN_IN), .B(keyinput_167), .ZN(n6362) );
  NOR4_X1 U7122 ( .A1(n6365), .A2(n6364), .A3(n6363), .A4(n6362), .ZN(n6368)
         );
  INV_X1 U7123 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n7541) );
  XNOR2_X1 U7124 ( .A(n7541), .B(keyinput_168), .ZN(n6367) );
  XNOR2_X1 U7125 ( .A(D_C_N_REG_SCAN_IN), .B(keyinput_169), .ZN(n6366) );
  NOR3_X1 U7126 ( .A1(n6368), .A2(n6367), .A3(n6366), .ZN(n6372) );
  XOR2_X1 U7127 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(keyinput_170), .Z(n6371)
         );
  XNOR2_X1 U7128 ( .A(n7520), .B(keyinput_171), .ZN(n6370) );
  XOR2_X1 U7129 ( .A(MORE_REG_SCAN_IN), .B(keyinput_172), .Z(n6369) );
  OAI211_X1 U7130 ( .C1(n6372), .C2(n6371), .A(n6370), .B(n6369), .ZN(n6375)
         );
  XOR2_X1 U7131 ( .A(W_R_N_REG_SCAN_IN), .B(keyinput_174), .Z(n6374) );
  XOR2_X1 U7132 ( .A(FLUSH_REG_SCAN_IN), .B(keyinput_173), .Z(n6373) );
  NAND3_X1 U7133 ( .A1(n6375), .A2(n6374), .A3(n6373), .ZN(n6386) );
  XOR2_X1 U7134 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_175), .Z(n6379)
         );
  XNOR2_X1 U7135 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(keyinput_177), .ZN(n6378)
         );
  XNOR2_X1 U7136 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(keyinput_176), .ZN(n6377)
         );
  XNOR2_X1 U7137 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_178), .ZN(n6376)
         );
  NOR4_X1 U7138 ( .A1(n6379), .A2(n6378), .A3(n6377), .A4(n6376), .ZN(n6385)
         );
  XOR2_X1 U7139 ( .A(REIP_REG_29__SCAN_IN), .B(keyinput_181), .Z(n6383) );
  XOR2_X1 U7140 ( .A(REIP_REG_28__SCAN_IN), .B(keyinput_182), .Z(n6382) );
  XOR2_X1 U7141 ( .A(REIP_REG_30__SCAN_IN), .B(keyinput_180), .Z(n6381) );
  XNOR2_X1 U7142 ( .A(REIP_REG_31__SCAN_IN), .B(keyinput_179), .ZN(n6380) );
  NAND4_X1 U7143 ( .A1(n6383), .A2(n6382), .A3(n6381), .A4(n6380), .ZN(n6384)
         );
  AOI21_X1 U7144 ( .B1(n6386), .B2(n6385), .A(n6384), .ZN(n6398) );
  XNOR2_X1 U7145 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_188), .ZN(n6388) );
  XNOR2_X1 U7146 ( .A(REIP_REG_23__SCAN_IN), .B(keyinput_187), .ZN(n6387) );
  NOR2_X1 U7147 ( .A1(n6388), .A2(n6387), .ZN(n6394) );
  XNOR2_X1 U7148 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_186), .ZN(n6390) );
  XNOR2_X1 U7149 ( .A(REIP_REG_26__SCAN_IN), .B(keyinput_184), .ZN(n6389) );
  NOR2_X1 U7150 ( .A1(n6390), .A2(n6389), .ZN(n6393) );
  XNOR2_X1 U7151 ( .A(REIP_REG_27__SCAN_IN), .B(keyinput_183), .ZN(n6392) );
  XNOR2_X1 U7152 ( .A(REIP_REG_25__SCAN_IN), .B(keyinput_185), .ZN(n6391) );
  NAND4_X1 U7153 ( .A1(n6394), .A2(n6393), .A3(n6392), .A4(n6391), .ZN(n6397)
         );
  XOR2_X1 U7154 ( .A(REIP_REG_21__SCAN_IN), .B(keyinput_189), .Z(n6396) );
  XOR2_X1 U7155 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_190), .Z(n6395) );
  OAI211_X1 U7156 ( .C1(n6398), .C2(n6397), .A(n6396), .B(n6395), .ZN(n6402)
         );
  XOR2_X1 U7157 ( .A(REIP_REG_19__SCAN_IN), .B(keyinput_191), .Z(n6401) );
  XOR2_X1 U7158 ( .A(REIP_REG_18__SCAN_IN), .B(keyinput_192), .Z(n6400) );
  XNOR2_X1 U7159 ( .A(REIP_REG_17__SCAN_IN), .B(keyinput_193), .ZN(n6399) );
  AOI211_X1 U7160 ( .C1(n6402), .C2(n6401), .A(n6400), .B(n6399), .ZN(n6407)
         );
  INV_X1 U7161 ( .A(keyinput_196), .ZN(n6403) );
  XNOR2_X1 U7162 ( .A(n6403), .B(BE_N_REG_2__SCAN_IN), .ZN(n6406) );
  XNOR2_X1 U7163 ( .A(BE_N_REG_3__SCAN_IN), .B(keyinput_195), .ZN(n6405) );
  XNOR2_X1 U7164 ( .A(REIP_REG_16__SCAN_IN), .B(keyinput_194), .ZN(n6404) );
  NOR4_X1 U7165 ( .A1(n6407), .A2(n6406), .A3(n6405), .A4(n6404), .ZN(n6414)
         );
  XNOR2_X1 U7166 ( .A(BE_N_REG_1__SCAN_IN), .B(keyinput_197), .ZN(n6413) );
  INV_X1 U7167 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n7069) );
  XNOR2_X1 U7168 ( .A(n7069), .B(keyinput_199), .ZN(n6411) );
  INV_X1 U7169 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n7065) );
  XNOR2_X1 U7170 ( .A(n7065), .B(keyinput_200), .ZN(n6410) );
  INV_X1 U7171 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n7102) );
  XNOR2_X1 U7172 ( .A(n7102), .B(keyinput_198), .ZN(n6409) );
  XNOR2_X1 U7173 ( .A(ADDRESS_REG_27__SCAN_IN), .B(keyinput_201), .ZN(n6408)
         );
  NOR4_X1 U7174 ( .A1(n6411), .A2(n6410), .A3(n6409), .A4(n6408), .ZN(n6412)
         );
  OAI21_X1 U7175 ( .B1(n6414), .B2(n6413), .A(n6412), .ZN(n6417) );
  XNOR2_X1 U7176 ( .A(ADDRESS_REG_26__SCAN_IN), .B(keyinput_202), .ZN(n6416)
         );
  XNOR2_X1 U7177 ( .A(ADDRESS_REG_25__SCAN_IN), .B(keyinput_203), .ZN(n6415)
         );
  NAND3_X1 U7178 ( .A1(n6417), .A2(n6416), .A3(n6415), .ZN(n6420) );
  XNOR2_X1 U7179 ( .A(ADDRESS_REG_24__SCAN_IN), .B(keyinput_204), .ZN(n6419)
         );
  XNOR2_X1 U7180 ( .A(ADDRESS_REG_23__SCAN_IN), .B(keyinput_205), .ZN(n6418)
         );
  AOI21_X1 U7181 ( .B1(n6420), .B2(n6419), .A(n6418), .ZN(n6424) );
  XNOR2_X1 U7182 ( .A(n7054), .B(keyinput_206), .ZN(n6423) );
  XNOR2_X1 U7183 ( .A(ADDRESS_REG_20__SCAN_IN), .B(keyinput_208), .ZN(n6422)
         );
  XNOR2_X1 U7184 ( .A(ADDRESS_REG_21__SCAN_IN), .B(keyinput_207), .ZN(n6421)
         );
  OAI211_X1 U7185 ( .C1(n6424), .C2(n6423), .A(n6422), .B(n6421), .ZN(n6428)
         );
  INV_X1 U7186 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n7047) );
  XNOR2_X1 U7187 ( .A(n7047), .B(keyinput_211), .ZN(n6427) );
  XNOR2_X1 U7188 ( .A(ADDRESS_REG_19__SCAN_IN), .B(keyinput_209), .ZN(n6426)
         );
  XNOR2_X1 U7189 ( .A(ADDRESS_REG_18__SCAN_IN), .B(keyinput_210), .ZN(n6425)
         );
  NAND4_X1 U7190 ( .A1(n6428), .A2(n6427), .A3(n6426), .A4(n6425), .ZN(n6432)
         );
  XNOR2_X1 U7191 ( .A(ADDRESS_REG_16__SCAN_IN), .B(keyinput_212), .ZN(n6431)
         );
  XNOR2_X1 U7192 ( .A(n7043), .B(keyinput_214), .ZN(n6430) );
  XNOR2_X1 U7193 ( .A(ADDRESS_REG_15__SCAN_IN), .B(keyinput_213), .ZN(n6429)
         );
  AOI211_X1 U7194 ( .C1(n6432), .C2(n6431), .A(n6430), .B(n6429), .ZN(n6435)
         );
  XNOR2_X1 U7195 ( .A(ADDRESS_REG_13__SCAN_IN), .B(keyinput_215), .ZN(n6434)
         );
  XNOR2_X1 U7196 ( .A(ADDRESS_REG_12__SCAN_IN), .B(keyinput_216), .ZN(n6433)
         );
  NOR3_X1 U7197 ( .A1(n6435), .A2(n6434), .A3(n6433), .ZN(n6439) );
  XNOR2_X1 U7198 ( .A(n7039), .B(keyinput_217), .ZN(n6438) );
  XNOR2_X1 U7199 ( .A(ADDRESS_REG_9__SCAN_IN), .B(keyinput_219), .ZN(n6437) );
  XNOR2_X1 U7200 ( .A(ADDRESS_REG_10__SCAN_IN), .B(keyinput_218), .ZN(n6436)
         );
  NOR4_X1 U7201 ( .A1(n6439), .A2(n6438), .A3(n6437), .A4(n6436), .ZN(n6442)
         );
  INV_X1 U7202 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n7034) );
  XNOR2_X1 U7203 ( .A(n7034), .B(keyinput_221), .ZN(n6441) );
  INV_X1 U7204 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n7036) );
  XNOR2_X1 U7205 ( .A(n7036), .B(keyinput_220), .ZN(n6440) );
  NOR3_X1 U7206 ( .A1(n6442), .A2(n6441), .A3(n6440), .ZN(n6445) );
  XNOR2_X1 U7207 ( .A(ADDRESS_REG_6__SCAN_IN), .B(keyinput_222), .ZN(n6444) );
  XNOR2_X1 U7208 ( .A(ADDRESS_REG_5__SCAN_IN), .B(keyinput_223), .ZN(n6443) );
  NOR3_X1 U7209 ( .A1(n6445), .A2(n6444), .A3(n6443), .ZN(n6448) );
  INV_X1 U7210 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n7030) );
  XNOR2_X1 U7211 ( .A(n7030), .B(keyinput_224), .ZN(n6447) );
  XNOR2_X1 U7212 ( .A(n7029), .B(keyinput_225), .ZN(n6446) );
  OAI21_X1 U7213 ( .B1(n6448), .B2(n6447), .A(n6446), .ZN(n6451) );
  XOR2_X1 U7214 ( .A(ADDRESS_REG_2__SCAN_IN), .B(keyinput_226), .Z(n6450) );
  XNOR2_X1 U7215 ( .A(ADDRESS_REG_1__SCAN_IN), .B(keyinput_227), .ZN(n6449) );
  NAND3_X1 U7216 ( .A1(n6451), .A2(n6450), .A3(n6449), .ZN(n6454) );
  XNOR2_X1 U7217 ( .A(n7533), .B(keyinput_229), .ZN(n6453) );
  XNOR2_X1 U7218 ( .A(ADDRESS_REG_0__SCAN_IN), .B(keyinput_228), .ZN(n6452) );
  NAND3_X1 U7219 ( .A1(n6454), .A2(n6453), .A3(n6452), .ZN(n6457) );
  XNOR2_X1 U7220 ( .A(STATE_REG_1__SCAN_IN), .B(keyinput_230), .ZN(n6456) );
  XNOR2_X1 U7221 ( .A(n7535), .B(keyinput_231), .ZN(n6455) );
  AOI21_X1 U7222 ( .B1(n6457), .B2(n6456), .A(n6455), .ZN(n6460) );
  XNOR2_X1 U7223 ( .A(DATAWIDTH_REG_0__SCAN_IN), .B(keyinput_232), .ZN(n6459)
         );
  XNOR2_X1 U7224 ( .A(DATAWIDTH_REG_1__SCAN_IN), .B(keyinput_233), .ZN(n6458)
         );
  OAI21_X1 U7225 ( .B1(n6460), .B2(n6459), .A(n6458), .ZN(n6463) );
  XOR2_X1 U7226 ( .A(DATAWIDTH_REG_3__SCAN_IN), .B(keyinput_235), .Z(n6462) );
  XOR2_X1 U7227 ( .A(DATAWIDTH_REG_2__SCAN_IN), .B(keyinput_234), .Z(n6461) );
  NAND3_X1 U7228 ( .A1(n6463), .A2(n6462), .A3(n6461), .ZN(n6469) );
  XNOR2_X1 U7229 ( .A(DATAWIDTH_REG_4__SCAN_IN), .B(keyinput_236), .ZN(n6468)
         );
  XOR2_X1 U7230 ( .A(DATAWIDTH_REG_7__SCAN_IN), .B(keyinput_239), .Z(n6466) );
  XNOR2_X1 U7231 ( .A(DATAWIDTH_REG_5__SCAN_IN), .B(keyinput_237), .ZN(n6465)
         );
  XNOR2_X1 U7232 ( .A(DATAWIDTH_REG_6__SCAN_IN), .B(keyinput_238), .ZN(n6464)
         );
  NAND3_X1 U7233 ( .A1(n6466), .A2(n6465), .A3(n6464), .ZN(n6467) );
  AOI21_X1 U7234 ( .B1(n6469), .B2(n6468), .A(n6467), .ZN(n6472) );
  INV_X1 U7235 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6985) );
  XNOR2_X1 U7236 ( .A(n6985), .B(keyinput_241), .ZN(n6471) );
  XNOR2_X1 U7237 ( .A(DATAWIDTH_REG_8__SCAN_IN), .B(keyinput_240), .ZN(n6470)
         );
  NOR3_X1 U7238 ( .A1(n6472), .A2(n6471), .A3(n6470), .ZN(n6480) );
  XOR2_X1 U7239 ( .A(DATAWIDTH_REG_13__SCAN_IN), .B(keyinput_245), .Z(n6476)
         );
  XOR2_X1 U7240 ( .A(DATAWIDTH_REG_11__SCAN_IN), .B(keyinput_243), .Z(n6475)
         );
  XOR2_X1 U7241 ( .A(DATAWIDTH_REG_12__SCAN_IN), .B(keyinput_244), .Z(n6474)
         );
  XNOR2_X1 U7242 ( .A(DATAWIDTH_REG_10__SCAN_IN), .B(keyinput_242), .ZN(n6473)
         );
  NAND4_X1 U7243 ( .A1(n6476), .A2(n6475), .A3(n6474), .A4(n6473), .ZN(n6479)
         );
  XOR2_X1 U7244 ( .A(DATAWIDTH_REG_15__SCAN_IN), .B(keyinput_247), .Z(n6478)
         );
  XNOR2_X1 U7245 ( .A(DATAWIDTH_REG_14__SCAN_IN), .B(keyinput_246), .ZN(n6477)
         );
  OAI211_X1 U7246 ( .C1(n6480), .C2(n6479), .A(n6478), .B(n6477), .ZN(n6484)
         );
  XOR2_X1 U7247 ( .A(DATAWIDTH_REG_18__SCAN_IN), .B(keyinput_250), .Z(n6483)
         );
  XNOR2_X1 U7248 ( .A(DATAWIDTH_REG_16__SCAN_IN), .B(keyinput_248), .ZN(n6482)
         );
  XNOR2_X1 U7249 ( .A(DATAWIDTH_REG_17__SCAN_IN), .B(keyinput_249), .ZN(n6481)
         );
  NAND4_X1 U7250 ( .A1(n6484), .A2(n6483), .A3(n6482), .A4(n6481), .ZN(n6487)
         );
  XNOR2_X1 U7251 ( .A(DATAWIDTH_REG_19__SCAN_IN), .B(keyinput_251), .ZN(n6486)
         );
  XNOR2_X1 U7252 ( .A(DATAWIDTH_REG_20__SCAN_IN), .B(keyinput_252), .ZN(n6485)
         );
  AOI21_X1 U7253 ( .B1(n6487), .B2(n6486), .A(n6485), .ZN(n6491) );
  XNOR2_X1 U7254 ( .A(n6990), .B(keyinput_254), .ZN(n6490) );
  INV_X1 U7255 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6989) );
  XNOR2_X1 U7256 ( .A(n6989), .B(keyinput_253), .ZN(n6489) );
  XNOR2_X1 U7257 ( .A(DATAWIDTH_REG_23__SCAN_IN), .B(keyinput_255), .ZN(n6488)
         );
  NOR4_X1 U7258 ( .A1(n6491), .A2(n6490), .A3(n6489), .A4(n6488), .ZN(n6492)
         );
  NAND2_X1 U7259 ( .A1(n6493), .A2(n6492), .ZN(n6494) );
  XOR2_X1 U7260 ( .A(n6495), .B(n6494), .Z(U2798) );
  OR2_X1 U7261 ( .A1(n6518), .A2(n6496), .ZN(n6497) );
  NAND2_X1 U7262 ( .A1(n6498), .A2(n6497), .ZN(n6808) );
  OAI21_X1 U7263 ( .B1(n6499), .B2(n6501), .A(n6500), .ZN(n6658) );
  INV_X1 U7264 ( .A(n6658), .ZN(n6695) );
  NAND2_X1 U7265 ( .A1(n6695), .A2(n7442), .ZN(n6510) );
  INV_X1 U7266 ( .A(n6502), .ZN(n6693) );
  OAI22_X1 U7267 ( .A1(n6503), .A2(n7429), .B1(n7445), .B2(n6693), .ZN(n6508)
         );
  INV_X1 U7268 ( .A(REIP_REG_28__SCAN_IN), .ZN(n7063) );
  INV_X1 U7269 ( .A(n6504), .ZN(n6506) );
  AOI21_X1 U7270 ( .B1(n7063), .B2(n6506), .A(n6505), .ZN(n6507) );
  AOI211_X1 U7271 ( .C1(EBX_REG_28__SCAN_IN), .C2(n7419), .A(n6508), .B(n6507), 
        .ZN(n6509) );
  OAI211_X1 U7272 ( .C1(n7421), .C2(n6808), .A(n6510), .B(n6509), .ZN(U2799)
         );
  INV_X1 U7273 ( .A(n6511), .ZN(n6528) );
  AOI21_X1 U7274 ( .B1(n6512), .B2(n6528), .A(n6499), .ZN(n6705) );
  INV_X1 U7275 ( .A(n6705), .ZN(n6661) );
  OAI22_X1 U7276 ( .A1(n6513), .A2(n7429), .B1(n7445), .B2(n6703), .ZN(n6517)
         );
  NOR2_X1 U7277 ( .A1(n7324), .A2(n6514), .ZN(n6515) );
  MUX2_X1 U7278 ( .A(n6515), .B(n6532), .S(REIP_REG_27__SCAN_IN), .Z(n6516) );
  AOI211_X1 U7279 ( .C1(EBX_REG_27__SCAN_IN), .C2(n7419), .A(n6517), .B(n6516), 
        .ZN(n6521) );
  AOI21_X1 U7280 ( .B1(n6519), .B2(n6525), .A(n6518), .ZN(n6821) );
  NAND2_X1 U7281 ( .A1(n6821), .A2(n7441), .ZN(n6520) );
  OAI211_X1 U7282 ( .C1(n6661), .C2(n7422), .A(n6521), .B(n6520), .ZN(U2800)
         );
  NAND2_X1 U7283 ( .A1(n6555), .A2(n6523), .ZN(n6524) );
  NAND2_X1 U7284 ( .A1(n6525), .A2(n6524), .ZN(n6828) );
  AOI21_X1 U7285 ( .B1(n6529), .B2(n6543), .A(n6511), .ZN(n6713) );
  NAND2_X1 U7286 ( .A1(n6713), .A2(n7442), .ZN(n6539) );
  INV_X1 U7287 ( .A(n6530), .ZN(n6711) );
  OAI22_X1 U7288 ( .A1(n6531), .A2(n7429), .B1(n7445), .B2(n6711), .ZN(n6537)
         );
  INV_X1 U7289 ( .A(n6532), .ZN(n6535) );
  AOI21_X1 U7290 ( .B1(n7372), .B2(n6533), .A(REIP_REG_26__SCAN_IN), .ZN(n6534) );
  NOR2_X1 U7291 ( .A1(n6535), .A2(n6534), .ZN(n6536) );
  AOI211_X1 U7292 ( .C1(EBX_REG_26__SCAN_IN), .C2(n7419), .A(n6537), .B(n6536), 
        .ZN(n6538) );
  OAI211_X1 U7293 ( .C1(n6828), .C2(n7421), .A(n6539), .B(n6538), .ZN(U2801)
         );
  INV_X1 U7294 ( .A(n6541), .ZN(n6545) );
  INV_X1 U7295 ( .A(n6542), .ZN(n6544) );
  OAI21_X1 U7296 ( .B1(n6545), .B2(n6544), .A(n6543), .ZN(n6723) );
  OAI21_X1 U7297 ( .B1(n7324), .B2(n6563), .A(n7301), .ZN(n6580) );
  INV_X1 U7298 ( .A(n6546), .ZN(n6547) );
  INV_X1 U7299 ( .A(REIP_REG_24__SCAN_IN), .ZN(n7055) );
  MUX2_X1 U7300 ( .A(n6547), .B(n7055), .S(REIP_REG_25__SCAN_IN), .Z(n6550) );
  OAI22_X1 U7301 ( .A1(n6548), .A2(n7429), .B1(n7445), .B2(n6716), .ZN(n6549)
         );
  AOI21_X1 U7302 ( .B1(n7372), .B2(n6550), .A(n6549), .ZN(n6551) );
  OAI21_X1 U7303 ( .B1(n7435), .B2(n6634), .A(n6551), .ZN(n6557) );
  OR2_X1 U7304 ( .A1(n6552), .A2(n6553), .ZN(n6554) );
  NAND2_X1 U7305 ( .A1(n6555), .A2(n6554), .ZN(n6840) );
  NOR2_X1 U7306 ( .A1(n6840), .A2(n7421), .ZN(n6556) );
  AOI211_X1 U7307 ( .C1(REIP_REG_25__SCAN_IN), .C2(n6580), .A(n6557), .B(n6556), .ZN(n6558) );
  OAI21_X1 U7308 ( .B1(n6723), .B2(n7422), .A(n6558), .ZN(U2802) );
  OAI21_X1 U7309 ( .B1(n6573), .B2(n6560), .A(n6541), .ZN(n6737) );
  NOR2_X1 U7310 ( .A1(n6577), .A2(n6561), .ZN(n6562) );
  OR2_X1 U7311 ( .A1(n6552), .A2(n6562), .ZN(n6635) );
  INV_X1 U7312 ( .A(n6635), .ZN(n6852) );
  INV_X1 U7313 ( .A(n6563), .ZN(n6564) );
  NOR2_X1 U7314 ( .A1(n7324), .A2(n6564), .ZN(n6565) );
  MUX2_X1 U7315 ( .A(n6565), .B(n6580), .S(REIP_REG_24__SCAN_IN), .Z(n6569) );
  AOI22_X1 U7316 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n7439), .B1(n7425), 
        .B2(n6736), .ZN(n6566) );
  OAI21_X1 U7317 ( .B1(n7435), .B2(n6567), .A(n6566), .ZN(n6568) );
  AOI211_X1 U7318 ( .C1(n6852), .C2(n7441), .A(n6569), .B(n6568), .ZN(n6570)
         );
  OAI21_X1 U7319 ( .B1(n6737), .B2(n7422), .A(n6570), .ZN(U2803) );
  AOI21_X1 U7320 ( .B1(n6574), .B2(n6589), .A(n6573), .ZN(n6749) );
  INV_X1 U7321 ( .A(n6749), .ZN(n6638) );
  AND2_X1 U7322 ( .A1(n6593), .A2(n6575), .ZN(n6576) );
  NOR2_X1 U7323 ( .A1(n6577), .A2(n6576), .ZN(n6856) );
  INV_X1 U7324 ( .A(n6578), .ZN(n6595) );
  NAND2_X1 U7325 ( .A1(n7372), .A2(n6595), .ZN(n7416) );
  NOR2_X1 U7326 ( .A1(n7416), .A2(n6579), .ZN(n6581) );
  OAI21_X1 U7327 ( .B1(n6581), .B2(REIP_REG_23__SCAN_IN), .A(n6580), .ZN(n6583) );
  AOI22_X1 U7328 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n7439), .B1(n7425), 
        .B2(n6745), .ZN(n6582) );
  OAI211_X1 U7329 ( .C1(n7435), .C2(n4846), .A(n6583), .B(n6582), .ZN(n6584)
         );
  AOI21_X1 U7330 ( .B1(n6856), .B2(n7441), .A(n6584), .ZN(n6585) );
  OAI21_X1 U7331 ( .B1(n6638), .B2(n7422), .A(n6585), .ZN(U2804) );
  NAND2_X1 U7332 ( .A1(n6586), .A2(n6587), .ZN(n6588) );
  INV_X1 U7333 ( .A(REIP_REG_21__SCAN_IN), .ZN(n7434) );
  INV_X1 U7334 ( .A(REIP_REG_20__SCAN_IN), .ZN(n7417) );
  NOR4_X1 U7335 ( .A1(REIP_REG_22__SCAN_IN), .A2(n7434), .A3(n7417), .A4(n7416), .ZN(n6604) );
  NAND2_X1 U7336 ( .A1(n6590), .A2(n6591), .ZN(n6592) );
  AND2_X1 U7337 ( .A1(n6593), .A2(n6592), .ZN(n6870) );
  NAND2_X1 U7338 ( .A1(n6870), .A2(n7441), .ZN(n6602) );
  INV_X1 U7339 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6755) );
  OAI22_X1 U7340 ( .A1(n6755), .A2(n7429), .B1(n6641), .B2(n7435), .ZN(n6594)
         );
  AOI21_X1 U7341 ( .B1(n7425), .B2(n6757), .A(n6594), .ZN(n6601) );
  NAND2_X1 U7342 ( .A1(n6595), .A2(REIP_REG_20__SCAN_IN), .ZN(n7431) );
  INV_X1 U7343 ( .A(n7431), .ZN(n6596) );
  NAND2_X1 U7344 ( .A1(n7301), .A2(n6596), .ZN(n6597) );
  NAND2_X1 U7345 ( .A1(n6598), .A2(n6597), .ZN(n7433) );
  OR2_X1 U7346 ( .A1(n7324), .A2(REIP_REG_21__SCAN_IN), .ZN(n7432) );
  NAND2_X1 U7347 ( .A1(n7433), .A2(n7432), .ZN(n6599) );
  NAND2_X1 U7348 ( .A1(n6599), .A2(REIP_REG_22__SCAN_IN), .ZN(n6600) );
  NAND3_X1 U7349 ( .A1(n6602), .A2(n6601), .A3(n6600), .ZN(n6603) );
  AOI211_X1 U7350 ( .C1(n6758), .C2(n7442), .A(n6604), .B(n6603), .ZN(n6605)
         );
  INV_X1 U7351 ( .A(n6605), .ZN(U2805) );
  OAI22_X1 U7352 ( .A1(n6607), .A2(n7429), .B1(n7445), .B2(n6606), .ZN(n6611)
         );
  OAI22_X1 U7353 ( .A1(n7435), .A2(n6609), .B1(n6608), .B2(n6618), .ZN(n6610)
         );
  AOI211_X1 U7354 ( .C1(n7441), .C2(n6612), .A(n6611), .B(n6610), .ZN(n6616)
         );
  NOR2_X1 U7355 ( .A1(n6626), .A2(n6613), .ZN(n6614) );
  OAI21_X1 U7356 ( .B1(n7324), .B2(n7286), .A(n7301), .ZN(n7294) );
  OAI21_X1 U7357 ( .B1(REIP_REG_3__SCAN_IN), .B2(n6614), .A(n7294), .ZN(n6615)
         );
  OAI211_X1 U7358 ( .C1(n7290), .C2(n6617), .A(n6616), .B(n6615), .ZN(U2824)
         );
  NOR2_X1 U7359 ( .A1(n6618), .A2(n3648), .ZN(n6624) );
  AOI22_X1 U7360 ( .A1(n7439), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n7425), 
        .B2(n6619), .ZN(n6622) );
  NAND2_X1 U7361 ( .A1(n7305), .A2(n6620), .ZN(n6621) );
  OAI211_X1 U7362 ( .C1(n7324), .C2(REIP_REG_1__SCAN_IN), .A(n6622), .B(n6621), 
        .ZN(n6623) );
  AOI211_X1 U7363 ( .C1(n7441), .C2(n6625), .A(n6624), .B(n6623), .ZN(n6628)
         );
  AOI22_X1 U7364 ( .A1(EBX_REG_1__SCAN_IN), .A2(n7419), .B1(n6626), .B2(
        REIP_REG_1__SCAN_IN), .ZN(n6627) );
  NAND2_X1 U7365 ( .A1(n6628), .A2(n6627), .ZN(U2826) );
  INV_X1 U7366 ( .A(n6629), .ZN(n6655) );
  INV_X1 U7367 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6630) );
  OAI222_X1 U7368 ( .A1(n6648), .A2(n6655), .B1(n6630), .B2(n7126), .C1(n6798), 
        .C2(n6647), .ZN(U2830) );
  OAI222_X1 U7369 ( .A1(n6648), .A2(n6658), .B1(n6631), .B2(n7126), .C1(n6808), 
        .C2(n6647), .ZN(U2831) );
  AOI22_X1 U7370 ( .A1(n6821), .A2(n7124), .B1(EBX_REG_27__SCAN_IN), .B2(n6636), .ZN(n6632) );
  OAI21_X1 U7371 ( .B1(n6661), .B2(n6648), .A(n6632), .ZN(U2832) );
  INV_X1 U7372 ( .A(n6713), .ZN(n6664) );
  OAI222_X1 U7373 ( .A1(n6664), .A2(n6648), .B1(n6633), .B2(n7126), .C1(n6828), 
        .C2(n6647), .ZN(U2833) );
  OAI222_X1 U7374 ( .A1(n6723), .A2(n6648), .B1(n6634), .B2(n7126), .C1(n6840), 
        .C2(n6647), .ZN(U2834) );
  OAI222_X1 U7375 ( .A1(n6648), .A2(n6737), .B1(n7126), .B2(n6567), .C1(n6635), 
        .C2(n6647), .ZN(U2835) );
  AOI22_X1 U7376 ( .A1(n6856), .A2(n7124), .B1(EBX_REG_23__SCAN_IN), .B2(n6636), .ZN(n6637) );
  OAI21_X1 U7377 ( .B1(n6638), .B2(n6648), .A(n6637), .ZN(U2836) );
  NAND2_X1 U7378 ( .A1(n6758), .A2(n4916), .ZN(n6640) );
  NAND2_X1 U7379 ( .A1(n6870), .A2(n7124), .ZN(n6639) );
  OAI211_X1 U7380 ( .C1(n6641), .C2(n7126), .A(n6640), .B(n6639), .ZN(U2837)
         );
  INV_X1 U7381 ( .A(n6642), .ZN(n6645) );
  INV_X1 U7382 ( .A(n6643), .ZN(n6776) );
  AOI21_X1 U7383 ( .B1(n6645), .B2(n6776), .A(n6644), .ZN(n6772) );
  INV_X1 U7384 ( .A(n6772), .ZN(n7423) );
  AOI21_X1 U7385 ( .B1(n6646), .B2(n6896), .A(n6877), .ZN(n6887) );
  INV_X1 U7386 ( .A(n6887), .ZN(n7420) );
  OAI222_X1 U7387 ( .A1(n6648), .A2(n7423), .B1(n7126), .B2(n4836), .C1(n7420), 
        .C2(n6647), .ZN(U2839) );
  INV_X1 U7388 ( .A(n6649), .ZN(n6652) );
  AOI22_X1 U7389 ( .A1(n7550), .A2(DATAI_30_), .B1(n7553), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6651) );
  NAND2_X1 U7390 ( .A1(n7554), .A2(DATAI_14_), .ZN(n6650) );
  OAI211_X1 U7391 ( .C1(n6652), .C2(n6669), .A(n6651), .B(n6650), .ZN(U2861)
         );
  AOI22_X1 U7392 ( .A1(n7550), .A2(DATAI_29_), .B1(n7553), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6654) );
  NAND2_X1 U7393 ( .A1(n7554), .A2(DATAI_13_), .ZN(n6653) );
  OAI211_X1 U7394 ( .C1(n6655), .C2(n6669), .A(n6654), .B(n6653), .ZN(U2862)
         );
  AOI22_X1 U7395 ( .A1(n7550), .A2(DATAI_28_), .B1(n7553), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6657) );
  NAND2_X1 U7396 ( .A1(n7554), .A2(DATAI_12_), .ZN(n6656) );
  OAI211_X1 U7397 ( .C1(n6658), .C2(n6669), .A(n6657), .B(n6656), .ZN(U2863)
         );
  AOI22_X1 U7398 ( .A1(n7550), .A2(DATAI_27_), .B1(n7553), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6660) );
  NAND2_X1 U7399 ( .A1(n7554), .A2(DATAI_11_), .ZN(n6659) );
  OAI211_X1 U7400 ( .C1(n6661), .C2(n6669), .A(n6660), .B(n6659), .ZN(U2864)
         );
  AOI22_X1 U7401 ( .A1(n7550), .A2(DATAI_26_), .B1(n7553), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U7402 ( .A1(n7554), .A2(DATAI_10_), .ZN(n6662) );
  OAI211_X1 U7403 ( .C1(n6664), .C2(n6669), .A(n6663), .B(n6662), .ZN(U2865)
         );
  AOI22_X1 U7404 ( .A1(n7550), .A2(DATAI_25_), .B1(n7553), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U7405 ( .A1(n7554), .A2(DATAI_9_), .ZN(n6665) );
  OAI211_X1 U7406 ( .C1(n6723), .C2(n6669), .A(n6666), .B(n6665), .ZN(U2866)
         );
  AOI22_X1 U7407 ( .A1(n7550), .A2(DATAI_24_), .B1(n7553), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n6668) );
  NAND2_X1 U7408 ( .A1(n7554), .A2(DATAI_8_), .ZN(n6667) );
  OAI211_X1 U7409 ( .C1(n6737), .C2(n6669), .A(n6668), .B(n6667), .ZN(U2867)
         );
  INV_X1 U7410 ( .A(n7554), .ZN(n6679) );
  NAND2_X1 U7411 ( .A1(n6749), .A2(n7551), .ZN(n6671) );
  AOI22_X1 U7412 ( .A1(n7550), .A2(DATAI_23_), .B1(n7553), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6670) );
  OAI211_X1 U7413 ( .C1(n6679), .C2(n6672), .A(n6671), .B(n6670), .ZN(U2868)
         );
  NAND2_X1 U7414 ( .A1(n6758), .A2(n7551), .ZN(n6674) );
  AOI22_X1 U7415 ( .A1(n7550), .A2(DATAI_22_), .B1(n7553), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6673) );
  OAI211_X1 U7416 ( .C1(n6679), .C2(n6675), .A(n6674), .B(n6673), .ZN(U2869)
         );
  NAND2_X1 U7417 ( .A1(n6772), .A2(n7551), .ZN(n6677) );
  AOI22_X1 U7418 ( .A1(n7550), .A2(DATAI_20_), .B1(n7553), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6676) );
  OAI211_X1 U7419 ( .C1(n6679), .C2(n6678), .A(n6677), .B(n6676), .ZN(U2871)
         );
  AOI21_X1 U7420 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n6751), .A(n6680), 
        .ZN(n6684) );
  XOR2_X1 U7421 ( .A(n6684), .B(n6683), .Z(n6807) );
  NOR2_X1 U7422 ( .A1(n7211), .A2(n7066), .ZN(n6804) );
  AOI21_X1 U7423 ( .B1(n7158), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n6804), 
        .ZN(n6685) );
  OAI21_X1 U7424 ( .B1(n7169), .B2(n6686), .A(n6685), .ZN(n6687) );
  AOI21_X1 U7425 ( .B1(n6629), .B2(n7165), .A(n6687), .ZN(n6688) );
  OAI21_X1 U7426 ( .B1(n7447), .B2(n6807), .A(n6688), .ZN(U2957) );
  AOI22_X1 U7427 ( .A1(n6698), .A2(n6689), .B1(n6751), .B2(n6812), .ZN(n6691)
         );
  XNOR2_X1 U7428 ( .A(n6751), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6690)
         );
  XNOR2_X1 U7429 ( .A(n6691), .B(n6690), .ZN(n6819) );
  NOR2_X1 U7430 ( .A1(n7211), .A2(n7063), .ZN(n6814) );
  AOI21_X1 U7431 ( .B1(n7158), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n6814), 
        .ZN(n6692) );
  OAI21_X1 U7432 ( .B1(n7169), .B2(n6693), .A(n6692), .ZN(n6694) );
  AOI21_X1 U7433 ( .B1(n6695), .B2(n7165), .A(n6694), .ZN(n6696) );
  OAI21_X1 U7434 ( .B1(n7447), .B2(n6819), .A(n6696), .ZN(U2958) );
  XNOR2_X1 U7435 ( .A(n6701), .B(n6812), .ZN(n6827) );
  NOR2_X1 U7436 ( .A1(n7211), .A2(n7061), .ZN(n6820) );
  AOI21_X1 U7437 ( .B1(n7158), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n6820), 
        .ZN(n6702) );
  OAI21_X1 U7438 ( .B1(n7169), .B2(n6703), .A(n6702), .ZN(n6704) );
  AOI21_X1 U7439 ( .B1(n6705), .B2(n7165), .A(n6704), .ZN(n6706) );
  OAI21_X1 U7440 ( .B1(n7447), .B2(n6827), .A(n6706), .ZN(U2959) );
  XNOR2_X1 U7441 ( .A(n6751), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6707)
         );
  XNOR2_X1 U7442 ( .A(n6708), .B(n6707), .ZN(n6838) );
  INV_X1 U7443 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6709) );
  NOR2_X1 U7444 ( .A1(n7211), .A2(n6709), .ZN(n6829) );
  AOI21_X1 U7445 ( .B1(n7158), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n6829), 
        .ZN(n6710) );
  OAI21_X1 U7446 ( .B1(n7169), .B2(n6711), .A(n6710), .ZN(n6712) );
  AOI21_X1 U7447 ( .B1(n6713), .B2(n7165), .A(n6712), .ZN(n6714) );
  OAI21_X1 U7448 ( .B1(n6838), .B2(n7447), .A(n6714), .ZN(U2960) );
  NOR2_X1 U7449 ( .A1(n7211), .A2(n7058), .ZN(n6841) );
  AOI21_X1 U7450 ( .B1(n7158), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n6841), 
        .ZN(n6715) );
  OAI21_X1 U7451 ( .B1(n7169), .B2(n6716), .A(n6715), .ZN(n6717) );
  INV_X1 U7452 ( .A(n6717), .ZN(n6722) );
  NAND2_X1 U7453 ( .A1(n6720), .A2(n6719), .ZN(n6839) );
  NAND3_X1 U7454 ( .A1(n6718), .A2(n6839), .A3(n7166), .ZN(n6721) );
  OAI211_X1 U7455 ( .C1(n6723), .C2(n6797), .A(n6722), .B(n6721), .ZN(U2961)
         );
  XNOR2_X1 U7456 ( .A(n6751), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6778)
         );
  NAND2_X2 U7457 ( .A1(n6741), .A2(n6778), .ZN(n6777) );
  AOI21_X1 U7458 ( .B1(n6769), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n6777), 
        .ZN(n6725) );
  XNOR2_X1 U7459 ( .A(n6751), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6762)
         );
  NAND2_X1 U7460 ( .A1(n6763), .A2(n6762), .ZN(n6874) );
  INV_X1 U7461 ( .A(n6777), .ZN(n6730) );
  NAND4_X1 U7462 ( .A1(n6730), .A2(n6769), .A3(n6729), .A4(n6884), .ZN(n6742)
         );
  NAND2_X1 U7463 ( .A1(n6732), .A2(n6731), .ZN(n6733) );
  XNOR2_X1 U7464 ( .A(n6733), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6854)
         );
  NOR2_X1 U7465 ( .A1(n7211), .A2(n7055), .ZN(n6851) );
  INV_X1 U7466 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6734) );
  NOR2_X1 U7467 ( .A1(n6791), .A2(n6734), .ZN(n6735) );
  AOI211_X1 U7468 ( .C1(n7154), .C2(n6736), .A(n6851), .B(n6735), .ZN(n6740)
         );
  INV_X1 U7469 ( .A(n6737), .ZN(n6738) );
  NAND2_X1 U7470 ( .A1(n6738), .A2(n7165), .ZN(n6739) );
  OAI211_X1 U7471 ( .C1(n6854), .C2(n7447), .A(n6740), .B(n6739), .ZN(U2962)
         );
  NAND2_X1 U7472 ( .A1(n6751), .A2(n6857), .ZN(n6743) );
  OAI21_X1 U7473 ( .B1(n6779), .B2(n6743), .A(n6742), .ZN(n6744) );
  XNOR2_X1 U7474 ( .A(n6744), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6863)
         );
  INV_X1 U7475 ( .A(n6745), .ZN(n6747) );
  INV_X1 U7476 ( .A(REIP_REG_23__SCAN_IN), .ZN(n7053) );
  NOR2_X1 U7477 ( .A1(n7211), .A2(n7053), .ZN(n6855) );
  AOI21_X1 U7478 ( .B1(n7158), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n6855), 
        .ZN(n6746) );
  OAI21_X1 U7479 ( .B1(n7169), .B2(n6747), .A(n6746), .ZN(n6748) );
  AOI21_X1 U7480 ( .B1(n6749), .B2(n7165), .A(n6748), .ZN(n6750) );
  OAI21_X1 U7481 ( .B1(n6863), .B2(n7447), .A(n6750), .ZN(U2963) );
  XNOR2_X1 U7482 ( .A(n6751), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6752)
         );
  XNOR2_X1 U7483 ( .A(n6753), .B(n6752), .ZN(n6872) );
  INV_X1 U7484 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6754) );
  NOR2_X1 U7485 ( .A1(n7211), .A2(n6754), .ZN(n6869) );
  NOR2_X1 U7486 ( .A1(n6791), .A2(n6755), .ZN(n6756) );
  AOI211_X1 U7487 ( .C1(n7154), .C2(n6757), .A(n6869), .B(n6756), .ZN(n6760)
         );
  NAND2_X1 U7488 ( .A1(n6758), .A2(n7165), .ZN(n6759) );
  OAI211_X1 U7489 ( .C1(n6872), .C2(n7447), .A(n6760), .B(n6759), .ZN(U2964)
         );
  OAI21_X1 U7490 ( .B1(n6644), .B2(n6761), .A(n6586), .ZN(n7117) );
  OR2_X1 U7491 ( .A1(n6763), .A2(n6762), .ZN(n6875) );
  NAND3_X1 U7492 ( .A1(n6875), .A2(n6874), .A3(n7166), .ZN(n6766) );
  NOR2_X1 U7493 ( .A1(n7211), .A2(n7434), .ZN(n6879) );
  NOR2_X1 U7494 ( .A1(n7169), .A2(n7446), .ZN(n6764) );
  AOI211_X1 U7495 ( .C1(n7158), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n6879), 
        .B(n6764), .ZN(n6765) );
  OAI211_X1 U7496 ( .C1(n6797), .C2(n7117), .A(n6766), .B(n6765), .ZN(U2965)
         );
  NOR2_X1 U7497 ( .A1(n6769), .A2(n6767), .ZN(n6768) );
  MUX2_X1 U7498 ( .A(n6769), .B(n6768), .S(n6777), .Z(n6770) );
  XNOR2_X1 U7499 ( .A(n6770), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6893)
         );
  NOR2_X1 U7500 ( .A1(n7211), .A2(n7417), .ZN(n6886) );
  NOR2_X1 U7501 ( .A1(n6791), .A2(n7430), .ZN(n6771) );
  AOI211_X1 U7502 ( .C1(n7154), .C2(n7426), .A(n6886), .B(n6771), .ZN(n6774)
         );
  NAND2_X1 U7503 ( .A1(n6772), .A2(n7165), .ZN(n6773) );
  OAI211_X1 U7504 ( .C1(n6893), .C2(n7447), .A(n6774), .B(n6773), .ZN(U2966)
         );
  OAI21_X1 U7505 ( .B1(n3662), .B2(n5987), .A(n6776), .ZN(n7120) );
  OAI21_X1 U7506 ( .B1(n6779), .B2(n6778), .A(n6777), .ZN(n6894) );
  NAND2_X1 U7507 ( .A1(n6894), .A2(n7166), .ZN(n6784) );
  NAND2_X1 U7508 ( .A1(n7276), .A2(REIP_REG_19__SCAN_IN), .ZN(n6900) );
  OAI21_X1 U7509 ( .B1(n6791), .B2(n6780), .A(n6900), .ZN(n6781) );
  AOI21_X1 U7510 ( .B1(n6782), .B2(n7154), .A(n6781), .ZN(n6783) );
  OAI211_X1 U7511 ( .C1(n6797), .C2(n7120), .A(n6784), .B(n6783), .ZN(U2967)
         );
  NAND2_X1 U7512 ( .A1(n6751), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n7162) );
  INV_X1 U7513 ( .A(n6787), .ZN(n6788) );
  NOR2_X1 U7514 ( .A1(n6751), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n7159)
         );
  NAND2_X1 U7515 ( .A1(n6788), .A2(n7159), .ZN(n7163) );
  OAI21_X1 U7516 ( .B1(n6785), .B2(n7162), .A(n7163), .ZN(n6789) );
  XNOR2_X1 U7517 ( .A(n6789), .B(n6907), .ZN(n6916) );
  NAND2_X1 U7518 ( .A1(n6916), .A2(n7166), .ZN(n6795) );
  INV_X1 U7519 ( .A(REIP_REG_18__SCAN_IN), .ZN(n7048) );
  NOR2_X1 U7520 ( .A1(n7211), .A2(n7048), .ZN(n6908) );
  NOR2_X1 U7521 ( .A1(n6791), .A2(n6790), .ZN(n6792) );
  AOI211_X1 U7522 ( .C1(n7154), .C2(n6793), .A(n6908), .B(n6792), .ZN(n6794)
         );
  OAI211_X1 U7523 ( .C1(n6797), .C2(n6796), .A(n6795), .B(n6794), .ZN(U2968)
         );
  INV_X1 U7524 ( .A(n6798), .ZN(n6805) );
  INV_X1 U7525 ( .A(n6799), .ZN(n6800) );
  AOI21_X1 U7526 ( .B1(n6802), .B2(n6801), .A(n6800), .ZN(n6803) );
  AOI211_X1 U7527 ( .C1(n7269), .C2(n6805), .A(n6804), .B(n6803), .ZN(n6806)
         );
  OAI21_X1 U7528 ( .B1(n6807), .B2(n6892), .A(n6806), .ZN(U2989) );
  INV_X1 U7529 ( .A(n6808), .ZN(n6815) );
  INV_X1 U7530 ( .A(n6809), .ZN(n6823) );
  AOI211_X1 U7531 ( .C1(n6812), .C2(n6811), .A(n6810), .B(n6823), .ZN(n6813)
         );
  AOI211_X1 U7532 ( .C1(n7269), .C2(n6815), .A(n6814), .B(n6813), .ZN(n6818)
         );
  INV_X1 U7533 ( .A(n6816), .ZN(n6825) );
  NAND2_X1 U7534 ( .A1(n6825), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6817) );
  OAI211_X1 U7535 ( .C1(n6819), .C2(n6892), .A(n6818), .B(n6817), .ZN(U2990)
         );
  AOI21_X1 U7536 ( .B1(n6821), .B2(n7269), .A(n6820), .ZN(n6822) );
  OAI21_X1 U7537 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n6823), .A(n6822), 
        .ZN(n6824) );
  AOI21_X1 U7538 ( .B1(n6825), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n6824), 
        .ZN(n6826) );
  OAI21_X1 U7539 ( .B1(n6827), .B2(n6892), .A(n6826), .ZN(U2991) );
  INV_X1 U7540 ( .A(n6828), .ZN(n6830) );
  AOI21_X1 U7541 ( .B1(n6830), .B2(n7269), .A(n6829), .ZN(n6834) );
  INV_X1 U7542 ( .A(n6831), .ZN(n6843) );
  OAI211_X1 U7543 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A(n6843), .B(n6832), .ZN(n6833) );
  OAI211_X1 U7544 ( .C1(n6847), .C2(n6835), .A(n6834), .B(n6833), .ZN(n6836)
         );
  INV_X1 U7545 ( .A(n6836), .ZN(n6837) );
  OAI21_X1 U7546 ( .B1(n6838), .B2(n6892), .A(n6837), .ZN(U2992) );
  NAND3_X1 U7547 ( .A1(n6718), .A2(n6839), .A3(n7278), .ZN(n6845) );
  NOR2_X1 U7548 ( .A1(n6840), .A2(n7212), .ZN(n6842) );
  AOI211_X1 U7549 ( .C1(n6843), .C2(n6846), .A(n6842), .B(n6841), .ZN(n6844)
         );
  OAI211_X1 U7550 ( .C1(n6847), .C2(n6846), .A(n6845), .B(n6844), .ZN(U2993)
         );
  NAND3_X1 U7551 ( .A1(n6864), .A2(n6857), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6848) );
  AOI21_X1 U7552 ( .B1(n6849), .B2(n6848), .A(n6847), .ZN(n6850) );
  AOI211_X1 U7553 ( .C1(n7269), .C2(n6852), .A(n6851), .B(n6850), .ZN(n6853)
         );
  OAI21_X1 U7554 ( .B1(n6854), .B2(n6892), .A(n6853), .ZN(U2994) );
  AOI21_X1 U7555 ( .B1(n6856), .B2(n7269), .A(n6855), .ZN(n6859) );
  NAND3_X1 U7556 ( .A1(n6864), .A2(n6857), .A3(n6860), .ZN(n6858) );
  OAI211_X1 U7557 ( .C1(n6865), .C2(n6860), .A(n6859), .B(n6858), .ZN(n6861)
         );
  INV_X1 U7558 ( .A(n6861), .ZN(n6862) );
  OAI21_X1 U7559 ( .B1(n6863), .B2(n6892), .A(n6862), .ZN(U2995) );
  NAND3_X1 U7560 ( .A1(n6864), .A2(n6888), .A3(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6866) );
  AOI21_X1 U7561 ( .B1(n6867), .B2(n6866), .A(n6865), .ZN(n6868) );
  AOI211_X1 U7562 ( .C1(n7269), .C2(n6870), .A(n6869), .B(n6868), .ZN(n6871)
         );
  OAI21_X1 U7563 ( .B1(n6872), .B2(n6892), .A(n6871), .ZN(U2996) );
  INV_X1 U7564 ( .A(n6873), .ZN(n6883) );
  NAND3_X1 U7565 ( .A1(n6875), .A2(n6874), .A3(n7278), .ZN(n6882) );
  OAI21_X1 U7566 ( .B1(n6877), .B2(n6876), .A(n6590), .ZN(n7118) );
  NOR2_X1 U7567 ( .A1(n7118), .A2(n7212), .ZN(n6878) );
  AOI211_X1 U7568 ( .C1(n6880), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n6879), .B(n6878), .ZN(n6881) );
  OAI211_X1 U7569 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n6883), .A(n6882), .B(n6881), .ZN(U2997) );
  NOR2_X1 U7570 ( .A1(n6895), .A2(n6884), .ZN(n6885) );
  AOI211_X1 U7571 ( .C1(n7269), .C2(n6887), .A(n6886), .B(n6885), .ZN(n6891)
         );
  OR3_X1 U7572 ( .A1(n6906), .A2(n6889), .A3(n6888), .ZN(n6890) );
  OAI211_X1 U7573 ( .C1(n6893), .C2(n6892), .A(n6891), .B(n6890), .ZN(U2998)
         );
  NAND2_X1 U7574 ( .A1(n6894), .A2(n7278), .ZN(n6905) );
  INV_X1 U7575 ( .A(n6895), .ZN(n6903) );
  INV_X1 U7576 ( .A(n6896), .ZN(n6897) );
  AOI21_X1 U7577 ( .B1(n6899), .B2(n6898), .A(n6897), .ZN(n7412) );
  INV_X1 U7578 ( .A(n7412), .ZN(n6901) );
  OAI21_X1 U7579 ( .B1(n6901), .B2(n7212), .A(n6900), .ZN(n6902) );
  AOI21_X1 U7580 ( .B1(n6903), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n6902), 
        .ZN(n6904) );
  OAI211_X1 U7581 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6906), .A(n6905), .B(n6904), .ZN(U2999) );
  NAND2_X1 U7582 ( .A1(n6907), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6914) );
  AOI21_X1 U7583 ( .B1(n6909), .B2(n7269), .A(n6908), .ZN(n6913) );
  NOR2_X1 U7584 ( .A1(n6910), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6911)
         );
  OAI21_X1 U7585 ( .B1(n7277), .B2(n6911), .A(INSTADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n6912) );
  OAI211_X1 U7586 ( .C1(n7282), .C2(n6914), .A(n6913), .B(n6912), .ZN(n6915)
         );
  AOI21_X1 U7587 ( .B1(n6916), .B2(n7278), .A(n6915), .ZN(n6917) );
  INV_X1 U7588 ( .A(n6917), .ZN(U3000) );
  OAI22_X1 U7589 ( .A1(n6919), .A2(n7459), .B1(n6918), .B2(n7513), .ZN(n6921)
         );
  MUX2_X1 U7590 ( .A(n6921), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6920), 
        .Z(U3456) );
  NOR2_X1 U7591 ( .A1(n6923), .A2(n6922), .ZN(n6975) );
  INV_X1 U7592 ( .A(n6975), .ZN(n6925) );
  AOI211_X1 U7593 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6925), .A(n6924), .B(
        n7565), .ZN(n6930) );
  OAI21_X1 U7594 ( .B1(n6976), .B2(n6974), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6926) );
  OAI21_X1 U7595 ( .B1(n6928), .B2(n6927), .A(n6926), .ZN(n6929) );
  NAND2_X1 U7596 ( .A1(n6930), .A2(n6929), .ZN(n6971) );
  NAND2_X1 U7597 ( .A1(n6971), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n6940) );
  INV_X1 U7598 ( .A(n6931), .ZN(n7561) );
  NAND2_X1 U7599 ( .A1(n6932), .A2(n7561), .ZN(n6933) );
  OAI21_X1 U7600 ( .B1(n6935), .B2(n6934), .A(n6933), .ZN(n6972) );
  AOI22_X1 U7601 ( .A1(n6974), .A2(n7583), .B1(n6936), .B2(n6972), .ZN(n6939)
         );
  NAND2_X1 U7602 ( .A1(n7582), .A2(n6975), .ZN(n6938) );
  NAND2_X1 U7603 ( .A1(n6976), .A2(n7591), .ZN(n6937) );
  NAND4_X1 U7604 ( .A1(n6940), .A2(n6939), .A3(n6938), .A4(n6937), .ZN(U3020)
         );
  NAND2_X1 U7605 ( .A1(n6971), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n6945) );
  AOI22_X1 U7606 ( .A1(n6974), .A2(n7598), .B1(n6941), .B2(n6972), .ZN(n6944)
         );
  NAND2_X1 U7607 ( .A1(n7597), .A2(n6975), .ZN(n6943) );
  NAND2_X1 U7608 ( .A1(n6976), .A2(n7599), .ZN(n6942) );
  NAND4_X1 U7609 ( .A1(n6945), .A2(n6944), .A3(n6943), .A4(n6942), .ZN(U3021)
         );
  NAND2_X1 U7610 ( .A1(n6971), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n6950) );
  AOI22_X1 U7611 ( .A1(n6974), .A2(n7607), .B1(n6946), .B2(n6972), .ZN(n6949)
         );
  NAND2_X1 U7612 ( .A1(n7605), .A2(n6975), .ZN(n6948) );
  NAND2_X1 U7613 ( .A1(n6976), .A2(n7606), .ZN(n6947) );
  NAND4_X1 U7614 ( .A1(n6950), .A2(n6949), .A3(n6948), .A4(n6947), .ZN(U3022)
         );
  NAND2_X1 U7615 ( .A1(n6971), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6955) );
  AOI22_X1 U7616 ( .A1(n6974), .A2(n7614), .B1(n6951), .B2(n6972), .ZN(n6954)
         );
  NAND2_X1 U7617 ( .A1(n7613), .A2(n6975), .ZN(n6953) );
  NAND2_X1 U7618 ( .A1(n6976), .A2(n7615), .ZN(n6952) );
  NAND4_X1 U7619 ( .A1(n6955), .A2(n6954), .A3(n6953), .A4(n6952), .ZN(U3023)
         );
  NAND2_X1 U7620 ( .A1(n6971), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n6960) );
  AOI22_X1 U7621 ( .A1(n6974), .A2(n7623), .B1(n6956), .B2(n6972), .ZN(n6959)
         );
  NAND2_X1 U7622 ( .A1(n7621), .A2(n6975), .ZN(n6958) );
  NAND2_X1 U7623 ( .A1(n6976), .A2(n7622), .ZN(n6957) );
  NAND4_X1 U7624 ( .A1(n6960), .A2(n6959), .A3(n6958), .A4(n6957), .ZN(U3024)
         );
  NAND2_X1 U7625 ( .A1(n6971), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n6965) );
  AOI22_X1 U7626 ( .A1(n6974), .A2(n7631), .B1(n6961), .B2(n6972), .ZN(n6964)
         );
  NAND2_X1 U7627 ( .A1(n7629), .A2(n6975), .ZN(n6963) );
  NAND2_X1 U7628 ( .A1(n6976), .A2(n7630), .ZN(n6962) );
  NAND4_X1 U7629 ( .A1(n6965), .A2(n6964), .A3(n6963), .A4(n6962), .ZN(U3025)
         );
  NAND2_X1 U7630 ( .A1(n6971), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n6970) );
  AOI22_X1 U7631 ( .A1(n6974), .A2(n7639), .B1(n6966), .B2(n6972), .ZN(n6969)
         );
  NAND2_X1 U7632 ( .A1(n7637), .A2(n6975), .ZN(n6968) );
  NAND2_X1 U7633 ( .A1(n6976), .A2(n7638), .ZN(n6967) );
  NAND4_X1 U7634 ( .A1(n6970), .A2(n6969), .A3(n6968), .A4(n6967), .ZN(U3026)
         );
  NAND2_X1 U7635 ( .A1(n6971), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n6980) );
  AOI22_X1 U7636 ( .A1(n6974), .A2(n7651), .B1(n6973), .B2(n6972), .ZN(n6979)
         );
  NAND2_X1 U7637 ( .A1(n7650), .A2(n6975), .ZN(n6978) );
  NAND2_X1 U7638 ( .A1(n6976), .A2(n7654), .ZN(n6977) );
  NAND4_X1 U7639 ( .A1(n6980), .A2(n6979), .A3(n6978), .A4(n6977), .ZN(U3027)
         );
  INV_X1 U7640 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6982) );
  OR2_X1 U7641 ( .A1(n7524), .A2(STATE_REG_0__SCAN_IN), .ZN(n7540) );
  INV_X1 U7642 ( .A(n3628), .ZN(n6993) );
  INV_X1 U7643 ( .A(BS16_N), .ZN(n6981) );
  NAND2_X1 U7644 ( .A1(n7533), .A2(n7535), .ZN(n7173) );
  AOI21_X1 U7645 ( .B1(n6981), .B2(n7173), .A(n6993), .ZN(n7519) );
  AOI21_X1 U7646 ( .B1(n6982), .B2(n6993), .A(n7519), .ZN(U3451) );
  INV_X1 U7647 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n7079) );
  NOR2_X1 U7648 ( .A1(n3628), .A2(n7079), .ZN(U3180) );
  AND2_X1 U7649 ( .A1(n6993), .A2(DATAWIDTH_REG_3__SCAN_IN), .ZN(U3179) );
  INV_X1 U7650 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n7078) );
  NOR2_X1 U7651 ( .A1(n3628), .A2(n7078), .ZN(U3178) );
  NOR2_X1 U7652 ( .A1(n3628), .A2(n6983), .ZN(U3177) );
  NOR2_X1 U7653 ( .A1(n3628), .A2(n6984), .ZN(U3176) );
  INV_X1 U7654 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n7080) );
  NOR2_X1 U7655 ( .A1(n3628), .A2(n7080), .ZN(U3175) );
  AND2_X1 U7656 ( .A1(n6993), .A2(DATAWIDTH_REG_8__SCAN_IN), .ZN(U3174) );
  NOR2_X1 U7657 ( .A1(n3628), .A2(n6985), .ZN(U3173) );
  NOR2_X1 U7658 ( .A1(n3628), .A2(n6986), .ZN(U3172) );
  AND2_X1 U7659 ( .A1(n6993), .A2(DATAWIDTH_REG_11__SCAN_IN), .ZN(U3171) );
  INV_X1 U7660 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n7077) );
  NOR2_X1 U7661 ( .A1(n3628), .A2(n7077), .ZN(U3170) );
  INV_X1 U7662 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n7075) );
  NOR2_X1 U7663 ( .A1(n3628), .A2(n7075), .ZN(U3169) );
  NOR2_X1 U7664 ( .A1(n3628), .A2(n6987), .ZN(U3168) );
  INV_X1 U7665 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n7074) );
  NOR2_X1 U7666 ( .A1(n3628), .A2(n7074), .ZN(U3167) );
  INV_X1 U7667 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n7076) );
  NOR2_X1 U7668 ( .A1(n3628), .A2(n7076), .ZN(U3166) );
  AND2_X1 U7669 ( .A1(n6993), .A2(DATAWIDTH_REG_17__SCAN_IN), .ZN(U3165) );
  AND2_X1 U7670 ( .A1(n6993), .A2(DATAWIDTH_REG_18__SCAN_IN), .ZN(U3164) );
  INV_X1 U7671 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n7073) );
  NOR2_X1 U7672 ( .A1(n3628), .A2(n7073), .ZN(U3163) );
  INV_X1 U7673 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6988) );
  NOR2_X1 U7674 ( .A1(n3628), .A2(n6988), .ZN(U3162) );
  NOR2_X1 U7675 ( .A1(n3628), .A2(n6989), .ZN(U3161) );
  NOR2_X1 U7676 ( .A1(n3628), .A2(n6990), .ZN(U3160) );
  INV_X1 U7677 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6991) );
  NOR2_X1 U7678 ( .A1(n3628), .A2(n6991), .ZN(U3159) );
  AND2_X1 U7679 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6993), .ZN(U3158) );
  AND2_X1 U7680 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6993), .ZN(U3157) );
  AND2_X1 U7681 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6993), .ZN(U3156) );
  AND2_X1 U7682 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6993), .ZN(U3155) );
  AND2_X1 U7683 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6993), .ZN(U3154) );
  AND2_X1 U7684 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6993), .ZN(U3153) );
  AND2_X1 U7685 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6993), .ZN(U3152) );
  AND2_X1 U7686 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6993), .ZN(U3151) );
  AND2_X1 U7687 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6992), .ZN(U3019)
         );
  AND2_X1 U7688 ( .A1(n7003), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  OAI21_X1 U7689 ( .B1(n7174), .B2(n6994), .A(n6993), .ZN(U2789) );
  AOI22_X1 U7690 ( .A1(n7192), .A2(LWORD_REG_0__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6995) );
  OAI21_X1 U7691 ( .B1(n6996), .B2(n7024), .A(n6995), .ZN(U2923) );
  AOI22_X1 U7692 ( .A1(n7192), .A2(LWORD_REG_1__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6997) );
  OAI21_X1 U7693 ( .B1(n6998), .B2(n7024), .A(n6997), .ZN(U2922) );
  AOI22_X1 U7694 ( .A1(n7192), .A2(LWORD_REG_2__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6999) );
  OAI21_X1 U7695 ( .B1(n7000), .B2(n7024), .A(n6999), .ZN(U2921) );
  AOI22_X1 U7696 ( .A1(n7192), .A2(LWORD_REG_3__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n7001) );
  OAI21_X1 U7697 ( .B1(n7002), .B2(n7024), .A(n7001), .ZN(U2920) );
  AOI22_X1 U7698 ( .A1(n7192), .A2(LWORD_REG_4__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n7004) );
  OAI21_X1 U7699 ( .B1(n7005), .B2(n7024), .A(n7004), .ZN(U2919) );
  AOI22_X1 U7700 ( .A1(n7192), .A2(LWORD_REG_5__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n7006) );
  OAI21_X1 U7701 ( .B1(n4246), .B2(n7024), .A(n7006), .ZN(U2918) );
  AOI22_X1 U7702 ( .A1(n7192), .A2(LWORD_REG_6__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n7007) );
  OAI21_X1 U7703 ( .B1(n4234), .B2(n7024), .A(n7007), .ZN(U2917) );
  AOI22_X1 U7704 ( .A1(n7192), .A2(LWORD_REG_7__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n7008) );
  OAI21_X1 U7705 ( .B1(n4250), .B2(n7024), .A(n7008), .ZN(U2916) );
  AOI22_X1 U7706 ( .A1(n7192), .A2(LWORD_REG_8__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n7009) );
  OAI21_X1 U7707 ( .B1(n7010), .B2(n7024), .A(n7009), .ZN(U2915) );
  AOI22_X1 U7708 ( .A1(n7192), .A2(LWORD_REG_9__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n7011) );
  OAI21_X1 U7709 ( .B1(n7012), .B2(n7024), .A(n7011), .ZN(U2914) );
  AOI22_X1 U7710 ( .A1(n7192), .A2(LWORD_REG_10__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n7013) );
  OAI21_X1 U7711 ( .B1(n7014), .B2(n7024), .A(n7013), .ZN(U2913) );
  AOI22_X1 U7712 ( .A1(n7192), .A2(LWORD_REG_11__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n7015) );
  OAI21_X1 U7713 ( .B1(n7016), .B2(n7024), .A(n7015), .ZN(U2912) );
  AOI22_X1 U7714 ( .A1(n7192), .A2(LWORD_REG_12__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n7017) );
  OAI21_X1 U7715 ( .B1(n7018), .B2(n7024), .A(n7017), .ZN(U2911) );
  AOI22_X1 U7716 ( .A1(n7492), .A2(LWORD_REG_13__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n7019) );
  OAI21_X1 U7717 ( .B1(n7020), .B2(n7024), .A(n7019), .ZN(U2910) );
  AOI22_X1 U7718 ( .A1(n7492), .A2(LWORD_REG_14__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n7021) );
  OAI21_X1 U7719 ( .B1(n7022), .B2(n7024), .A(n7021), .ZN(U2909) );
  AOI22_X1 U7720 ( .A1(n7492), .A2(LWORD_REG_15__SCAN_IN), .B1(n7003), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n7023) );
  OAI21_X1 U7721 ( .B1(n4924), .B2(n7024), .A(n7023), .ZN(U2908) );
  INV_X1 U7722 ( .A(n7540), .ZN(n7543) );
  NAND2_X1 U7723 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7174), .ZN(n7064) );
  CLKBUF_X1 U7724 ( .A(n7064), .Z(n7067) );
  OAI222_X1 U7725 ( .A1(n7071), .A2(n7026), .B1(n7025), .B2(n7543), .C1(n5013), 
        .C2(n7067), .ZN(U3184) );
  INV_X1 U7726 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n7027) );
  OAI222_X1 U7727 ( .A1(n7071), .A2(n5074), .B1(n7027), .B2(n7174), .C1(n7026), 
        .C2(n7067), .ZN(U3185) );
  INV_X1 U7728 ( .A(REIP_REG_4__SCAN_IN), .ZN(n7285) );
  INV_X1 U7729 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n7028) );
  OAI222_X1 U7730 ( .A1(n7071), .A2(n7285), .B1(n7028), .B2(n7543), .C1(n5074), 
        .C2(n7064), .ZN(U3186) );
  OAI222_X1 U7731 ( .A1(n7071), .A2(n7302), .B1(n7029), .B2(n7174), .C1(n7285), 
        .C2(n7067), .ZN(U3187) );
  INV_X1 U7732 ( .A(REIP_REG_6__SCAN_IN), .ZN(n7311) );
  OAI222_X1 U7733 ( .A1(n7071), .A2(n7311), .B1(n7030), .B2(n7543), .C1(n7302), 
        .C2(n7067), .ZN(U3188) );
  INV_X1 U7734 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n7031) );
  OAI222_X1 U7735 ( .A1(n7071), .A2(n5363), .B1(n7031), .B2(n7174), .C1(n7311), 
        .C2(n7064), .ZN(U3189) );
  INV_X1 U7736 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n7032) );
  OAI222_X1 U7737 ( .A1(n7071), .A2(n7033), .B1(n7032), .B2(n7543), .C1(n5363), 
        .C2(n7067), .ZN(U3190) );
  OAI222_X1 U7738 ( .A1(n7071), .A2(n7035), .B1(n7034), .B2(n7543), .C1(n7033), 
        .C2(n7064), .ZN(U3191) );
  OAI222_X1 U7739 ( .A1(n7071), .A2(n5831), .B1(n7036), .B2(n7543), .C1(n7035), 
        .C2(n7064), .ZN(U3192) );
  INV_X1 U7740 ( .A(REIP_REG_11__SCAN_IN), .ZN(n7354) );
  INV_X1 U7741 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n7037) );
  OAI222_X1 U7742 ( .A1(n7071), .A2(n7354), .B1(n7037), .B2(n7543), .C1(n5831), 
        .C2(n7064), .ZN(U3193) );
  INV_X1 U7743 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n7038) );
  OAI222_X1 U7744 ( .A1(n7071), .A2(n7366), .B1(n7038), .B2(n7543), .C1(n7354), 
        .C2(n7064), .ZN(U3194) );
  INV_X1 U7745 ( .A(REIP_REG_13__SCAN_IN), .ZN(n7040) );
  OAI222_X1 U7746 ( .A1(n7064), .A2(n7366), .B1(n7039), .B2(n7543), .C1(n7040), 
        .C2(n7071), .ZN(U3195) );
  OAI222_X1 U7747 ( .A1(n7071), .A2(n5970), .B1(n7041), .B2(n7543), .C1(n7040), 
        .C2(n7067), .ZN(U3196) );
  INV_X1 U7748 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n7042) );
  OAI222_X1 U7749 ( .A1(n7071), .A2(n7044), .B1(n7042), .B2(n7543), .C1(n5970), 
        .C2(n7067), .ZN(U3197) );
  OAI222_X1 U7750 ( .A1(n7064), .A2(n7044), .B1(n7043), .B2(n7543), .C1(n6017), 
        .C2(n7071), .ZN(U3198) );
  INV_X1 U7751 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n7045) );
  OAI222_X1 U7752 ( .A1(n7071), .A2(n7392), .B1(n7045), .B2(n7543), .C1(n6017), 
        .C2(n7067), .ZN(U3199) );
  INV_X1 U7753 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n7046) );
  OAI222_X1 U7754 ( .A1(n7071), .A2(n7048), .B1(n7046), .B2(n7543), .C1(n7392), 
        .C2(n7067), .ZN(U3200) );
  INV_X1 U7755 ( .A(REIP_REG_19__SCAN_IN), .ZN(n7405) );
  OAI222_X1 U7756 ( .A1(n7067), .A2(n7048), .B1(n7047), .B2(n7543), .C1(n7405), 
        .C2(n7071), .ZN(U3201) );
  OAI222_X1 U7757 ( .A1(n7071), .A2(n7417), .B1(n7049), .B2(n7543), .C1(n7405), 
        .C2(n7067), .ZN(U3202) );
  OAI222_X1 U7758 ( .A1(n7071), .A2(n7434), .B1(n7050), .B2(n7543), .C1(n7417), 
        .C2(n7067), .ZN(U3203) );
  INV_X1 U7759 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n7051) );
  OAI222_X1 U7760 ( .A1(n7071), .A2(n6754), .B1(n7051), .B2(n7543), .C1(n7434), 
        .C2(n7067), .ZN(U3204) );
  INV_X1 U7761 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n7052) );
  OAI222_X1 U7762 ( .A1(n7071), .A2(n7053), .B1(n7052), .B2(n7543), .C1(n6754), 
        .C2(n7067), .ZN(U3205) );
  OAI222_X1 U7763 ( .A1(n7071), .A2(n7055), .B1(n7054), .B2(n7543), .C1(n7053), 
        .C2(n7067), .ZN(U3206) );
  INV_X1 U7764 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n7056) );
  OAI222_X1 U7765 ( .A1(n7071), .A2(n7058), .B1(n7056), .B2(n7174), .C1(n7055), 
        .C2(n7067), .ZN(U3207) );
  OAI222_X1 U7766 ( .A1(n7067), .A2(n7058), .B1(n7057), .B2(n7174), .C1(n6709), 
        .C2(n7071), .ZN(U3208) );
  INV_X1 U7767 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n7059) );
  OAI222_X1 U7768 ( .A1(n7064), .A2(n6709), .B1(n7059), .B2(n7174), .C1(n7061), 
        .C2(n7071), .ZN(U3209) );
  OAI222_X1 U7769 ( .A1(n7064), .A2(n7061), .B1(n7060), .B2(n7174), .C1(n7063), 
        .C2(n7071), .ZN(U3210) );
  INV_X1 U7770 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n7062) );
  OAI222_X1 U7771 ( .A1(n7064), .A2(n7063), .B1(n7062), .B2(n7174), .C1(n7066), 
        .C2(n7071), .ZN(U3211) );
  OAI222_X1 U7772 ( .A1(n7067), .A2(n7066), .B1(n7065), .B2(n7174), .C1(n7068), 
        .C2(n7071), .ZN(U3212) );
  OAI222_X1 U7773 ( .A1(n7071), .A2(n7070), .B1(n7069), .B2(n7174), .C1(n7068), 
        .C2(n7067), .ZN(U3213) );
  INV_X1 U7774 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n7093) );
  INV_X1 U7775 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n7072) );
  AOI22_X1 U7776 ( .A1(n7543), .A2(n7093), .B1(n7072), .B2(n7540), .ZN(U3445)
         );
  NOR4_X1 U7777 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(n7090) );
  AOI211_X1 U7778 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_6__SCAN_IN), .B(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n7089) );
  NAND4_X1 U7779 ( .A1(n7076), .A2(n7075), .A3(n7074), .A4(n7073), .ZN(n7087)
         );
  NAND4_X1 U7780 ( .A1(n7080), .A2(n7079), .A3(n7078), .A4(n7077), .ZN(n7086)
         );
  NOR4_X1 U7781 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n7084) );
  NOR4_X1 U7782 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_31__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n7083) );
  NOR4_X1 U7783 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(
        DATAWIDTH_REG_8__SCAN_IN), .ZN(n7082) );
  NOR4_X1 U7784 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n7081) );
  NAND4_X1 U7785 ( .A1(n7084), .A2(n7083), .A3(n7082), .A4(n7081), .ZN(n7085)
         );
  NOR3_X1 U7786 ( .A1(n7087), .A2(n7086), .A3(n7085), .ZN(n7088) );
  NAND3_X1 U7787 ( .A1(n7090), .A2(n7089), .A3(n7088), .ZN(n7103) );
  INV_X1 U7788 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7522) );
  NAND2_X1 U7789 ( .A1(n5013), .A2(n7522), .ZN(n7092) );
  NOR3_X1 U7790 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(REIP_REG_0__SCAN_IN), .ZN(n7099) );
  NOR2_X1 U7791 ( .A1(n7103), .A2(n7099), .ZN(n7091) );
  AOI22_X1 U7792 ( .A1(n7093), .A2(n7103), .B1(n7092), .B2(n7091), .ZN(U2795)
         );
  INV_X1 U7793 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n7096) );
  INV_X1 U7794 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n7094) );
  AOI22_X1 U7795 ( .A1(n7174), .A2(n7096), .B1(n7094), .B2(n7540), .ZN(U3446)
         );
  INV_X1 U7796 ( .A(n7103), .ZN(n7106) );
  AOI211_X1 U7797 ( .C1(REIP_REG_0__SCAN_IN), .C2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(REIP_REG_1__SCAN_IN), .B(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7095) );
  AOI21_X1 U7798 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n7095), .ZN(n7097) );
  AOI22_X1 U7799 ( .A1(n7106), .A2(n7097), .B1(n7096), .B2(n7103), .ZN(U3468)
         );
  INV_X1 U7800 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n7101) );
  INV_X1 U7801 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n7098) );
  AOI22_X1 U7802 ( .A1(n7543), .A2(n7101), .B1(n7098), .B2(n7540), .ZN(U3447)
         );
  OAI21_X1 U7803 ( .B1(REIP_REG_1__SCAN_IN), .B2(n7099), .A(n7106), .ZN(n7100)
         );
  OAI21_X1 U7804 ( .B1(n7106), .B2(n7101), .A(n7100), .ZN(U2794) );
  INV_X1 U7805 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n7104) );
  AOI22_X1 U7806 ( .A1(n7174), .A2(n7104), .B1(n7102), .B2(n7540), .ZN(U3448)
         );
  NOR2_X1 U7807 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n7105) );
  AOI22_X1 U7808 ( .A1(n7106), .A2(n7105), .B1(n7104), .B2(n7103), .ZN(U3469)
         );
  AOI22_X1 U7809 ( .A1(n7351), .A2(n4916), .B1(n7124), .B2(n7345), .ZN(n7107)
         );
  OAI21_X1 U7810 ( .B1(n7126), .B2(n7108), .A(n7107), .ZN(U2848) );
  OR2_X1 U7811 ( .A1(n5876), .A2(n7109), .ZN(n7110) );
  AND2_X1 U7812 ( .A1(n7110), .A2(n5984), .ZN(n7544) );
  AND2_X1 U7813 ( .A1(n7112), .A2(n7111), .ZN(n7113) );
  NOR2_X1 U7814 ( .A1(n7114), .A2(n7113), .ZN(n7398) );
  AOI22_X1 U7815 ( .A1(n7544), .A2(n4916), .B1(n7124), .B2(n7398), .ZN(n7115)
         );
  OAI21_X1 U7816 ( .B1(n7126), .B2(n7116), .A(n7115), .ZN(U2842) );
  INV_X1 U7817 ( .A(n7117), .ZN(n7552) );
  INV_X1 U7818 ( .A(n7118), .ZN(n7440) );
  AOI22_X1 U7819 ( .A1(n7552), .A2(n4916), .B1(n7124), .B2(n7440), .ZN(n7119)
         );
  OAI21_X1 U7820 ( .B1(n7126), .B2(n7436), .A(n7119), .ZN(U2838) );
  INV_X1 U7821 ( .A(n7120), .ZN(n7547) );
  AOI22_X1 U7822 ( .A1(n7547), .A2(n4916), .B1(n7124), .B2(n7412), .ZN(n7121)
         );
  OAI21_X1 U7823 ( .B1(n7126), .B2(n7409), .A(n7121), .ZN(U2840) );
  XNOR2_X1 U7824 ( .A(n7123), .B(n7122), .ZN(n7284) );
  AOI22_X1 U7825 ( .A1(n7139), .A2(n4916), .B1(n7124), .B2(n7284), .ZN(n7125)
         );
  OAI21_X1 U7826 ( .B1(n7126), .B2(n7297), .A(n7125), .ZN(U2855) );
  AOI22_X1 U7827 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n7158), .B1(n7276), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n7133) );
  INV_X1 U7828 ( .A(n7127), .ZN(n7131) );
  XNOR2_X1 U7829 ( .A(n7129), .B(n7234), .ZN(n7130) );
  XNOR2_X1 U7830 ( .A(n7128), .B(n7130), .ZN(n7230) );
  AOI22_X1 U7831 ( .A1(n7131), .A2(n7165), .B1(n7230), .B2(n7166), .ZN(n7132)
         );
  OAI211_X1 U7832 ( .C1(n7169), .C2(n7134), .A(n7133), .B(n7132), .ZN(U2984)
         );
  AOI22_X1 U7833 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n7158), .B1(n7276), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n7141) );
  OAI21_X1 U7834 ( .B1(n7137), .B2(n3640), .A(n3642), .ZN(n7138) );
  INV_X1 U7835 ( .A(n7138), .ZN(n7204) );
  AOI22_X1 U7836 ( .A1(n7165), .A2(n7139), .B1(n7204), .B2(n7166), .ZN(n7140)
         );
  OAI211_X1 U7837 ( .C1(n7169), .C2(n7289), .A(n7141), .B(n7140), .ZN(U2982)
         );
  AOI22_X1 U7838 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n7158), .B1(n7276), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n7147) );
  OAI21_X1 U7839 ( .B1(n7142), .B2(n7144), .A(n7143), .ZN(n7145) );
  INV_X1 U7840 ( .A(n7145), .ZN(n7222) );
  AOI22_X1 U7841 ( .A1(n7222), .A2(n7166), .B1(n7165), .B2(n7306), .ZN(n7146)
         );
  OAI211_X1 U7842 ( .C1(n7169), .C2(n7309), .A(n7147), .B(n7146), .ZN(U2981)
         );
  AOI22_X1 U7843 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n7158), .B1(n7276), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n7153) );
  CLKBUF_X1 U7844 ( .A(n7148), .Z(n7149) );
  XNOR2_X1 U7845 ( .A(n7150), .B(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n7151)
         );
  XNOR2_X1 U7846 ( .A(n7149), .B(n7151), .ZN(n7216) );
  AOI22_X1 U7847 ( .A1(n7216), .A2(n7166), .B1(n7165), .B2(n7318), .ZN(n7152)
         );
  OAI211_X1 U7848 ( .C1(n7169), .C2(n7321), .A(n7153), .B(n7152), .ZN(U2980)
         );
  AOI22_X1 U7849 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n7158), .B1(n7276), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n7156) );
  AOI22_X1 U7850 ( .A1(n7351), .A2(n7165), .B1(n7154), .B2(n7350), .ZN(n7155)
         );
  OAI211_X1 U7851 ( .C1(n7447), .C2(n7157), .A(n7156), .B(n7155), .ZN(U2975)
         );
  AOI22_X1 U7852 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n7158), .B1(n7276), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n7168) );
  INV_X1 U7853 ( .A(n7159), .ZN(n7160) );
  NAND2_X1 U7854 ( .A1(n7160), .A2(n7162), .ZN(n7161) );
  MUX2_X1 U7855 ( .A(n7162), .B(n7161), .S(n6787), .Z(n7164) );
  NAND2_X1 U7856 ( .A1(n7164), .A2(n7163), .ZN(n7279) );
  AOI22_X1 U7857 ( .A1(n7279), .A2(n7166), .B1(n7165), .B2(n7544), .ZN(n7167)
         );
  OAI211_X1 U7858 ( .C1(n7169), .C2(n7401), .A(n7168), .B(n7167), .ZN(U2969)
         );
  OAI21_X1 U7859 ( .B1(n7170), .B2(n7517), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n7171) );
  OAI21_X1 U7860 ( .B1(n7178), .B2(n3848), .A(n7171), .ZN(U2790) );
  OAI222_X1 U7861 ( .A1(n7174), .A2(n7173), .B1(n7174), .B2(n7172), .C1(
        CODEFETCH_REG_SCAN_IN), .C2(n7540), .ZN(U2791) );
  INV_X1 U7862 ( .A(n7175), .ZN(n7176) );
  NAND2_X1 U7863 ( .A1(n7190), .A2(n7176), .ZN(n7177) );
  OAI211_X1 U7864 ( .C1(n7190), .C2(n7179), .A(n7178), .B(n7177), .ZN(U3474)
         );
  OAI22_X1 U7865 ( .A1(n7540), .A2(n7179), .B1(W_R_N_REG_SCAN_IN), .B2(n7543), 
        .ZN(n7180) );
  INV_X1 U7866 ( .A(n7180), .ZN(U3470) );
  NAND2_X1 U7867 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .ZN(n7538) );
  INV_X1 U7868 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7526) );
  NOR2_X1 U7869 ( .A1(n7535), .A2(n7526), .ZN(n7528) );
  INV_X1 U7870 ( .A(HOLD), .ZN(n7531) );
  NOR2_X1 U7871 ( .A1(n7524), .A2(n7531), .ZN(n7181) );
  OAI22_X1 U7872 ( .A1(n7528), .A2(n7181), .B1(n7533), .B2(n7531), .ZN(n7182)
         );
  NAND3_X1 U7873 ( .A1(n7183), .A2(n7538), .A3(n7182), .ZN(U3182) );
  NOR2_X1 U7874 ( .A1(READY_N), .A2(n3848), .ZN(n7500) );
  OAI211_X1 U7875 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n7500), .A(n7507), .B(
        n7514), .ZN(n7184) );
  NAND2_X1 U7876 ( .A1(n7185), .A2(n7184), .ZN(U3150) );
  INV_X1 U7877 ( .A(n7186), .ZN(n7187) );
  AOI211_X1 U7878 ( .C1(n3915), .C2(n7520), .A(n7188), .B(n7187), .ZN(n7189)
         );
  OAI21_X1 U7879 ( .B1(n7189), .B2(n3848), .A(n7514), .ZN(n7194) );
  AOI211_X1 U7880 ( .C1(n7192), .C2(n7502), .A(n7191), .B(n7190), .ZN(n7193)
         );
  MUX2_X1 U7881 ( .A(n7194), .B(REQUESTPENDING_REG_SCAN_IN), .S(n7193), .Z(
        U3472) );
  AOI21_X1 U7882 ( .B1(n7269), .B2(n7196), .A(n7195), .ZN(n7202) );
  NOR4_X1 U7883 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n4801), .A3(n7198), 
        .A4(n7197), .ZN(n7199) );
  AOI21_X1 U7884 ( .B1(n7200), .B2(n7278), .A(n7199), .ZN(n7201) );
  OAI211_X1 U7885 ( .C1(n7203), .C2(n4096), .A(n7202), .B(n7201), .ZN(U3005)
         );
  OAI21_X1 U7886 ( .B1(INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n7219), .ZN(n7207) );
  AOI22_X1 U7887 ( .A1(n7269), .A2(n7284), .B1(n7276), .B2(REIP_REG_4__SCAN_IN), .ZN(n7206) );
  AOI22_X1 U7888 ( .A1(n7208), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .B1(n7278), 
        .B2(n7204), .ZN(n7205) );
  OAI211_X1 U7889 ( .C1(n7218), .C2(n7207), .A(n7206), .B(n7205), .ZN(U3014)
         );
  AND2_X1 U7890 ( .A1(n7219), .A2(n7260), .ZN(n7209) );
  AOI211_X1 U7891 ( .C1(n7213), .C2(n7210), .A(n7209), .B(n7208), .ZN(n7226)
         );
  OAI22_X1 U7892 ( .A1(n7212), .A2(n7314), .B1(n7311), .B2(n7211), .ZN(n7215)
         );
  NOR4_X1 U7893 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n7213), .A3(n7219), 
        .A4(n7218), .ZN(n7214) );
  AOI211_X1 U7894 ( .C1(n7216), .C2(n7278), .A(n7215), .B(n7214), .ZN(n7217)
         );
  OAI21_X1 U7895 ( .B1(n7226), .B2(n4771), .A(n7217), .ZN(U3012) );
  NOR2_X1 U7896 ( .A1(n7219), .A2(n7218), .ZN(n7220) );
  NOR2_X1 U7897 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n7220), .ZN(n7225)
         );
  INV_X1 U7898 ( .A(n7299), .ZN(n7221) );
  AOI22_X1 U7899 ( .A1(n7222), .A2(n7278), .B1(n7269), .B2(n7221), .ZN(n7224)
         );
  NAND2_X1 U7900 ( .A1(n7276), .A2(REIP_REG_5__SCAN_IN), .ZN(n7223) );
  OAI211_X1 U7901 ( .C1(n7226), .C2(n7225), .A(n7224), .B(n7223), .ZN(U3013)
         );
  AOI22_X1 U7902 ( .A1(n7269), .A2(n7227), .B1(n7276), .B2(REIP_REG_2__SCAN_IN), .ZN(n7239) );
  NAND2_X1 U7903 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n7229) );
  OAI21_X1 U7904 ( .B1(n7229), .B2(n7233), .A(n7228), .ZN(n7231) );
  AOI22_X1 U7905 ( .A1(n7231), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n7278), 
        .B2(n7230), .ZN(n7238) );
  OR2_X1 U7906 ( .A1(n7233), .A2(n7232), .ZN(n7237) );
  NAND3_X1 U7907 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n7235), .A3(n7234), 
        .ZN(n7236) );
  NAND4_X1 U7908 ( .A1(n7239), .A2(n7238), .A3(n7237), .A4(n7236), .ZN(U3016)
         );
  NAND2_X1 U7909 ( .A1(n7245), .A2(n7240), .ZN(n7258) );
  INV_X1 U7910 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n7241) );
  AOI22_X1 U7911 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n7241), .B1(
        INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n4790), .ZN(n7250) );
  AOI21_X1 U7912 ( .B1(n7269), .B2(n7243), .A(n7242), .ZN(n7249) );
  OAI21_X1 U7913 ( .B1(n7246), .B2(n7245), .A(n7244), .ZN(n7254) );
  AOI22_X1 U7914 ( .A1(n7247), .A2(n7278), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n7254), .ZN(n7248) );
  OAI211_X1 U7915 ( .C1(n7258), .C2(n7250), .A(n7249), .B(n7248), .ZN(U3008)
         );
  INV_X1 U7916 ( .A(n7251), .ZN(n7336) );
  INV_X1 U7917 ( .A(n7252), .ZN(n7253) );
  AOI21_X1 U7918 ( .B1(n7269), .B2(n7336), .A(n7253), .ZN(n7257) );
  AOI22_X1 U7919 ( .A1(n7255), .A2(n7278), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n7254), .ZN(n7256) );
  OAI211_X1 U7920 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n7258), .A(n7257), 
        .B(n7256), .ZN(U3009) );
  AOI21_X1 U7921 ( .B1(n7261), .B2(n7260), .A(n7259), .ZN(n7275) );
  INV_X1 U7922 ( .A(n7262), .ZN(n7263) );
  AOI21_X1 U7923 ( .B1(n7269), .B2(n7264), .A(n7263), .ZN(n7267) );
  AOI22_X1 U7924 ( .A1(n7265), .A2(n7278), .B1(n7272), .B2(n7268), .ZN(n7266)
         );
  OAI211_X1 U7925 ( .C1(n7275), .C2(n7268), .A(n7267), .B(n7266), .ZN(U3003)
         );
  AOI222_X1 U7926 ( .A1(n7270), .A2(n7278), .B1(n7269), .B2(n7384), .C1(
        REIP_REG_16__SCAN_IN), .C2(n7276), .ZN(n7274) );
  NAND2_X1 U7927 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n7271) );
  OAI211_X1 U7928 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A(n7272), .B(n7271), .ZN(n7273) );
  OAI211_X1 U7929 ( .C1(n7275), .C2(n4818), .A(n7274), .B(n7273), .ZN(U3002)
         );
  AOI22_X1 U7930 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n7277), .B1(n7276), .B2(REIP_REG_17__SCAN_IN), .ZN(n7281) );
  AOI22_X1 U7931 ( .A1(n7279), .A2(n7278), .B1(n7269), .B2(n7398), .ZN(n7280)
         );
  OAI211_X1 U7932 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n7282), .A(n7281), .B(n7280), .ZN(U3001) );
  AOI22_X1 U7933 ( .A1(n7441), .A2(n7284), .B1(n7283), .B2(n7461), .ZN(n7296)
         );
  INV_X1 U7934 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n7288) );
  NAND3_X1 U7935 ( .A1(n7372), .A2(n7286), .A3(n7285), .ZN(n7287) );
  OAI211_X1 U7936 ( .C1(n7429), .C2(n7288), .A(n7315), .B(n7287), .ZN(n7293)
         );
  OAI22_X1 U7937 ( .A1(n7291), .A2(n7290), .B1(n7289), .B2(n7445), .ZN(n7292)
         );
  AOI211_X1 U7938 ( .C1(REIP_REG_4__SCAN_IN), .C2(n7294), .A(n7293), .B(n7292), 
        .ZN(n7295) );
  OAI211_X1 U7939 ( .C1(n7297), .C2(n7435), .A(n7296), .B(n7295), .ZN(U2823)
         );
  OAI22_X1 U7940 ( .A1(n7421), .A2(n7299), .B1(n7429), .B2(n7298), .ZN(n7300)
         );
  AOI211_X1 U7941 ( .C1(n7419), .C2(EBX_REG_5__SCAN_IN), .A(n7411), .B(n7300), 
        .ZN(n7308) );
  OAI21_X1 U7942 ( .B1(n7324), .B2(n7310), .A(n7301), .ZN(n7329) );
  OAI21_X1 U7943 ( .B1(n7324), .B2(n7303), .A(n7302), .ZN(n7304) );
  AOI22_X1 U7944 ( .A1(n7306), .A2(n7305), .B1(n7329), .B2(n7304), .ZN(n7307)
         );
  OAI211_X1 U7945 ( .C1(n7309), .C2(n7445), .A(n7308), .B(n7307), .ZN(U2822)
         );
  AND3_X1 U7946 ( .A1(n7372), .A2(n7311), .A3(n7310), .ZN(n7330) );
  NOR2_X1 U7947 ( .A1(n7312), .A2(n7435), .ZN(n7313) );
  AOI211_X1 U7948 ( .C1(REIP_REG_6__SCAN_IN), .C2(n7329), .A(n7330), .B(n7313), 
        .ZN(n7320) );
  NOR2_X1 U7949 ( .A1(n7421), .A2(n7314), .ZN(n7317) );
  OAI21_X1 U7950 ( .B1(n7429), .B2(n4233), .A(n7315), .ZN(n7316) );
  AOI211_X1 U7951 ( .C1(n7318), .C2(n7442), .A(n7317), .B(n7316), .ZN(n7319)
         );
  OAI211_X1 U7952 ( .C1(n7321), .C2(n7445), .A(n7320), .B(n7319), .ZN(U2821)
         );
  AOI22_X1 U7953 ( .A1(n7441), .A2(n7322), .B1(n7419), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n7334) );
  NOR3_X1 U7954 ( .A1(n7324), .A2(REIP_REG_7__SCAN_IN), .A3(n7323), .ZN(n7325)
         );
  AOI211_X1 U7955 ( .C1(n7439), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n7411), 
        .B(n7325), .ZN(n7333) );
  INV_X1 U7956 ( .A(n7326), .ZN(n7327) );
  AOI22_X1 U7957 ( .A1(n7328), .A2(n7442), .B1(n7327), .B2(n7425), .ZN(n7332)
         );
  OAI21_X1 U7958 ( .B1(n7330), .B2(n7329), .A(REIP_REG_7__SCAN_IN), .ZN(n7331)
         );
  NAND4_X1 U7959 ( .A1(n7334), .A2(n7333), .A3(n7332), .A4(n7331), .ZN(U2820)
         );
  AOI21_X1 U7960 ( .B1(n7336), .B2(n7441), .A(n7335), .ZN(n7344) );
  AOI22_X1 U7961 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n7439), .B1(
        EBX_REG_9__SCAN_IN), .B2(n7419), .ZN(n7343) );
  AOI21_X1 U7962 ( .B1(REIP_REG_9__SCAN_IN), .B2(n7337), .A(n7411), .ZN(n7342)
         );
  INV_X1 U7963 ( .A(n7338), .ZN(n7340) );
  AOI22_X1 U7964 ( .A1(n7340), .A2(n7442), .B1(n7425), .B2(n7339), .ZN(n7341)
         );
  NAND4_X1 U7965 ( .A1(n7344), .A2(n7343), .A3(n7342), .A4(n7341), .ZN(U2818)
         );
  NAND3_X1 U7966 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        n7354), .ZN(n7347) );
  AOI22_X1 U7967 ( .A1(n7441), .A2(n7345), .B1(n7419), .B2(EBX_REG_11__SCAN_IN), .ZN(n7346) );
  OAI21_X1 U7968 ( .B1(n7348), .B2(n7347), .A(n7346), .ZN(n7349) );
  AOI211_X1 U7969 ( .C1(n7439), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n7411), 
        .B(n7349), .ZN(n7353) );
  AOI22_X1 U7970 ( .A1(n7351), .A2(n7442), .B1(n7425), .B2(n7350), .ZN(n7352)
         );
  OAI211_X1 U7971 ( .C1(n7367), .C2(n7354), .A(n7353), .B(n7352), .ZN(U2816)
         );
  INV_X1 U7972 ( .A(n7355), .ZN(n7358) );
  NAND2_X1 U7973 ( .A1(n7419), .A2(EBX_REG_12__SCAN_IN), .ZN(n7357) );
  AOI21_X1 U7974 ( .B1(n7439), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n7411), 
        .ZN(n7356) );
  OAI211_X1 U7975 ( .C1(n7358), .C2(n7421), .A(n7357), .B(n7356), .ZN(n7359)
         );
  INV_X1 U7976 ( .A(n7359), .ZN(n7360) );
  OAI211_X1 U7977 ( .C1(n7362), .C2(n7422), .A(n7361), .B(n7360), .ZN(n7363)
         );
  AOI21_X1 U7978 ( .B1(n7364), .B2(n7425), .A(n7363), .ZN(n7365) );
  OAI21_X1 U7979 ( .B1(n7367), .B2(n7366), .A(n7365), .ZN(U2815) );
  INV_X1 U7980 ( .A(n7368), .ZN(n7369) );
  OAI22_X1 U7981 ( .A1(n7382), .A2(n5970), .B1(n7421), .B2(n7369), .ZN(n7370)
         );
  AOI211_X1 U7982 ( .C1(n7439), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n7411), 
        .B(n7370), .ZN(n7379) );
  NAND2_X1 U7983 ( .A1(n7372), .A2(n7371), .ZN(n7373) );
  OAI22_X1 U7984 ( .A1(n7375), .A2(n7422), .B1(n7374), .B2(n7373), .ZN(n7376)
         );
  AOI21_X1 U7985 ( .B1(n7377), .B2(n7425), .A(n7376), .ZN(n7378) );
  OAI211_X1 U7986 ( .C1(n7380), .C2(n7435), .A(n7379), .B(n7378), .ZN(U2813)
         );
  OAI21_X1 U7987 ( .B1(REIP_REG_16__SCAN_IN), .B2(REIP_REG_15__SCAN_IN), .A(
        n7394), .ZN(n7381) );
  OAI22_X1 U7988 ( .A1(n7382), .A2(n6017), .B1(n7393), .B2(n7381), .ZN(n7383)
         );
  AOI211_X1 U7989 ( .C1(n7439), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n7411), 
        .B(n7383), .ZN(n7390) );
  INV_X1 U7990 ( .A(n7384), .ZN(n7385) );
  OAI22_X1 U7991 ( .A1(n7386), .A2(n7422), .B1(n7421), .B2(n7385), .ZN(n7387)
         );
  AOI21_X1 U7992 ( .B1(n7388), .B2(n7425), .A(n7387), .ZN(n7389) );
  OAI211_X1 U7993 ( .C1(n7391), .C2(n7435), .A(n7390), .B(n7389), .ZN(U2811)
         );
  OAI21_X1 U7994 ( .B1(n7394), .B2(n7393), .A(n7392), .ZN(n7397) );
  AOI22_X1 U7995 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n7439), .B1(
        EBX_REG_17__SCAN_IN), .B2(n7419), .ZN(n7395) );
  INV_X1 U7996 ( .A(n7395), .ZN(n7396) );
  AOI211_X1 U7997 ( .C1(n7402), .C2(n7397), .A(n7411), .B(n7396), .ZN(n7400)
         );
  AOI22_X1 U7998 ( .A1(n7544), .A2(n7442), .B1(n7441), .B2(n7398), .ZN(n7399)
         );
  OAI211_X1 U7999 ( .C1(n7401), .C2(n7445), .A(n7400), .B(n7399), .ZN(U2810)
         );
  OAI21_X1 U8000 ( .B1(n7403), .B2(n7402), .A(REIP_REG_19__SCAN_IN), .ZN(n7408) );
  INV_X1 U8001 ( .A(n7404), .ZN(n7406) );
  NAND3_X1 U8002 ( .A1(n7406), .A2(REIP_REG_18__SCAN_IN), .A3(n7405), .ZN(
        n7407) );
  OAI211_X1 U8003 ( .C1(n7435), .C2(n7409), .A(n7408), .B(n7407), .ZN(n7410)
         );
  AOI211_X1 U8004 ( .C1(n7439), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n7411), 
        .B(n7410), .ZN(n7414) );
  AOI22_X1 U8005 ( .A1(n7547), .A2(n7442), .B1(n7441), .B2(n7412), .ZN(n7413)
         );
  OAI211_X1 U8006 ( .C1(n7415), .C2(n7445), .A(n7414), .B(n7413), .ZN(U2808)
         );
  AOI21_X1 U8007 ( .B1(n7417), .B2(n7416), .A(n7433), .ZN(n7418) );
  AOI21_X1 U8008 ( .B1(n7419), .B2(EBX_REG_20__SCAN_IN), .A(n7418), .ZN(n7428)
         );
  OAI22_X1 U8009 ( .A1(n7423), .A2(n7422), .B1(n7421), .B2(n7420), .ZN(n7424)
         );
  AOI21_X1 U8010 ( .B1(n7426), .B2(n7425), .A(n7424), .ZN(n7427) );
  OAI211_X1 U8011 ( .C1(n7430), .C2(n7429), .A(n7428), .B(n7427), .ZN(U2807)
         );
  NOR2_X1 U8012 ( .A1(n7432), .A2(n7431), .ZN(n7438) );
  OAI22_X1 U8013 ( .A1(n7436), .A2(n7435), .B1(n7434), .B2(n7433), .ZN(n7437)
         );
  AOI211_X1 U8014 ( .C1(n7439), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n7438), 
        .B(n7437), .ZN(n7444) );
  AOI22_X1 U8015 ( .A1(n7552), .A2(n7442), .B1(n7441), .B2(n7440), .ZN(n7443)
         );
  OAI211_X1 U8016 ( .C1(n7446), .C2(n7445), .A(n7444), .B(n7443), .ZN(U2806)
         );
  OAI21_X1 U8017 ( .B1(n7449), .B2(n7448), .A(n7447), .ZN(U2793) );
  NAND2_X1 U8018 ( .A1(n7450), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n7468) );
  AOI22_X1 U8019 ( .A1(n7454), .A2(n7453), .B1(n7452), .B2(n7451), .ZN(n7469)
         );
  OAI22_X1 U8020 ( .A1(n7469), .A2(n7459), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n7455), .ZN(n7457) );
  OAI22_X1 U8021 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n7466), .B1(n7457), .B2(n7456), .ZN(n7458) );
  OAI21_X1 U8022 ( .B1(n7468), .B2(n7459), .A(n7458), .ZN(U3461) );
  INV_X1 U8023 ( .A(n7460), .ZN(n7462) );
  NAND4_X1 U8024 ( .A1(n7463), .A2(n7462), .A3(n7501), .A4(n7461), .ZN(n7464)
         );
  OAI21_X1 U8025 ( .B1(n7466), .B2(n7465), .A(n7464), .ZN(U3455) );
  INV_X1 U8026 ( .A(n7467), .ZN(n7477) );
  AND3_X1 U8027 ( .A1(n7469), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n7468), 
        .ZN(n7470) );
  INV_X1 U8028 ( .A(n7470), .ZN(n7475) );
  OAI22_X1 U8029 ( .A1(n7472), .A2(n7471), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n7470), .ZN(n7473) );
  OAI21_X1 U8030 ( .B1(n7475), .B2(n7474), .A(n7473), .ZN(n7476) );
  AOI222_X1 U8031 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7477), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n7476), .C1(n7477), .C2(n7476), 
        .ZN(n7478) );
  AOI222_X1 U8032 ( .A1(n7480), .A2(n7479), .B1(n7480), .B2(n7478), .C1(n7479), 
        .C2(n7478), .ZN(n7481) );
  OR2_X1 U8033 ( .A1(n7481), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n7491)
         );
  NOR2_X1 U8034 ( .A1(MORE_REG_SCAN_IN), .A2(FLUSH_REG_SCAN_IN), .ZN(n7486) );
  INV_X1 U8035 ( .A(n7482), .ZN(n7485) );
  INV_X1 U8036 ( .A(n7483), .ZN(n7484) );
  OAI211_X1 U8037 ( .C1(n7487), .C2(n7486), .A(n7485), .B(n7484), .ZN(n7488)
         );
  NOR2_X1 U8038 ( .A1(n7489), .A2(n7488), .ZN(n7490) );
  NAND2_X1 U8039 ( .A1(n7518), .A2(n7499), .ZN(n7494) );
  NAND2_X1 U8040 ( .A1(READY_N), .A2(n7492), .ZN(n7493) );
  NAND2_X1 U8041 ( .A1(n7494), .A2(n7493), .ZN(n7498) );
  OR2_X1 U8042 ( .A1(n7496), .A2(n7495), .ZN(n7497) );
  AOI21_X1 U8043 ( .B1(n7501), .B2(n7500), .A(n7499), .ZN(n7505) );
  OAI21_X1 U8044 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7502), .A(n7512), .ZN(
        n7510) );
  OAI211_X1 U8045 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n7510), .ZN(n7503) );
  OAI211_X1 U8046 ( .C1(n7506), .C2(n7505), .A(n7504), .B(n7503), .ZN(U3149)
         );
  OAI221_X1 U8047 ( .B1(n7508), .B2(STATE2_REG_0__SCAN_IN), .C1(n7508), .C2(
        n7512), .A(n7507), .ZN(U3453) );
  AOI221_X1 U8048 ( .B1(n7511), .B2(STATE2_REG_0__SCAN_IN), .C1(n7510), .C2(
        STATE2_REG_0__SCAN_IN), .A(n7509), .ZN(n7516) );
  OAI211_X1 U8049 ( .C1(n7514), .C2(n7513), .A(n3848), .B(n7512), .ZN(n7515)
         );
  OAI211_X1 U8050 ( .C1(n7518), .C2(n7517), .A(n7516), .B(n7515), .ZN(U3148)
         );
  INV_X1 U8051 ( .A(n7519), .ZN(n7521) );
  OAI21_X1 U8052 ( .B1(n3628), .B2(n7520), .A(n7521), .ZN(U2792) );
  OAI21_X1 U8053 ( .B1(n3628), .B2(n7522), .A(n7521), .ZN(U3452) );
  OAI221_X1 U8054 ( .B1(n7533), .B2(NA_N), .C1(n7533), .C2(n7524), .A(n7535), 
        .ZN(n7534) );
  AOI21_X1 U8055 ( .B1(n7524), .B2(n7533), .A(n7531), .ZN(n7525) );
  OAI21_X1 U8056 ( .B1(n7526), .B2(n7525), .A(n7540), .ZN(n7527) );
  OAI211_X1 U8057 ( .C1(STATE_REG_2__SCAN_IN), .C2(n7538), .A(n7534), .B(n7527), .ZN(U3181) );
  INV_X1 U8058 ( .A(NA_N), .ZN(n7530) );
  AOI21_X1 U8059 ( .B1(n7528), .B2(n7530), .A(STATE_REG_2__SCAN_IN), .ZN(n7539) );
  AOI21_X1 U8060 ( .B1(READY_N), .B2(n7530), .A(n7529), .ZN(n7532) );
  AOI211_X1 U8061 ( .C1(REQUESTPENDING_REG_SCAN_IN), .C2(n7533), .A(n7532), 
        .B(n7531), .ZN(n7536) );
  OAI21_X1 U8062 ( .B1(n7536), .B2(n7535), .A(n7534), .ZN(n7537) );
  OAI21_X1 U8063 ( .B1(n7539), .B2(n7538), .A(n7537), .ZN(U3183) );
  AOI22_X1 U8064 ( .A1(n7543), .A2(n7542), .B1(n7541), .B2(n7540), .ZN(U3473)
         );
  AOI22_X1 U8065 ( .A1(n7544), .A2(n7551), .B1(n7550), .B2(DATAI_17_), .ZN(
        n7546) );
  AOI22_X1 U8066 ( .A1(n7554), .A2(DATAI_1_), .B1(n7553), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n7545) );
  NAND2_X1 U8067 ( .A1(n7546), .A2(n7545), .ZN(U2874) );
  AOI22_X1 U8068 ( .A1(n7547), .A2(n7551), .B1(n7550), .B2(DATAI_19_), .ZN(
        n7549) );
  AOI22_X1 U8069 ( .A1(n7554), .A2(DATAI_3_), .B1(n7553), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n7548) );
  NAND2_X1 U8070 ( .A1(n7549), .A2(n7548), .ZN(U2872) );
  AOI22_X1 U8071 ( .A1(n7552), .A2(n7551), .B1(n7550), .B2(DATAI_21_), .ZN(
        n7556) );
  AOI22_X1 U8072 ( .A1(n7554), .A2(DATAI_5_), .B1(n7553), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n7555) );
  NAND2_X1 U8073 ( .A1(n7556), .A2(n7555), .ZN(U2870) );
  NOR2_X1 U8074 ( .A1(n7644), .A2(n7580), .ZN(n7559) );
  NAND2_X1 U8075 ( .A1(n7581), .A2(n7557), .ZN(n7563) );
  INV_X1 U8076 ( .A(n7579), .ZN(n7558) );
  AOI21_X1 U8077 ( .B1(n7559), .B2(n7563), .A(n7558), .ZN(n7569) );
  INV_X1 U8078 ( .A(n7569), .ZN(n7562) );
  AOI22_X1 U8079 ( .A1(n7562), .A2(n7570), .B1(n7561), .B2(n7560), .ZN(n7648)
         );
  NOR2_X1 U8080 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7564), .ZN(n7643)
         );
  AOI22_X1 U8081 ( .A1(n7653), .A2(n7583), .B1(n7582), .B2(n7643), .ZN(n7572)
         );
  INV_X1 U8082 ( .A(n7643), .ZN(n7567) );
  AOI211_X1 U8083 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n7567), .A(n7566), .B(
        n7565), .ZN(n7568) );
  OAI21_X1 U8084 ( .B1(n7570), .B2(n7569), .A(n7568), .ZN(n7645) );
  AOI22_X1 U8085 ( .A1(n7645), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n7591), 
        .B2(n7644), .ZN(n7571) );
  OAI211_X1 U8086 ( .C1(n7648), .C2(n7594), .A(n7572), .B(n7571), .ZN(U3100)
         );
  NOR2_X1 U8087 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n7575), .ZN(n7589)
         );
  NAND2_X1 U8088 ( .A1(n7574), .A2(n7573), .ZN(n7578) );
  NOR3_X2 U8089 ( .A1(n7576), .A2(n7575), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n7649) );
  INV_X1 U8090 ( .A(n7649), .ZN(n7577) );
  NAND2_X1 U8091 ( .A1(n7578), .A2(n7577), .ZN(n7584) );
  OAI21_X1 U8092 ( .B1(n7581), .B2(n7580), .A(n7579), .ZN(n7586) );
  AOI22_X1 U8093 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7589), .B1(n7584), .B2(
        n7586), .ZN(n7659) );
  AOI22_X1 U8094 ( .A1(n7652), .A2(n7583), .B1(n7582), .B2(n7649), .ZN(n7593)
         );
  INV_X1 U8095 ( .A(n7584), .ZN(n7585) );
  NAND2_X1 U8096 ( .A1(n7586), .A2(n7585), .ZN(n7588) );
  OAI211_X1 U8097 ( .C1(n7590), .C2(n7589), .A(n7588), .B(n7587), .ZN(n7655)
         );
  AOI22_X1 U8098 ( .A1(n7655), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n7591), 
        .B2(n7653), .ZN(n7592) );
  OAI211_X1 U8099 ( .C1(n7659), .C2(n7594), .A(n7593), .B(n7592), .ZN(U3092)
         );
  AOI22_X1 U8100 ( .A1(n7653), .A2(n7598), .B1(n7597), .B2(n7643), .ZN(n7596)
         );
  AOI22_X1 U8101 ( .A1(n7645), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n7599), 
        .B2(n7644), .ZN(n7595) );
  OAI211_X1 U8102 ( .C1(n7648), .C2(n7602), .A(n7596), .B(n7595), .ZN(U3101)
         );
  AOI22_X1 U8103 ( .A1(n7652), .A2(n7598), .B1(n7597), .B2(n7649), .ZN(n7601)
         );
  AOI22_X1 U8104 ( .A1(n7655), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n7599), 
        .B2(n7653), .ZN(n7600) );
  OAI211_X1 U8105 ( .C1(n7659), .C2(n7602), .A(n7601), .B(n7600), .ZN(U3093)
         );
  AOI22_X1 U8106 ( .A1(n7653), .A2(n7607), .B1(n7605), .B2(n7643), .ZN(n7604)
         );
  AOI22_X1 U8107 ( .A1(n7645), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n7606), 
        .B2(n7644), .ZN(n7603) );
  OAI211_X1 U8108 ( .C1(n7648), .C2(n7610), .A(n7604), .B(n7603), .ZN(U3102)
         );
  AOI22_X1 U8109 ( .A1(n7653), .A2(n7606), .B1(n7605), .B2(n7649), .ZN(n7609)
         );
  AOI22_X1 U8110 ( .A1(n7655), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n7607), 
        .B2(n7652), .ZN(n7608) );
  OAI211_X1 U8111 ( .C1(n7659), .C2(n7610), .A(n7609), .B(n7608), .ZN(U3094)
         );
  AOI22_X1 U8112 ( .A1(n7653), .A2(n7614), .B1(n7613), .B2(n7643), .ZN(n7612)
         );
  AOI22_X1 U8113 ( .A1(n7645), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n7615), 
        .B2(n7644), .ZN(n7611) );
  OAI211_X1 U8114 ( .C1(n7648), .C2(n7618), .A(n7612), .B(n7611), .ZN(U3103)
         );
  AOI22_X1 U8115 ( .A1(n7652), .A2(n7614), .B1(n7613), .B2(n7649), .ZN(n7617)
         );
  AOI22_X1 U8116 ( .A1(n7655), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n7615), 
        .B2(n7653), .ZN(n7616) );
  OAI211_X1 U8117 ( .C1(n7659), .C2(n7618), .A(n7617), .B(n7616), .ZN(U3095)
         );
  AOI22_X1 U8118 ( .A1(n7653), .A2(n7623), .B1(n7621), .B2(n7643), .ZN(n7620)
         );
  AOI22_X1 U8119 ( .A1(n7645), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n7622), 
        .B2(n7644), .ZN(n7619) );
  OAI211_X1 U8120 ( .C1(n7648), .C2(n7626), .A(n7620), .B(n7619), .ZN(U3104)
         );
  AOI22_X1 U8121 ( .A1(n7653), .A2(n7622), .B1(n7621), .B2(n7649), .ZN(n7625)
         );
  AOI22_X1 U8122 ( .A1(n7655), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n7623), 
        .B2(n7652), .ZN(n7624) );
  OAI211_X1 U8123 ( .C1(n7659), .C2(n7626), .A(n7625), .B(n7624), .ZN(U3096)
         );
  AOI22_X1 U8124 ( .A1(n7653), .A2(n7631), .B1(n7629), .B2(n7643), .ZN(n7628)
         );
  AOI22_X1 U8125 ( .A1(n7645), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n7630), 
        .B2(n7644), .ZN(n7627) );
  OAI211_X1 U8126 ( .C1(n7648), .C2(n7634), .A(n7628), .B(n7627), .ZN(U3105)
         );
  AOI22_X1 U8127 ( .A1(n7653), .A2(n7630), .B1(n7629), .B2(n7649), .ZN(n7633)
         );
  AOI22_X1 U8128 ( .A1(n7655), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n7631), 
        .B2(n7652), .ZN(n7632) );
  OAI211_X1 U8129 ( .C1(n7659), .C2(n7634), .A(n7633), .B(n7632), .ZN(U3097)
         );
  AOI22_X1 U8130 ( .A1(n7653), .A2(n7639), .B1(n7637), .B2(n7643), .ZN(n7636)
         );
  AOI22_X1 U8131 ( .A1(n7645), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n7638), 
        .B2(n7644), .ZN(n7635) );
  OAI211_X1 U8132 ( .C1(n7648), .C2(n7642), .A(n7636), .B(n7635), .ZN(U3106)
         );
  AOI22_X1 U8133 ( .A1(n7653), .A2(n7638), .B1(n7637), .B2(n7649), .ZN(n7641)
         );
  AOI22_X1 U8134 ( .A1(n7655), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n7639), 
        .B2(n7652), .ZN(n7640) );
  OAI211_X1 U8135 ( .C1(n7659), .C2(n7642), .A(n7641), .B(n7640), .ZN(U3098)
         );
  AOI22_X1 U8136 ( .A1(n7653), .A2(n7651), .B1(n7650), .B2(n7643), .ZN(n7647)
         );
  AOI22_X1 U8137 ( .A1(n7645), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n7654), 
        .B2(n7644), .ZN(n7646) );
  OAI211_X1 U8138 ( .C1(n7648), .C2(n7658), .A(n7647), .B(n7646), .ZN(U3107)
         );
  AOI22_X1 U8139 ( .A1(n7652), .A2(n7651), .B1(n7650), .B2(n7649), .ZN(n7657)
         );
  AOI22_X1 U8140 ( .A1(n7655), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n7654), 
        .B2(n7653), .ZN(n7656) );
  OAI211_X1 U8141 ( .C1(n7659), .C2(n7658), .A(n7657), .B(n7656), .ZN(U3099)
         );
  AND2_X1 U3672 ( .A1(n4978), .A2(n3676), .ZN(n3772) );
  CLKBUF_X2 U3670 ( .A(n3772), .Z(n3936) );
  AND2_X1 U3673 ( .A1(n5128), .A2(n5163), .ZN(n3980) );
  AND2_X2 U3686 ( .A1(n3669), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4974)
         );
  OR2_X1 U3690 ( .A1(n6590), .A2(n6591), .ZN(n6593) );
  CLKBUF_X1 U3986 ( .A(n7192), .Z(n7492) );
  CLKBUF_X1 U5406 ( .A(n4110), .Z(n6708) );
endmodule

