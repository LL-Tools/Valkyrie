

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740;

  INV_X2 U7174 ( .A(n15691), .ZN(n9345) );
  XNOR2_X1 U7175 ( .A(n9474), .B(n13958), .ZN(n9531) );
  OAI21_X1 U7176 ( .B1(n8831), .B2(n12957), .A(n8830), .ZN(n7455) );
  INV_X1 U7177 ( .A(n11914), .ZN(n7628) );
  NAND2_X1 U7178 ( .A1(n10136), .A2(n10135), .ZN(n11818) );
  INV_X1 U7179 ( .A(n10527), .ZN(n6434) );
  CLKBUF_X2 U7180 ( .A(n8137), .Z(n12880) );
  NAND4_X2 U7181 ( .A1(n8988), .A2(n8987), .A3(n8986), .A4(n8985), .ZN(n13978)
         );
  INV_X1 U7182 ( .A(n10616), .ZN(n10506) );
  INV_X1 U7183 ( .A(n11545), .ZN(n15523) );
  OR2_X1 U7184 ( .A1(n11156), .A2(n11151), .ZN(n11150) );
  INV_X1 U7185 ( .A(n8137), .ZN(n8179) );
  NAND4_X1 U7186 ( .A1(n9641), .A2(n9640), .A3(n9639), .A4(n9638), .ZN(n14819)
         );
  XNOR2_X1 U7188 ( .A(n10041), .B(P1_IR_REG_26__SCAN_IN), .ZN(n10050) );
  AND2_X1 U7189 ( .A1(n10777), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10775) );
  INV_X1 U7190 ( .A(n10527), .ZN(n6435) );
  NOR2_X1 U7191 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n9575) );
  OAI21_X1 U7192 ( .B1(n12373), .B2(n10397), .A(n10396), .ZN(n12403) );
  INV_X1 U7193 ( .A(n10252), .ZN(n10287) );
  CLKBUF_X2 U7194 ( .A(n12935), .Z(n12932) );
  INV_X1 U7195 ( .A(n9321), .ZN(n9328) );
  INV_X1 U7196 ( .A(n11804), .ZN(n9552) );
  INV_X2 U7197 ( .A(n8969), .ZN(n7406) );
  INV_X1 U7198 ( .A(n11042), .ZN(n8768) );
  CLKBUF_X2 U7199 ( .A(n10292), .Z(n10283) );
  AND2_X1 U7200 ( .A1(n10083), .A2(n9989), .ZN(n10297) );
  NAND2_X1 U7201 ( .A1(n9600), .A2(n9601), .ZN(n9587) );
  NAND2_X1 U7202 ( .A1(n7893), .A2(n13430), .ZN(n10714) );
  INV_X1 U7203 ( .A(n12988), .ZN(n8346) );
  INV_X1 U7204 ( .A(n13172), .ZN(n13168) );
  INV_X1 U7205 ( .A(n14310), .ZN(n8989) );
  INV_X1 U7206 ( .A(n8996), .ZN(n9262) );
  INV_X1 U7207 ( .A(n9614), .ZN(n9959) );
  AND2_X2 U7208 ( .A1(n6937), .A2(n6936), .ZN(n11498) );
  OR2_X1 U7209 ( .A1(n9600), .A2(n15422), .ZN(n9602) );
  INV_X1 U7210 ( .A(n8346), .ZN(n12985) );
  NAND2_X1 U7211 ( .A1(n12944), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6958) );
  NAND2_X1 U7212 ( .A1(n7250), .A2(n8780), .ZN(n14393) );
  NAND2_X1 U7214 ( .A1(n8747), .A2(n8746), .ZN(n14275) );
  AND2_X1 U7215 ( .A1(n8872), .A2(n8871), .ZN(n10453) );
  NAND2_X1 U7216 ( .A1(n9659), .A2(n9658), .ZN(n11868) );
  NAND4_X2 U7218 ( .A1(n9696), .A2(n9695), .A3(n9694), .A4(n9693), .ZN(n14815)
         );
  INV_X1 U7219 ( .A(n15023), .ZN(n15383) );
  OR2_X1 U7220 ( .A1(n7887), .A2(n10850), .ZN(n6426) );
  AND2_X1 U7221 ( .A1(n12343), .A2(n13383), .ZN(n6427) );
  OR2_X1 U7222 ( .A1(n14085), .A2(n6922), .ZN(n6428) );
  INV_X2 U7223 ( .A(n10299), .ZN(n10292) );
  NAND2_X2 U7225 ( .A1(n10018), .A2(n10016), .ZN(n7278) );
  AND2_X2 U7226 ( .A1(n13479), .A2(n7315), .ZN(n7961) );
  INV_X1 U7227 ( .A(n8153), .ZN(n8126) );
  NOR2_X2 U7228 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7350) );
  OR2_X2 U7229 ( .A1(n9631), .A2(n10797), .ZN(n9628) );
  AOI22_X2 U7230 ( .A1(n13219), .A2(n13218), .B1(n12939), .B2(n12934), .ZN(
        n12937) );
  INV_X1 U7231 ( .A(n11830), .ZN(n11564) );
  NOR2_X1 U7232 ( .A1(n15171), .A2(n10567), .ZN(n15138) );
  NAND2_X4 U7233 ( .A1(n8885), .A2(n14647), .ZN(n11042) );
  XNOR2_X2 U7234 ( .A(n10886), .B(n10885), .ZN(n10884) );
  NAND2_X2 U7235 ( .A1(n10805), .A2(n10804), .ZN(n10886) );
  BUF_X4 U7236 ( .A(n9854), .Z(n6429) );
  NAND2_X1 U7237 ( .A1(n9590), .A2(n9589), .ZN(n9854) );
  NAND2_X2 U7238 ( .A1(n15127), .A2(n10021), .ZN(n15110) );
  OAI211_X4 U7239 ( .C1(n6857), .C2(n6854), .A(n15128), .B(n6853), .ZN(n15127)
         );
  OAI21_X2 U7240 ( .B1(n13259), .B2(n7446), .A(n7442), .ZN(n13282) );
  NAND2_X2 U7241 ( .A1(n13316), .A2(n12913), .ZN(n13259) );
  NOR2_X2 U7242 ( .A1(n6432), .A2(n11390), .ZN(n13716) );
  CLKBUF_X2 U7243 ( .A(n13723), .Z(n6432) );
  XNOR2_X2 U7244 ( .A(n7855), .B(P3_IR_REG_1__SCAN_IN), .ZN(n8113) );
  AOI21_X2 U7245 ( .B1(n7481), .B2(n7482), .A(n6524), .ZN(n7479) );
  INV_X2 U7246 ( .A(n13054), .ZN(n13059) );
  XNOR2_X2 U7247 ( .A(n15523), .B(n14819), .ZN(n11321) );
  OAI21_X2 U7248 ( .B1(n8826), .B2(n8825), .A(n8824), .ZN(n8831) );
  INV_X4 U7249 ( .A(n11365), .ZN(n13188) );
  XNOR2_X2 U7250 ( .A(n8781), .B(n8788), .ZN(n11774) );
  XNOR2_X2 U7251 ( .A(n8792), .B(SI_20_), .ZN(n8781) );
  XNOR2_X2 U7252 ( .A(n10991), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n10896) );
  NAND2_X2 U7253 ( .A1(n10889), .A2(n10888), .ZN(n10991) );
  XNOR2_X1 U7254 ( .A(n15548), .B(n14815), .ZN(n12028) );
  AOI21_X2 U7255 ( .B1(n6427), .B2(n7441), .A(n6562), .ZN(n7440) );
  OAI21_X2 U7256 ( .B1(n11329), .B2(n11212), .A(n11211), .ZN(n11214) );
  AOI21_X2 U7257 ( .B1(n11332), .B2(n11331), .A(n11330), .ZN(n11329) );
  INV_X1 U7258 ( .A(n11458), .ZN(n14993) );
  AND2_X4 U7259 ( .A1(n8471), .A2(n6978), .ZN(n12988) );
  OAI21_X2 U7260 ( .B1(n6741), .B2(n7990), .A(n6738), .ZN(n7991) );
  MUX2_X1 U7261 ( .A(n15378), .B(n15377), .S(n15550), .Z(n15379) );
  AND2_X1 U7262 ( .A1(n15315), .A2(n6819), .ZN(n15401) );
  MUX2_X1 U7263 ( .A(n15281), .B(n15377), .S(n15554), .Z(n15282) );
  CLKBUF_X1 U7264 ( .A(n13459), .Z(n7093) );
  AND2_X1 U7265 ( .A1(n15121), .A2(n10017), .ZN(n15158) );
  NAND2_X1 U7266 ( .A1(n12145), .A2(n10004), .ZN(n12188) );
  NAND2_X1 U7267 ( .A1(n6946), .A2(n6944), .ZN(n8773) );
  NAND2_X1 U7268 ( .A1(n11575), .A2(n11576), .ZN(n11574) );
  CLKBUF_X1 U7269 ( .A(n6430), .Z(n7063) );
  INV_X1 U7270 ( .A(n13974), .ZN(n12372) );
  INV_X2 U7271 ( .A(n10294), .ZN(n10105) );
  AOI21_X1 U7272 ( .B1(n11982), .B2(n9478), .A(n12264), .ZN(n9370) );
  INV_X1 U7273 ( .A(n11979), .ZN(n15649) );
  INV_X2 U7274 ( .A(n10616), .ZN(n10582) );
  NAND4_X2 U7275 ( .A1(n9608), .A2(n9610), .A3(n9606), .A4(n9607), .ZN(n10096)
         );
  CLKBUF_X2 U7276 ( .A(n9328), .Z(n12875) );
  BUF_X2 U7277 ( .A(n9691), .Z(n10615) );
  NAND2_X2 U7278 ( .A1(n8471), .A2(n10817), .ZN(n8110) );
  NAND2_X1 U7279 ( .A1(n13214), .A2(n15428), .ZN(n9691) );
  NAND2_X2 U7280 ( .A1(n8950), .A2(n8949), .ZN(n9464) );
  XNOR2_X1 U7281 ( .A(n7915), .B(n7914), .ZN(n7966) );
  NOR2_X1 U7282 ( .A1(n6967), .A2(n6968), .ZN(n8084) );
  OR2_X1 U7283 ( .A1(n9845), .A2(n9844), .ZN(n9979) );
  INV_X1 U7284 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7866) );
  INV_X1 U7285 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7094) );
  INV_X1 U7286 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7854) );
  INV_X1 U7287 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7448) );
  AND2_X1 U7288 ( .A1(n9352), .A2(n7633), .ZN(n7002) );
  OAI211_X1 U7289 ( .C1(n10608), .C2(n6835), .A(n7790), .B(n6833), .ZN(n10694)
         );
  OR2_X1 U7290 ( .A1(n10076), .A2(n15552), .ZN(n10079) );
  AND3_X1 U7291 ( .A1(n6686), .A2(n6713), .A3(n6685), .ZN(n15381) );
  NAND2_X1 U7292 ( .A1(n6642), .A2(n10271), .ZN(n14699) );
  AOI21_X1 U7293 ( .B1(n13672), .B2(n13718), .A(n13545), .ZN(n13674) );
  OAI211_X1 U7294 ( .C1(n15096), .C2(n15354), .A(n15095), .B(n15094), .ZN(
        n15307) );
  AND2_X1 U7295 ( .A1(n15280), .A2(n15279), .ZN(n15377) );
  AND2_X1 U7296 ( .A1(n10631), .A2(n10630), .ZN(n10635) );
  INV_X1 U7297 ( .A(n15014), .ZN(n7730) );
  NAND2_X1 U7298 ( .A1(n6890), .A2(n6887), .ZN(n15448) );
  AND2_X1 U7299 ( .A1(n9484), .A2(n9483), .ZN(n9494) );
  NAND2_X1 U7300 ( .A1(n6964), .A2(n6963), .ZN(n13257) );
  AND2_X1 U7301 ( .A1(n10379), .A2(n8853), .ZN(n14078) );
  OR2_X1 U7302 ( .A1(n6893), .A2(n6590), .ZN(n6890) );
  NAND2_X1 U7303 ( .A1(n14146), .A2(n10366), .ZN(n14131) );
  XNOR2_X1 U7304 ( .A(n9214), .B(n9204), .ZN(n13811) );
  AND2_X1 U7305 ( .A1(n10641), .A2(n10640), .ZN(n15376) );
  NAND2_X1 U7306 ( .A1(n13318), .A2(n13317), .ZN(n13316) );
  XNOR2_X1 U7307 ( .A(n8861), .B(n8856), .ZN(n13212) );
  NAND2_X1 U7308 ( .A1(n10212), .A2(n10211), .ZN(n14782) );
  OAI21_X1 U7309 ( .B1(n10578), .B2(n10577), .A(n10576), .ZN(n10580) );
  CLKBUF_X1 U7310 ( .A(n13634), .Z(n6988) );
  NAND2_X1 U7311 ( .A1(n8850), .A2(n8855), .ZN(n14634) );
  OR2_X1 U7312 ( .A1(n8849), .A2(n8848), .ZN(n8850) );
  NAND2_X1 U7313 ( .A1(n9952), .A2(n9951), .ZN(n15023) );
  AND2_X1 U7314 ( .A1(n7741), .A2(n6919), .ZN(n6918) );
  NAND2_X1 U7315 ( .A1(n9943), .A2(n9942), .ZN(n15042) );
  NAND2_X1 U7316 ( .A1(n8836), .A2(n8835), .ZN(n14356) );
  XNOR2_X1 U7317 ( .A(n8843), .B(n8842), .ZN(n12890) );
  NOR2_X1 U7318 ( .A1(n10718), .A2(n6995), .ZN(n7957) );
  NAND2_X1 U7319 ( .A1(n8395), .A2(n8394), .ZN(n13756) );
  NAND2_X1 U7320 ( .A1(n8786), .A2(n8785), .ZN(n14196) );
  NAND2_X2 U7321 ( .A1(n8800), .A2(n8799), .ZN(n14378) );
  NAND2_X2 U7322 ( .A1(n6638), .A2(n9860), .ZN(n15151) );
  NAND2_X1 U7323 ( .A1(n8363), .A2(n8362), .ZN(n13775) );
  NAND2_X1 U7324 ( .A1(n8384), .A2(n8383), .ZN(n13762) );
  XNOR2_X1 U7325 ( .A(n8798), .B(n8797), .ZN(n12045) );
  XNOR2_X1 U7326 ( .A(n6639), .B(n8784), .ZN(n11823) );
  NAND2_X1 U7327 ( .A1(n12146), .A2(n12152), .ZN(n12145) );
  NAND2_X1 U7328 ( .A1(n9795), .A2(n9794), .ZN(n15271) );
  NAND2_X1 U7329 ( .A1(n9815), .A2(n9814), .ZN(n15345) );
  XNOR2_X1 U7330 ( .A(n12720), .B(n7287), .ZN(n12710) );
  NAND2_X1 U7331 ( .A1(n7012), .A2(n10002), .ZN(n7701) );
  AND2_X1 U7332 ( .A1(n7304), .A2(n7303), .ZN(n13387) );
  NAND2_X1 U7333 ( .A1(n8675), .A2(n8674), .ZN(n12609) );
  XNOR2_X1 U7334 ( .A(n8748), .B(n8749), .ZN(n11195) );
  NAND2_X1 U7335 ( .A1(n8731), .A2(n8730), .ZN(n14546) );
  OR2_X1 U7336 ( .A1(n11842), .A2(n11845), .ZN(n7304) );
  NAND2_X1 U7337 ( .A1(n7697), .A2(n9745), .ZN(n12423) );
  OAI22_X1 U7338 ( .A1(n7354), .A2(n7353), .B1(n10493), .B2(n7352), .ZN(n10496) );
  OR2_X1 U7339 ( .A1(n12251), .A2(n12445), .ZN(n12401) );
  NAND2_X1 U7340 ( .A1(n11290), .A2(n11291), .ZN(n11553) );
  NAND2_X1 U7341 ( .A1(n8644), .A2(n8643), .ZN(n12409) );
  NAND2_X1 U7342 ( .A1(n8632), .A2(n8631), .ZN(n12445) );
  NOR2_X1 U7343 ( .A1(n7626), .A2(n11937), .ZN(n12252) );
  AND2_X1 U7344 ( .A1(n6924), .A2(n10101), .ZN(n7794) );
  NAND2_X1 U7345 ( .A1(n8623), .A2(n8622), .ZN(n15624) );
  NAND2_X1 U7346 ( .A1(n9687), .A2(n9686), .ZN(n15548) );
  INV_X1 U7347 ( .A(n12064), .ZN(n12104) );
  NAND2_X1 U7348 ( .A1(n8612), .A2(n8613), .ZN(n12064) );
  INV_X1 U7349 ( .A(n12935), .ZN(n6430) );
  NAND4_X1 U7350 ( .A1(n9000), .A2(n8999), .A3(n8998), .A4(n8997), .ZN(n13977)
         );
  NAND2_X1 U7351 ( .A1(n8586), .A2(n8585), .ZN(n15657) );
  NAND2_X1 U7352 ( .A1(n6804), .A2(n8618), .ZN(n6645) );
  NAND2_X1 U7353 ( .A1(n6789), .A2(n8164), .ZN(n15699) );
  NAND2_X1 U7354 ( .A1(n7591), .A2(n7589), .ZN(n8254) );
  NAND2_X1 U7355 ( .A1(n8616), .A2(n8615), .ZN(n6804) );
  AND4_X2 U7356 ( .A1(n9593), .A2(n9594), .A3(n9595), .A4(n9592), .ZN(n11156)
         );
  OR2_X1 U7357 ( .A1(n11394), .A2(n6644), .ZN(n11396) );
  INV_X1 U7360 ( .A(n10453), .ZN(n9533) );
  NAND2_X1 U7361 ( .A1(n15653), .A2(n10453), .ZN(n9401) );
  NAND2_X1 U7362 ( .A1(n10084), .A2(n10083), .ZN(n10252) );
  OAI211_X1 U7363 ( .C1(n8866), .C2(n10806), .A(n8576), .B(n8575), .ZN(n13827)
         );
  NAND2_X1 U7364 ( .A1(n10621), .A2(n7388), .ZN(n10527) );
  AND3_X1 U7365 ( .A1(n8686), .A2(n8687), .A3(n8688), .ZN(n8708) );
  INV_X2 U7366 ( .A(n8983), .ZN(n9259) );
  AND2_X1 U7367 ( .A1(n8634), .A2(n6987), .ZN(n7481) );
  INV_X1 U7368 ( .A(n11924), .ZN(n10430) );
  MUX2_X1 U7369 ( .A(P2_IR_REG_0__SCAN_IN), .B(n14648), .S(n11042), .Z(n11485)
         );
  XNOR2_X1 U7370 ( .A(n7892), .B(n7891), .ZN(n13430) );
  OAI211_X1 U7371 ( .C1(n8880), .C2(n8879), .A(n8878), .B(n8877), .ZN(n11924)
         );
  NAND2_X1 U7372 ( .A1(n10472), .A2(n11825), .ZN(n10617) );
  AND2_X1 U7373 ( .A1(n7912), .A2(n6473), .ZN(n13054) );
  XNOR2_X1 U7374 ( .A(n8547), .B(n8548), .ZN(n10875) );
  MUX2_X1 U7375 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7812), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n7825) );
  NAND2_X1 U7376 ( .A1(n10043), .A2(n10044), .ZN(n12109) );
  INV_X1 U7377 ( .A(n10031), .ZN(n11825) );
  INV_X1 U7378 ( .A(n8614), .ZN(n8615) );
  AND2_X1 U7379 ( .A1(n7704), .A2(n6826), .ZN(n9590) );
  XNOR2_X1 U7380 ( .A(n6683), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8949) );
  XNOR2_X1 U7381 ( .A(n8463), .B(n8462), .ZN(n11804) );
  MUX2_X1 U7382 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7911), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n7912) );
  AOI21_X1 U7383 ( .B1(n8571), .B2(n8570), .A(n8569), .ZN(n8600) );
  XNOR2_X1 U7384 ( .A(n8617), .B(SI_6_), .ZN(n8614) );
  OAI21_X1 U7385 ( .B1(n8650), .B2(P2_DATAO_REG_3__SCAN_IN), .A(n7028), .ZN(
        n8582) );
  INV_X1 U7386 ( .A(n8684), .ZN(n6431) );
  INV_X2 U7387 ( .A(n14640), .ZN(n14646) );
  XNOR2_X1 U7388 ( .A(n8085), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8087) );
  OR2_X1 U7389 ( .A1(n14629), .A2(n14630), .ZN(n8890) );
  OR2_X1 U7390 ( .A1(n8084), .A2(n8083), .ZN(n8085) );
  XNOR2_X1 U7391 ( .A(n8543), .B(n8541), .ZN(n14647) );
  NAND2_X1 U7392 ( .A1(n8145), .A2(n8144), .ZN(n8147) );
  NOR2_X1 U7393 ( .A1(n6764), .A2(n7820), .ZN(n7826) );
  NOR2_X1 U7394 ( .A1(n9587), .A2(n7707), .ZN(n7703) );
  AND3_X1 U7395 ( .A1(n7833), .A2(n7805), .A3(n6594), .ZN(n8460) );
  NAND2_X1 U7396 ( .A1(n9603), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9605) );
  NAND2_X1 U7397 ( .A1(n9979), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9981) );
  OAI21_X1 U7398 ( .B1(n10818), .B2(n10797), .A(n7020), .ZN(n8567) );
  XNOR2_X1 U7399 ( .A(n7094), .B(n7862), .ZN(n11344) );
  INV_X4 U7400 ( .A(n10818), .ZN(n10786) );
  BUF_X1 U7401 ( .A(n7973), .Z(n11122) );
  AND2_X1 U7402 ( .A1(n8744), .A2(n8743), .ZN(n8765) );
  OR2_X1 U7403 ( .A1(n9845), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n9843) );
  NAND3_X1 U7404 ( .A1(n7824), .A2(n7913), .A3(n7821), .ZN(n6968) );
  XNOR2_X1 U7405 ( .A(n7866), .B(n7867), .ZN(n11219) );
  NAND2_X1 U7406 ( .A1(n8556), .A2(n8573), .ZN(n8577) );
  OAI211_X1 U7407 ( .C1(n6731), .C2(n15422), .A(n9622), .B(n6730), .ZN(n14828)
         );
  AND2_X1 U7408 ( .A1(n8544), .A2(n14413), .ZN(n8556) );
  AND2_X1 U7409 ( .A1(n7975), .A2(n7854), .ZN(n7846) );
  INV_X1 U7410 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9699) );
  INV_X4 U7411 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7412 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9841) );
  INV_X1 U7413 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7816) );
  INV_X1 U7414 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9839) );
  INV_X1 U7415 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7809) );
  NOR2_X1 U7416 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n9571) );
  INV_X1 U7417 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n7452) );
  INV_X1 U7418 ( .A(P1_RD_REG_SCAN_IN), .ZN(n8061) );
  INV_X1 U7419 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n14072) );
  NOR2_X2 U7420 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7975) );
  INV_X1 U7421 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9633) );
  INV_X1 U7422 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7879) );
  INV_X4 U7423 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7424 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8544) );
  INV_X4 U7425 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7426 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9656) );
  INV_X1 U7427 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9769) );
  NOR2_X1 U7428 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9580) );
  INV_X1 U7429 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7869) );
  INV_X1 U7430 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9766) );
  NOR2_X1 U7431 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7351) );
  INV_X1 U7432 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7837) );
  INV_X1 U7433 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8764) );
  INV_X1 U7434 ( .A(n10527), .ZN(n6433) );
  OR2_X1 U7435 ( .A1(n13194), .A2(n8087), .ZN(n8137) );
  OAI222_X1 U7436 ( .A1(n13805), .A2(n13197), .B1(P3_U3151), .B2(n13194), .C1(
        n13808), .C2(n13196), .ZN(P3_U3265) );
  NAND2_X1 U7437 ( .A1(n13194), .A2(n8087), .ZN(n9321) );
  OAI21_X2 U7438 ( .B1(n7083), .B2(n11778), .A(n6969), .ZN(n11781) );
  NOR2_X4 U7439 ( .A1(n12422), .A2(n12423), .ZN(n12565) );
  OR2_X2 U7440 ( .A1(n12334), .A2(n14674), .ZN(n12422) );
  INV_X1 U7441 ( .A(n8328), .ZN(n7205) );
  INV_X1 U7442 ( .A(n8138), .ZN(n9318) );
  NAND2_X1 U7443 ( .A1(n13216), .A2(n8949), .ZN(n8983) );
  OAI21_X1 U7444 ( .B1(n9424), .B2(n9423), .A(n9422), .ZN(n9426) );
  AOI21_X1 U7445 ( .B1(n6762), .B2(n13133), .A(n13134), .ZN(n13138) );
  NOR2_X1 U7446 ( .A1(n8403), .A2(n7218), .ZN(n7217) );
  OAI21_X1 U7447 ( .B1(n7743), .B2(n7744), .A(n10361), .ZN(n7269) );
  NAND2_X1 U7448 ( .A1(n6897), .A2(n6896), .ZN(n10771) );
  AND2_X1 U7449 ( .A1(n13516), .A2(n12997), .ZN(n13180) );
  OR2_X1 U7450 ( .A1(n9309), .A2(n9308), .ZN(n13171) );
  NAND2_X1 U7451 ( .A1(n7201), .A2(n6453), .ZN(n13634) );
  NOR2_X1 U7452 ( .A1(n8032), .A2(n7180), .ZN(n7179) );
  INV_X1 U7453 ( .A(n8029), .ZN(n7180) );
  NOR2_X1 U7454 ( .A1(n14393), .A2(n13964), .ZN(n10359) );
  NAND2_X1 U7455 ( .A1(n7751), .A2(n7749), .ZN(n14258) );
  NOR2_X1 U7456 ( .A1(n9523), .A2(n7750), .ZN(n7749) );
  INV_X1 U7457 ( .A(n10353), .ZN(n7750) );
  NOR2_X1 U7458 ( .A1(n6480), .A2(n7754), .ZN(n7753) );
  INV_X1 U7459 ( .A(n10347), .ZN(n7754) );
  INV_X1 U7460 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8882) );
  NOR2_X1 U7461 ( .A1(n12720), .A2(n12567), .ZN(n7763) );
  NAND2_X1 U7462 ( .A1(n6979), .A2(n6512), .ZN(n8715) );
  NAND2_X1 U7463 ( .A1(n8708), .A2(n8702), .ZN(n6979) );
  INV_X1 U7464 ( .A(n8699), .ZN(n8701) );
  AND4_X1 U7465 ( .A1(n8263), .A2(n8262), .A3(n8261), .A4(n8260), .ZN(n13275)
         );
  NAND2_X1 U7466 ( .A1(n7214), .A2(n7212), .ZN(n13554) );
  AND2_X1 U7467 ( .A1(n7213), .A2(n7641), .ZN(n7212) );
  NOR2_X1 U7468 ( .A1(n6545), .A2(n7670), .ZN(n7669) );
  INV_X1 U7469 ( .A(n8315), .ZN(n7670) );
  NAND2_X1 U7470 ( .A1(n7747), .A2(n6472), .ZN(n7255) );
  NAND2_X1 U7471 ( .A1(n10444), .A2(n9512), .ZN(n10432) );
  OR2_X1 U7472 ( .A1(n14087), .A2(n14093), .ZN(n9512) );
  XNOR2_X1 U7473 ( .A(n14149), .B(n14160), .ZN(n14143) );
  NAND2_X1 U7474 ( .A1(n6865), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6683) );
  OR2_X1 U7475 ( .A1(n9965), .A2(n6517), .ZN(n7528) );
  INV_X1 U7476 ( .A(n7526), .ZN(n7525) );
  OAI22_X1 U7477 ( .A1(n9965), .A2(n7527), .B1(n15023), .B2(n12964), .ZN(n7526) );
  OR2_X1 U7478 ( .A1(n9927), .A2(n9926), .ZN(n9957) );
  OR2_X1 U7479 ( .A1(n6856), .A2(n6491), .ZN(n6854) );
  OR2_X1 U7480 ( .A1(n6858), .A2(n6491), .ZN(n6853) );
  NAND2_X1 U7481 ( .A1(n7100), .A2(n13859), .ZN(n9363) );
  NAND2_X1 U7482 ( .A1(n9478), .A2(n10330), .ZN(n7101) );
  NAND2_X1 U7483 ( .A1(n9359), .A2(n9361), .ZN(n7102) );
  NAND2_X1 U7484 ( .A1(n9367), .A2(n11710), .ZN(n9368) );
  MUX2_X1 U7485 ( .A(n10488), .B(n10487), .S(n6433), .Z(n10489) );
  INV_X1 U7486 ( .A(n10559), .ZN(n10541) );
  AND2_X1 U7487 ( .A1(n6502), .A2(n7070), .ZN(n6677) );
  INV_X1 U7488 ( .A(n9428), .ZN(n7070) );
  AND2_X1 U7489 ( .A1(n7358), .A2(n7076), .ZN(n7075) );
  INV_X1 U7490 ( .A(n9429), .ZN(n7076) );
  NAND2_X1 U7491 ( .A1(n7357), .A2(n9429), .ZN(n7356) );
  NAND2_X1 U7492 ( .A1(n7359), .A2(n7358), .ZN(n7357) );
  XNOR2_X1 U7493 ( .A(n14993), .B(n11127), .ZN(n10472) );
  NAND2_X1 U7494 ( .A1(n6659), .A2(n9444), .ZN(n9448) );
  NAND2_X1 U7495 ( .A1(n9446), .A2(n9445), .ZN(n6659) );
  INV_X1 U7496 ( .A(n9445), .ZN(n7073) );
  NAND2_X1 U7497 ( .A1(n10617), .A2(n10471), .ZN(n10621) );
  NAND3_X1 U7498 ( .A1(n6650), .A2(n6649), .A3(n6648), .ZN(n7814) );
  INV_X1 U7499 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n6649) );
  INV_X1 U7500 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n6648) );
  NAND2_X1 U7501 ( .A1(n10419), .A2(n7548), .ZN(n7547) );
  INV_X1 U7502 ( .A(n10418), .ZN(n7548) );
  INV_X1 U7503 ( .A(n6478), .ZN(n6906) );
  AND2_X1 U7504 ( .A1(n8742), .A2(n7779), .ZN(n8744) );
  NAND2_X1 U7505 ( .A1(n6832), .A2(n7386), .ZN(n10604) );
  NAND2_X1 U7506 ( .A1(n10599), .A2(n7387), .ZN(n7386) );
  OAI21_X1 U7507 ( .B1(n10596), .B2(n6831), .A(n6829), .ZN(n6832) );
  NOR2_X1 U7508 ( .A1(n10598), .A2(n10595), .ZN(n6831) );
  INV_X1 U7509 ( .A(n7520), .ZN(n6818) );
  NAND2_X1 U7510 ( .A1(n8668), .A2(n10872), .ZN(n8687) );
  OAI21_X1 U7511 ( .B1(n8650), .B2(n10862), .A(n7033), .ZN(n8636) );
  NAND2_X1 U7512 ( .A1(n8650), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7033) );
  NAND2_X1 U7513 ( .A1(n11206), .A2(n7982), .ZN(n7983) );
  OAI21_X1 U7514 ( .B1(n7507), .B2(n7508), .A(n7500), .ZN(n7503) );
  NAND2_X1 U7515 ( .A1(n11027), .A2(n6526), .ZN(n7502) );
  AND2_X1 U7516 ( .A1(n7501), .A2(n11352), .ZN(n7500) );
  AND2_X1 U7517 ( .A1(n10845), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7990) );
  NAND2_X1 U7518 ( .A1(n13463), .A2(n7518), .ZN(n7900) );
  INV_X1 U7519 ( .A(n9317), .ZN(n9350) );
  NAND2_X1 U7520 ( .A1(n7223), .A2(n8079), .ZN(n8464) );
  NAND2_X1 U7521 ( .A1(n13540), .A2(n8456), .ZN(n7672) );
  NOR2_X1 U7522 ( .A1(n8447), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n7223) );
  AOI21_X1 U7523 ( .B1(n7217), .B2(n13003), .A(n6522), .ZN(n7216) );
  NAND2_X1 U7524 ( .A1(n13603), .A2(n7217), .ZN(n7215) );
  OR2_X1 U7525 ( .A1(n13789), .A2(n13373), .ZN(n13037) );
  NOR2_X1 U7526 ( .A1(n12203), .A2(n7640), .ZN(n7639) );
  INV_X1 U7527 ( .A(n12201), .ZN(n7640) );
  OR2_X1 U7528 ( .A1(n13278), .A2(n13270), .ZN(n13117) );
  INV_X1 U7529 ( .A(n6968), .ZN(n6966) );
  NAND2_X1 U7530 ( .A1(n6654), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7916) );
  AOI21_X1 U7531 ( .B1(n7190), .B2(n7192), .A(n6627), .ZN(n7188) );
  NAND2_X1 U7532 ( .A1(n8460), .A2(n6494), .ZN(n7909) );
  AND2_X1 U7533 ( .A1(n8018), .A2(n8015), .ZN(n7614) );
  INV_X1 U7534 ( .A(n8191), .ZN(n8018) );
  NAND2_X1 U7535 ( .A1(n10806), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8009) );
  NAND2_X1 U7536 ( .A1(n8852), .A2(n8851), .ZN(n14352) );
  AND2_X1 U7537 ( .A1(n6688), .A2(n6438), .ZN(n7553) );
  OR2_X1 U7538 ( .A1(n14111), .A2(n7558), .ZN(n7557) );
  AND2_X1 U7539 ( .A1(n6463), .A2(n14099), .ZN(n6797) );
  OR2_X1 U7540 ( .A1(n9243), .A2(n9241), .ZN(n9256) );
  INV_X1 U7541 ( .A(n10337), .ZN(n6901) );
  NAND2_X1 U7542 ( .A1(n10330), .A2(n13859), .ZN(n10384) );
  INV_X1 U7543 ( .A(n11044), .ZN(n9288) );
  INV_X1 U7544 ( .A(n8853), .ZN(n7611) );
  NOR2_X1 U7545 ( .A1(n12817), .A2(n14562), .ZN(n14311) );
  INV_X1 U7546 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8887) );
  AOI21_X1 U7547 ( .B1(n7761), .B2(n10283), .A(n10203), .ZN(n10205) );
  AND2_X1 U7548 ( .A1(n9671), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9688) );
  INV_X1 U7549 ( .A(n9673), .ZN(n9671) );
  OR2_X1 U7550 ( .A1(n10637), .A2(n10636), .ZN(n7784) );
  NOR2_X1 U7551 ( .A1(n9872), .A2(n14694), .ZN(n6675) );
  OR2_X1 U7552 ( .A1(n15345), .A2(n15242), .ZN(n10546) );
  OR2_X1 U7553 ( .A1(n12770), .A2(n14788), .ZN(n10531) );
  OR2_X1 U7554 ( .A1(n15199), .A2(n10225), .ZN(n10562) );
  INV_X1 U7555 ( .A(n11253), .ZN(n7049) );
  NAND2_X1 U7556 ( .A1(n8832), .A2(n7455), .ZN(n8838) );
  NAND2_X1 U7557 ( .A1(n7260), .A2(n7261), .ZN(n6640) );
  AND2_X1 U7558 ( .A1(n8716), .A2(n7262), .ZN(n7261) );
  AOI21_X1 U7559 ( .B1(n8715), .B2(n8714), .A(n8713), .ZN(n8716) );
  NAND2_X1 U7560 ( .A1(n8714), .A2(n8694), .ZN(n8699) );
  XNOR2_X1 U7561 ( .A(n8689), .B(SI_13_), .ZN(n8688) );
  OR2_X1 U7562 ( .A1(n9755), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9756) );
  NAND2_X1 U7563 ( .A1(n8659), .A2(n10848), .ZN(n8684) );
  INV_X1 U7564 ( .A(n6717), .ZN(n7457) );
  XNOR2_X1 U7565 ( .A(n8636), .B(SI_8_), .ZN(n8633) );
  XNOR2_X1 U7566 ( .A(n8625), .B(SI_7_), .ZN(n8624) );
  NOR2_X1 U7567 ( .A1(n8568), .A2(n10839), .ZN(n8569) );
  INV_X1 U7568 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10765) );
  INV_X1 U7569 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7295) );
  NAND2_X1 U7570 ( .A1(n10771), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n7121) );
  OAI21_X1 U7571 ( .B1(n12923), .B2(n13238), .A(n12922), .ZN(n12924) );
  INV_X1 U7572 ( .A(n7171), .ZN(n7170) );
  NAND2_X1 U7573 ( .A1(n9350), .A2(n9318), .ZN(n12883) );
  AOI21_X1 U7574 ( .B1(n13525), .B2(n9318), .A(n8469), .ZN(n9308) );
  AND2_X1 U7575 ( .A1(n8380), .A2(n8379), .ZN(n13251) );
  NAND2_X1 U7576 ( .A1(n8126), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8107) );
  AND2_X1 U7577 ( .A1(n8109), .A2(n8106), .ZN(n6962) );
  OR2_X1 U7578 ( .A1(n8137), .A2(n15689), .ZN(n8106) );
  AND2_X1 U7579 ( .A1(n7984), .A2(n10734), .ZN(n11030) );
  NAND2_X1 U7580 ( .A1(n7032), .A2(n7054), .ZN(n7984) );
  INV_X1 U7581 ( .A(n7983), .ZN(n7032) );
  INV_X1 U7582 ( .A(n13388), .ZN(n7303) );
  NAND2_X1 U7583 ( .A1(n11839), .A2(n13398), .ZN(n6741) );
  INV_X1 U7584 ( .A(n6739), .ZN(n6738) );
  OAI21_X1 U7585 ( .B1(n6740), .B2(n7990), .A(n10850), .ZN(n6739) );
  NOR2_X1 U7586 ( .A1(n7885), .A2(n12659), .ZN(n7511) );
  OAI211_X1 U7587 ( .C1(n7343), .C2(n7341), .A(n7340), .B(n7996), .ZN(n7997)
         );
  NAND2_X1 U7588 ( .A1(n7345), .A2(n7337), .ZN(n7340) );
  AND2_X1 U7589 ( .A1(n7969), .A2(n7918), .ZN(n8002) );
  INV_X1 U7590 ( .A(n7642), .ZN(n7641) );
  NAND2_X1 U7591 ( .A1(n7645), .A2(n8417), .ZN(n7644) );
  NAND2_X1 U7592 ( .A1(n7047), .A2(n7204), .ZN(n7201) );
  OAI21_X1 U7593 ( .B1(n12613), .B2(n6786), .A(n6783), .ZN(n12758) );
  AOI21_X1 U7594 ( .B1(n6787), .B2(n6785), .A(n6784), .ZN(n6783) );
  INV_X1 U7595 ( .A(n6787), .ZN(n6786) );
  INV_X1 U7596 ( .A(n13135), .ZN(n6784) );
  AND3_X1 U7597 ( .A1(n8116), .A2(n8115), .A3(n8114), .ZN(n13732) );
  OR2_X1 U7598 ( .A1(n8110), .A2(n10842), .ZN(n8116) );
  OAI211_X1 U7599 ( .C1(n12992), .C2(n12991), .A(n12990), .B(n12989), .ZN(
        n13516) );
  OR2_X1 U7600 ( .A1(n13702), .A2(n13249), .ZN(n13043) );
  NAND2_X1 U7601 ( .A1(n8320), .A2(n8319), .ZN(n13712) );
  AOI21_X1 U7602 ( .B1(n7665), .B2(n7209), .A(n6529), .ZN(n7208) );
  INV_X1 U7603 ( .A(n7795), .ZN(n7209) );
  NAND2_X1 U7604 ( .A1(n7211), .A2(n7795), .ZN(n7666) );
  INV_X1 U7605 ( .A(n12276), .ZN(n7211) );
  AND2_X1 U7606 ( .A1(n13168), .A2(n8472), .ZN(n13724) );
  AND2_X1 U7607 ( .A1(n13168), .A2(n11281), .ZN(n13722) );
  NAND2_X1 U7608 ( .A1(n8344), .A2(n8343), .ZN(n8342) );
  NAND2_X1 U7609 ( .A1(n7175), .A2(n7173), .ZN(n8306) );
  AOI21_X1 U7610 ( .B1(n7176), .B2(n7178), .A(n7174), .ZN(n7173) );
  INV_X1 U7611 ( .A(n8033), .ZN(n7174) );
  INV_X1 U7612 ( .A(n7593), .ZN(n7592) );
  OAI21_X1 U7613 ( .B1(n8210), .B2(n7594), .A(n8234), .ZN(n7593) );
  NAND2_X1 U7614 ( .A1(n10830), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8019) );
  INV_X1 U7615 ( .A(n7587), .ZN(n7586) );
  OAI21_X1 U7616 ( .B1(n8159), .B2(n7588), .A(n8173), .ZN(n7587) );
  NAND2_X1 U7617 ( .A1(n8147), .A2(n8009), .ZN(n8160) );
  AND2_X1 U7618 ( .A1(n9129), .A2(n9128), .ZN(n12805) );
  AND2_X1 U7619 ( .A1(n9214), .A2(n9213), .ZN(n13812) );
  NAND2_X1 U7620 ( .A1(n7396), .A2(n6484), .ZN(n7395) );
  NAND2_X1 U7621 ( .A1(n6806), .A2(n11748), .ZN(n7396) );
  NAND2_X1 U7622 ( .A1(n6807), .A2(n9030), .ZN(n6806) );
  NAND2_X1 U7623 ( .A1(n6484), .A2(n9030), .ZN(n7397) );
  NAND2_X1 U7624 ( .A1(n6802), .A2(n6800), .ZN(n7130) );
  AOI21_X1 U7625 ( .B1(n13927), .B2(n6803), .A(n6801), .ZN(n6800) );
  NAND2_X1 U7626 ( .A1(n13926), .A2(n6803), .ZN(n6802) );
  AND2_X1 U7627 ( .A1(n13905), .A2(n7129), .ZN(n7128) );
  NAND2_X1 U7628 ( .A1(n13833), .A2(n13832), .ZN(n7129) );
  OR2_X1 U7629 ( .A1(n9220), .A2(n13900), .ZN(n9243) );
  XNOR2_X1 U7630 ( .A(n14378), .B(n8969), .ZN(n13814) );
  NAND2_X1 U7631 ( .A1(n7405), .A2(n7404), .ZN(n11637) );
  AND2_X1 U7632 ( .A1(n9006), .A2(n8995), .ZN(n7404) );
  NAND2_X1 U7633 ( .A1(n13861), .A2(n13862), .ZN(n13860) );
  NOR2_X1 U7634 ( .A1(n7410), .A2(n7134), .ZN(n7132) );
  INV_X1 U7635 ( .A(n6471), .ZN(n7410) );
  INV_X1 U7636 ( .A(n8566), .ZN(n8592) );
  NAND2_X1 U7637 ( .A1(n6438), .A2(n10429), .ZN(n7556) );
  INV_X1 U7638 ( .A(n10432), .ZN(n10375) );
  NAND2_X1 U7639 ( .A1(n10369), .A2(n6577), .ZN(n7747) );
  INV_X1 U7640 ( .A(n10368), .ZN(n7748) );
  AND2_X1 U7641 ( .A1(n14130), .A2(n10424), .ZN(n10425) );
  OAI21_X1 U7642 ( .B1(n14176), .B2(n7265), .A(n7263), .ZN(n14146) );
  INV_X1 U7643 ( .A(n7264), .ZN(n7263) );
  OAI21_X1 U7644 ( .B1(n7265), .B2(n14177), .A(n6552), .ZN(n7264) );
  NOR2_X1 U7645 ( .A1(n7267), .A2(n10363), .ZN(n7266) );
  INV_X1 U7646 ( .A(n10362), .ZN(n7267) );
  NAND2_X1 U7647 ( .A1(n14176), .A2(n14177), .ZN(n7268) );
  NAND2_X1 U7648 ( .A1(n14187), .A2(n10420), .ZN(n10422) );
  NOR2_X1 U7649 ( .A1(n10359), .A2(n10358), .ZN(n7744) );
  NOR2_X1 U7650 ( .A1(n10359), .A2(n10360), .ZN(n7743) );
  NAND2_X1 U7651 ( .A1(n6791), .A2(n7615), .ZN(n14208) );
  NOR2_X1 U7652 ( .A1(n14393), .A2(n7617), .ZN(n7615) );
  INV_X1 U7653 ( .A(n14298), .ZN(n6791) );
  NAND2_X1 U7654 ( .A1(n10352), .A2(n6508), .ZN(n7751) );
  INV_X1 U7655 ( .A(n14305), .ZN(n7752) );
  NAND2_X1 U7656 ( .A1(n14319), .A2(n10346), .ZN(n7755) );
  XNOR2_X1 U7657 ( .A(n11914), .B(n13976), .ZN(n11911) );
  NAND2_X1 U7658 ( .A1(n10387), .A2(n6796), .ZN(n10337) );
  INV_X1 U7659 ( .A(n15657), .ZN(n6796) );
  NAND2_X1 U7660 ( .A1(n11042), .A2(n10817), .ZN(n8566) );
  XNOR2_X1 U7661 ( .A(n7611), .B(n13960), .ZN(n10456) );
  OR2_X1 U7662 ( .A1(n8870), .A2(n8873), .ZN(n8872) );
  NAND2_X1 U7663 ( .A1(n8880), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8870) );
  NOR2_X1 U7664 ( .A1(n7678), .A2(n7680), .ZN(n7677) );
  NAND2_X1 U7665 ( .A1(n9688), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9705) );
  OR2_X1 U7666 ( .A1(n11498), .A2(n10252), .ZN(n10093) );
  AND2_X1 U7667 ( .A1(n10098), .A2(n10097), .ZN(n10099) );
  INV_X1 U7668 ( .A(n14785), .ZN(n7245) );
  OAI21_X1 U7669 ( .B1(n7688), .B2(n14680), .A(n6643), .ZN(n14751) );
  OAI21_X1 U7670 ( .B1(n7687), .B2(n6930), .A(n6926), .ZN(n6643) );
  NAND2_X1 U7671 ( .A1(n6928), .A2(n6927), .ZN(n6926) );
  INV_X1 U7672 ( .A(n9688), .ZN(n6680) );
  AOI21_X1 U7673 ( .B1(n15133), .B2(n9944), .A(n9888), .ZN(n14691) );
  INV_X1 U7674 ( .A(n9660), .ZN(n9896) );
  INV_X1 U7675 ( .A(n9691), .ZN(n9929) );
  XNOR2_X1 U7676 ( .A(n14981), .B(n14974), .ZN(n14980) );
  OAI21_X1 U7677 ( .B1(n15059), .B2(n7271), .A(n7270), .ZN(n15014) );
  INV_X1 U7678 ( .A(n7272), .ZN(n7271) );
  AOI21_X1 U7679 ( .B1(n7272), .B2(n10662), .A(n6538), .ZN(n7270) );
  NOR2_X1 U7680 ( .A1(n10650), .A2(n7273), .ZN(n7272) );
  NAND2_X1 U7681 ( .A1(n9941), .A2(n9940), .ZN(n15030) );
  NAND2_X1 U7682 ( .A1(n9916), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9927) );
  OR2_X1 U7683 ( .A1(n15099), .A2(n9935), .ZN(n15070) );
  NAND2_X1 U7684 ( .A1(n15112), .A2(n15396), .ZN(n15079) );
  NAND2_X1 U7685 ( .A1(n6675), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9907) );
  NAND2_X1 U7686 ( .A1(n11823), .A2(n9902), .ZN(n6638) );
  NOR2_X1 U7687 ( .A1(n7761), .A2(n15271), .ZN(n7760) );
  INV_X1 U7688 ( .A(n9632), .ZN(n9847) );
  NAND2_X2 U7689 ( .A1(n9986), .A2(n15436), .ZN(n9632) );
  NAND2_X1 U7690 ( .A1(n9587), .A2(n7705), .ZN(n7704) );
  NOR2_X1 U7691 ( .A1(n7703), .A2(n7706), .ZN(n6826) );
  INV_X1 U7692 ( .A(n7710), .ZN(n7705) );
  XNOR2_X1 U7693 ( .A(n6827), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9589) );
  XNOR2_X1 U7694 ( .A(n6637), .B(n8571), .ZN(n9620) );
  INV_X1 U7695 ( .A(n8570), .ZN(n6637) );
  NAND2_X1 U7696 ( .A1(n15490), .A2(n9611), .ZN(n9622) );
  NAND2_X1 U7697 ( .A1(n11944), .A2(n11945), .ZN(n7113) );
  INV_X1 U7698 ( .A(n13582), .ZN(n13551) );
  AND3_X1 U7699 ( .A1(n8313), .A2(n8312), .A3(n8311), .ZN(n13293) );
  NAND2_X1 U7700 ( .A1(n13192), .A2(n13193), .ZN(n7171) );
  NAND2_X1 U7701 ( .A1(n13869), .A2(n13868), .ZN(n13867) );
  NAND2_X1 U7702 ( .A1(n9286), .A2(n9285), .ZN(n14093) );
  NAND2_X1 U7703 ( .A1(n14682), .A2(n14681), .ZN(n14680) );
  NAND2_X1 U7704 ( .A1(n9949), .A2(n9948), .ZN(n14801) );
  NAND2_X1 U7705 ( .A1(n11312), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n11650) );
  NAND2_X1 U7706 ( .A1(n9362), .A2(n9361), .ZN(n6662) );
  NAND2_X1 U7707 ( .A1(n11484), .A2(n6665), .ZN(n6664) );
  OAI21_X1 U7708 ( .B1(n9356), .B2(n6665), .A(n11690), .ZN(n6663) );
  INV_X1 U7709 ( .A(n10495), .ZN(n7021) );
  INV_X1 U7710 ( .A(n9389), .ZN(n7366) );
  AND2_X1 U7711 ( .A1(n12724), .A2(n7364), .ZN(n7363) );
  NAND2_X1 U7712 ( .A1(n9392), .A2(n9389), .ZN(n7364) );
  INV_X1 U7713 ( .A(n9395), .ZN(n7362) );
  NAND2_X1 U7714 ( .A1(n6840), .A2(n7380), .ZN(n10510) );
  NAND2_X1 U7715 ( .A1(n10503), .A2(n10505), .ZN(n7380) );
  NOR2_X1 U7716 ( .A1(n6838), .A2(n10500), .ZN(n6839) );
  INV_X1 U7717 ( .A(n9402), .ZN(n7383) );
  NAND2_X1 U7718 ( .A1(n10513), .A2(n10515), .ZN(n7372) );
  NAND2_X1 U7719 ( .A1(n7017), .A2(n6511), .ZN(n7016) );
  INV_X1 U7720 ( .A(n10560), .ZN(n7017) );
  AND2_X1 U7721 ( .A1(n7019), .A2(n7018), .ZN(n10559) );
  AND2_X1 U7722 ( .A1(n6956), .A2(n9427), .ZN(n7359) );
  INV_X1 U7723 ( .A(n9425), .ZN(n6956) );
  NAND2_X1 U7724 ( .A1(n6955), .A2(n9425), .ZN(n7358) );
  INV_X1 U7725 ( .A(n9427), .ZN(n6955) );
  INV_X1 U7726 ( .A(n13129), .ZN(n6761) );
  INV_X1 U7727 ( .A(n9432), .ZN(n7099) );
  NOR2_X1 U7728 ( .A1(n7378), .A2(n10579), .ZN(n7379) );
  NAND2_X1 U7729 ( .A1(n7392), .A2(n10586), .ZN(n7391) );
  INV_X1 U7730 ( .A(n10585), .ZN(n7392) );
  INV_X1 U7731 ( .A(n6953), .ZN(n6952) );
  OAI21_X1 U7732 ( .B1(n7384), .B2(n6954), .A(n9451), .ZN(n6953) );
  NAND2_X1 U7733 ( .A1(n9447), .A2(n7385), .ZN(n7384) );
  MUX2_X1 U7734 ( .A(n13960), .B(n14352), .S(n9478), .Z(n9481) );
  OAI21_X1 U7735 ( .B1(n14352), .B2(n9497), .A(n7103), .ZN(n9482) );
  OR2_X1 U7736 ( .A1(n13960), .A2(n9473), .ZN(n7103) );
  NAND2_X1 U7737 ( .A1(n10472), .A2(n11890), .ZN(n7388) );
  NAND2_X1 U7738 ( .A1(n7158), .A2(n13172), .ZN(n7157) );
  AOI21_X1 U7739 ( .B1(n7037), .B2(n8489), .A(n13158), .ZN(n13162) );
  OAI21_X1 U7740 ( .B1(n13149), .B2(n6539), .A(n7038), .ZN(n7037) );
  NAND2_X1 U7741 ( .A1(n13147), .A2(n13145), .ZN(n7664) );
  INV_X1 U7742 ( .A(n8046), .ZN(n7596) );
  NAND2_X1 U7743 ( .A1(n7199), .A2(n8042), .ZN(n7198) );
  INV_X1 U7744 ( .A(n8330), .ZN(n7199) );
  NAND2_X1 U7745 ( .A1(n6603), .A2(n7200), .ZN(n7196) );
  INV_X1 U7746 ( .A(n8042), .ZN(n7200) );
  NOR2_X1 U7747 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n7813) );
  NOR2_X1 U7748 ( .A1(n14177), .A2(n7570), .ZN(n7569) );
  INV_X1 U7749 ( .A(n10421), .ZN(n7570) );
  AOI21_X1 U7750 ( .B1(n9745), .B2(n9619), .A(n7699), .ZN(n7698) );
  INV_X1 U7751 ( .A(n10287), .ZN(n7699) );
  INV_X1 U7752 ( .A(n9745), .ZN(n7700) );
  INV_X1 U7753 ( .A(n15111), .ZN(n7145) );
  NOR2_X1 U7754 ( .A1(n7462), .A2(n8860), .ZN(n7461) );
  INV_X1 U7755 ( .A(n7465), .ZN(n7462) );
  INV_X1 U7756 ( .A(n8788), .ZN(n8787) );
  INV_X1 U7757 ( .A(n6949), .ZN(n6948) );
  OAI21_X1 U7758 ( .B1(n7792), .B2(n6950), .A(n8749), .ZN(n6949) );
  INV_X1 U7759 ( .A(n8733), .ZN(n6950) );
  OAI21_X1 U7760 ( .B1(n8812), .B2(P2_DATAO_REG_14__SCAN_IN), .A(n6977), .ZN(
        n8692) );
  NAND2_X1 U7761 ( .A1(n8812), .A2(n11021), .ZN(n6977) );
  INV_X1 U7762 ( .A(n8598), .ZN(n8608) );
  NAND2_X1 U7763 ( .A1(n8601), .A2(SI_3_), .ZN(n8599) );
  NAND2_X1 U7764 ( .A1(n10818), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7020) );
  AND2_X1 U7765 ( .A1(n8070), .A2(n7230), .ZN(n7229) );
  INV_X1 U7766 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n7230) );
  INV_X1 U7767 ( .A(n8286), .ZN(n8071) );
  OAI21_X1 U7768 ( .B1(n11365), .B2(P3_REG1_REG_1__SCAN_IN), .A(n6993), .ZN(
        n7919) );
  NAND2_X1 U7769 ( .A1(n11365), .A2(n15689), .ZN(n6993) );
  INV_X1 U7770 ( .A(n11355), .ZN(n7314) );
  NAND2_X1 U7771 ( .A1(n6744), .A2(n6742), .ZN(n6746) );
  AND2_X1 U7772 ( .A1(n6743), .A2(n6568), .ZN(n6742) );
  AND2_X1 U7773 ( .A1(n6746), .A2(n11849), .ZN(n7989) );
  NAND2_X1 U7774 ( .A1(n7348), .A2(n7346), .ZN(n7992) );
  AND2_X1 U7775 ( .A1(n7347), .A2(n7774), .ZN(n7346) );
  NOR2_X1 U7776 ( .A1(n10713), .A2(n7057), .ZN(n7896) );
  AND2_X1 U7777 ( .A1(n10977), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7057) );
  OR2_X1 U7778 ( .A1(n8464), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9317) );
  AND2_X1 U7779 ( .A1(n7225), .A2(n8457), .ZN(n7671) );
  NAND2_X1 U7780 ( .A1(n7159), .A2(n13371), .ZN(n13163) );
  OR2_X1 U7781 ( .A1(n13675), .A2(n13570), .ZN(n13159) );
  NAND2_X1 U7782 ( .A1(n8074), .A2(n6622), .ZN(n8421) );
  INV_X1 U7783 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n7235) );
  OR2_X1 U7784 ( .A1(n13243), .A2(n13569), .ZN(n13151) );
  INV_X1 U7785 ( .A(n8385), .ZN(n8074) );
  NOR2_X1 U7786 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(P3_REG3_REG_8__SCAN_IN), 
        .ZN(n7227) );
  INV_X1 U7787 ( .A(n8197), .ZN(n8066) );
  OR2_X1 U7788 ( .A1(n13383), .A2(n8204), .ZN(n13090) );
  OR2_X1 U7789 ( .A1(n13385), .A2(n11731), .ZN(n13073) );
  NAND2_X1 U7790 ( .A1(n6974), .A2(n6973), .ZN(n13065) );
  NAND2_X1 U7791 ( .A1(n13191), .A2(n13054), .ZN(n13172) );
  AND2_X1 U7792 ( .A1(n13001), .A2(n13145), .ZN(n13144) );
  OR2_X1 U7793 ( .A1(n13768), .A2(n13251), .ZN(n13034) );
  OR2_X1 U7794 ( .A1(n13366), .A2(n13374), .ZN(n13135) );
  AND2_X1 U7795 ( .A1(n8247), .A2(n12076), .ZN(n8248) );
  NOR2_X1 U7796 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n7810) );
  AND2_X1 U7797 ( .A1(n7452), .A2(n7809), .ZN(n6771) );
  AND2_X1 U7798 ( .A1(n8462), .A2(n7806), .ZN(n7453) );
  NAND2_X1 U7799 ( .A1(n8268), .A2(n8029), .ZN(n8280) );
  NAND2_X1 U7800 ( .A1(n10812), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8007) );
  INV_X1 U7801 ( .A(n12136), .ZN(n7401) );
  INV_X1 U7802 ( .A(n9064), .ZN(n7402) );
  NOR2_X1 U7803 ( .A1(n9153), .A2(n7413), .ZN(n7412) );
  INV_X1 U7804 ( .A(n9129), .ZN(n7413) );
  INV_X1 U7805 ( .A(n7266), .ZN(n7265) );
  INV_X1 U7806 ( .A(n12398), .ZN(n7737) );
  NOR2_X1 U7807 ( .A1(n7738), .A2(n6906), .ZN(n6903) );
  AND2_X1 U7808 ( .A1(n10343), .A2(n10342), .ZN(n7738) );
  NOR2_X1 U7809 ( .A1(n6906), .A2(n10339), .ZN(n6904) );
  INV_X1 U7810 ( .A(n9032), .ZN(n8941) );
  NOR2_X1 U7811 ( .A1(n7563), .A2(n7560), .ZN(n7559) );
  INV_X1 U7812 ( .A(n10388), .ZN(n7560) );
  INV_X1 U7813 ( .A(n7559), .ZN(n6873) );
  NAND2_X1 U7814 ( .A1(n12049), .A2(n12053), .ZN(n12051) );
  NAND2_X1 U7815 ( .A1(n10453), .A2(n11815), .ZN(n10377) );
  OR2_X1 U7816 ( .A1(n10755), .A2(n10747), .ZN(n10749) );
  NAND2_X1 U7817 ( .A1(n9355), .A2(n11485), .ZN(n10754) );
  INV_X1 U7818 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8531) );
  INV_X1 U7819 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8532) );
  INV_X1 U7820 ( .A(n8619), .ZN(n8726) );
  INV_X1 U7821 ( .A(n10271), .ZN(n6943) );
  INV_X1 U7822 ( .A(n14970), .ZN(n6722) );
  OR2_X1 U7823 ( .A1(n14970), .A2(n7023), .ZN(n6721) );
  INV_X1 U7824 ( .A(n10021), .ZN(n7715) );
  NOR2_X1 U7825 ( .A1(n14803), .A2(n15404), .ZN(n7146) );
  AND2_X1 U7826 ( .A1(n9890), .A2(n7536), .ZN(n7535) );
  NAND2_X1 U7827 ( .A1(n9880), .A2(n7539), .ZN(n7536) );
  INV_X1 U7828 ( .A(n15158), .ZN(n10018) );
  OR2_X1 U7829 ( .A1(n15271), .A2(n15240), .ZN(n10530) );
  OR2_X1 U7830 ( .A1(n9785), .A2(n9784), .ZN(n9798) );
  AOI21_X1 U7831 ( .B1(n12710), .B2(n7719), .A(n6533), .ZN(n7718) );
  INV_X1 U7832 ( .A(n10007), .ZN(n7719) );
  NAND2_X1 U7833 ( .A1(n12430), .A2(n10006), .ZN(n6849) );
  INV_X1 U7834 ( .A(n10006), .ZN(n6850) );
  AOI21_X1 U7835 ( .B1(n11876), .B2(n7141), .A(n6523), .ZN(n7140) );
  INV_X1 U7836 ( .A(n9670), .ZN(n7141) );
  OR2_X1 U7837 ( .A1(n12028), .A2(n12024), .ZN(n9999) );
  NOR2_X1 U7838 ( .A1(n11876), .A2(n12028), .ZN(n10000) );
  NAND2_X1 U7839 ( .A1(n7712), .A2(n7711), .ZN(n15059) );
  AOI21_X1 U7840 ( .B1(n7713), .B2(n7716), .A(n6546), .ZN(n7711) );
  NAND2_X1 U7841 ( .A1(n15191), .A2(n7538), .ZN(n15120) );
  NAND2_X1 U7842 ( .A1(n15193), .A2(n15192), .ZN(n15191) );
  NOR2_X1 U7843 ( .A1(n7152), .A2(n15213), .ZN(n7150) );
  NAND2_X1 U7844 ( .A1(n6816), .A2(n6818), .ZN(n6814) );
  AND2_X1 U7845 ( .A1(n7153), .A2(n6811), .ZN(n6816) );
  NOR2_X1 U7846 ( .A1(n7531), .A2(n7154), .ZN(n7153) );
  NAND2_X1 U7847 ( .A1(n7520), .A2(n6817), .ZN(n6811) );
  INV_X1 U7848 ( .A(n10531), .ZN(n7154) );
  OR2_X1 U7849 ( .A1(n6818), .A2(n12559), .ZN(n6812) );
  INV_X1 U7850 ( .A(n10083), .ZN(n10645) );
  NAND2_X1 U7851 ( .A1(n7542), .A2(n7540), .ZN(n12149) );
  NOR2_X1 U7852 ( .A1(n12152), .A2(n7541), .ZN(n7540) );
  INV_X1 U7853 ( .A(n9697), .ZN(n7541) );
  NAND2_X1 U7854 ( .A1(n7709), .A2(n7708), .ZN(n7707) );
  INV_X1 U7855 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n7709) );
  INV_X1 U7856 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9574) );
  INV_X1 U7857 ( .A(n8816), .ZN(n7478) );
  AOI21_X1 U7858 ( .B1(n7474), .B2(n7477), .A(n7472), .ZN(n7471) );
  INV_X1 U7859 ( .A(n8791), .ZN(n7472) );
  NAND2_X1 U7860 ( .A1(n9586), .A2(n9792), .ZN(n9982) );
  OAI21_X1 U7861 ( .B1(n9979), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9973) );
  INV_X1 U7862 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9572) );
  NAND2_X1 U7863 ( .A1(n8734), .A2(n14461), .ZN(n8755) );
  NAND2_X1 U7864 ( .A1(n8722), .A2(n8706), .ZN(n8713) );
  NAND2_X1 U7865 ( .A1(n8692), .A2(n10975), .ZN(n8714) );
  XNOR2_X1 U7866 ( .A(n8657), .B(SI_10_), .ZN(n8654) );
  NAND2_X1 U7867 ( .A1(n6645), .A2(n6518), .ZN(n7015) );
  NAND2_X1 U7868 ( .A1(n8563), .A2(n8562), .ZN(n8570) );
  XNOR2_X1 U7869 ( .A(n10891), .B(n10800), .ZN(n10890) );
  NAND2_X1 U7870 ( .A1(n13260), .A2(n13237), .ZN(n7447) );
  INV_X1 U7871 ( .A(n13237), .ZN(n7444) );
  NAND2_X1 U7872 ( .A1(n7061), .A2(n13239), .ZN(n13307) );
  NAND2_X1 U7873 ( .A1(n13257), .A2(n7062), .ZN(n7061) );
  AND2_X1 U7874 ( .A1(n13238), .A2(n13237), .ZN(n7062) );
  OR2_X1 U7875 ( .A1(n7439), .A2(n6479), .ZN(n6444) );
  AND2_X1 U7876 ( .A1(n13247), .A2(n7428), .ZN(n7427) );
  OR2_X1 U7877 ( .A1(n13336), .A2(n7429), .ZN(n7428) );
  INV_X1 U7878 ( .A(n12908), .ZN(n7429) );
  OAI211_X1 U7879 ( .C1(n8346), .C2(n10838), .A(n8135), .B(n8134), .ZN(n11448)
         );
  AND2_X1 U7880 ( .A1(n12164), .A2(n12163), .ZN(n12342) );
  AND2_X1 U7881 ( .A1(n8355), .A2(n8354), .ZN(n13249) );
  OR2_X1 U7882 ( .A1(n8153), .A2(n8154), .ZN(n8155) );
  OR2_X1 U7883 ( .A1(n8138), .A2(n11366), .ZN(n8120) );
  NAND2_X1 U7884 ( .A1(n8113), .A2(n7974), .ZN(n7336) );
  OR2_X1 U7885 ( .A1(n11344), .A2(n7498), .ZN(n7496) );
  NAND2_X1 U7886 ( .A1(n7983), .A2(n6492), .ZN(n7330) );
  NAND2_X1 U7887 ( .A1(n11030), .A2(n6483), .ZN(n7328) );
  AND2_X1 U7888 ( .A1(n6647), .A2(n11356), .ZN(n10740) );
  NAND2_X1 U7889 ( .A1(n7942), .A2(n10820), .ZN(n6647) );
  NAND2_X1 U7890 ( .A1(n7312), .A2(n7314), .ZN(n7311) );
  NAND2_X1 U7891 ( .A1(n6646), .A2(n11356), .ZN(n7312) );
  NAND2_X1 U7892 ( .A1(n10740), .A2(n10741), .ZN(n6646) );
  AND3_X1 U7893 ( .A1(n7504), .A2(n7505), .A3(n7506), .ZN(n7876) );
  OAI21_X1 U7894 ( .B1(n7331), .B2(n7332), .A(n7323), .ZN(n7327) );
  NAND2_X1 U7895 ( .A1(n11030), .A2(n6525), .ZN(n7326) );
  AND2_X1 U7896 ( .A1(n7324), .A2(n11352), .ZN(n7323) );
  INV_X1 U7897 ( .A(n11521), .ZN(n7307) );
  AOI21_X1 U7898 ( .B1(n11214), .B2(n11036), .A(n11035), .ZN(n11038) );
  NAND2_X1 U7899 ( .A1(n7311), .A2(n7946), .ZN(n7309) );
  NAND2_X1 U7900 ( .A1(n11849), .A2(n7495), .ZN(n7491) );
  NOR2_X1 U7901 ( .A1(n11520), .A2(n6651), .ZN(n11843) );
  AND2_X1 U7902 ( .A1(n7948), .A2(n11529), .ZN(n6651) );
  NOR2_X1 U7903 ( .A1(n11843), .A2(n11844), .ZN(n11842) );
  NAND3_X1 U7904 ( .A1(n7486), .A2(P3_REG1_REG_9__SCAN_IN), .A3(n7487), .ZN(
        n13395) );
  NOR2_X1 U7905 ( .A1(n13387), .A2(n7302), .ZN(n12658) );
  AND2_X1 U7906 ( .A1(n7952), .A2(n13393), .ZN(n7302) );
  NAND3_X1 U7907 ( .A1(n6426), .A2(n7886), .A3(n6465), .ZN(n7512) );
  NAND2_X1 U7908 ( .A1(n7511), .A2(n13416), .ZN(n7510) );
  NOR2_X1 U7909 ( .A1(n13406), .A2(n7305), .ZN(n13427) );
  NOR2_X1 U7910 ( .A1(n7306), .A2(n13412), .ZN(n7305) );
  INV_X1 U7911 ( .A(n7954), .ZN(n7306) );
  NAND2_X1 U7912 ( .A1(n7992), .A2(n13430), .ZN(n10709) );
  NAND2_X1 U7913 ( .A1(n7003), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n13434) );
  INV_X1 U7914 ( .A(n13432), .ZN(n7003) );
  NAND2_X1 U7915 ( .A1(n13427), .A2(n13426), .ZN(n13425) );
  NAND2_X1 U7916 ( .A1(n7896), .A2(n7993), .ZN(n7517) );
  NAND2_X1 U7917 ( .A1(n7517), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7515) );
  NOR2_X1 U7918 ( .A1(n7896), .A2(n7993), .ZN(n13459) );
  NOR2_X1 U7919 ( .A1(n7093), .A2(n7515), .ZN(n13460) );
  NAND2_X1 U7920 ( .A1(n13466), .A2(n13465), .ZN(n13464) );
  NAND2_X1 U7921 ( .A1(n7997), .A2(n13485), .ZN(n13503) );
  NAND2_X1 U7922 ( .A1(n7485), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n13478) );
  NAND2_X1 U7923 ( .A1(n6779), .A2(n6778), .ZN(n7673) );
  AOI21_X1 U7924 ( .B1(n6780), .B2(n6782), .A(n7225), .ZN(n6778) );
  NAND2_X1 U7925 ( .A1(n13556), .A2(n6780), .ZN(n6779) );
  NAND2_X1 U7926 ( .A1(n7672), .A2(n7671), .ZN(n9302) );
  AND2_X1 U7927 ( .A1(n9302), .A2(n9301), .ZN(n13521) );
  AOI21_X1 U7928 ( .B1(n13163), .B2(n6781), .A(n7158), .ZN(n6780) );
  INV_X1 U7929 ( .A(n13160), .ZN(n6781) );
  INV_X1 U7930 ( .A(n13163), .ZN(n6782) );
  NAND2_X1 U7931 ( .A1(n13554), .A2(n8442), .ZN(n13540) );
  NAND2_X1 U7932 ( .A1(n8078), .A2(n8077), .ZN(n8447) );
  INV_X1 U7933 ( .A(n8434), .ZN(n8078) );
  NAND2_X1 U7934 ( .A1(n7215), .A2(n6452), .ZN(n7214) );
  INV_X1 U7935 ( .A(n8417), .ZN(n7646) );
  NAND2_X1 U7936 ( .A1(n8074), .A2(n7236), .ZN(n8408) );
  AOI21_X1 U7937 ( .B1(n7204), .B2(n7203), .A(n6555), .ZN(n7202) );
  INV_X1 U7938 ( .A(n7669), .ZN(n7203) );
  NAND2_X1 U7939 ( .A1(n6998), .A2(n13104), .ZN(n12070) );
  NAND2_X1 U7940 ( .A1(n13099), .A2(n13100), .ZN(n13015) );
  NAND2_X1 U7941 ( .A1(n11732), .A2(n8063), .ZN(n8167) );
  INV_X1 U7942 ( .A(n11554), .ZN(n11782) );
  AND2_X1 U7943 ( .A1(n13066), .A2(n13065), .ZN(n13007) );
  NAND2_X1 U7944 ( .A1(n13802), .A2(n12985), .ZN(n9307) );
  NAND2_X1 U7945 ( .A1(n8525), .A2(n8524), .ZN(n12933) );
  INV_X1 U7946 ( .A(n13144), .ZN(n13593) );
  AOI21_X1 U7947 ( .B1(n6437), .B2(n13005), .A(n6531), .ZN(n7648) );
  INV_X1 U7948 ( .A(n7655), .ZN(n7654) );
  OAI21_X1 U7949 ( .B1(n13611), .B2(n7658), .A(n13034), .ZN(n7655) );
  NAND2_X1 U7950 ( .A1(n7659), .A2(n13038), .ZN(n7658) );
  INV_X1 U7951 ( .A(n7660), .ZN(n7659) );
  NOR2_X1 U7952 ( .A1(n13006), .A2(n7653), .ZN(n7652) );
  INV_X1 U7953 ( .A(n8356), .ZN(n7653) );
  NOR2_X1 U7954 ( .A1(n13046), .A2(n7661), .ZN(n7660) );
  INV_X1 U7955 ( .A(n13043), .ZN(n7661) );
  NAND2_X1 U7956 ( .A1(n12758), .A2(n7667), .ZN(n8487) );
  AND2_X1 U7957 ( .A1(n13037), .A2(n13040), .ZN(n13653) );
  AND2_X1 U7958 ( .A1(n7638), .A2(n8482), .ZN(n7637) );
  NAND2_X1 U7959 ( .A1(n13018), .A2(n6506), .ZN(n7638) );
  AND2_X1 U7960 ( .A1(n8279), .A2(n8264), .ZN(n7665) );
  NAND2_X1 U7961 ( .A1(n7666), .A2(n8264), .ZN(n12205) );
  AND2_X1 U7962 ( .A1(n13117), .A2(n13118), .ZN(n13018) );
  NAND2_X1 U7963 ( .A1(n9551), .A2(n13000), .ZN(n13728) );
  OAI21_X1 U7964 ( .B1(n12874), .B2(n12873), .A(n12872), .ZN(n12948) );
  NAND2_X1 U7965 ( .A1(n7600), .A2(n7601), .ZN(n9311) );
  AOI21_X1 U7966 ( .B1(n7603), .B2(n7602), .A(n6625), .ZN(n7601) );
  NAND2_X1 U7967 ( .A1(n8081), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7915) );
  NAND2_X1 U7968 ( .A1(n6966), .A2(n6965), .ZN(n8081) );
  NAND2_X1 U7969 ( .A1(n7605), .A2(n8060), .ZN(n9304) );
  NAND2_X1 U7970 ( .A1(n7606), .A2(n6616), .ZN(n7605) );
  INV_X1 U7971 ( .A(n8444), .ZN(n7606) );
  NOR2_X1 U7972 ( .A1(n8392), .A2(n7194), .ZN(n7193) );
  INV_X1 U7973 ( .A(n8052), .ZN(n7194) );
  NAND2_X1 U7974 ( .A1(n8382), .A2(n8051), .ZN(n8053) );
  OAI21_X1 U7975 ( .B1(n8371), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n8049), .ZN(
        n8382) );
  INV_X1 U7976 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n6763) );
  NAND2_X1 U7977 ( .A1(n8048), .A2(n8049), .ZN(n8371) );
  OR2_X1 U7978 ( .A1(n8047), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8048) );
  INV_X1 U7979 ( .A(n7598), .ZN(n7597) );
  OAI21_X1 U7980 ( .B1(n8343), .B2(n7599), .A(n8358), .ZN(n7598) );
  INV_X1 U7981 ( .A(n8044), .ZN(n7599) );
  NAND2_X1 U7982 ( .A1(n8329), .A2(n8042), .ZN(n8344) );
  NAND2_X1 U7983 ( .A1(n7833), .A2(n7805), .ZN(n7449) );
  XNOR2_X1 U7984 ( .A(n7836), .B(P3_IR_REG_16__SCAN_IN), .ZN(n11017) );
  AOI21_X1 U7985 ( .B1(n7177), .B2(n7179), .A(n6560), .ZN(n7176) );
  INV_X1 U7986 ( .A(n8265), .ZN(n7177) );
  INV_X1 U7987 ( .A(n7179), .ZN(n7178) );
  OR2_X1 U7988 ( .A1(n8282), .A2(n11025), .ZN(n8295) );
  NAND2_X1 U7989 ( .A1(n8252), .A2(n8027), .ZN(n8266) );
  NAND2_X1 U7990 ( .A1(n8266), .A2(n8265), .ZN(n8268) );
  NAND2_X1 U7991 ( .A1(n8254), .A2(n8253), .ZN(n8252) );
  INV_X1 U7992 ( .A(n8023), .ZN(n7594) );
  AND2_X1 U7993 ( .A1(n8023), .A2(n8022), .ZN(n8210) );
  NAND2_X1 U7994 ( .A1(n7183), .A2(n7181), .ZN(n8211) );
  AOI21_X1 U7995 ( .B1(n7184), .B2(n7186), .A(n7182), .ZN(n7181) );
  INV_X1 U7996 ( .A(n8021), .ZN(n7182) );
  NAND2_X1 U7997 ( .A1(n8211), .A2(n8210), .ZN(n8209) );
  AND2_X1 U7998 ( .A1(n8021), .A2(n8020), .ZN(n8221) );
  NOR2_X1 U7999 ( .A1(n7851), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n7849) );
  NAND2_X1 U8000 ( .A1(n8019), .A2(n8017), .ZN(n8191) );
  NAND2_X1 U8001 ( .A1(n8016), .A2(n7614), .ZN(n8194) );
  NAND2_X1 U8002 ( .A1(n7585), .A2(n7583), .ZN(n8187) );
  AOI21_X1 U8003 ( .B1(n7586), .B2(n7588), .A(n7584), .ZN(n7583) );
  INV_X1 U8004 ( .A(n8013), .ZN(n7584) );
  NAND2_X1 U8005 ( .A1(n8131), .A2(n8007), .ZN(n8145) );
  NAND2_X1 U8006 ( .A1(n7135), .A2(n7133), .ZN(n12803) );
  NAND2_X1 U8007 ( .A1(n7395), .A2(n7397), .ZN(n7393) );
  NAND2_X1 U8008 ( .A1(n8947), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9220) );
  INV_X1 U8009 ( .A(n9207), .ZN(n8947) );
  OAI21_X1 U8010 ( .B1(n7130), .B2(n7416), .A(n7126), .ZN(n9214) );
  AOI21_X1 U8011 ( .B1(n7415), .B2(n7127), .A(n6559), .ZN(n7126) );
  INV_X1 U8012 ( .A(n7128), .ZN(n7127) );
  NAND2_X1 U8013 ( .A1(n8943), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9072) );
  INV_X1 U8014 ( .A(n9066), .ZN(n8943) );
  INV_X1 U8015 ( .A(n7412), .ZN(n7409) );
  INV_X1 U8016 ( .A(n13888), .ZN(n7414) );
  NAND2_X1 U8017 ( .A1(n13867), .A2(n7419), .ZN(n7418) );
  NOR2_X1 U8018 ( .A1(n13936), .A2(n9239), .ZN(n7419) );
  AOI211_X1 U8019 ( .C1(n9480), .C2(n9479), .A(n9494), .B(n9490), .ZN(n9502)
         );
  NAND2_X1 U8020 ( .A1(n8970), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8959) );
  OR2_X1 U8021 ( .A1(n8983), .A2(n11049), .ZN(n8958) );
  NOR3_X1 U8022 ( .A1(n13990), .A2(n11049), .A3(n13991), .ZN(n13989) );
  OR2_X1 U8023 ( .A1(n13989), .A2(n6705), .ZN(n6704) );
  NOR2_X1 U8024 ( .A1(n13983), .A2(n8964), .ZN(n6705) );
  AND2_X1 U8025 ( .A1(n6704), .A2(n6703), .ZN(n11072) );
  INV_X1 U8026 ( .A(n11050), .ZN(n6703) );
  AND2_X1 U8027 ( .A1(n11464), .A2(n11463), .ZN(n11466) );
  OAI22_X1 U8028 ( .A1(n15578), .A2(n15577), .B1(n15580), .B2(
        P2_REG1_REG_12__SCAN_IN), .ZN(n15598) );
  INV_X1 U8029 ( .A(n12457), .ZN(n15586) );
  OR2_X1 U8030 ( .A1(n14046), .A2(n14062), .ZN(n14065) );
  AND2_X1 U8031 ( .A1(n7610), .A2(n7609), .ZN(n7608) );
  INV_X1 U8032 ( .A(n10427), .ZN(n6880) );
  AOI21_X1 U8033 ( .B1(n6918), .B2(n6916), .A(n6915), .ZN(n6914) );
  INV_X1 U8034 ( .A(n6918), .ZN(n6917) );
  INV_X1 U8035 ( .A(n10357), .ZN(n6916) );
  NAND2_X1 U8036 ( .A1(n6875), .A2(n6874), .ZN(n14187) );
  NAND2_X1 U8037 ( .A1(n6877), .A2(n6544), .ZN(n6874) );
  NAND2_X1 U8038 ( .A1(n14246), .A2(n7550), .ZN(n14221) );
  OAI21_X1 U8039 ( .B1(n14258), .B2(n14261), .A(n10357), .ZN(n14213) );
  NOR3_X1 U8040 ( .A1(n14298), .A2(n14537), .A3(n14275), .ZN(n14252) );
  NAND2_X1 U8041 ( .A1(n6907), .A2(n6911), .ZN(n10352) );
  AND2_X1 U8042 ( .A1(n12813), .A2(n6912), .ZN(n6911) );
  NAND2_X1 U8043 ( .A1(n12669), .A2(n10350), .ZN(n6912) );
  INV_X1 U8044 ( .A(n10350), .ZN(n6913) );
  INV_X1 U8045 ( .A(n10408), .ZN(n7577) );
  NAND2_X1 U8046 ( .A1(n12574), .A2(n10407), .ZN(n7578) );
  NAND2_X1 U8047 ( .A1(n10349), .A2(n10348), .ZN(n12670) );
  NAND2_X1 U8048 ( .A1(n6486), .A2(n6798), .ZN(n12817) );
  NOR3_X1 U8049 ( .A1(n12401), .A2(n12409), .A3(n12678), .ZN(n6798) );
  AND2_X1 U8050 ( .A1(n7561), .A2(n6871), .ZN(n6870) );
  INV_X1 U8051 ( .A(n7562), .ZN(n7561) );
  NAND2_X1 U8052 ( .A1(n7559), .A2(n6872), .ZN(n6871) );
  OAI21_X1 U8053 ( .B1(n11911), .B2(n7563), .A(n10390), .ZN(n7562) );
  OR2_X1 U8054 ( .A1(n11932), .A2(n6873), .ZN(n6869) );
  NAND2_X1 U8055 ( .A1(n11930), .A2(n10388), .ZN(n11912) );
  NAND2_X1 U8056 ( .A1(n11911), .A2(n11912), .ZN(n12054) );
  OAI211_X1 U8057 ( .C1(n6901), .C2(n6872), .A(n6898), .B(n11908), .ZN(n11907)
         );
  NOR2_X1 U8058 ( .A1(n6901), .A2(n6900), .ZN(n6899) );
  INV_X1 U8059 ( .A(n10336), .ZN(n6900) );
  NAND2_X1 U8060 ( .A1(n11707), .A2(n10336), .ZN(n11927) );
  NAND2_X1 U8061 ( .A1(n11927), .A2(n6872), .ZN(n11928) );
  AND2_X1 U8062 ( .A1(n9288), .A2(n9287), .ZN(n14285) );
  NAND2_X1 U8063 ( .A1(n13856), .A2(n11485), .ZN(n10747) );
  OR2_X1 U8064 ( .A1(n9464), .A2(n13980), .ZN(n8966) );
  INV_X1 U8065 ( .A(n14286), .ZN(n14192) );
  NAND2_X1 U8066 ( .A1(n14643), .A2(n8834), .ZN(n8836) );
  NAND2_X1 U8067 ( .A1(n8814), .A2(n8813), .ZN(n14149) );
  NAND2_X1 U8068 ( .A1(n8794), .A2(n8793), .ZN(n14180) );
  AND2_X1 U8069 ( .A1(n10707), .A2(n10706), .ZN(n9293) );
  AND2_X1 U8070 ( .A1(n7580), .A2(n8887), .ZN(n7579) );
  INV_X1 U8071 ( .A(n7582), .ZN(n7580) );
  INV_X1 U8072 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8541) );
  NAND2_X1 U8073 ( .A1(n7423), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8883) );
  OR2_X1 U8074 ( .A1(n8672), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8680) );
  AND2_X1 U8075 ( .A1(n14774), .A2(n7685), .ZN(n7684) );
  OR2_X1 U8076 ( .A1(n14700), .A2(n7686), .ZN(n7685) );
  INV_X1 U8077 ( .A(n10278), .ZN(n7686) );
  AND2_X1 U8078 ( .A1(n7684), .A2(n6942), .ZN(n6941) );
  OR2_X1 U8079 ( .A1(n14722), .A2(n6943), .ZN(n6942) );
  NAND2_X1 U8080 ( .A1(n6941), .A2(n6943), .ZN(n6939) );
  AND2_X1 U8081 ( .A1(n10199), .A2(n14650), .ZN(n7691) );
  OR2_X1 U8082 ( .A1(n12583), .A2(n10181), .ZN(n7696) );
  AND2_X1 U8083 ( .A1(n6570), .A2(n10159), .ZN(n7693) );
  OAI21_X1 U8084 ( .B1(n10105), .B2(n11156), .A(n10086), .ZN(n11146) );
  INV_X1 U8085 ( .A(n9870), .ZN(n9861) );
  AND2_X1 U8086 ( .A1(n14733), .A2(n14734), .ZN(n14731) );
  INV_X1 U8087 ( .A(n10240), .ZN(n6932) );
  NAND2_X1 U8088 ( .A1(n14689), .A2(n7690), .ZN(n7689) );
  INV_X1 U8089 ( .A(n10247), .ZN(n7690) );
  NAND2_X2 U8090 ( .A1(n10084), .A2(n10645), .ZN(n10299) );
  NAND2_X1 U8091 ( .A1(n10627), .A2(n6834), .ZN(n6833) );
  NAND2_X1 U8092 ( .A1(n10627), .A2(n6836), .ZN(n6835) );
  NAND2_X1 U8093 ( .A1(n10612), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9618) );
  OR2_X1 U8094 ( .A1(n6429), .A2(n14822), .ZN(n9608) );
  AND2_X1 U8095 ( .A1(n15505), .A2(n10920), .ZN(n14877) );
  INV_X1 U8096 ( .A(n7058), .ZN(n14941) );
  XNOR2_X1 U8097 ( .A(n10626), .B(n10625), .ZN(n10665) );
  NAND2_X1 U8098 ( .A1(n15298), .A2(n14724), .ZN(n15048) );
  NAND2_X1 U8099 ( .A1(n15093), .A2(n15092), .ZN(n15091) );
  INV_X1 U8100 ( .A(n7146), .ZN(n9891) );
  INV_X1 U8101 ( .A(n6675), .ZN(n9884) );
  OR2_X1 U8102 ( .A1(n15125), .A2(n15124), .ZN(n6823) );
  NAND2_X1 U8103 ( .A1(n7147), .A2(n7535), .ZN(n15123) );
  NAND2_X1 U8104 ( .A1(n15193), .A2(n7148), .ZN(n7147) );
  NAND2_X1 U8105 ( .A1(n7281), .A2(n10016), .ZN(n15156) );
  OR2_X1 U8106 ( .A1(n15178), .A2(n7736), .ZN(n7281) );
  INV_X1 U8107 ( .A(n7278), .ZN(n7280) );
  NAND2_X1 U8108 ( .A1(n9829), .A2(n9828), .ZN(n15199) );
  NOR2_X1 U8109 ( .A1(n15236), .A2(n7533), .ZN(n7532) );
  INV_X1 U8110 ( .A(n10530), .ZN(n7533) );
  NAND2_X1 U8111 ( .A1(n15263), .A2(n15262), .ZN(n15261) );
  NAND2_X1 U8112 ( .A1(n12767), .A2(n10531), .ZN(n15263) );
  AOI21_X1 U8113 ( .B1(n7733), .B2(n7735), .A(n6535), .ZN(n7732) );
  AND2_X1 U8114 ( .A1(n7734), .A2(n12332), .ZN(n7733) );
  OR2_X1 U8115 ( .A1(n12189), .A2(n7735), .ZN(n7734) );
  INV_X1 U8116 ( .A(n10005), .ZN(n7735) );
  NAND2_X1 U8117 ( .A1(n12188), .A2(n12189), .ZN(n12187) );
  NAND2_X1 U8118 ( .A1(n12149), .A2(n6824), .ZN(n12192) );
  NOR2_X1 U8119 ( .A1(n12189), .A2(n6825), .ZN(n6824) );
  INV_X1 U8120 ( .A(n9713), .ZN(n6825) );
  NAND2_X1 U8121 ( .A1(n7051), .A2(n7050), .ZN(n12334) );
  NAND2_X1 U8122 ( .A1(n7701), .A2(n10003), .ZN(n12146) );
  NAND3_X1 U8123 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n9673) );
  NAND2_X1 U8124 ( .A1(n6845), .A2(n9996), .ZN(n11507) );
  INV_X1 U8125 ( .A(n10488), .ZN(n9612) );
  INV_X1 U8126 ( .A(n15241), .ZN(n15258) );
  AND2_X1 U8127 ( .A1(n13200), .A2(n13203), .ZN(n10038) );
  NAND2_X1 U8128 ( .A1(n9850), .A2(n9849), .ZN(n15332) );
  NAND2_X1 U8129 ( .A1(n9783), .A2(n9782), .ZN(n12770) );
  NAND2_X1 U8130 ( .A1(n10982), .A2(n9902), .ZN(n6716) );
  NAND2_X1 U8131 ( .A1(n7463), .A2(n7465), .ZN(n8861) );
  XNOR2_X1 U8132 ( .A(n8826), .B(n8825), .ZN(n12241) );
  AND2_X1 U8133 ( .A1(n14416), .A2(n10047), .ZN(n7248) );
  XNOR2_X1 U8134 ( .A(n8815), .B(n8816), .ZN(n12108) );
  NAND2_X1 U8135 ( .A1(n7467), .A2(n7471), .ZN(n8803) );
  OR2_X1 U8136 ( .A1(n8773), .A2(n7473), .ZN(n7467) );
  XNOR2_X1 U8137 ( .A(n8803), .B(n8804), .ZN(n9882) );
  XNOR2_X1 U8138 ( .A(n8678), .B(n8688), .ZN(n11024) );
  AOI21_X1 U8139 ( .B1(n7285), .B2(n6431), .A(n7284), .ZN(n7283) );
  AND2_X1 U8140 ( .A1(n9771), .A2(n9780), .ZN(n11663) );
  NAND2_X1 U8141 ( .A1(n7480), .A2(n8626), .ZN(n8635) );
  INV_X1 U8142 ( .A(n8624), .ZN(n6957) );
  NAND2_X1 U8143 ( .A1(n10769), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n6897) );
  NAND2_X1 U8144 ( .A1(n10896), .A2(n6448), .ZN(n6884) );
  OR2_X1 U8145 ( .A1(n10993), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6885) );
  NOR2_X1 U8146 ( .A1(n11944), .A2(n11945), .ZN(n7112) );
  NOR2_X1 U8147 ( .A1(n7112), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7111) );
  NAND2_X1 U8148 ( .A1(n7294), .A2(n15451), .ZN(n7293) );
  NAND2_X1 U8149 ( .A1(n6961), .A2(n6960), .ZN(n11379) );
  NAND2_X1 U8150 ( .A1(n13064), .A2(n12935), .ZN(n6960) );
  INV_X1 U8151 ( .A(n13604), .ZN(n13263) );
  AOI21_X1 U8152 ( .B1(n7434), .B2(n7432), .A(n6505), .ZN(n7431) );
  INV_X1 U8153 ( .A(n7434), .ZN(n7433) );
  NOR2_X1 U8154 ( .A1(n11781), .A2(n11780), .ZN(n12161) );
  NAND2_X1 U8155 ( .A1(n11581), .A2(n13385), .ZN(n11582) );
  NAND2_X1 U8156 ( .A1(n11553), .A2(n11552), .ZN(n11583) );
  NAND2_X1 U8157 ( .A1(n11179), .A2(n11178), .ZN(n13362) );
  NAND2_X1 U8158 ( .A1(n6769), .A2(n6768), .ZN(n6770) );
  AOI21_X1 U8159 ( .B1(n6436), .B2(n6458), .A(n6566), .ZN(n6768) );
  NOR2_X1 U8160 ( .A1(n7170), .A2(n13000), .ZN(n7167) );
  AOI21_X1 U8161 ( .B1(n13179), .B2(n13178), .A(n7034), .ZN(n13182) );
  NAND2_X1 U8162 ( .A1(n7036), .A2(n7035), .ZN(n7034) );
  NAND2_X1 U8163 ( .A1(n7161), .A2(n7160), .ZN(n13179) );
  AOI21_X1 U8164 ( .B1(n6504), .B2(n7169), .A(n7168), .ZN(n7166) );
  NOR2_X1 U8165 ( .A1(n7170), .A2(n13186), .ZN(n7169) );
  NOR2_X1 U8166 ( .A1(n7170), .A2(n13192), .ZN(n7168) );
  NAND2_X1 U8167 ( .A1(n12883), .A2(n9324), .ZN(n13522) );
  NAND2_X1 U8168 ( .A1(n8093), .A2(n8092), .ZN(n13542) );
  NAND2_X1 U8169 ( .A1(n13531), .A2(n9318), .ZN(n8093) );
  NAND2_X1 U8170 ( .A1(n8428), .A2(n8427), .ZN(n13582) );
  INV_X1 U8171 ( .A(n13251), .ZN(n13623) );
  INV_X1 U8172 ( .A(n13249), .ZN(n13655) );
  NAND2_X1 U8173 ( .A1(n8327), .A2(n8326), .ZN(n13654) );
  NAND2_X1 U8174 ( .A1(n7991), .A2(n7349), .ZN(n12661) );
  NOR2_X1 U8175 ( .A1(n10719), .A2(n10720), .ZN(n10718) );
  NOR2_X1 U8176 ( .A1(n7994), .A2(n7993), .ZN(n13455) );
  OR2_X1 U8177 ( .A1(n13476), .A2(n13657), .ZN(n13474) );
  XNOR2_X1 U8178 ( .A(n7907), .B(n7962), .ZN(n7499) );
  NOR2_X1 U8179 ( .A1(n13511), .A2(n6454), .ZN(n7965) );
  NAND2_X1 U8180 ( .A1(n6749), .A2(n6632), .ZN(n7316) );
  AND2_X1 U8181 ( .A1(n8002), .A2(n8001), .ZN(n13504) );
  OR2_X1 U8182 ( .A1(n8474), .A2(n13638), .ZN(n7044) );
  NAND2_X1 U8183 ( .A1(n8348), .A2(n8347), .ZN(n13702) );
  OR2_X1 U8184 ( .A1(n11221), .A2(n8346), .ZN(n8348) );
  INV_X1 U8185 ( .A(n6790), .ZN(n6789) );
  OAI21_X1 U8186 ( .B1(n8346), .B2(n10866), .A(n8163), .ZN(n6790) );
  OR2_X1 U8187 ( .A1(n11989), .A2(n15715), .ZN(n13588) );
  INV_X1 U8188 ( .A(n12933), .ZN(n13744) );
  OR2_X1 U8189 ( .A1(n11435), .A2(n8346), .ZN(n8363) );
  NAND2_X1 U8190 ( .A1(n8299), .A2(n8298), .ZN(n13236) );
  NAND2_X1 U8191 ( .A1(n8239), .A2(n8238), .ZN(n13110) );
  OR2_X1 U8192 ( .A1(n15721), .A2(n15715), .ZN(n13790) );
  OAI21_X1 U8193 ( .B1(n8160), .B2(n7588), .A(n7586), .ZN(n8176) );
  NAND2_X1 U8194 ( .A1(n8162), .A2(n8011), .ZN(n8174) );
  NAND2_X1 U8195 ( .A1(n12045), .A2(n8834), .ZN(n8800) );
  NAND2_X1 U8196 ( .A1(n6799), .A2(n6803), .ZN(n13835) );
  OR2_X1 U8197 ( .A1(n13926), .A2(n13927), .ZN(n6799) );
  NAND2_X1 U8198 ( .A1(n8771), .A2(n8770), .ZN(n14232) );
  NAND2_X1 U8199 ( .A1(n12890), .A2(n8592), .ZN(n8841) );
  NAND2_X1 U8200 ( .A1(n7418), .A2(n6805), .ZN(n13854) );
  AND2_X1 U8201 ( .A1(n9270), .A2(n6498), .ZN(n6805) );
  AND2_X1 U8202 ( .A1(n7621), .A2(n6569), .ZN(n7619) );
  NAND2_X1 U8203 ( .A1(n11042), .A2(n7620), .ZN(n7621) );
  NAND2_X1 U8204 ( .A1(n13896), .A2(n9230), .ZN(n13869) );
  OAI211_X1 U8205 ( .C1(n13860), .C2(n8991), .A(n8990), .B(n13825), .ZN(n7405)
         );
  AOI21_X1 U8206 ( .B1(n11471), .B2(n11473), .A(n13822), .ZN(n8990) );
  AOI21_X1 U8207 ( .B1(n8768), .B2(n14000), .A(n6456), .ZN(n8586) );
  NAND2_X1 U8208 ( .A1(n11774), .A2(n8834), .ZN(n7250) );
  NAND2_X1 U8209 ( .A1(n8665), .A2(n8664), .ZN(n14571) );
  NAND2_X1 U8210 ( .A1(n12543), .A2(n8834), .ZN(n8829) );
  NAND2_X1 U8211 ( .A1(n8721), .A2(n8720), .ZN(n14313) );
  NAND2_X1 U8212 ( .A1(n9265), .A2(n9264), .ZN(n13961) );
  NAND2_X1 U8213 ( .A1(n6695), .A2(n9250), .ZN(n14125) );
  NAND2_X1 U8214 ( .A1(n14114), .A2(n9258), .ZN(n6695) );
  OR2_X1 U8215 ( .A1(n14150), .A2(n9464), .ZN(n9226) );
  OR2_X1 U8216 ( .A1(n9135), .A2(n9134), .ZN(n13966) );
  OAI21_X1 U8217 ( .B1(n6476), .B2(n14006), .A(n11074), .ZN(n14009) );
  AOI21_X1 U8218 ( .B1(n14009), .B2(n11133), .A(n11132), .ZN(n14019) );
  NOR2_X1 U8219 ( .A1(n11418), .A2(n7082), .ZN(n11459) );
  OR2_X1 U8220 ( .A1(n11420), .A2(n11417), .ZN(n7082) );
  NOR2_X1 U8221 ( .A1(n11459), .A2(n7081), .ZN(n12465) );
  AND2_X1 U8222 ( .A1(n11462), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7081) );
  NAND2_X1 U8223 ( .A1(n6984), .A2(n9170), .ZN(n14066) );
  INV_X1 U8224 ( .A(n14049), .ZN(n6984) );
  XNOR2_X1 U8225 ( .A(n10447), .B(n10446), .ZN(n14355) );
  INV_X1 U8226 ( .A(n10456), .ZN(n10446) );
  AOI21_X1 U8227 ( .B1(n6472), .B2(n7258), .A(n7254), .ZN(n7253) );
  AOI21_X1 U8228 ( .B1(n14351), .B2(n14344), .A(n10467), .ZN(n10468) );
  NAND2_X1 U8229 ( .A1(n10437), .A2(n13847), .ZN(n14085) );
  OR2_X1 U8230 ( .A1(n10434), .A2(n10455), .ZN(n10437) );
  OAI21_X1 U8231 ( .B1(n14107), .B2(n7556), .A(n7552), .ZN(n10433) );
  OAI21_X1 U8232 ( .B1(n7747), .B2(n7258), .A(n6472), .ZN(n10445) );
  NAND2_X1 U8233 ( .A1(n14103), .A2(n7053), .ZN(n10376) );
  NOR2_X1 U8234 ( .A1(n10375), .A2(n7258), .ZN(n7053) );
  INV_X1 U8235 ( .A(n14356), .ZN(n14099) );
  NAND2_X1 U8236 ( .A1(n8698), .A2(n8697), .ZN(n14562) );
  OR2_X1 U8237 ( .A1(n14312), .A2(n10454), .ZN(n14346) );
  INV_X1 U8238 ( .A(n15627), .ZN(n14344) );
  INV_X1 U8239 ( .A(n14346), .ZN(n15630) );
  OR2_X1 U8240 ( .A1(n8866), .A2(n10812), .ZN(n8564) );
  OR2_X1 U8241 ( .A1(n14341), .A2(n14070), .ZN(n15627) );
  AOI21_X1 U8242 ( .B1(n7545), .B2(n14339), .A(n6614), .ZN(n14354) );
  INV_X1 U8243 ( .A(n14353), .ZN(n6992) );
  AOI21_X1 U8244 ( .B1(n6457), .B2(n14579), .A(n6428), .ZN(n10441) );
  INV_X1 U8245 ( .A(n14089), .ZN(n6922) );
  NAND2_X1 U8246 ( .A1(n6680), .A2(n9689), .ZN(n9690) );
  AND2_X1 U8247 ( .A1(n9964), .A2(n9963), .ZN(n12964) );
  OR2_X1 U8248 ( .A1(n10313), .A2(n6429), .ZN(n9964) );
  NAND2_X2 U8249 ( .A1(n9893), .A2(n9892), .ZN(n15113) );
  NAND2_X1 U8250 ( .A1(n12045), .A2(n9902), .ZN(n9893) );
  NOR2_X1 U8251 ( .A1(n7677), .A2(n7676), .ZN(n7675) );
  NAND2_X1 U8252 ( .A1(n12890), .A2(n9902), .ZN(n9952) );
  AOI21_X1 U8253 ( .B1(n11901), .B2(n6934), .A(n6537), .ZN(n6933) );
  INV_X1 U8254 ( .A(n11901), .ZN(n6935) );
  NAND2_X1 U8255 ( .A1(n9806), .A2(n9805), .ZN(n15351) );
  INV_X1 U8256 ( .A(n10096), .ZN(n9991) );
  INV_X1 U8257 ( .A(n14812), .ZN(n12590) );
  AND2_X1 U8258 ( .A1(n10312), .A2(n11490), .ZN(n14766) );
  NAND2_X1 U8259 ( .A1(n6641), .A2(n10278), .ZN(n7240) );
  NAND2_X1 U8260 ( .A1(n14699), .A2(n14700), .ZN(n6641) );
  INV_X1 U8261 ( .A(n14774), .ZN(n7239) );
  NAND2_X1 U8262 ( .A1(n12543), .A2(n9902), .ZN(n9925) );
  INV_X1 U8263 ( .A(n15256), .ZN(n14788) );
  NAND2_X1 U8264 ( .A1(n9913), .A2(n9912), .ZN(n14802) );
  OR2_X1 U8265 ( .A1(n15100), .A2(n6429), .ZN(n9913) );
  NAND2_X1 U8266 ( .A1(n9899), .A2(n9898), .ZN(n15089) );
  OAI211_X1 U8267 ( .C1(n14828), .C2(n10912), .A(n10913), .B(n7029), .ZN(
        n14831) );
  NAND2_X1 U8268 ( .A1(n14828), .A2(n10912), .ZN(n7029) );
  NAND2_X1 U8269 ( .A1(n6728), .A2(n10924), .ZN(n14910) );
  NAND2_X1 U8270 ( .A1(n14908), .A2(n14907), .ZN(n6728) );
  OR2_X1 U8271 ( .A1(n14917), .A2(n14918), .ZN(n6734) );
  AND2_X1 U8272 ( .A1(n6733), .A2(n6732), .ZN(n11264) );
  NOR2_X1 U8273 ( .A1(n11000), .A2(n11002), .ZN(n6732) );
  XNOR2_X1 U8274 ( .A(n7090), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14992) );
  NAND2_X1 U8275 ( .A1(n7092), .A2(n7091), .ZN(n7090) );
  NAND2_X1 U8276 ( .A1(n14980), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7092) );
  OAI21_X1 U8277 ( .B1(n15019), .B2(n15160), .A(n15018), .ZN(n15285) );
  XNOR2_X1 U8278 ( .A(n6682), .B(n15017), .ZN(n15019) );
  AOI21_X1 U8279 ( .B1(n15030), .B2(n10650), .A(n6517), .ZN(n6682) );
  AND2_X1 U8280 ( .A1(n15016), .A2(n15015), .ZN(n15284) );
  NAND2_X1 U8281 ( .A1(n15014), .A2(n15017), .ZN(n15015) );
  NAND2_X1 U8282 ( .A1(n7730), .A2(n7729), .ZN(n15016) );
  NAND2_X1 U8283 ( .A1(n7071), .A2(n7072), .ZN(n15040) );
  NAND2_X1 U8284 ( .A1(n15036), .A2(n10650), .ZN(n7071) );
  AND2_X1 U8285 ( .A1(n9957), .A2(n9928), .ZN(n15052) );
  NAND2_X1 U8286 ( .A1(n6852), .A2(n6851), .ZN(n15129) );
  AND2_X1 U8287 ( .A1(n6821), .A2(n6820), .ZN(n15315) );
  INV_X1 U8288 ( .A(n15126), .ZN(n6820) );
  NAND2_X1 U8289 ( .A1(n6822), .A2(n15260), .ZN(n6821) );
  NAND2_X1 U8290 ( .A1(n6823), .A2(n15123), .ZN(n6822) );
  NAND2_X1 U8291 ( .A1(n14643), .A2(n9902), .ZN(n9943) );
  OR2_X1 U8292 ( .A1(n10076), .A2(n15549), .ZN(n10069) );
  AND2_X1 U8293 ( .A1(n15040), .A2(n6861), .ZN(n15384) );
  NOR2_X1 U8294 ( .A1(n15289), .A2(n7137), .ZN(n6861) );
  INV_X1 U8295 ( .A(n15039), .ZN(n7137) );
  AOI22_X1 U8296 ( .A1(n9848), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n15507), .B2(
        n9847), .ZN(n7519) );
  AND2_X1 U8297 ( .A1(n6864), .A2(n6863), .ZN(n6936) );
  OR2_X1 U8298 ( .A1(n9619), .A2(n10875), .ZN(n6937) );
  NAND2_X1 U8299 ( .A1(n9632), .A2(n6449), .ZN(n6864) );
  NOR2_X1 U8300 ( .A1(n9843), .A2(n9842), .ZN(n9846) );
  NAND2_X1 U8301 ( .A1(n10896), .A2(n10895), .ZN(n10994) );
  NAND2_X1 U8302 ( .A1(n11650), .A2(n11649), .ZN(n11793) );
  NAND2_X1 U8303 ( .A1(n11650), .A2(n6894), .ZN(n11794) );
  NOR2_X1 U8304 ( .A1(n6895), .A2(n11792), .ZN(n6894) );
  INV_X1 U8305 ( .A(n11649), .ZN(n6895) );
  XNOR2_X1 U8306 ( .A(n12498), .B(n12496), .ZN(n12495) );
  INV_X1 U8307 ( .A(n6889), .ZN(n6887) );
  NOR2_X1 U8308 ( .A1(n10330), .A2(n9401), .ZN(n6665) );
  INV_X1 U8309 ( .A(n10493), .ZN(n10494) );
  OAI21_X1 U8310 ( .B1(n6434), .B2(n11865), .A(n6985), .ZN(n10492) );
  NAND2_X1 U8311 ( .A1(n6434), .A2(n11830), .ZN(n6985) );
  NAND2_X1 U8312 ( .A1(n6670), .A2(n9372), .ZN(n6667) );
  OAI21_X1 U8313 ( .B1(n6670), .B2(n9372), .A(n11911), .ZN(n6669) );
  AND2_X1 U8314 ( .A1(n9375), .A2(n10390), .ZN(n9376) );
  NAND2_X1 U8315 ( .A1(n10498), .A2(n7370), .ZN(n7369) );
  AOI21_X1 U8316 ( .B1(n10496), .B2(n10497), .A(n7021), .ZN(n7368) );
  NAND2_X1 U8317 ( .A1(n6838), .A2(n10500), .ZN(n6837) );
  AOI21_X1 U8318 ( .B1(n13071), .B2(n13070), .A(n13069), .ZN(n13081) );
  NAND2_X1 U8319 ( .A1(n7360), .A2(n7361), .ZN(n6658) );
  AOI21_X1 U8320 ( .B1(n7363), .B2(n7365), .A(n7362), .ZN(n7361) );
  AND2_X1 U8321 ( .A1(n9391), .A2(n7366), .ZN(n7365) );
  INV_X1 U8322 ( .A(n10509), .ZN(n7010) );
  NOR2_X1 U8323 ( .A1(n10541), .A2(n7799), .ZN(n10542) );
  AND2_X1 U8324 ( .A1(n10559), .A2(n7016), .ZN(n7087) );
  OAI211_X1 U8325 ( .C1(n13125), .C2(n6760), .A(n13130), .B(n6759), .ZN(n6762)
         );
  OR2_X1 U8326 ( .A1(n6761), .A2(n13126), .ZN(n6760) );
  OR2_X1 U8327 ( .A1(n6576), .A2(n6761), .ZN(n6759) );
  NAND2_X1 U8328 ( .A1(n9431), .A2(n7099), .ZN(n7098) );
  NAND2_X1 U8329 ( .A1(n9430), .A2(n6677), .ZN(n6676) );
  NAND2_X1 U8330 ( .A1(n7390), .A2(n10585), .ZN(n7389) );
  INV_X1 U8331 ( .A(n10586), .ZN(n7390) );
  NAND2_X1 U8332 ( .A1(n6758), .A2(n6757), .ZN(n6756) );
  INV_X1 U8333 ( .A(n13140), .ZN(n6757) );
  INV_X1 U8334 ( .A(n13141), .ZN(n7067) );
  INV_X1 U8335 ( .A(n13142), .ZN(n7066) );
  NAND2_X1 U8336 ( .A1(n6661), .A2(n6660), .ZN(n9446) );
  NAND2_X1 U8337 ( .A1(n9441), .A2(n9443), .ZN(n6660) );
  AOI21_X1 U8338 ( .B1(n6755), .B2(n7065), .A(n6754), .ZN(n13149) );
  NOR2_X1 U8339 ( .A1(n13024), .A2(n7066), .ZN(n7065) );
  NAND2_X1 U8340 ( .A1(n13144), .A2(n13143), .ZN(n6754) );
  NAND2_X1 U8341 ( .A1(n6756), .A2(n6532), .ZN(n6755) );
  NAND2_X1 U8342 ( .A1(n13243), .A2(n7039), .ZN(n7038) );
  NOR2_X1 U8343 ( .A1(n13595), .A2(n13172), .ZN(n7039) );
  AND2_X1 U8344 ( .A1(n6587), .A2(n6830), .ZN(n6829) );
  NAND2_X1 U8345 ( .A1(n10595), .A2(n10598), .ZN(n6830) );
  AOI21_X1 U8346 ( .B1(n7471), .B2(n7473), .A(n7469), .ZN(n7468) );
  INV_X1 U8347 ( .A(n8802), .ZN(n7469) );
  NAND2_X1 U8348 ( .A1(n7505), .A2(n10738), .ZN(n7501) );
  INV_X1 U8349 ( .A(n7191), .ZN(n7190) );
  OAI21_X1 U8350 ( .B1(n7193), .B2(n7192), .A(n8404), .ZN(n7191) );
  INV_X1 U8351 ( .A(n8054), .ZN(n7192) );
  INV_X1 U8352 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n6753) );
  INV_X1 U8353 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n6751) );
  AND2_X1 U8354 ( .A1(n7384), .A2(n6954), .ZN(n6951) );
  NOR2_X1 U8355 ( .A1(n14244), .A2(n10382), .ZN(n10411) );
  INV_X1 U8356 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7421) );
  INV_X1 U8357 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8533) );
  INV_X1 U8358 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8741) );
  NOR2_X1 U8359 ( .A1(n7777), .A2(n9879), .ZN(n9880) );
  NOR2_X1 U8360 ( .A1(n9808), .A2(n9807), .ZN(n7000) );
  NAND2_X1 U8361 ( .A1(n15271), .A2(n15240), .ZN(n10533) );
  INV_X1 U8362 ( .A(n7522), .ZN(n6817) );
  INV_X1 U8363 ( .A(n7532), .ZN(n7531) );
  AND2_X1 U8364 ( .A1(n6591), .A2(n8779), .ZN(n7474) );
  INV_X1 U8365 ( .A(n8708), .ZN(n8710) );
  INV_X1 U8366 ( .A(n8654), .ZN(n8655) );
  AOI21_X1 U8367 ( .B1(n7440), .B2(n12355), .A(n7438), .ZN(n7437) );
  INV_X1 U8368 ( .A(n12529), .ZN(n7438) );
  NOR2_X1 U8369 ( .A1(n7226), .A2(n7225), .ZN(n7224) );
  OAI21_X1 U8370 ( .B1(n13163), .B2(n13172), .A(n7157), .ZN(n7226) );
  INV_X1 U8371 ( .A(n10737), .ZN(n7507) );
  INV_X1 U8372 ( .A(n11525), .ZN(n6747) );
  NAND2_X1 U8373 ( .A1(n7329), .A2(n10735), .ZN(n7324) );
  AND2_X1 U8374 ( .A1(n10977), .A2(n7956), .ZN(n6995) );
  INV_X1 U8375 ( .A(n13454), .ZN(n7341) );
  NOR2_X1 U8376 ( .A1(n7341), .A2(n7338), .ZN(n7337) );
  NAND2_X1 U8377 ( .A1(n7960), .A2(n13485), .ZN(n7315) );
  INV_X1 U8378 ( .A(n13502), .ZN(n7322) );
  AND2_X1 U8379 ( .A1(n8073), .A2(n7237), .ZN(n7236) );
  INV_X1 U8380 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n7237) );
  AND2_X1 U8381 ( .A1(n14485), .A2(n7234), .ZN(n7233) );
  INV_X1 U8382 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n7234) );
  INV_X1 U8383 ( .A(n8335), .ZN(n8072) );
  AOI21_X1 U8384 ( .B1(n8483), .B2(n13127), .A(n6788), .ZN(n6787) );
  INV_X1 U8385 ( .A(n13130), .ZN(n6788) );
  INV_X1 U8386 ( .A(n13127), .ZN(n6785) );
  INV_X1 U8387 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8064) );
  OR2_X1 U8388 ( .A1(n13384), .A2(n11779), .ZN(n13082) );
  INV_X1 U8389 ( .A(n15699), .ZN(n11584) );
  INV_X1 U8390 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n8063) );
  CLKBUF_X1 U8391 ( .A(n11441), .Z(n13719) );
  AOI21_X1 U8392 ( .B1(n7221), .B2(n7220), .A(n6551), .ZN(n7219) );
  INV_X1 U8393 ( .A(n7671), .ZN(n7220) );
  NAND2_X1 U8394 ( .A1(n7651), .A2(n13004), .ZN(n7650) );
  INV_X1 U8395 ( .A(n7652), .ZN(n7651) );
  INV_X1 U8396 ( .A(n13021), .ZN(n7668) );
  INV_X1 U8397 ( .A(n8060), .ZN(n7604) );
  INV_X1 U8398 ( .A(n6616), .ZN(n7602) );
  INV_X1 U8399 ( .A(n7814), .ZN(n6772) );
  NAND2_X1 U8400 ( .A1(n7197), .A2(n7195), .ZN(n8047) );
  AND2_X1 U8401 ( .A1(n7196), .A2(n7595), .ZN(n7195) );
  AOI21_X1 U8402 ( .B1(n7597), .B2(n7599), .A(n7596), .ZN(n7595) );
  NAND2_X1 U8403 ( .A1(n8047), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8049) );
  INV_X1 U8404 ( .A(n7185), .ZN(n7184) );
  OAI21_X1 U8405 ( .B1(n7614), .B2(n7186), .A(n8221), .ZN(n7185) );
  INV_X1 U8406 ( .A(n8019), .ZN(n7186) );
  NAND2_X1 U8407 ( .A1(n7846), .A2(n7094), .ZN(n7863) );
  NOR2_X1 U8408 ( .A1(n9192), .A2(n6624), .ZN(n6694) );
  NAND2_X1 U8409 ( .A1(n9486), .A2(n9485), .ZN(n7042) );
  NAND2_X1 U8410 ( .A1(n9498), .A2(n9497), .ZN(n6982) );
  NAND2_X1 U8411 ( .A1(n9499), .A2(n9473), .ZN(n6981) );
  INV_X1 U8412 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8530) );
  INV_X1 U8413 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8529) );
  NAND2_X1 U8414 ( .A1(n15594), .A2(n12458), .ZN(n12459) );
  NOR2_X1 U8415 ( .A1(n15607), .A2(n12467), .ZN(n6706) );
  NOR2_X1 U8416 ( .A1(n15604), .A2(n15605), .ZN(n6707) );
  INV_X1 U8417 ( .A(n9256), .ZN(n9254) );
  AOI21_X1 U8418 ( .B1(n7566), .B2(n7565), .A(n6565), .ZN(n7564) );
  INV_X1 U8419 ( .A(n7569), .ZN(n7565) );
  AND2_X1 U8420 ( .A1(n7632), .A2(n7631), .ZN(n7630) );
  NOR2_X1 U8421 ( .A1(n14378), .A2(n14149), .ZN(n7632) );
  NAND2_X1 U8422 ( .A1(n6694), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U8423 ( .A1(n10357), .A2(n14261), .ZN(n6919) );
  INV_X1 U8424 ( .A(n7739), .ZN(n6915) );
  AOI21_X1 U8425 ( .B1(n7741), .B2(n7743), .A(n6520), .ZN(n7739) );
  INV_X1 U8426 ( .A(n10419), .ZN(n7549) );
  NOR2_X1 U8427 ( .A1(n6878), .A2(n7546), .ZN(n6876) );
  NAND2_X1 U8428 ( .A1(n6461), .A2(n14257), .ZN(n7617) );
  NOR2_X1 U8429 ( .A1(n9139), .A2(n9130), .ZN(n6693) );
  NOR2_X1 U8430 ( .A1(n6913), .A2(n6909), .ZN(n6908) );
  INV_X1 U8431 ( .A(n10348), .ZN(n6909) );
  INV_X1 U8432 ( .A(n10407), .ZN(n7574) );
  NOR2_X1 U8433 ( .A1(n14571), .A2(n12735), .ZN(n7613) );
  INV_X1 U8434 ( .A(n12052), .ZN(n7563) );
  INV_X1 U8435 ( .A(n9008), .ZN(n6689) );
  NAND2_X1 U8436 ( .A1(n10330), .A2(n11690), .ZN(n11705) );
  NAND2_X1 U8437 ( .A1(n6487), .A2(n10384), .ZN(n10755) );
  NAND2_X1 U8438 ( .A1(n10422), .A2(n7569), .ZN(n7568) );
  NAND2_X1 U8439 ( .A1(n7568), .A2(n7566), .ZN(n14120) );
  NAND2_X1 U8440 ( .A1(n6868), .A2(n6867), .ZN(n12373) );
  AOI21_X1 U8441 ( .B1(n6870), .B2(n6873), .A(n6548), .ZN(n6867) );
  AND2_X1 U8442 ( .A1(n9533), .A2(n11924), .ZN(n9274) );
  NAND2_X1 U8443 ( .A1(n6496), .A2(n8541), .ZN(n7582) );
  INV_X1 U8444 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8898) );
  INV_X1 U8445 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8896) );
  INV_X1 U8446 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8932) );
  NOR2_X1 U8447 ( .A1(n9831), .A2(n9830), .ZN(n6681) );
  INV_X1 U8448 ( .A(n14753), .ZN(n6930) );
  NOR2_X1 U8449 ( .A1(n6930), .A2(n6932), .ZN(n6928) );
  INV_X1 U8450 ( .A(n7689), .ZN(n6927) );
  OAI21_X1 U8451 ( .B1(n10904), .B2(n7700), .A(n7698), .ZN(n10171) );
  NAND2_X1 U8452 ( .A1(n10607), .A2(n10609), .ZN(n6836) );
  NOR2_X1 U8453 ( .A1(n10609), .A2(n10607), .ZN(n6834) );
  INV_X1 U8454 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9734) );
  OR2_X1 U8455 ( .A1(n10650), .A2(n6517), .ZN(n7527) );
  NAND2_X1 U8456 ( .A1(n6561), .A2(n7758), .ZN(n7757) );
  INV_X1 U8457 ( .A(n10029), .ZN(n7273) );
  OR2_X1 U8458 ( .A1(n7535), .A2(n7146), .ZN(n7143) );
  NOR2_X1 U8459 ( .A1(n7537), .A2(n7149), .ZN(n7148) );
  INV_X1 U8460 ( .A(n9880), .ZN(n7537) );
  NOR2_X1 U8461 ( .A1(n15199), .A2(n15345), .ZN(n7771) );
  NAND2_X1 U8462 ( .A1(n7000), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9831) );
  INV_X1 U8463 ( .A(n7000), .ZN(n9817) );
  AOI21_X1 U8464 ( .B1(n6474), .B2(n6850), .A(n6847), .ZN(n6846) );
  INV_X1 U8465 ( .A(n7718), .ZN(n6847) );
  AOI21_X1 U8466 ( .B1(n7718), .B2(n12714), .A(n6554), .ZN(n7276) );
  NAND2_X1 U8467 ( .A1(n15252), .A2(n15251), .ZN(n15226) );
  NAND2_X1 U8468 ( .A1(n9796), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9808) );
  INV_X1 U8469 ( .A(n9798), .ZN(n9796) );
  AOI21_X1 U8470 ( .B1(n12714), .B2(n7524), .A(n7523), .ZN(n7522) );
  INV_X1 U8471 ( .A(n12765), .ZN(n7523) );
  INV_X1 U8472 ( .A(n9765), .ZN(n7524) );
  NAND2_X1 U8473 ( .A1(n6679), .A2(n6610), .ZN(n9785) );
  INV_X1 U8474 ( .A(n9759), .ZN(n6679) );
  INV_X1 U8475 ( .A(n9705), .ZN(n6673) );
  NAND2_X1 U8476 ( .A1(n11879), .A2(n9669), .ZN(n10652) );
  NAND2_X1 U8477 ( .A1(n11865), .A2(n11564), .ZN(n11761) );
  AND2_X1 U8478 ( .A1(n7724), .A2(n15370), .ZN(n7720) );
  NAND2_X1 U8479 ( .A1(n7763), .A2(n12565), .ZN(n12769) );
  NAND2_X1 U8480 ( .A1(n11498), .A2(n11151), .ZN(n11253) );
  AOI21_X1 U8481 ( .B1(n7461), .B2(n7459), .A(n6626), .ZN(n7458) );
  INV_X1 U8482 ( .A(n8848), .ZN(n7459) );
  INV_X1 U8483 ( .A(n7461), .ZN(n7460) );
  NAND2_X1 U8484 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), 
        .ZN(n7710) );
  AOI21_X1 U8485 ( .B1(n7466), .B2(n8848), .A(n6613), .ZN(n7465) );
  INV_X1 U8486 ( .A(n8846), .ZN(n7466) );
  INV_X1 U8487 ( .A(n7474), .ZN(n7473) );
  AOI21_X1 U8488 ( .B1(n6948), .B2(n6950), .A(n6945), .ZN(n6944) );
  INV_X1 U8489 ( .A(n8755), .ZN(n6945) );
  INV_X1 U8490 ( .A(n7286), .ZN(n7285) );
  OAI21_X1 U8491 ( .B1(n7456), .B2(n6431), .A(n8676), .ZN(n7286) );
  INV_X1 U8492 ( .A(n8687), .ZN(n7284) );
  OR2_X1 U8493 ( .A1(n9714), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9741) );
  NAND2_X1 U8494 ( .A1(n8624), .A2(n8626), .ZN(n6987) );
  AND2_X1 U8495 ( .A1(n8605), .A2(n8608), .ZN(n6997) );
  INV_X1 U8496 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n14414) );
  NAND3_X1 U8497 ( .A1(n6636), .A2(n6635), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n6634) );
  INV_X1 U8498 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n6635) );
  XNOR2_X1 U8499 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n10774) );
  NAND2_X1 U8500 ( .A1(n7119), .A2(n7121), .ZN(n10891) );
  AND2_X1 U8501 ( .A1(n10988), .A2(n10987), .ZN(n11308) );
  OR2_X1 U8502 ( .A1(n10985), .A2(n10984), .ZN(n10988) );
  INV_X1 U8503 ( .A(n15441), .ZN(n6892) );
  INV_X1 U8504 ( .A(n12899), .ZN(n7432) );
  XNOR2_X1 U8505 ( .A(n12935), .B(n11584), .ZN(n11585) );
  NAND2_X1 U8506 ( .A1(n12531), .A2(n12532), .ZN(n12700) );
  NAND2_X1 U8507 ( .A1(n8071), .A2(n8070), .ZN(n8300) );
  INV_X1 U8508 ( .A(n13260), .ZN(n6963) );
  INV_X1 U8509 ( .A(n13259), .ZN(n6964) );
  AND2_X1 U8510 ( .A1(n8190), .A2(n8189), .ZN(n8204) );
  AOI21_X1 U8511 ( .B1(n13225), .B2(n12899), .A(n7435), .ZN(n7434) );
  INV_X1 U8512 ( .A(n13355), .ZN(n7435) );
  NAND2_X1 U8513 ( .A1(n8071), .A2(n6468), .ZN(n8321) );
  INV_X1 U8514 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n7228) );
  NAND2_X1 U8515 ( .A1(n8071), .A2(n7229), .ZN(n8309) );
  NAND2_X1 U8516 ( .A1(n7163), .A2(n7162), .ZN(n7161) );
  NAND2_X1 U8517 ( .A1(n13173), .A2(n7164), .ZN(n7163) );
  NAND2_X1 U8518 ( .A1(n13744), .A2(n13542), .ZN(n7164) );
  AND2_X1 U8519 ( .A1(n13170), .A2(n13171), .ZN(n7160) );
  INV_X1 U8520 ( .A(n6458), .ZN(n7035) );
  AND2_X1 U8521 ( .A1(n12883), .A2(n12882), .ZN(n12997) );
  AND4_X1 U8522 ( .A1(n8278), .A2(n8277), .A3(n8276), .A4(n8275), .ZN(n13270)
         );
  NAND2_X1 U8523 ( .A1(n7921), .A2(n11108), .ZN(n6644) );
  OR2_X1 U8524 ( .A1(n11402), .A2(n11401), .ZN(n11404) );
  NAND2_X1 U8525 ( .A1(n7055), .A2(n7054), .ZN(n7872) );
  INV_X1 U8526 ( .A(n7871), .ZN(n7055) );
  NAND2_X1 U8527 ( .A1(n11027), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n11026) );
  NAND2_X1 U8528 ( .A1(n11027), .A2(n6482), .ZN(n7504) );
  NAND2_X1 U8529 ( .A1(n7507), .A2(n7509), .ZN(n7506) );
  NAND2_X1 U8530 ( .A1(n11030), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n11029) );
  AND2_X1 U8531 ( .A1(n7325), .A2(n7328), .ZN(n7987) );
  AND2_X1 U8532 ( .A1(n7330), .A2(n7329), .ZN(n7325) );
  NAND2_X1 U8533 ( .A1(n7941), .A2(n8188), .ZN(n11356) );
  NAND2_X1 U8534 ( .A1(n7313), .A2(n10740), .ZN(n11357) );
  OR2_X1 U8535 ( .A1(n6994), .A2(n10741), .ZN(n7313) );
  NAND2_X1 U8536 ( .A1(n7988), .A2(n6747), .ZN(n6743) );
  NAND2_X1 U8537 ( .A1(n6994), .A2(n6485), .ZN(n7310) );
  CLKBUF_X1 U8538 ( .A(n11346), .Z(n11532) );
  NOR2_X1 U8539 ( .A1(n7989), .A2(n6745), .ZN(n11840) );
  INV_X1 U8540 ( .A(n13399), .ZN(n6740) );
  NAND2_X1 U8541 ( .A1(n11840), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n11839) );
  NOR2_X1 U8542 ( .A1(n13397), .A2(n7043), .ZN(n7885) );
  AND2_X1 U8543 ( .A1(n10845), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7043) );
  NOR2_X1 U8544 ( .A1(n13408), .A2(n13409), .ZN(n13406) );
  INV_X1 U8545 ( .A(n7991), .ZN(n13414) );
  NAND3_X1 U8546 ( .A1(n7991), .A2(n6467), .A3(n7349), .ZN(n7348) );
  OAI21_X1 U8547 ( .B1(n7992), .B2(n13430), .A(n10709), .ZN(n13432) );
  NAND3_X1 U8548 ( .A1(n7512), .A2(n7510), .A3(n7773), .ZN(n7893) );
  AND2_X1 U8549 ( .A1(n10977), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7004) );
  NAND2_X1 U8550 ( .A1(n13464), .A2(n7060), .ZN(n13481) );
  OR2_X1 U8551 ( .A1(n7959), .A2(n11017), .ZN(n7060) );
  NAND2_X1 U8552 ( .A1(n7320), .A2(n7322), .ZN(n7319) );
  INV_X1 U8553 ( .A(n13503), .ZN(n7320) );
  NAND2_X1 U8554 ( .A1(n6749), .A2(n6470), .ZN(n7318) );
  NAND2_X1 U8555 ( .A1(n9317), .A2(n8465), .ZN(n13525) );
  NAND2_X1 U8556 ( .A1(n8080), .A2(n8464), .ZN(n13531) );
  NAND2_X1 U8557 ( .A1(n7672), .A2(n8457), .ZN(n8459) );
  INV_X1 U8558 ( .A(n7223), .ZN(n8449) );
  AND2_X1 U8559 ( .A1(n13163), .A2(n13164), .ZN(n13537) );
  NAND2_X1 U8560 ( .A1(n8076), .A2(n8075), .ZN(n8434) );
  INV_X1 U8561 ( .A(n8421), .ZN(n8076) );
  NAND2_X1 U8562 ( .A1(n7643), .A2(n8417), .ZN(n13566) );
  NAND2_X1 U8563 ( .A1(n13579), .A2(n13580), .ZN(n7643) );
  AND2_X1 U8564 ( .A1(n6774), .A2(n7662), .ZN(n13568) );
  AOI21_X1 U8565 ( .B1(n7645), .B2(n6455), .A(n7663), .ZN(n7662) );
  INV_X1 U8566 ( .A(n13151), .ZN(n7663) );
  INV_X1 U8567 ( .A(n13565), .ZN(n8489) );
  NAND2_X1 U8568 ( .A1(n7215), .A2(n7216), .ZN(n13579) );
  AND2_X1 U8569 ( .A1(n13756), .A2(n13263), .ZN(n13147) );
  OR2_X1 U8570 ( .A1(n8374), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8385) );
  NAND2_X1 U8571 ( .A1(n8072), .A2(n7231), .ZN(n8374) );
  AND2_X1 U8572 ( .A1(n7233), .A2(n7232), .ZN(n7231) );
  INV_X1 U8573 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n7232) );
  NAND2_X1 U8574 ( .A1(n8072), .A2(n7233), .ZN(n8364) );
  OR2_X1 U8575 ( .A1(n8321), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8335) );
  NAND2_X1 U8576 ( .A1(n8072), .A2(n14485), .ZN(n8349) );
  NAND2_X1 U8577 ( .A1(n12758), .A2(n13021), .ZN(n13630) );
  NAND2_X1 U8578 ( .A1(n8069), .A2(n8068), .ZN(n8286) );
  INV_X1 U8579 ( .A(n8271), .ZN(n8069) );
  OR2_X1 U8580 ( .A1(n8258), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8271) );
  INV_X1 U8581 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8067) );
  OR2_X1 U8582 ( .A1(n8241), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8258) );
  NAND2_X1 U8583 ( .A1(n8480), .A2(n8479), .ZN(n12202) );
  NAND2_X1 U8584 ( .A1(n8066), .A2(n8065), .ZN(n8226) );
  NAND4_X1 U8585 ( .A1(n8063), .A2(n11732), .A3(n7238), .A4(n8064), .ZN(n8197)
         );
  INV_X1 U8586 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n7238) );
  NAND2_X1 U8587 ( .A1(n11694), .A2(n13074), .ZN(n6766) );
  INV_X1 U8588 ( .A(n8476), .ZN(n13079) );
  INV_X1 U8589 ( .A(n11697), .ZN(n13074) );
  NAND2_X1 U8590 ( .A1(n13077), .A2(n13076), .ZN(n11697) );
  NAND2_X1 U8591 ( .A1(n9316), .A2(n9315), .ZN(n12994) );
  AND2_X1 U8592 ( .A1(n13135), .A2(n13131), .ZN(n13130) );
  OAI21_X1 U8593 ( .B1(n12070), .B2(n7635), .A(n6542), .ZN(n12613) );
  NAND3_X1 U8594 ( .A1(n13121), .A2(n7637), .A3(n6477), .ZN(n7636) );
  AND2_X1 U8595 ( .A1(n12280), .A2(n13275), .ZN(n13049) );
  OAI21_X1 U8596 ( .B1(n12013), .B2(n8249), .A(n8248), .ZN(n8251) );
  NAND2_X1 U8597 ( .A1(n12948), .A2(n12947), .ZN(n12992) );
  NAND2_X1 U8598 ( .A1(n9314), .A2(n9313), .ZN(n12874) );
  OR2_X1 U8599 ( .A1(n9311), .A2(n9310), .ZN(n9314) );
  NAND2_X1 U8600 ( .A1(n8059), .A2(n8058), .ZN(n8444) );
  NAND2_X1 U8601 ( .A1(n8431), .A2(n8057), .ZN(n8059) );
  INV_X1 U8602 ( .A(n7821), .ZN(n7820) );
  NAND2_X1 U8603 ( .A1(n8055), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7624) );
  AND2_X1 U8604 ( .A1(n7910), .A2(n7909), .ZN(n13191) );
  AOI21_X1 U8605 ( .B1(n7592), .B2(n7594), .A(n7590), .ZN(n7589) );
  INV_X1 U8606 ( .A(n8025), .ZN(n7590) );
  OR2_X1 U8607 ( .A1(n7843), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n7882) );
  INV_X1 U8608 ( .A(n8011), .ZN(n7588) );
  AND2_X1 U8609 ( .A1(n8011), .A2(n8010), .ZN(n8159) );
  NAND2_X1 U8610 ( .A1(n8160), .A2(n8159), .ZN(n8162) );
  AND2_X1 U8611 ( .A1(n8009), .A2(n8008), .ZN(n8144) );
  NAND2_X1 U8612 ( .A1(n10797), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8006) );
  NAND2_X1 U8613 ( .A1(n10876), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8005) );
  XNOR2_X1 U8614 ( .A(n6748), .B(n7854), .ZN(n7973) );
  NAND2_X1 U8615 ( .A1(n7853), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6748) );
  XNOR2_X1 U8616 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n8112) );
  OR2_X1 U8617 ( .A1(n7400), .A2(n11627), .ZN(n6807) );
  INV_X1 U8618 ( .A(n9019), .ZN(n7400) );
  OR2_X1 U8619 ( .A1(n9172), .A2(n9171), .ZN(n6803) );
  AND2_X1 U8620 ( .A1(n6978), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7620) );
  OR2_X1 U8621 ( .A1(n11483), .A2(n8963), .ZN(n13861) );
  OR2_X1 U8622 ( .A1(n9174), .A2(n9173), .ZN(n9192) );
  INV_X1 U8623 ( .A(n6694), .ZN(n9205) );
  AOI21_X1 U8624 ( .B1(n6810), .B2(n6475), .A(n6808), .ZN(n12507) );
  OAI21_X1 U8625 ( .B1(n9090), .B2(n9091), .A(n6809), .ZN(n6808) );
  INV_X1 U8626 ( .A(n12135), .ZN(n6810) );
  AND2_X1 U8627 ( .A1(n9105), .A2(n9104), .ZN(n12508) );
  NAND2_X1 U8628 ( .A1(n12803), .A2(n7412), .ZN(n7411) );
  NOR2_X1 U8629 ( .A1(n9228), .A2(n9227), .ZN(n9229) );
  NAND2_X1 U8630 ( .A1(n12002), .A2(n9050), .ZN(n12135) );
  NAND2_X1 U8631 ( .A1(n12135), .A2(n12136), .ZN(n12134) );
  NAND2_X1 U8632 ( .A1(n8977), .A2(n8976), .ZN(n11473) );
  AND2_X1 U8633 ( .A1(n8982), .A2(n8981), .ZN(n13822) );
  NAND2_X1 U8634 ( .A1(n6693), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9166) );
  NAND2_X1 U8635 ( .A1(n8946), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9174) );
  INV_X1 U8636 ( .A(n9166), .ZN(n8946) );
  XNOR2_X1 U8637 ( .A(n14113), .B(n8969), .ZN(n9251) );
  NOR2_X1 U8638 ( .A1(n11072), .A2(n6541), .ZN(n15565) );
  AND2_X1 U8639 ( .A1(n11239), .A2(n11094), .ZN(n11096) );
  OR2_X1 U8640 ( .A1(n11428), .A2(n11427), .ZN(n11464) );
  XNOR2_X1 U8641 ( .A(n12459), .B(n15607), .ZN(n15612) );
  XNOR2_X1 U8642 ( .A(n7079), .B(n12640), .ZN(n12636) );
  AOI21_X1 U8643 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n12636), .A(n7078), .ZN(
        n14036) );
  NOR2_X1 U8644 ( .A1(n7079), .A2(n12469), .ZN(n7078) );
  AOI22_X1 U8645 ( .A1(n14052), .A2(n14051), .B1(n14050), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n14060) );
  INV_X1 U8646 ( .A(n10461), .ZN(n10379) );
  INV_X1 U8647 ( .A(n10444), .ZN(n7254) );
  INV_X1 U8648 ( .A(n7553), .ZN(n7552) );
  NAND2_X1 U8649 ( .A1(n10432), .A2(n7555), .ZN(n7554) );
  NAND2_X1 U8650 ( .A1(n7553), .A2(n10432), .ZN(n6687) );
  INV_X1 U8651 ( .A(n7556), .ZN(n7555) );
  NAND2_X1 U8652 ( .A1(n6797), .A2(n14178), .ZN(n14096) );
  NAND2_X1 U8653 ( .A1(n7257), .A2(n10374), .ZN(n7256) );
  INV_X1 U8654 ( .A(n7745), .ZN(n7257) );
  NOR2_X1 U8655 ( .A1(n14102), .A2(n7746), .ZN(n7745) );
  INV_X1 U8656 ( .A(n10371), .ZN(n7746) );
  AND2_X1 U8657 ( .A1(n9256), .A2(n9244), .ZN(n14114) );
  NAND2_X1 U8658 ( .A1(n10428), .A2(n10427), .ZN(n14107) );
  NAND2_X1 U8659 ( .A1(n14178), .A2(n7630), .ZN(n14132) );
  NAND2_X1 U8660 ( .A1(n14178), .A2(n7632), .ZN(n14147) );
  NAND2_X1 U8661 ( .A1(n14178), .A2(n14168), .ZN(n14164) );
  INV_X1 U8662 ( .A(n14297), .ZN(n6793) );
  INV_X1 U8663 ( .A(n6693), .ZN(n9155) );
  OR2_X1 U8664 ( .A1(n9117), .A2(n8944), .ZN(n9137) );
  NAND2_X1 U8665 ( .A1(n8945), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9139) );
  INV_X1 U8666 ( .A(n9137), .ZN(n8945) );
  OAI21_X1 U8667 ( .B1(n12574), .B2(n7575), .A(n7572), .ZN(n12814) );
  AOI21_X1 U8668 ( .B1(n7576), .B2(n7574), .A(n7573), .ZN(n7572) );
  INV_X1 U8669 ( .A(n7576), .ZN(n7575) );
  INV_X1 U8670 ( .A(n10409), .ZN(n7573) );
  NAND2_X1 U8671 ( .A1(n6486), .A2(n12732), .ZN(n12677) );
  OR2_X1 U8672 ( .A1(n9072), .A2(n11460), .ZN(n9094) );
  OR2_X1 U8673 ( .A1(n9094), .A2(n9093), .ZN(n9117) );
  OAI21_X1 U8674 ( .B1(n12051), .B2(n6905), .A(n6902), .ZN(n12726) );
  NAND2_X1 U8675 ( .A1(n6440), .A2(n6478), .ZN(n6905) );
  AOI21_X1 U8676 ( .B1(n6440), .B2(n6904), .A(n6903), .ZN(n6902) );
  NAND2_X1 U8677 ( .A1(n12726), .A2(n10344), .ZN(n12725) );
  NAND2_X1 U8678 ( .A1(n8941), .A2(n6530), .ZN(n9066) );
  AND2_X1 U8679 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n8942) );
  NAND2_X1 U8680 ( .A1(n8941), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9053) );
  NOR2_X1 U8681 ( .A1(n12401), .A2(n12409), .ZN(n12732) );
  NAND2_X1 U8682 ( .A1(n12051), .A2(n10339), .ZN(n12247) );
  NAND2_X1 U8683 ( .A1(n12247), .A2(n12248), .ZN(n12369) );
  NAND2_X1 U8684 ( .A1(n6690), .A2(n6689), .ZN(n9032) );
  NOR2_X1 U8685 ( .A1(n6692), .A2(n6691), .ZN(n6690) );
  NOR2_X1 U8686 ( .A1(n11937), .A2(n7625), .ZN(n12062) );
  NAND2_X1 U8687 ( .A1(n7628), .A2(n6796), .ZN(n7625) );
  NAND2_X1 U8688 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9008) );
  NAND2_X1 U8689 ( .A1(n6689), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9020) );
  NAND2_X1 U8690 ( .A1(n11932), .A2(n11931), .ZN(n11930) );
  NAND2_X1 U8691 ( .A1(n7627), .A2(n6796), .ZN(n11938) );
  INV_X1 U8692 ( .A(n11937), .ZN(n7627) );
  NOR2_X1 U8693 ( .A1(n11971), .A2(n11979), .ZN(n11972) );
  OR2_X1 U8694 ( .A1(n13859), .A2(n11485), .ZN(n11971) );
  INV_X1 U8695 ( .A(n15648), .ZN(n15656) );
  NAND2_X1 U8696 ( .A1(n8881), .A2(n8882), .ZN(n8880) );
  INV_X1 U8697 ( .A(n8807), .ZN(n8805) );
  OR2_X1 U8698 ( .A1(n8680), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8718) );
  OR2_X1 U8699 ( .A1(n8627), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8629) );
  OR2_X1 U8700 ( .A1(n8629), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8638) );
  OR2_X1 U8701 ( .A1(n8594), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8619) );
  INV_X1 U8702 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8573) );
  INV_X1 U8703 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8550) );
  INV_X1 U8704 ( .A(n6681), .ZN(n9852) );
  INV_X1 U8705 ( .A(n14765), .ZN(n7676) );
  INV_X1 U8706 ( .A(n10144), .ZN(n6934) );
  NAND2_X1 U8707 ( .A1(n7001), .A2(n9905), .ZN(n9917) );
  INV_X1 U8708 ( .A(n9907), .ZN(n7001) );
  OR2_X1 U8709 ( .A1(n10270), .A2(n10269), .ZN(n10271) );
  CLKBUF_X1 U8710 ( .A(n11826), .Z(n11827) );
  NAND2_X1 U8711 ( .A1(n10091), .A2(n6923), .ZN(n11144) );
  NAND2_X1 U8712 ( .A1(n6681), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9870) );
  OR2_X1 U8713 ( .A1(n9735), .A2(n9734), .ZN(n9747) );
  AND2_X1 U8714 ( .A1(n12587), .A2(n12582), .ZN(n12583) );
  INV_X1 U8715 ( .A(n14819), .ZN(n9995) );
  NOR2_X1 U8716 ( .A1(n14715), .A2(n7681), .ZN(n7680) );
  INV_X1 U8717 ( .A(n14708), .ZN(n7681) );
  OAI22_X1 U8718 ( .A1(n14715), .A2(n7679), .B1(n10223), .B2(n10224), .ZN(
        n7678) );
  AND2_X1 U8719 ( .A1(n10207), .A2(n7244), .ZN(n7243) );
  INV_X1 U8720 ( .A(n10211), .ZN(n7244) );
  NAND2_X1 U8721 ( .A1(n14842), .A2(n7006), .ZN(n14866) );
  AND2_X1 U8722 ( .A1(n7008), .A2(n7007), .ZN(n7006) );
  NAND2_X1 U8723 ( .A1(n14843), .A2(n10915), .ZN(n7007) );
  OR2_X1 U8724 ( .A1(n14843), .A2(n10915), .ZN(n7008) );
  OR2_X1 U8725 ( .A1(n11274), .A2(n11273), .ZN(n11611) );
  OR2_X1 U8726 ( .A1(n11613), .A2(n11612), .ZN(n11669) );
  AND2_X1 U8727 ( .A1(n6737), .A2(n6736), .ZN(n11658) );
  NOR2_X1 U8728 ( .A1(n11604), .A2(n11605), .ZN(n6736) );
  INV_X1 U8729 ( .A(n11606), .ZN(n6737) );
  OR2_X1 U8730 ( .A1(n12121), .A2(n7059), .ZN(n7058) );
  NOR2_X1 U8731 ( .A1(n12124), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7059) );
  NAND2_X1 U8732 ( .A1(n6719), .A2(n6720), .ZN(n14981) );
  AND2_X1 U8733 ( .A1(n6721), .A2(n6629), .ZN(n6720) );
  INV_X1 U8734 ( .A(n10030), .ZN(n7727) );
  AND2_X1 U8735 ( .A1(n10028), .A2(n7714), .ZN(n7713) );
  NAND2_X1 U8736 ( .A1(n10024), .A2(n7715), .ZN(n7714) );
  INV_X1 U8737 ( .A(n10024), .ZN(n7716) );
  NAND2_X1 U8738 ( .A1(n10025), .A2(n15048), .ZN(n15071) );
  INV_X1 U8739 ( .A(n15047), .ZN(n15093) );
  NOR2_X2 U8740 ( .A1(n15230), .A2(n7770), .ZN(n15183) );
  NAND2_X1 U8741 ( .A1(n15186), .A2(n7771), .ZN(n7770) );
  NOR2_X1 U8742 ( .A1(n15230), .A2(n7769), .ZN(n15198) );
  INV_X1 U8743 ( .A(n7771), .ZN(n7769) );
  NAND2_X1 U8744 ( .A1(n15211), .A2(n10012), .ZN(n15190) );
  NAND2_X1 U8745 ( .A1(n6815), .A2(n7520), .ZN(n12767) );
  NAND2_X1 U8746 ( .A1(n12559), .A2(n7522), .ZN(n6815) );
  NAND2_X1 U8747 ( .A1(n12559), .A2(n9765), .ZN(n12713) );
  OR2_X1 U8748 ( .A1(n9747), .A2(n9746), .ZN(n9759) );
  NAND2_X1 U8749 ( .A1(n6679), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9774) );
  NAND2_X1 U8750 ( .A1(n12419), .A2(n10006), .ZN(n12556) );
  NAND2_X1 U8751 ( .A1(n7534), .A2(n6528), .ZN(n12561) );
  NAND2_X1 U8752 ( .A1(n12421), .A2(n12420), .ZN(n12419) );
  NAND2_X1 U8753 ( .A1(n12192), .A2(n9726), .ZN(n12328) );
  NAND2_X1 U8754 ( .A1(n6673), .A2(n6671), .ZN(n9735) );
  NOR2_X1 U8755 ( .A1(n6674), .A2(n6672), .ZN(n6671) );
  NAND2_X1 U8756 ( .A1(n6673), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9718) );
  NAND2_X1 U8757 ( .A1(n12149), .A2(n9713), .ZN(n12190) );
  OR2_X1 U8758 ( .A1(n10001), .A2(n10000), .ZN(n10002) );
  NAND2_X1 U8759 ( .A1(n11509), .A2(n11770), .ZN(n11871) );
  INV_X1 U8760 ( .A(n10651), .ZN(n11512) );
  AND2_X1 U8761 ( .A1(n15191), .A2(n10562), .ZN(n15179) );
  AND2_X1 U8762 ( .A1(n15195), .A2(n15194), .ZN(n15340) );
  AND2_X1 U8763 ( .A1(n7151), .A2(n7530), .ZN(n15215) );
  NAND2_X1 U8764 ( .A1(n6812), .A2(n6816), .ZN(n7151) );
  NAND2_X1 U8765 ( .A1(n7542), .A2(n9697), .ZN(n12151) );
  NAND2_X1 U8766 ( .A1(n9986), .A2(n6862), .ZN(n6863) );
  AND2_X1 U8767 ( .A1(n15436), .A2(n14825), .ZN(n6862) );
  AND2_X1 U8768 ( .A1(n9585), .A2(n9604), .ZN(n7077) );
  INV_X1 U8769 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U8770 ( .A1(n8849), .A2(n8848), .ZN(n8855) );
  XNOR2_X1 U8771 ( .A(n8838), .B(n8833), .ZN(n14643) );
  NAND2_X1 U8772 ( .A1(n7249), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10041) );
  AND2_X1 U8773 ( .A1(n6501), .A2(n9581), .ZN(n7247) );
  NAND2_X1 U8774 ( .A1(n9982), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9983) );
  NOR2_X1 U8775 ( .A1(n9976), .A2(n9975), .ZN(n9977) );
  OR2_X1 U8776 ( .A1(n9973), .A2(n9572), .ZN(n9978) );
  NOR2_X1 U8777 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n9975) );
  NAND2_X1 U8778 ( .A1(n8783), .A2(n8782), .ZN(n6639) );
  INV_X1 U8779 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9980) );
  XNOR2_X1 U8780 ( .A(n8763), .B(n8762), .ZN(n11453) );
  NAND2_X1 U8781 ( .A1(n6947), .A2(n8733), .ZN(n8748) );
  NAND2_X1 U8782 ( .A1(n8717), .A2(n6640), .ZN(n10978) );
  INV_X1 U8783 ( .A(n8715), .ZN(n8712) );
  OAI21_X1 U8784 ( .B1(n7122), .B2(n8702), .A(n8708), .ZN(n8691) );
  XNOR2_X1 U8785 ( .A(n8677), .B(n8676), .ZN(n10982) );
  OR2_X1 U8786 ( .A1(n9684), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9698) );
  INV_X1 U8787 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10777) );
  AND2_X1 U8788 ( .A1(n10768), .A2(n10767), .ZN(n10772) );
  XNOR2_X1 U8789 ( .A(n10799), .B(n15496), .ZN(n10803) );
  NAND2_X1 U8790 ( .A1(n11305), .A2(n11304), .ZN(n11648) );
  INV_X1 U8791 ( .A(n7299), .ZN(n7298) );
  NOR2_X1 U8792 ( .A1(n6446), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7300) );
  NOR2_X1 U8793 ( .A1(n6892), .A2(n15443), .ZN(n6889) );
  INV_X1 U8794 ( .A(n7292), .ZN(n7291) );
  NOR2_X1 U8795 ( .A1(n7291), .A2(n6889), .ZN(n6888) );
  INV_X1 U8796 ( .A(n13381), .ZN(n12537) );
  NOR2_X1 U8797 ( .A1(n12342), .A2(n6427), .ZN(n12354) );
  OR2_X1 U8798 ( .A1(n13226), .A2(n13225), .ZN(n13227) );
  INV_X1 U8799 ( .A(n13380), .ZN(n12702) );
  NAND2_X1 U8800 ( .A1(n13335), .A2(n12908), .ZN(n13248) );
  OAI21_X1 U8801 ( .B1(n13337), .B2(n7429), .A(n7427), .ZN(n13246) );
  NAND2_X1 U8802 ( .A1(n7436), .A2(n7440), .ZN(n12530) );
  NAND2_X1 U8803 ( .A1(n12342), .A2(n7441), .ZN(n7436) );
  AND2_X1 U8804 ( .A1(n12925), .A2(n7443), .ZN(n7442) );
  NAND2_X1 U8805 ( .A1(n7445), .A2(n7444), .ZN(n7443) );
  NAND2_X1 U8806 ( .A1(n8433), .A2(n8432), .ZN(n13675) );
  AOI22_X1 U8807 ( .A1(n13307), .A2(n6970), .B1(n13308), .B2(n13595), .ZN(
        n6972) );
  NAND2_X1 U8808 ( .A1(n12918), .A2(n13569), .ZN(n6970) );
  NAND2_X1 U8809 ( .A1(n8420), .A2(n8419), .ZN(n8488) );
  AND2_X1 U8810 ( .A1(n11180), .A2(n11281), .ZN(n13357) );
  AOI21_X1 U8811 ( .B1(n7427), .B2(n7429), .A(n6513), .ZN(n7425) );
  NAND2_X1 U8812 ( .A1(n13257), .A2(n13237), .ZN(n13327) );
  NAND2_X1 U8813 ( .A1(n6509), .A2(n7085), .ZN(n7084) );
  INV_X1 U8814 ( .A(n11181), .ZN(n7085) );
  NAND2_X1 U8815 ( .A1(n13337), .A2(n13336), .ZN(n13335) );
  NOR2_X1 U8816 ( .A1(n12161), .A2(n7787), .ZN(n12164) );
  AND2_X1 U8817 ( .A1(n8441), .A2(n8440), .ZN(n13570) );
  NAND2_X1 U8818 ( .A1(n13227), .A2(n12899), .ZN(n13356) );
  NAND2_X1 U8819 ( .A1(n7430), .A2(n7434), .ZN(n13354) );
  NAND2_X1 U8820 ( .A1(n13226), .A2(n12899), .ZN(n7430) );
  INV_X1 U8821 ( .A(n13351), .ZN(n13353) );
  INV_X1 U8822 ( .A(n12997), .ZN(n13368) );
  NAND2_X1 U8823 ( .A1(n8402), .A2(n8401), .ZN(n13604) );
  INV_X1 U8824 ( .A(P3_U3897), .ZN(n13372) );
  NAND4_X1 U8825 ( .A1(n8158), .A2(n8157), .A3(n8156), .A4(n8155), .ZN(n11554)
         );
  OR2_X1 U8826 ( .A1(n8138), .A2(n11696), .ZN(n8156) );
  OR2_X1 U8827 ( .A1(n8138), .A2(n11295), .ZN(n8129) );
  OR2_X1 U8828 ( .A1(n8153), .A2(n8117), .ZN(n8119) );
  INV_X1 U8829 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7802) );
  NAND2_X1 U8830 ( .A1(n7336), .A2(n7334), .ZN(n11393) );
  NOR2_X1 U8831 ( .A1(n7335), .A2(n15689), .ZN(n7334) );
  INV_X1 U8832 ( .A(n7976), .ZN(n7335) );
  NAND2_X1 U8833 ( .A1(n7336), .A2(n7976), .ZN(n11391) );
  CLKBUF_X1 U8834 ( .A(n11038), .Z(n6994) );
  NAND2_X1 U8835 ( .A1(n6653), .A2(n6652), .ZN(n11520) );
  NAND2_X1 U8836 ( .A1(n7309), .A2(n7307), .ZN(n6653) );
  NAND2_X1 U8837 ( .A1(n6564), .A2(n11038), .ZN(n6652) );
  AND2_X1 U8838 ( .A1(n7310), .A2(n7308), .ZN(n11522) );
  INV_X1 U8839 ( .A(n7309), .ZN(n7308) );
  NAND2_X1 U8840 ( .A1(n7492), .A2(n7095), .ZN(n7486) );
  NOR2_X1 U8841 ( .A1(n11346), .A2(n11531), .ZN(n7490) );
  NAND2_X1 U8842 ( .A1(n7489), .A2(n11849), .ZN(n7488) );
  INV_X1 U8843 ( .A(n7304), .ZN(n13389) );
  AND2_X1 U8844 ( .A1(n6741), .A2(n6740), .ZN(n13401) );
  AOI21_X1 U8845 ( .B1(n13395), .B2(n7487), .A(n13394), .ZN(n13397) );
  NAND2_X1 U8846 ( .A1(n13425), .A2(n6604), .ZN(n10719) );
  INV_X1 U8847 ( .A(n7345), .ZN(n7344) );
  NOR2_X1 U8848 ( .A1(n7093), .A2(n7516), .ZN(n13442) );
  INV_X1 U8849 ( .A(n7517), .ZN(n7516) );
  NOR2_X1 U8850 ( .A1(n13455), .A2(n7342), .ZN(n13440) );
  NAND2_X1 U8851 ( .A1(n7514), .A2(n13458), .ZN(n13463) );
  NAND2_X1 U8852 ( .A1(n7339), .A2(n13454), .ZN(n13457) );
  OR2_X1 U8853 ( .A1(n7997), .A2(n13485), .ZN(n6750) );
  NAND2_X1 U8854 ( .A1(n7318), .A2(n7319), .ZN(n13506) );
  NAND2_X1 U8855 ( .A1(n13478), .A2(n7901), .ZN(n7484) );
  XNOR2_X1 U8856 ( .A(n7104), .B(n7162), .ZN(n13668) );
  NAND2_X1 U8857 ( .A1(n9302), .A2(n7221), .ZN(n13519) );
  NAND2_X1 U8858 ( .A1(n6777), .A2(n6780), .ZN(n9346) );
  OR2_X1 U8859 ( .A1(n13556), .A2(n6782), .ZN(n6777) );
  XNOR2_X1 U8860 ( .A(n13538), .B(n13537), .ZN(n13672) );
  NAND2_X1 U8861 ( .A1(n13556), .A2(n13160), .ZN(n13538) );
  NAND2_X1 U8862 ( .A1(n7214), .A2(n7641), .ZN(n13550) );
  NAND2_X1 U8863 ( .A1(n7201), .A2(n7202), .ZN(n13636) );
  NAND2_X1 U8864 ( .A1(n8316), .A2(n8315), .ZN(n12756) );
  INV_X1 U8865 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11732) );
  INV_X1 U8866 ( .A(n13645), .ZN(n15685) );
  INV_X1 U8867 ( .A(n13588), .ZN(n13659) );
  AOI21_X1 U8868 ( .B1(n13195), .B2(n12985), .A(n7789), .ZN(n12996) );
  INV_X1 U8869 ( .A(n9309), .ZN(n13741) );
  OAI21_X1 U8870 ( .B1(n13603), .B2(n13003), .A(n13002), .ZN(n13594) );
  OAI21_X1 U8871 ( .B1(n13632), .B2(n6447), .A(n7654), .ZN(n13601) );
  NAND2_X1 U8872 ( .A1(n8373), .A2(n8372), .ZN(n13768) );
  NAND2_X1 U8873 ( .A1(n7649), .A2(n13004), .ZN(n13612) );
  NAND2_X1 U8874 ( .A1(n6988), .A2(n7652), .ZN(n7649) );
  NAND2_X1 U8875 ( .A1(n7657), .A2(n13038), .ZN(n13610) );
  NAND2_X1 U8876 ( .A1(n13632), .A2(n7660), .ZN(n7657) );
  NAND2_X1 U8877 ( .A1(n6988), .A2(n8356), .ZN(n13622) );
  NAND2_X1 U8878 ( .A1(n13632), .A2(n13043), .ZN(n13620) );
  NAND2_X1 U8879 ( .A1(n8334), .A2(n8333), .ZN(n13789) );
  NAND2_X1 U8880 ( .A1(n7206), .A2(n8328), .ZN(n13652) );
  NAND2_X1 U8881 ( .A1(n8316), .A2(n7669), .ZN(n7206) );
  NAND2_X1 U8882 ( .A1(n8308), .A2(n8307), .ZN(n13366) );
  NAND2_X1 U8883 ( .A1(n8285), .A2(n8284), .ZN(n12790) );
  OAI21_X1 U8884 ( .B1(n8480), .B2(n6477), .A(n7637), .ZN(n12389) );
  NAND2_X1 U8885 ( .A1(n7666), .A2(n7665), .ZN(n12207) );
  NAND2_X1 U8886 ( .A1(n8270), .A2(n8269), .ZN(n13278) );
  OR2_X1 U8887 ( .A1(n10873), .A2(n8346), .ZN(n8270) );
  AND2_X1 U8888 ( .A1(n11169), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13797) );
  XNOR2_X1 U8889 ( .A(n9311), .B(n9305), .ZN(n13802) );
  AND2_X1 U8890 ( .A1(n6494), .A2(n7452), .ZN(n7451) );
  NAND2_X1 U8891 ( .A1(n7189), .A2(n8054), .ZN(n8405) );
  INV_X1 U8892 ( .A(n13191), .ZN(n11964) );
  OAI21_X1 U8893 ( .B1(n8344), .B2(n7599), .A(n7597), .ZN(n8357) );
  NAND2_X1 U8894 ( .A1(n8342), .A2(n8044), .ZN(n8359) );
  OAI21_X1 U8895 ( .B1(n8266), .B2(n7178), .A(n7176), .ZN(n8296) );
  OAI21_X1 U8896 ( .B1(n8211), .B2(n7594), .A(n7592), .ZN(n8237) );
  NAND2_X1 U8897 ( .A1(n8209), .A2(n8023), .ZN(n8235) );
  NAND2_X1 U8898 ( .A1(n8194), .A2(n8019), .ZN(n8223) );
  INV_X1 U8899 ( .A(n7849), .ZN(n7873) );
  NAND2_X1 U8900 ( .A1(n8016), .A2(n8015), .ZN(n8192) );
  INV_X1 U8901 ( .A(n7846), .ZN(n7861) );
  XNOR2_X1 U8902 ( .A(n9040), .B(n9038), .ZN(n11748) );
  NAND2_X1 U8903 ( .A1(n7398), .A2(n9030), .ZN(n11749) );
  NAND2_X1 U8904 ( .A1(n11574), .A2(n7399), .ZN(n7398) );
  INV_X1 U8905 ( .A(n6807), .ZN(n7399) );
  AND2_X1 U8906 ( .A1(n7135), .A2(n6493), .ZN(n12804) );
  NAND2_X1 U8907 ( .A1(n12134), .A2(n9064), .ZN(n12483) );
  OAI21_X1 U8908 ( .B1(n11574), .B2(n7397), .A(n7395), .ZN(n12004) );
  NAND2_X1 U8909 ( .A1(n7417), .A2(n9191), .ZN(n10727) );
  NAND2_X1 U8910 ( .A1(n7130), .A2(n7128), .ZN(n7417) );
  OR2_X1 U8911 ( .A1(n9216), .A2(n9215), .ZN(n7786) );
  OAI21_X1 U8912 ( .B1(n13835), .B2(n13833), .A(n13832), .ZN(n13906) );
  NAND2_X1 U8913 ( .A1(n12506), .A2(n9105), .ZN(n12550) );
  NAND2_X1 U8914 ( .A1(n8683), .A2(n8682), .ZN(n12678) );
  AOI21_X1 U8915 ( .B1(n6471), .B2(n7409), .A(n7408), .ZN(n7407) );
  INV_X1 U8916 ( .A(n9164), .ZN(n7408) );
  NAND2_X1 U8917 ( .A1(n11574), .A2(n9019), .ZN(n11628) );
  AND2_X1 U8918 ( .A1(n9295), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13938) );
  NAND2_X1 U8919 ( .A1(n13867), .A2(n9240), .ZN(n13935) );
  INV_X1 U8920 ( .A(n13938), .ZN(n13952) );
  NAND2_X1 U8921 ( .A1(n7793), .A2(n9533), .ZN(n9534) );
  OR2_X1 U8922 ( .A1(n9464), .A2(n11975), .ZN(n8973) );
  OR2_X1 U8923 ( .A1(n9464), .A2(n11599), .ZN(n8960) );
  INV_X1 U8924 ( .A(n6704), .ZN(n11051) );
  OAI21_X1 U8925 ( .B1(n14019), .B2(n14014), .A(n11076), .ZN(n14017) );
  AND2_X1 U8926 ( .A1(n6709), .A2(n6708), .ZN(n11236) );
  INV_X1 U8927 ( .A(n11223), .ZN(n6708) );
  NAND2_X1 U8928 ( .A1(n14017), .A2(n11224), .ZN(n6709) );
  NOR2_X1 U8929 ( .A1(n11236), .A2(n7080), .ZN(n11238) );
  AND2_X1 U8930 ( .A1(n11228), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7080) );
  OAI21_X1 U8931 ( .B1(n12465), .B2(n12464), .A(n6553), .ZN(n15578) );
  AND2_X1 U8932 ( .A1(n8673), .A2(n8680), .ZN(n15580) );
  OR2_X1 U8933 ( .A1(n15593), .A2(n15592), .ZN(n15594) );
  OAI22_X1 U8934 ( .A1(n14036), .A2(n14035), .B1(n14043), .B2(n12637), .ZN(
        n14052) );
  NAND2_X1 U8935 ( .A1(n14065), .A2(n14047), .ZN(n14049) );
  OAI21_X1 U8936 ( .B1(n14069), .B2(n15597), .A(n6462), .ZN(n6700) );
  OAI21_X1 U8937 ( .B1(n14068), .B2(n15591), .A(n15608), .ZN(n6702) );
  NOR2_X1 U8938 ( .A1(n15618), .A2(n14072), .ZN(n6698) );
  INV_X1 U8939 ( .A(n14071), .ZN(n6697) );
  NOR2_X1 U8940 ( .A1(n8884), .A2(n14320), .ZN(n14073) );
  NAND2_X1 U8941 ( .A1(n7747), .A2(n10371), .ZN(n10372) );
  OAI21_X1 U8942 ( .B1(n10428), .B2(n14106), .A(n6879), .ZN(n6881) );
  AOI21_X1 U8943 ( .B1(n6880), .B2(n14111), .A(n7558), .ZN(n6879) );
  NAND2_X1 U8944 ( .A1(n12241), .A2(n8834), .ZN(n8823) );
  NAND2_X1 U8945 ( .A1(n7756), .A2(n10364), .ZN(n14144) );
  NAND2_X1 U8946 ( .A1(n7268), .A2(n7266), .ZN(n7756) );
  NAND2_X1 U8947 ( .A1(n7268), .A2(n10362), .ZN(n14158) );
  NAND2_X1 U8948 ( .A1(n10422), .A2(n10421), .ZN(n14172) );
  NAND2_X1 U8949 ( .A1(n7740), .A2(n7742), .ZN(n14194) );
  NAND2_X1 U8950 ( .A1(n14213), .A2(n7744), .ZN(n7740) );
  NAND2_X1 U8951 ( .A1(n14221), .A2(n10418), .ZN(n14204) );
  NAND2_X1 U8952 ( .A1(n14246), .A2(n10417), .ZN(n14223) );
  NAND2_X1 U8953 ( .A1(n7751), .A2(n10353), .ZN(n14296) );
  NAND2_X1 U8954 ( .A1(n10352), .A2(n10351), .ZN(n14304) );
  INV_X1 U8955 ( .A(n6910), .ZN(n12812) );
  AOI21_X1 U8956 ( .B1(n12670), .B2(n12672), .A(n6913), .ZN(n6910) );
  NAND2_X1 U8957 ( .A1(n7578), .A2(n10408), .ZN(n12671) );
  NAND2_X1 U8958 ( .A1(n7755), .A2(n10347), .ZN(n12572) );
  NAND2_X1 U8959 ( .A1(n10827), .A2(n8834), .ZN(n8623) );
  NAND2_X1 U8960 ( .A1(n6869), .A2(n6870), .ZN(n12056) );
  NAND2_X1 U8961 ( .A1(n11928), .A2(n10337), .ZN(n11909) );
  NAND2_X1 U8962 ( .A1(n6795), .A2(n6794), .ZN(n11941) );
  NAND2_X1 U8963 ( .A1(n14323), .A2(n11641), .ZN(n6794) );
  OR2_X1 U8964 ( .A1(n14326), .A2(n6796), .ZN(n6795) );
  OAI22_X1 U8965 ( .A1(n14192), .A2(n11982), .B1(n10330), .B2(n14190), .ZN(
        n11983) );
  OAI21_X1 U8966 ( .B1(n14192), .B2(n10330), .A(n11597), .ZN(n11620) );
  INV_X1 U8967 ( .A(n14180), .ZN(n14599) );
  INV_X1 U8968 ( .A(n14313), .ZN(n14617) );
  INV_X1 U8969 ( .A(n15624), .ZN(n12375) );
  AND2_X1 U8970 ( .A1(n7579), .A2(n8888), .ZN(n6866) );
  INV_X1 U8971 ( .A(n8949), .ZN(n14635) );
  NAND2_X1 U8972 ( .A1(n8901), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8543) );
  INV_X1 U8973 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11021) );
  INV_X1 U8974 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n11025) );
  XNOR2_X1 U8975 ( .A(n8651), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11462) );
  INV_X1 U8976 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10880) );
  INV_X1 U8977 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10828) );
  INV_X1 U8978 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10814) );
  INV_X1 U8979 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10810) );
  INV_X1 U8980 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10806) );
  INV_X1 U8981 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10812) );
  NAND2_X1 U8982 ( .A1(n8557), .A2(n8572), .ZN(n11071) );
  NAND2_X1 U8983 ( .A1(n8554), .A2(n6710), .ZN(n13983) );
  INV_X1 U8984 ( .A(n6711), .ZN(n6710) );
  OAI21_X1 U8985 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(P2_IR_REG_1__SCAN_IN), .A(
        n6712), .ZN(n6711) );
  NAND2_X1 U8986 ( .A1(n11902), .A2(n11901), .ZN(n11900) );
  NAND2_X1 U8987 ( .A1(n11816), .A2(n10144), .ZN(n11902) );
  NAND2_X1 U8988 ( .A1(n6940), .A2(n6938), .ZN(n12961) );
  AND2_X1 U8989 ( .A1(n6939), .A2(n7683), .ZN(n6938) );
  AOI21_X1 U8990 ( .B1(n7684), .B2(n7686), .A(n6527), .ZN(n7683) );
  AND3_X2 U8991 ( .A1(n9637), .A2(n9636), .A3(n9635), .ZN(n11545) );
  NAND2_X1 U8992 ( .A1(n12968), .A2(n10109), .ZN(n11538) );
  NAND2_X1 U8993 ( .A1(n6925), .A2(n7056), .ZN(n6924) );
  INV_X1 U8994 ( .A(n10099), .ZN(n7056) );
  OR2_X1 U8995 ( .A1(n14731), .A2(n7689), .ZN(n14688) );
  INV_X1 U8996 ( .A(n12624), .ZN(n7694) );
  INV_X1 U8997 ( .A(n7695), .ZN(n12625) );
  NAND2_X1 U8998 ( .A1(n7242), .A2(n14782), .ZN(n14707) );
  NAND2_X1 U8999 ( .A1(n9904), .A2(n9903), .ZN(n15099) );
  NAND2_X1 U9000 ( .A1(n12108), .A2(n9902), .ZN(n9904) );
  NAND2_X1 U9001 ( .A1(n14680), .A2(n10240), .ZN(n14733) );
  INV_X1 U9002 ( .A(n6929), .ZN(n14752) );
  AOI21_X1 U9003 ( .B1(n14680), .B2(n6931), .A(n7688), .ZN(n6929) );
  NOR2_X1 U9004 ( .A1(n7689), .A2(n6932), .ZN(n6931) );
  INV_X1 U9005 ( .A(n7674), .ZN(n14764) );
  AOI21_X1 U9006 ( .B1(n14707), .B2(n7680), .A(n7678), .ZN(n7674) );
  NAND2_X1 U9007 ( .A1(n6680), .A2(n9674), .ZN(n11886) );
  INV_X1 U9008 ( .A(n14776), .ZN(n14792) );
  AND2_X1 U9009 ( .A1(n10314), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11490) );
  NAND2_X1 U9010 ( .A1(n10694), .A2(n10649), .ZN(n10685) );
  INV_X1 U9011 ( .A(n10683), .ZN(n10684) );
  NAND2_X1 U9012 ( .A1(n9934), .A2(n9933), .ZN(n15037) );
  NAND2_X1 U9013 ( .A1(n9923), .A2(n9922), .ZN(n15090) );
  OR2_X1 U9014 ( .A1(n15078), .A2(n6429), .ZN(n9923) );
  NAND2_X1 U9015 ( .A1(n9867), .A2(n9866), .ZN(n15122) );
  OR2_X1 U9016 ( .A1(n15149), .A2(n6429), .ZN(n9867) );
  NAND2_X1 U9017 ( .A1(n9878), .A2(n9877), .ZN(n14804) );
  OR2_X1 U9018 ( .A1(n15169), .A2(n6429), .ZN(n9878) );
  OR2_X1 U9019 ( .A1(n9790), .A2(n9789), .ZN(n15256) );
  OR2_X1 U9020 ( .A1(n9614), .A2(n10936), .ZN(n9615) );
  OR2_X1 U9021 ( .A1(n9691), .A2(n9609), .ZN(n9610) );
  NAND2_X1 U9022 ( .A1(n6726), .A2(n10916), .ZN(n15503) );
  NAND2_X1 U9023 ( .A1(n14866), .A2(n14865), .ZN(n6726) );
  NAND2_X1 U9024 ( .A1(n14875), .A2(n6727), .ZN(n14908) );
  AND2_X1 U9025 ( .A1(n6729), .A2(n10921), .ZN(n6727) );
  INV_X1 U9026 ( .A(n10922), .ZN(n6729) );
  AND2_X1 U9027 ( .A1(n14910), .A2(n10927), .ZN(n10958) );
  NOR2_X1 U9028 ( .A1(n10960), .A2(n10959), .ZN(n14919) );
  NOR2_X1 U9029 ( .A1(n11264), .A2(n11263), .ZN(n11266) );
  NOR2_X1 U9030 ( .A1(n11658), .A2(n6735), .ZN(n12121) );
  OR2_X1 U9031 ( .A1(n11660), .A2(n11657), .ZN(n6735) );
  XNOR2_X1 U9032 ( .A(n7058), .B(n12127), .ZN(n14939) );
  NOR2_X1 U9033 ( .A1(n14954), .A2(n7022), .ZN(n14971) );
  NAND2_X1 U9034 ( .A1(n10611), .A2(n10610), .ZN(n15012) );
  XNOR2_X1 U9035 ( .A(n7529), .B(n10665), .ZN(n9985) );
  NAND2_X1 U9036 ( .A1(n7730), .A2(n7723), .ZN(n7721) );
  AND2_X1 U9037 ( .A1(n10665), .A2(n7729), .ZN(n7723) );
  OAI21_X1 U9038 ( .B1(n10665), .B2(n7726), .A(n7725), .ZN(n7724) );
  NAND2_X1 U9039 ( .A1(n10665), .A2(n10030), .ZN(n7725) );
  NOR2_X1 U9040 ( .A1(n7729), .A2(n7727), .ZN(n7726) );
  NOR2_X1 U9041 ( .A1(n15050), .A2(n15160), .ZN(n15295) );
  NAND2_X1 U9042 ( .A1(n9915), .A2(n9914), .ZN(n15298) );
  NAND2_X1 U9043 ( .A1(n12241), .A2(n9902), .ZN(n9915) );
  NAND2_X1 U9044 ( .A1(n15123), .A2(n9891), .ZN(n15106) );
  AND2_X1 U9045 ( .A1(n9885), .A2(n9907), .ZN(n15133) );
  OAI21_X1 U9046 ( .B1(n15178), .B2(n6441), .A(n7277), .ZN(n15145) );
  NAND2_X1 U9047 ( .A1(n7281), .A2(n7280), .ZN(n15165) );
  NAND2_X1 U9048 ( .A1(n15261), .A2(n7532), .ZN(n15237) );
  NAND2_X1 U9049 ( .A1(n12711), .A2(n12710), .ZN(n12709) );
  NAND2_X1 U9050 ( .A1(n12555), .A2(n10007), .ZN(n12711) );
  NAND2_X1 U9051 ( .A1(n11024), .A2(n9902), .ZN(n7288) );
  AND2_X1 U9052 ( .A1(n7534), .A2(n6495), .ZN(n12429) );
  OAI21_X1 U9053 ( .B1(n12188), .B2(n7735), .A(n7733), .ZN(n12331) );
  NAND2_X1 U9054 ( .A1(n12187), .A2(n10005), .ZN(n12333) );
  CLKBUF_X1 U9055 ( .A(n12147), .Z(n12196) );
  INV_X1 U9056 ( .A(n15234), .ZN(n15524) );
  OR2_X1 U9057 ( .A1(n15533), .A2(n15354), .ZN(n15248) );
  NAND2_X1 U9058 ( .A1(n15284), .A2(n15370), .ZN(n6686) );
  INV_X1 U9059 ( .A(n15285), .ZN(n6685) );
  INV_X1 U9060 ( .A(n15099), .ZN(n15396) );
  AOI21_X1 U9061 ( .B1(n15317), .B2(n15370), .A(n15316), .ZN(n6819) );
  NAND2_X1 U9062 ( .A1(n9732), .A2(n9731), .ZN(n14674) );
  NAND2_X1 U9063 ( .A1(n9703), .A2(n9702), .ZN(n12220) );
  INV_X1 U9064 ( .A(n9589), .ZN(n15428) );
  CLKBUF_X1 U9065 ( .A(n9986), .Z(n14836) );
  NAND2_X1 U9066 ( .A1(n6990), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10042) );
  NAND2_X1 U9067 ( .A1(n9976), .A2(n7248), .ZN(n6990) );
  NAND2_X1 U9068 ( .A1(n8796), .A2(n8795), .ZN(n8798) );
  XNOR2_X1 U9069 ( .A(n9883), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15437) );
  INV_X1 U9070 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n11103) );
  INV_X1 U9071 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10878) );
  INV_X1 U9072 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10830) );
  INV_X1 U9073 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10792) );
  XNOR2_X1 U9074 ( .A(n9644), .B(P1_IR_REG_4__SCAN_IN), .ZN(n15507) );
  OAI21_X1 U9075 ( .B1(n10817), .B2(n10798), .A(n7052), .ZN(n8547) );
  NAND2_X1 U9076 ( .A1(n10817), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7052) );
  NAND2_X1 U9077 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6731) );
  NAND2_X1 U9078 ( .A1(n9611), .A2(n15422), .ZN(n6730) );
  NAND2_X1 U9079 ( .A1(n6897), .A2(n10770), .ZN(n10782) );
  XNOR2_X1 U9080 ( .A(n10803), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n10802) );
  NAND2_X1 U9081 ( .A1(n10994), .A2(n6882), .ZN(n6886) );
  AND2_X1 U9082 ( .A1(n6885), .A2(n6884), .ZN(n6883) );
  AND2_X1 U9083 ( .A1(n10993), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6882) );
  NAND2_X1 U9084 ( .A1(n10995), .A2(n10996), .ZN(n11305) );
  XNOR2_X1 U9085 ( .A(n11648), .B(n11646), .ZN(n11312) );
  NAND2_X1 U9086 ( .A1(n11790), .A2(n7111), .ZN(n7110) );
  INV_X1 U9087 ( .A(n7112), .ZN(n7108) );
  NOR2_X1 U9088 ( .A1(n12838), .A2(n12837), .ZN(n12839) );
  NAND2_X1 U9089 ( .A1(n6891), .A2(n7289), .ZN(n15462) );
  INV_X1 U9090 ( .A(n7290), .ZN(n7289) );
  NAND2_X1 U9091 ( .A1(n6890), .A2(n6888), .ZN(n6891) );
  OAI21_X1 U9092 ( .B1(n7293), .B2(n7291), .A(n15459), .ZN(n7290) );
  NAND2_X1 U9093 ( .A1(n7118), .A2(n7292), .ZN(n7117) );
  INV_X1 U9094 ( .A(n15459), .ZN(n7118) );
  OR2_X1 U9095 ( .A1(n12864), .A2(n12863), .ZN(n6893) );
  NAND2_X1 U9096 ( .A1(n11583), .A2(n11582), .ZN(n11588) );
  NAND2_X1 U9097 ( .A1(n13184), .A2(n7171), .ZN(n6765) );
  NAND2_X1 U9098 ( .A1(n6426), .A2(n7886), .ZN(n12655) );
  AOI21_X1 U9099 ( .B1(n7972), .B2(n13509), .A(n7971), .ZN(n7005) );
  NAND2_X1 U9100 ( .A1(n7499), .A2(n13495), .ZN(n7089) );
  NAND2_X1 U9101 ( .A1(n7634), .A2(n7002), .ZN(P3_U3204) );
  OR2_X1 U9102 ( .A1(n9566), .A2(n13663), .ZN(n7634) );
  INV_X1 U9103 ( .A(n9351), .ZN(n7633) );
  OAI21_X1 U9104 ( .B1(n13742), .B2(n15731), .A(n8528), .ZN(P3_U3486) );
  OAI22_X1 U9105 ( .A1(n13744), .A2(n13709), .B1(n15734), .B2(n8526), .ZN(
        n8527) );
  OAI21_X1 U9106 ( .B1(n13742), .B2(n15721), .A(n7013), .ZN(P3_U3454) );
  INV_X1 U9107 ( .A(n7014), .ZN(n7013) );
  OAI22_X1 U9108 ( .A1(n13744), .A2(n13790), .B1(n15722), .B2(n13743), .ZN(
        n7014) );
  OAI222_X1 U9109 ( .A1(P3_U3151), .A2(n11041), .B1(n13808), .B2(n10834), .C1(
        n10833), .C2(n13805), .ZN(P3_U3290) );
  OAI21_X1 U9110 ( .B1(n14099), .B2(n13925), .A(n9298), .ZN(n9299) );
  NAND2_X1 U9111 ( .A1(n7405), .A2(n8995), .ZN(n11640) );
  OAI211_X1 U9112 ( .C1(n6701), .C2(n11455), .A(n6699), .B(n6696), .ZN(
        P2_U3233) );
  NOR2_X1 U9113 ( .A1(n6698), .A2(n6697), .ZN(n6696) );
  AOI21_X1 U9114 ( .B1(n14069), .B2(n15610), .A(n6702), .ZN(n6701) );
  NAND2_X1 U9115 ( .A1(n6700), .A2(n11455), .ZN(n6699) );
  INV_X1 U9116 ( .A(n10469), .ZN(n10470) );
  OAI21_X1 U9117 ( .B1(n14354), .B2(n14312), .A(n10468), .ZN(n10469) );
  AOI21_X1 U9118 ( .B1(n6457), .B2(n15630), .A(n14090), .ZN(n14091) );
  NOR2_X1 U9119 ( .A1(n15670), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7025) );
  NAND2_X1 U9120 ( .A1(n6534), .A2(n6445), .ZN(n6976) );
  OAI21_X1 U9121 ( .B1(n10441), .B2(n15668), .A(n6920), .ZN(P2_U3527) );
  NOR2_X1 U9122 ( .A1(n6503), .A2(n6921), .ZN(n6920) );
  NOR2_X1 U9123 ( .A1(n15670), .A2(n10438), .ZN(n6921) );
  NOR2_X1 U9124 ( .A1(n15666), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7027) );
  NAND2_X1 U9125 ( .A1(n7543), .A2(n6611), .ZN(n7544) );
  NAND2_X1 U9126 ( .A1(n6445), .A2(n6991), .ZN(n7543) );
  XNOR2_X1 U9127 ( .A(n7240), .B(n7239), .ZN(n14781) );
  MUX2_X1 U9128 ( .A(n14995), .B(n14994), .S(n14993), .Z(n14997) );
  OAI21_X1 U9129 ( .B1(n15384), .B2(n15552), .A(n6859), .ZN(P1_U3555) );
  AOI21_X1 U9130 ( .B1(n15042), .B2(n12686), .A(n6860), .ZN(n6859) );
  NOR2_X1 U9131 ( .A1(n15554), .A2(n15290), .ZN(n6860) );
  NAND2_X1 U9132 ( .A1(n10626), .A2(n12478), .ZN(n10073) );
  OAI21_X1 U9133 ( .B1(n15381), .B2(n15549), .A(n7155), .ZN(P1_U3524) );
  INV_X1 U9134 ( .A(n7156), .ZN(n7155) );
  OAI22_X1 U9135 ( .A1(n15383), .A2(n10072), .B1(n15550), .B2(n15382), .ZN(
        n7156) );
  OAI21_X1 U9136 ( .B1(n15384), .B2(n15549), .A(n7138), .ZN(P1_U3523) );
  INV_X1 U9137 ( .A(n7139), .ZN(n7138) );
  OAI22_X1 U9138 ( .A1(n7759), .A2(n10072), .B1(n15550), .B2(n15385), .ZN(
        n7139) );
  NAND2_X1 U9139 ( .A1(n11794), .A2(n7114), .ZN(n11946) );
  NAND2_X1 U9140 ( .A1(n7301), .A2(n12499), .ZN(n12824) );
  NAND2_X1 U9141 ( .A1(n12495), .A2(n15584), .ZN(n7301) );
  AOI21_X1 U9142 ( .B1(n15474), .B2(n15473), .A(n15472), .ZN(n15482) );
  INV_X1 U9143 ( .A(n6893), .ZN(n15442) );
  NOR2_X1 U9144 ( .A1(n13181), .A2(n12995), .ZN(n6436) );
  AND2_X1 U9145 ( .A1(n13611), .A2(n7650), .ZN(n6437) );
  NAND2_X1 U9146 ( .A1(n13503), .A2(n6750), .ZN(n13476) );
  INV_X1 U9147 ( .A(n13476), .ZN(n6749) );
  OAI21_X1 U9148 ( .B1(n9846), .B2(n7791), .A(n9979), .ZN(n11458) );
  NAND2_X1 U9149 ( .A1(n7345), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7342) );
  NAND2_X1 U9150 ( .A1(n14356), .A2(n14110), .ZN(n6438) );
  OR2_X1 U9151 ( .A1(n12790), .A2(n13376), .ZN(n13121) );
  INV_X1 U9152 ( .A(n15042), .ZN(n7759) );
  AND2_X1 U9153 ( .A1(n8108), .A2(n8107), .ZN(n6439) );
  AND2_X1 U9154 ( .A1(n12248), .A2(n7737), .ZN(n6440) );
  NAND2_X1 U9155 ( .A1(n6489), .A2(n7488), .ZN(n7881) );
  OR2_X1 U9156 ( .A1(n7279), .A2(n7736), .ZN(n6441) );
  AND2_X1 U9157 ( .A1(n7319), .A2(n7999), .ZN(n6442) );
  OR2_X1 U9158 ( .A1(n10383), .A2(n14305), .ZN(n6443) );
  INV_X1 U9159 ( .A(n14157), .ZN(n7571) );
  OR2_X1 U9160 ( .A1(n14355), .A2(n14575), .ZN(n6445) );
  AND2_X1 U9161 ( .A1(n12825), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6446) );
  NAND2_X1 U9162 ( .A1(n7656), .A2(n13038), .ZN(n6447) );
  NAND2_X1 U9163 ( .A1(n8653), .A2(n8652), .ZN(n12735) );
  INV_X1 U9164 ( .A(n12710), .ZN(n12714) );
  AND2_X1 U9165 ( .A1(n10895), .A2(n11226), .ZN(n6448) );
  XNOR2_X1 U9166 ( .A(n15053), .B(n15037), .ZN(n10662) );
  NAND2_X1 U9167 ( .A1(n7411), .A2(n9152), .ZN(n13887) );
  AND2_X1 U9168 ( .A1(n10817), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6449) );
  NAND2_X1 U9169 ( .A1(n9925), .A2(n9924), .ZN(n15053) );
  INV_X1 U9170 ( .A(n15053), .ZN(n7758) );
  AND2_X1 U9171 ( .A1(n7578), .A2(n7576), .ZN(n6450) );
  AND2_X1 U9172 ( .A1(n6776), .A2(n13033), .ZN(n6451) );
  AND2_X1 U9173 ( .A1(n6558), .A2(n7216), .ZN(n6452) );
  AND2_X1 U9174 ( .A1(n7207), .A2(n7202), .ZN(n6453) );
  AND2_X1 U9175 ( .A1(n7961), .A2(n6599), .ZN(n6454) );
  AND2_X1 U9176 ( .A1(n7664), .A2(n13146), .ZN(n6455) );
  AND2_X1 U9177 ( .A1(n11042), .A2(n6507), .ZN(n6456) );
  AND2_X1 U9178 ( .A1(n10445), .A2(n10376), .ZN(n6457) );
  NOR2_X1 U9179 ( .A1(n12994), .A2(n12993), .ZN(n6458) );
  INV_X1 U9180 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n8065) );
  NAND2_X1 U9181 ( .A1(n11585), .A2(n11782), .ZN(n11777) );
  AND2_X1 U9182 ( .A1(n10113), .A2(n10109), .ZN(n6459) );
  AND2_X1 U9183 ( .A1(n6563), .A2(n6837), .ZN(n6460) );
  AND2_X1 U9184 ( .A1(n14608), .A2(n7618), .ZN(n6461) );
  NAND2_X1 U9185 ( .A1(n14068), .A2(n15613), .ZN(n6462) );
  AND2_X1 U9186 ( .A1(n7630), .A2(n7629), .ZN(n6463) );
  INV_X1 U9187 ( .A(n9450), .ZN(n7385) );
  INV_X1 U9188 ( .A(n15251), .ZN(n15262) );
  NAND2_X1 U9189 ( .A1(n10530), .A2(n10533), .ZN(n15251) );
  INV_X1 U9190 ( .A(n12609), .ZN(n7612) );
  AND3_X1 U9191 ( .A1(n6426), .A2(n7886), .A3(P3_REG1_REG_11__SCAN_IN), .ZN(
        n6464) );
  AND2_X1 U9192 ( .A1(n13416), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n6465) );
  AND3_X1 U9193 ( .A1(n7349), .A2(n7991), .A3(P3_REG2_REG_11__SCAN_IN), .ZN(
        n6466) );
  AND2_X1 U9194 ( .A1(n13413), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n6467) );
  INV_X1 U9195 ( .A(n13371), .ZN(n13552) );
  NAND2_X1 U9196 ( .A1(n8455), .A2(n8454), .ZN(n13371) );
  AND2_X1 U9197 ( .A1(n7229), .A2(n7228), .ZN(n6468) );
  AND2_X1 U9198 ( .A1(n14740), .A2(n10199), .ZN(n6469) );
  INV_X1 U9199 ( .A(n15548), .ZN(n7767) );
  INV_X1 U9200 ( .A(n13186), .ZN(n7172) );
  AND2_X1 U9201 ( .A1(n7322), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6470) );
  INV_X1 U9202 ( .A(n9464), .ZN(n9258) );
  NAND2_X1 U9203 ( .A1(n7498), .A2(n11344), .ZN(n11198) );
  INV_X1 U9204 ( .A(n14809), .ZN(n7287) );
  OAI21_X1 U9205 ( .B1(n14258), .B2(n6917), .A(n6914), .ZN(n14176) );
  INV_X1 U9206 ( .A(n11931), .ZN(n6872) );
  AND2_X1 U9207 ( .A1(n7414), .A2(n9152), .ZN(n6471) );
  AND2_X1 U9208 ( .A1(n10375), .A2(n7256), .ZN(n6472) );
  NAND4_X1 U9209 ( .A1(n8121), .A2(n8120), .A3(n8118), .A4(n8119), .ZN(n13723)
         );
  NAND2_X1 U9210 ( .A1(n6775), .A2(n6451), .ZN(n13592) );
  NAND2_X1 U9211 ( .A1(n12803), .A2(n9129), .ZN(n13878) );
  CLKBUF_X3 U9212 ( .A(n10786), .Z(n6978) );
  NOR2_X1 U9213 ( .A1(n14298), .A2(n14275), .ZN(n14251) );
  OR2_X1 U9214 ( .A1(n15054), .A2(n7757), .ZN(n10032) );
  NAND2_X1 U9215 ( .A1(n7747), .A2(n7745), .ZN(n14103) );
  NAND2_X2 U9216 ( .A1(n8950), .A2(n14635), .ZN(n8984) );
  NAND2_X1 U9217 ( .A1(n12713), .A2(n12714), .ZN(n12712) );
  NAND2_X1 U9218 ( .A1(n8460), .A2(n7453), .ZN(n6473) );
  AND2_X1 U9219 ( .A1(n12557), .A2(n6849), .ZN(n6474) );
  NOR2_X1 U9220 ( .A1(n7403), .A2(n7402), .ZN(n6475) );
  NOR2_X1 U9221 ( .A1(n15565), .A2(n15566), .ZN(n6476) );
  NAND2_X1 U9222 ( .A1(n13018), .A2(n7639), .ZN(n6477) );
  NAND2_X1 U9223 ( .A1(n8754), .A2(n8753), .ZN(n14537) );
  NAND2_X1 U9224 ( .A1(n12409), .A2(n13971), .ZN(n6478) );
  NAND4_X1 U9225 ( .A1(n9650), .A2(n9649), .A3(n9648), .A4(n9647), .ZN(n14818)
         );
  AND2_X1 U9226 ( .A1(n12528), .A2(n13381), .ZN(n6479) );
  NOR2_X1 U9227 ( .A1(n12609), .A2(n13969), .ZN(n6480) );
  AND2_X1 U9228 ( .A1(n10232), .A2(n10231), .ZN(n6481) );
  AND2_X1 U9229 ( .A1(n9274), .A2(n11815), .ZN(n14310) );
  AND2_X1 U9230 ( .A1(n7509), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n6482) );
  AND2_X1 U9231 ( .A1(n7333), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U9232 ( .A1(n9040), .A2(n9039), .ZN(n6484) );
  AND2_X1 U9233 ( .A1(n7314), .A2(n10740), .ZN(n6485) );
  XNOR2_X1 U9234 ( .A(n14113), .B(n14125), .ZN(n14111) );
  INV_X1 U9235 ( .A(n7688), .ZN(n7687) );
  OAI21_X1 U9236 ( .B1(n7689), .B2(n14734), .A(n10251), .ZN(n7688) );
  AND2_X1 U9237 ( .A1(n9178), .A2(n9179), .ZN(n13833) );
  INV_X1 U9238 ( .A(n9355), .ZN(n13856) );
  NAND2_X1 U9239 ( .A1(n6488), .A2(n8960), .ZN(n9355) );
  AND2_X1 U9240 ( .A1(n7613), .A2(n7612), .ZN(n6486) );
  OR2_X1 U9241 ( .A1(n10330), .A2(n13859), .ZN(n6487) );
  AND3_X1 U9242 ( .A1(n8959), .A2(n8958), .A3(n8961), .ZN(n6488) );
  OR2_X1 U9243 ( .A1(n11346), .A2(n7491), .ZN(n6489) );
  NAND2_X1 U9244 ( .A1(n8597), .A2(n8596), .ZN(n11914) );
  XNOR2_X1 U9245 ( .A(n9981), .B(n9980), .ZN(n11775) );
  NAND2_X1 U9246 ( .A1(n8066), .A2(n7227), .ZN(n6490) );
  NOR2_X1 U9247 ( .A1(n15151), .A2(n15122), .ZN(n6491) );
  AND2_X1 U9248 ( .A1(n7333), .A2(n11041), .ZN(n6492) );
  NAND2_X1 U9249 ( .A1(n14751), .A2(n10256), .ZN(n14658) );
  NAND2_X1 U9250 ( .A1(n9113), .A2(n9112), .ZN(n6493) );
  AND2_X1 U9251 ( .A1(n7453), .A2(n7807), .ZN(n6494) );
  INV_X1 U9252 ( .A(n15192), .ZN(n7149) );
  OR2_X1 U9253 ( .A1(n12420), .A2(n12427), .ZN(n6495) );
  INV_X1 U9254 ( .A(n15177), .ZN(n7736) );
  INV_X1 U9255 ( .A(n10330), .ZN(n9353) );
  XNOR2_X1 U9256 ( .A(n7850), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11529) );
  XNOR2_X1 U9257 ( .A(n15023), .B(n15038), .ZN(n15017) );
  INV_X1 U9258 ( .A(n15017), .ZN(n7729) );
  AND4_X1 U9259 ( .A1(n8932), .A2(n8898), .A3(n8896), .A4(n8540), .ZN(n6496)
         );
  INV_X1 U9260 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7708) );
  NAND4_X1 U9261 ( .A1(n9580), .A2(n15490), .A3(n9633), .A4(n14414), .ZN(n9974) );
  INV_X1 U9262 ( .A(n9974), .ZN(n9792) );
  NAND3_X2 U9263 ( .A1(n9628), .A2(n9627), .A3(n9626), .ZN(n11259) );
  INV_X1 U9264 ( .A(n10374), .ZN(n7258) );
  NAND2_X1 U9265 ( .A1(n13171), .A2(n13169), .ZN(n13520) );
  INV_X1 U9266 ( .A(n13520), .ZN(n7162) );
  OR2_X1 U9267 ( .A1(n13762), .A2(n13320), .ZN(n6497) );
  NAND2_X1 U9268 ( .A1(n13034), .A2(n13035), .ZN(n13611) );
  NAND2_X1 U9269 ( .A1(n13151), .A2(n8416), .ZN(n13580) );
  INV_X1 U9270 ( .A(n13580), .ZN(n7645) );
  INV_X1 U9271 ( .A(n9452), .ZN(n6954) );
  NAND2_X1 U9272 ( .A1(n9307), .A2(n9306), .ZN(n9309) );
  XNOR2_X1 U9273 ( .A(n15042), .B(n14801), .ZN(n10650) );
  INV_X1 U9274 ( .A(n12355), .ZN(n7441) );
  INV_X1 U9275 ( .A(n13002), .ZN(n7218) );
  NAND2_X1 U9276 ( .A1(n9253), .A2(n9252), .ZN(n6498) );
  INV_X1 U9277 ( .A(n10499), .ZN(n7370) );
  INV_X1 U9278 ( .A(n10600), .ZN(n7387) );
  XNOR2_X1 U9279 ( .A(n8817), .B(SI_24_), .ZN(n8815) );
  AND2_X1 U9280 ( .A1(n15040), .A2(n15039), .ZN(n6499) );
  OR2_X1 U9281 ( .A1(n13455), .A2(n7344), .ZN(n6500) );
  INV_X1 U9282 ( .A(n10735), .ZN(n7333) );
  AND2_X1 U9283 ( .A1(n7248), .A2(n10040), .ZN(n6501) );
  INV_X1 U9284 ( .A(n13859), .ZN(n11690) );
  NAND2_X1 U9285 ( .A1(n8549), .A2(n7619), .ZN(n13859) );
  NAND2_X1 U9286 ( .A1(n8829), .A2(n8828), .ZN(n14113) );
  INV_X1 U9287 ( .A(n14113), .ZN(n7629) );
  NAND2_X1 U9288 ( .A1(n9432), .A2(n7371), .ZN(n6502) );
  NOR2_X1 U9289 ( .A1(n7609), .A2(n14582), .ZN(n6503) );
  XOR2_X1 U9290 ( .A(n13032), .B(n13031), .Z(n6504) );
  INV_X1 U9291 ( .A(n14102), .ZN(n10373) );
  XNOR2_X1 U9292 ( .A(n14356), .B(n13961), .ZN(n14102) );
  AND2_X1 U9293 ( .A1(n12900), .A2(n13374), .ZN(n6505) );
  AND2_X1 U9294 ( .A1(n7639), .A2(n12076), .ZN(n6506) );
  AND2_X1 U9295 ( .A1(n6978), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6507) );
  AND2_X1 U9296 ( .A1(n10351), .A2(n7752), .ZN(n6508) );
  INV_X1 U9297 ( .A(n12567), .ZN(n12755) );
  NAND2_X1 U9298 ( .A1(n6716), .A2(n9757), .ZN(n12567) );
  XNOR2_X1 U9299 ( .A(n8647), .B(SI_9_), .ZN(n8645) );
  XOR2_X1 U9300 ( .A(n13732), .B(n12935), .Z(n6509) );
  AND2_X1 U9301 ( .A1(n7568), .A2(n10423), .ZN(n6510) );
  OR2_X1 U9302 ( .A1(n10555), .A2(n10554), .ZN(n6511) );
  INV_X1 U9303 ( .A(n8626), .ZN(n7482) );
  AND2_X1 U9304 ( .A1(n8701), .A2(n8700), .ZN(n6512) );
  INV_X1 U9305 ( .A(n7477), .ZN(n7476) );
  AND2_X1 U9306 ( .A1(n12910), .A2(n13615), .ZN(n6513) );
  INV_X1 U9307 ( .A(n10429), .ZN(n7558) );
  NAND2_X1 U9308 ( .A1(n11485), .A2(n9357), .ZN(n6514) );
  AND2_X1 U9309 ( .A1(n15351), .A2(n14791), .ZN(n6515) );
  AND2_X1 U9310 ( .A1(n7417), .A2(n7415), .ZN(n6516) );
  INV_X1 U9311 ( .A(n10502), .ZN(n6838) );
  NOR2_X1 U9312 ( .A1(n15230), .A2(n15345), .ZN(n7772) );
  INV_X1 U9313 ( .A(n7616), .ZN(n14230) );
  NOR2_X1 U9314 ( .A1(n14298), .A2(n7617), .ZN(n7616) );
  AND2_X1 U9315 ( .A1(n15042), .A2(n9950), .ZN(n6517) );
  AND2_X1 U9316 ( .A1(n7481), .A2(n8645), .ZN(n6518) );
  OR2_X1 U9317 ( .A1(n9486), .A2(n9485), .ZN(n6519) );
  NAND2_X1 U9318 ( .A1(n13671), .A2(n13552), .ZN(n13164) );
  INV_X1 U9319 ( .A(n13164), .ZN(n7158) );
  AND2_X1 U9320 ( .A1(n14196), .A2(n14206), .ZN(n6520) );
  AND2_X1 U9321 ( .A1(n6982), .A2(n6981), .ZN(n6521) );
  AND2_X1 U9322 ( .A1(n13756), .A2(n13604), .ZN(n6522) );
  AND2_X1 U9323 ( .A1(n11903), .A2(n15543), .ZN(n6523) );
  INV_X1 U9324 ( .A(n11531), .ZN(n7495) );
  AND2_X1 U9325 ( .A1(n8636), .A2(SI_8_), .ZN(n6524) );
  NOR2_X1 U9326 ( .A1(n9238), .A2(n9237), .ZN(n9239) );
  AND2_X1 U9327 ( .A1(n6483), .A2(n11352), .ZN(n6525) );
  AND2_X1 U9328 ( .A1(n6482), .A2(n11352), .ZN(n6526) );
  AND2_X1 U9329 ( .A1(n10286), .A2(n10285), .ZN(n6527) );
  INV_X1 U9330 ( .A(n7225), .ZN(n13165) );
  OAI211_X1 U9331 ( .C1(n8096), .C2(n9304), .A(n8104), .B(n8103), .ZN(n7225)
         );
  OAI22_X1 U9332 ( .A1(n7710), .A2(n7708), .B1(P1_IR_REG_31__SCAN_IN), .B2(
        P1_IR_REG_30__SCAN_IN), .ZN(n7706) );
  AND2_X1 U9333 ( .A1(n6495), .A2(n9754), .ZN(n6528) );
  INV_X1 U9334 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n15422) );
  INV_X1 U9335 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8766) );
  AND2_X1 U9336 ( .A1(n13278), .A2(n13377), .ZN(n6529) );
  AND2_X1 U9337 ( .A1(n10004), .A2(n9712), .ZN(n12152) );
  AND2_X1 U9338 ( .A1(n8942), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6530) );
  AND2_X1 U9339 ( .A1(n13768), .A2(n13623), .ZN(n6531) );
  AND2_X1 U9340 ( .A1(n7067), .A2(n7656), .ZN(n6532) );
  INV_X1 U9341 ( .A(n10019), .ZN(n7279) );
  NOR2_X1 U9342 ( .A1(n12720), .A2(n14809), .ZN(n6533) );
  AND2_X1 U9343 ( .A1(n14354), .A2(n14353), .ZN(n6534) );
  NOR2_X1 U9344 ( .A1(n14674), .A2(n14812), .ZN(n6535) );
  AND2_X1 U9345 ( .A1(n7411), .A2(n6471), .ZN(n6536) );
  NOR2_X1 U9346 ( .A1(n10150), .A2(n10149), .ZN(n6537) );
  NOR2_X1 U9347 ( .A1(n15042), .A2(n14801), .ZN(n6538) );
  OR2_X1 U9348 ( .A1(n13148), .A2(n13580), .ZN(n6539) );
  INV_X1 U9349 ( .A(n7539), .ZN(n7538) );
  NAND2_X1 U9350 ( .A1(n7736), .A2(n10562), .ZN(n7539) );
  AND2_X1 U9351 ( .A1(n6952), .A2(n6954), .ZN(n6540) );
  AND2_X1 U9352 ( .A1(n11080), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6541) );
  AND2_X1 U9353 ( .A1(n7636), .A2(n13122), .ZN(n6542) );
  NOR2_X1 U9354 ( .A1(n14731), .A2(n10247), .ZN(n6543) );
  INV_X1 U9355 ( .A(n7551), .ZN(n7550) );
  NAND2_X1 U9356 ( .A1(n14229), .A2(n10417), .ZN(n7551) );
  NOR2_X1 U9357 ( .A1(n13653), .A2(n7205), .ZN(n7204) );
  OR2_X1 U9358 ( .A1(n7551), .A2(n7549), .ZN(n6544) );
  AND2_X1 U9359 ( .A1(n13712), .A2(n13654), .ZN(n6545) );
  AND2_X1 U9360 ( .A1(n15298), .A2(n15090), .ZN(n6546) );
  NAND2_X1 U9361 ( .A1(n8460), .A2(n8462), .ZN(n6547) );
  AND2_X1 U9362 ( .A1(n11571), .A2(n12064), .ZN(n6548) );
  OR2_X1 U9363 ( .A1(n14393), .A2(n14189), .ZN(n6549) );
  OR2_X1 U9364 ( .A1(n7437), .A2(n6479), .ZN(n6550) );
  INV_X1 U9365 ( .A(n7332), .ZN(n7329) );
  NOR2_X1 U9366 ( .A1(n8188), .A2(n7985), .ZN(n7332) );
  INV_X1 U9367 ( .A(n7508), .ZN(n7505) );
  NOR2_X1 U9368 ( .A1(n8188), .A2(n15729), .ZN(n7508) );
  AND2_X1 U9369 ( .A1(n9309), .A2(n13370), .ZN(n6551) );
  INV_X1 U9370 ( .A(n12764), .ZN(n7521) );
  AND2_X1 U9371 ( .A1(n10365), .A2(n10364), .ZN(n6552) );
  OR2_X1 U9372 ( .A1(n12462), .A2(n12463), .ZN(n6553) );
  INV_X1 U9373 ( .A(n7134), .ZN(n7133) );
  NAND2_X1 U9374 ( .A1(n12805), .A2(n6493), .ZN(n7134) );
  INV_X1 U9375 ( .A(n7546), .ZN(n6877) );
  NAND2_X1 U9376 ( .A1(n6549), .A2(n7547), .ZN(n7546) );
  NAND2_X1 U9377 ( .A1(n8407), .A2(n8406), .ZN(n13243) );
  NAND2_X1 U9378 ( .A1(n10009), .A2(n10008), .ZN(n6554) );
  NOR2_X1 U9379 ( .A1(n13789), .A2(n13640), .ZN(n6555) );
  NOR2_X1 U9380 ( .A1(n13401), .A2(n7990), .ZN(n6556) );
  AND2_X1 U9381 ( .A1(n10824), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n6557) );
  AND2_X1 U9382 ( .A1(n13159), .A2(n13160), .ZN(n13557) );
  AND2_X1 U9383 ( .A1(n13043), .A2(n13042), .ZN(n13637) );
  INV_X1 U9384 ( .A(n13637), .ZN(n7207) );
  INV_X1 U9385 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10797) );
  INV_X1 U9386 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10862) );
  NOR2_X1 U9387 ( .A1(n8429), .A2(n7646), .ZN(n6558) );
  INV_X1 U9388 ( .A(n7416), .ZN(n7415) );
  NAND2_X1 U9389 ( .A1(n9199), .A2(n9191), .ZN(n7416) );
  AND2_X1 U9390 ( .A1(n9203), .A2(n9202), .ZN(n6559) );
  INV_X1 U9391 ( .A(n11849), .ZN(n7492) );
  INV_X1 U9392 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10795) );
  INV_X1 U9393 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7913) );
  INV_X1 U9394 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10790) );
  OR2_X1 U9395 ( .A1(n8294), .A2(n8031), .ZN(n6560) );
  AND2_X1 U9396 ( .A1(n15383), .A2(n7759), .ZN(n6561) );
  AND2_X1 U9397 ( .A1(n12344), .A2(n13382), .ZN(n6562) );
  AND2_X1 U9398 ( .A1(n12996), .A2(n13369), .ZN(n13177) );
  INV_X1 U9399 ( .A(n13177), .ZN(n7036) );
  OR2_X1 U9400 ( .A1(n10505), .A2(n10503), .ZN(n6563) );
  AND2_X1 U9401 ( .A1(n14178), .A2(n6463), .ZN(n14095) );
  AND2_X1 U9402 ( .A1(n6485), .A2(n7307), .ZN(n6564) );
  NAND2_X1 U9403 ( .A1(n14122), .A2(n14121), .ZN(n6565) );
  NAND2_X1 U9404 ( .A1(n12999), .A2(n12998), .ZN(n6566) );
  NAND2_X1 U9405 ( .A1(n7327), .A2(n7326), .ZN(n7988) );
  INV_X1 U9406 ( .A(n9431), .ZN(n7371) );
  AOI21_X1 U9407 ( .B1(n15448), .B2(n7293), .A(n7117), .ZN(n15461) );
  INV_X1 U9408 ( .A(n15461), .ZN(n7116) );
  AOI21_X1 U9409 ( .B1(n7877), .B2(n7495), .A(n6557), .ZN(n7494) );
  OR2_X1 U9410 ( .A1(n13756), .A2(n13263), .ZN(n13145) );
  INV_X1 U9411 ( .A(n10584), .ZN(n7376) );
  OR2_X1 U9412 ( .A1(n7218), .A2(n13003), .ZN(n13602) );
  INV_X1 U9413 ( .A(n10581), .ZN(n7378) );
  OR2_X1 U9414 ( .A1(n7957), .A2(n7993), .ZN(n6567) );
  OR2_X1 U9415 ( .A1(n11529), .A2(n12116), .ZN(n6568) );
  OR2_X1 U9416 ( .A1(n11042), .A2(n13983), .ZN(n6569) );
  NOR2_X1 U9417 ( .A1(n12581), .A2(n10181), .ZN(n6570) );
  NOR2_X1 U9418 ( .A1(n12332), .A2(n12420), .ZN(n6571) );
  AND2_X1 U9419 ( .A1(n7148), .A2(n9891), .ZN(n6572) );
  AND2_X1 U9420 ( .A1(n13169), .A2(n13167), .ZN(n6573) );
  AND2_X1 U9421 ( .A1(n13105), .A2(n13099), .ZN(n6574) );
  AND2_X1 U9422 ( .A1(n10768), .A2(n7105), .ZN(n6575) );
  AND2_X1 U9423 ( .A1(n13124), .A2(n13123), .ZN(n6576) );
  NOR2_X1 U9424 ( .A1(n10370), .A2(n7748), .ZN(n6577) );
  NOR2_X1 U9425 ( .A1(n10665), .A2(n7727), .ZN(n6578) );
  AND2_X1 U9426 ( .A1(n7227), .A2(n8067), .ZN(n6579) );
  AND2_X1 U9427 ( .A1(n15448), .A2(n15449), .ZN(n6580) );
  AND2_X1 U9428 ( .A1(n7645), .A2(n7664), .ZN(n6581) );
  AND2_X1 U9429 ( .A1(n9114), .A2(n9105), .ZN(n6582) );
  AND2_X1 U9430 ( .A1(n6747), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n6583) );
  INV_X1 U9431 ( .A(n15404), .ZN(n15132) );
  NAND2_X1 U9432 ( .A1(n15437), .A2(n9632), .ZN(n15404) );
  AND2_X1 U9433 ( .A1(n15261), .A2(n10530), .ZN(n6584) );
  AND2_X1 U9434 ( .A1(n7096), .A2(n9368), .ZN(n6585) );
  INV_X1 U9435 ( .A(n14081), .ZN(n14585) );
  NAND2_X1 U9436 ( .A1(n8858), .A2(n8857), .ZN(n14081) );
  OR2_X1 U9437 ( .A1(n7370), .A2(n10498), .ZN(n6586) );
  OR2_X1 U9438 ( .A1(n10599), .A2(n7387), .ZN(n6587) );
  OR2_X1 U9439 ( .A1(n9443), .A2(n9441), .ZN(n6588) );
  NOR2_X1 U9440 ( .A1(n8710), .A2(n8709), .ZN(n8711) );
  NAND2_X2 U9441 ( .A1(n8841), .A2(n8840), .ZN(n14087) );
  INV_X1 U9442 ( .A(n14087), .ZN(n7609) );
  AND2_X1 U9443 ( .A1(n7654), .A2(n6497), .ZN(n6589) );
  AND2_X1 U9444 ( .A1(n6892), .A2(n15443), .ZN(n6590) );
  AND2_X1 U9445 ( .A1(n7796), .A2(n7778), .ZN(n6591) );
  OR2_X1 U9446 ( .A1(n10513), .A2(n10515), .ZN(n6592) );
  OR2_X1 U9447 ( .A1(n7385), .A2(n9447), .ZN(n6593) );
  AND2_X1 U9448 ( .A1(n7448), .A2(n6763), .ZN(n6594) );
  OR2_X1 U9449 ( .A1(n7383), .A2(n9403), .ZN(n6595) );
  INV_X1 U9450 ( .A(n8666), .ZN(n7456) );
  NAND2_X1 U9451 ( .A1(n8684), .A2(n8661), .ZN(n8666) );
  OR2_X1 U9452 ( .A1(n7675), .A2(n6481), .ZN(n6596) );
  NOR2_X1 U9453 ( .A1(n7678), .A2(n6481), .ZN(n6597) );
  INV_X1 U9454 ( .A(n7788), .ZN(n6878) );
  INV_X1 U9455 ( .A(n7222), .ZN(n7221) );
  NAND2_X1 U9456 ( .A1(n9301), .A2(n13520), .ZN(n7222) );
  INV_X1 U9457 ( .A(n7567), .ZN(n7566) );
  NAND2_X1 U9458 ( .A1(n7571), .A2(n10423), .ZN(n7567) );
  INV_X1 U9459 ( .A(n7446), .ZN(n7445) );
  NAND2_X1 U9460 ( .A1(n7776), .A2(n7447), .ZN(n7446) );
  AND2_X1 U9461 ( .A1(n8764), .A2(n8766), .ZN(n6598) );
  AND2_X1 U9462 ( .A1(n7903), .A2(n6764), .ZN(n6599) );
  NAND2_X1 U9463 ( .A1(n8487), .A2(n8486), .ZN(n13632) );
  INV_X1 U9464 ( .A(n14275), .ZN(n7618) );
  NAND2_X1 U9465 ( .A1(n12212), .A2(n10159), .ZN(n12517) );
  AND2_X1 U9466 ( .A1(n12732), .A2(n14628), .ZN(n12733) );
  NAND2_X1 U9467 ( .A1(n12700), .A2(n12697), .ZN(n12784) );
  NAND2_X1 U9468 ( .A1(n6828), .A2(n7140), .ZN(n12023) );
  NAND2_X1 U9469 ( .A1(n7142), .A2(n9670), .ZN(n11873) );
  NOR2_X1 U9470 ( .A1(n12672), .A2(n7577), .ZN(n7576) );
  AND2_X1 U9471 ( .A1(n8415), .A2(n8414), .ZN(n13569) );
  NAND2_X1 U9472 ( .A1(n8823), .A2(n8822), .ZN(n14135) );
  INV_X1 U9473 ( .A(n14135), .ZN(n7631) );
  AND2_X1 U9474 ( .A1(n12732), .A2(n7613), .ZN(n6600) );
  AND2_X1 U9475 ( .A1(n12565), .A2(n12755), .ZN(n6601) );
  AND2_X1 U9476 ( .A1(n15664), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6602) );
  INV_X1 U9477 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n6752) );
  INV_X1 U9478 ( .A(n14546), .ZN(n6792) );
  AND2_X1 U9479 ( .A1(n7597), .A2(n7198), .ZN(n6603) );
  INV_X1 U9480 ( .A(n13832), .ZN(n6801) );
  XNOR2_X1 U9481 ( .A(n11793), .B(n11791), .ZN(n11790) );
  OR2_X1 U9482 ( .A1(n7955), .A2(n13430), .ZN(n6604) );
  NAND2_X1 U9483 ( .A1(n8446), .A2(n8445), .ZN(n13671) );
  INV_X1 U9484 ( .A(n13671), .ZN(n7159) );
  OR2_X1 U9485 ( .A1(n13741), .A2(n13709), .ZN(n6605) );
  INV_X1 U9486 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8873) );
  INV_X1 U9487 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6691) );
  INV_X1 U9488 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6672) );
  OR2_X1 U9489 ( .A1(n15392), .A2(n10080), .ZN(n6606) );
  OR2_X1 U9490 ( .A1(n15396), .A2(n10080), .ZN(n6607) );
  NAND2_X1 U9491 ( .A1(n7512), .A2(n7510), .ZN(n6608) );
  NAND2_X1 U9492 ( .A1(n7347), .A2(n7348), .ZN(n6609) );
  AND2_X1 U9493 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_REG3_REG_13__SCAN_IN), 
        .ZN(n6610) );
  OR2_X1 U9494 ( .A1(n6602), .A2(n15666), .ZN(n6611) );
  NAND2_X1 U9495 ( .A1(n9976), .A2(n14416), .ZN(n6612) );
  AND2_X1 U9496 ( .A1(n8854), .A2(n14491), .ZN(n6613) );
  NAND2_X1 U9497 ( .A1(n10460), .A2(n10459), .ZN(n6614) );
  OR2_X1 U9498 ( .A1(n13741), .A2(n13790), .ZN(n6615) );
  INV_X1 U9499 ( .A(n7530), .ZN(n7152) );
  AOI21_X1 U9500 ( .B1(n7532), .B2(n15251), .A(n6515), .ZN(n7530) );
  INV_X1 U9501 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10876) );
  INV_X1 U9502 ( .A(n7762), .ZN(n7761) );
  INV_X1 U9503 ( .A(n12770), .ZN(n7762) );
  NAND2_X1 U9504 ( .A1(n9682), .A2(n9681), .ZN(n15543) );
  INV_X1 U9505 ( .A(n15543), .ZN(n7768) );
  AND2_X1 U9506 ( .A1(n11508), .A2(n11564), .ZN(n11509) );
  INV_X1 U9507 ( .A(n11448), .ZN(n6973) );
  NAND2_X1 U9508 ( .A1(n12547), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6616) );
  AND2_X1 U9509 ( .A1(n11058), .A2(n14647), .ZN(n15610) );
  OAI21_X1 U9510 ( .B1(n10483), .B2(n9612), .A(n10487), .ZN(n11254) );
  NAND2_X1 U9511 ( .A1(n9716), .A2(n9715), .ZN(n12516) );
  INV_X1 U9512 ( .A(n12516), .ZN(n7050) );
  XNOR2_X1 U9513 ( .A(n8542), .B(n8887), .ZN(n8885) );
  AND2_X1 U9514 ( .A1(n15691), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n6617) );
  OR2_X1 U9515 ( .A1(n15670), .A2(n9468), .ZN(n6618) );
  AND2_X1 U9516 ( .A1(n11986), .A2(n15660), .ZN(n14575) );
  INV_X1 U9517 ( .A(n14575), .ZN(n14579) );
  INV_X2 U9518 ( .A(n9401), .ZN(n9473) );
  INV_X1 U9519 ( .A(n9476), .ZN(n9497) );
  AND2_X1 U9520 ( .A1(n11064), .A2(n11048), .ZN(n15587) );
  AND2_X1 U9521 ( .A1(n6744), .A2(n6743), .ZN(n6619) );
  INV_X1 U9522 ( .A(n12147), .ZN(n7051) );
  AND2_X1 U9523 ( .A1(n7328), .A2(n7330), .ZN(n6620) );
  AND2_X1 U9524 ( .A1(n7504), .A2(n7506), .ZN(n6621) );
  AND2_X1 U9525 ( .A1(n7236), .A2(n7235), .ZN(n6622) );
  AND2_X1 U9526 ( .A1(n11583), .A2(n7083), .ZN(n6623) );
  NAND2_X1 U9527 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n6624) );
  AND2_X1 U9528 ( .A1(n15434), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6625) );
  AND2_X1 U9529 ( .A1(n8859), .A2(SI_30_), .ZN(n6626) );
  AND2_X1 U9530 ( .A1(n12043), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6627) );
  INV_X1 U9531 ( .A(n6733), .ZN(n14916) );
  OR2_X1 U9532 ( .A1(n14919), .A2(n6734), .ZN(n6733) );
  NAND2_X1 U9533 ( .A1(n7487), .A2(n7486), .ZN(n6628) );
  NOR2_X1 U9534 ( .A1(n9303), .A2(n7604), .ZN(n7603) );
  AOI21_X1 U9535 ( .B1(n11532), .B2(n11530), .A(n11531), .ZN(n7493) );
  OR2_X1 U9536 ( .A1(n14968), .A2(n14969), .ZN(n6629) );
  INV_X1 U9537 ( .A(n7023), .ZN(n7022) );
  NAND2_X1 U9538 ( .A1(n14955), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7023) );
  INV_X1 U9539 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n14413) );
  OR2_X1 U9540 ( .A1(n9587), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n6630) );
  AND2_X1 U9541 ( .A1(n6866), .A2(n7581), .ZN(n14629) );
  INV_X1 U9542 ( .A(n8000), .ZN(n7321) );
  AND2_X1 U9543 ( .A1(n14875), .A2(n10921), .ZN(n6631) );
  AND2_X1 U9544 ( .A1(n6470), .A2(n7321), .ZN(n6632) );
  NAND2_X1 U9545 ( .A1(n8511), .A2(n8512), .ZN(n13796) );
  AND2_X1 U9546 ( .A1(n7496), .A2(n11198), .ZN(n6633) );
  INV_X1 U9547 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n7338) );
  NAND2_X1 U9548 ( .A1(n7983), .A2(n11041), .ZN(n10734) );
  INV_X1 U9549 ( .A(n11041), .ZN(n7054) );
  INV_X2 U9550 ( .A(n13801), .ZN(n13808) );
  NAND2_X2 U9551 ( .A1(n10817), .A2(P3_U3151), .ZN(n13805) );
  INV_X4 U9552 ( .A(n6978), .ZN(n10817) );
  NAND2_X2 U9553 ( .A1(n6634), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n6714) );
  INV_X1 U9554 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6636) );
  XNOR2_X1 U9555 ( .A(n8567), .B(n10839), .ZN(n8571) );
  NAND2_X2 U9556 ( .A1(n6640), .A2(n8722), .ZN(n8732) );
  NAND2_X1 U9557 ( .A1(n14721), .A2(n14722), .ZN(n6642) );
  NAND2_X1 U9558 ( .A1(n14658), .A2(n14659), .ZN(n10264) );
  NAND2_X1 U9559 ( .A1(n6644), .A2(n11394), .ZN(n11395) );
  NAND2_X1 U9560 ( .A1(n6645), .A2(n6957), .ZN(n7480) );
  NAND2_X1 U9561 ( .A1(n6645), .A2(n7481), .ZN(n7251) );
  XNOR2_X1 U9562 ( .A(n6645), .B(n8624), .ZN(n10827) );
  INV_X1 U9563 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U9564 ( .A1(n13443), .A2(n6567), .ZN(n13466) );
  NAND2_X1 U9565 ( .A1(n13445), .A2(n13444), .ZN(n13443) );
  NAND2_X1 U9566 ( .A1(n7825), .A2(n6654), .ZN(n12959) );
  NAND4_X1 U9567 ( .A1(n7824), .A2(n7821), .A3(n7823), .A4(n7822), .ZN(n6654)
         );
  NAND2_X1 U9568 ( .A1(n6655), .A2(n6595), .ZN(n9414) );
  OAI21_X1 U9569 ( .B1(n6657), .B2(n6656), .A(n7381), .ZN(n6655) );
  AOI21_X1 U9570 ( .B1(n6658), .B2(n9397), .A(n9396), .ZN(n6656) );
  OAI21_X1 U9571 ( .B1(n6658), .B2(n9397), .A(n9522), .ZN(n6657) );
  NAND3_X1 U9572 ( .A1(n9440), .A2(n9439), .A3(n6588), .ZN(n6661) );
  NAND4_X1 U9573 ( .A1(n9363), .A2(n6664), .A3(n6663), .A4(n6662), .ZN(n6986)
         );
  NAND3_X1 U9574 ( .A1(n6668), .A2(n9380), .A3(n6666), .ZN(n9383) );
  NAND3_X1 U9575 ( .A1(n6667), .A2(n9376), .A3(n9371), .ZN(n6666) );
  NAND2_X1 U9576 ( .A1(n6669), .A2(n9376), .ZN(n6668) );
  NAND2_X1 U9577 ( .A1(n7097), .A2(n6585), .ZN(n6670) );
  INV_X1 U9578 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6674) );
  NAND3_X1 U9579 ( .A1(n6678), .A2(n7098), .A3(n6676), .ZN(n9435) );
  NAND3_X1 U9580 ( .A1(n9430), .A2(n7355), .A3(n6502), .ZN(n6678) );
  NAND2_X1 U9581 ( .A1(n9435), .A2(n9436), .ZN(n9434) );
  XNOR2_X2 U9582 ( .A(n8890), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8950) );
  NAND2_X1 U9583 ( .A1(n6684), .A2(n15287), .ZN(n15288) );
  NAND2_X1 U9584 ( .A1(n15381), .A2(n15554), .ZN(n6684) );
  OAI21_X1 U9585 ( .B1(n14107), .B2(n7554), .A(n6687), .ZN(n10455) );
  NAND2_X1 U9586 ( .A1(n7557), .A2(n14102), .ZN(n6688) );
  INV_X1 U9587 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6692) );
  NOR2_X1 U9588 ( .A1(n6707), .A2(n6706), .ZN(n7079) );
  NAND3_X1 U9589 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n6712) );
  INV_X1 U9590 ( .A(n15283), .ZN(n6713) );
  NAND2_X4 U9591 ( .A1(n6715), .A2(n6714), .ZN(n10818) );
  NAND3_X1 U9592 ( .A1(n6715), .A2(n6714), .A3(n8545), .ZN(n9599) );
  NAND2_X2 U9593 ( .A1(n8062), .A2(n7068), .ZN(n6715) );
  NAND2_X1 U9594 ( .A1(n7123), .A2(n8658), .ZN(n6717) );
  NAND2_X1 U9595 ( .A1(n6717), .A2(n8711), .ZN(n7260) );
  XNOR2_X1 U9596 ( .A(n7457), .B(n7456), .ZN(n10904) );
  INV_X1 U9597 ( .A(n6718), .ZN(n15146) );
  NOR2_X2 U9598 ( .A1(n15130), .A2(n15113), .ZN(n15112) );
  NAND2_X1 U9599 ( .A1(n6718), .A2(n15404), .ZN(n15130) );
  NOR2_X1 U9600 ( .A1(n15167), .A2(n15151), .ZN(n6718) );
  NAND2_X1 U9601 ( .A1(n14954), .A2(n6722), .ZN(n6719) );
  INV_X1 U9602 ( .A(n10916), .ZN(n6724) );
  NAND3_X1 U9603 ( .A1(n10919), .A2(n6725), .A3(n6723), .ZN(n15505) );
  NAND2_X1 U9604 ( .A1(n6724), .A2(n15502), .ZN(n6723) );
  NAND3_X1 U9605 ( .A1(n14865), .A2(n15502), .A3(n14866), .ZN(n6725) );
  NAND2_X1 U9606 ( .A1(n11349), .A2(n6583), .ZN(n6744) );
  NAND2_X1 U9607 ( .A1(n11349), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n11350) );
  NOR2_X1 U9608 ( .A1(n6746), .A2(n11849), .ZN(n6745) );
  NAND2_X1 U9609 ( .A1(n11113), .A2(n11114), .ZN(n11112) );
  XNOR2_X1 U9610 ( .A(n7973), .B(n15680), .ZN(n11114) );
  INV_X1 U9611 ( .A(n10734), .ZN(n7331) );
  NAND3_X1 U9612 ( .A1(n7979), .A2(P3_REG2_REG_3__SCAN_IN), .A3(n11203), .ZN(
        n11335) );
  NAND2_X1 U9613 ( .A1(n7979), .A2(n11203), .ZN(n11337) );
  NAND4_X1 U9614 ( .A1(n7094), .A2(n7874), .A3(n7869), .A4(n6751), .ZN(n7819)
         );
  INV_X2 U9615 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7874) );
  NAND3_X1 U9616 ( .A1(n7837), .A2(n6753), .A3(n6752), .ZN(n7818) );
  NAND3_X1 U9617 ( .A1(n13139), .A2(n13637), .A3(n13653), .ZN(n6758) );
  NAND3_X1 U9618 ( .A1(n7833), .A2(n7805), .A3(n7448), .ZN(n6764) );
  NAND2_X1 U9619 ( .A1(n6764), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7906) );
  NAND4_X1 U9620 ( .A1(n6765), .A2(n7166), .A3(n7165), .A4(n7031), .ZN(
        P3_U3296) );
  NAND2_X1 U9621 ( .A1(n6766), .A2(n13077), .ZN(n11737) );
  NAND2_X1 U9622 ( .A1(n6767), .A2(n13011), .ZN(n8477) );
  XNOR2_X1 U9623 ( .A(n6767), .B(n13011), .ZN(n15709) );
  NAND2_X1 U9624 ( .A1(n11739), .A2(n13082), .ZN(n6767) );
  NAND2_X1 U9625 ( .A1(n12981), .A2(n6436), .ZN(n6769) );
  XNOR2_X1 U9626 ( .A(n6770), .B(n11284), .ZN(n13187) );
  AND3_X2 U9627 ( .A1(n6771), .A2(n7811), .A3(n7810), .ZN(n7821) );
  AND3_X2 U9628 ( .A1(n6772), .A2(n7813), .A3(n7975), .ZN(n7824) );
  NOR2_X2 U9629 ( .A1(n7817), .A2(n6773), .ZN(n7823) );
  NAND4_X1 U9630 ( .A1(n7854), .A2(n7816), .A3(n7448), .A4(n7815), .ZN(n6773)
         );
  NAND3_X1 U9631 ( .A1(n7801), .A2(n7866), .A3(n7879), .ZN(n7817) );
  NOR2_X2 U9632 ( .A1(n7819), .A2(n7818), .ZN(n7822) );
  NAND3_X1 U9633 ( .A1(n6775), .A2(n6451), .A3(n6581), .ZN(n6774) );
  NAND2_X1 U9634 ( .A1(n13632), .A2(n6589), .ZN(n6775) );
  NAND3_X1 U9635 ( .A1(n7654), .A2(n6447), .A3(n6497), .ZN(n6776) );
  OAI21_X1 U9636 ( .B1(n12613), .B2(n8483), .A(n13127), .ZN(n12798) );
  NOR2_X2 U9637 ( .A1(n14208), .A2(n14196), .ZN(n14195) );
  NAND2_X2 U9638 ( .A1(n6793), .A2(n6792), .ZN(n14298) );
  NAND3_X1 U9639 ( .A1(n7628), .A2(n12104), .A3(n6796), .ZN(n7626) );
  INV_X2 U9640 ( .A(n8866), .ZN(n8769) );
  NAND2_X2 U9641 ( .A1(n11042), .A2(n6978), .ZN(n8866) );
  NAND3_X1 U9642 ( .A1(n6797), .A2(n14178), .A3(n7609), .ZN(n10461) );
  NAND2_X1 U9643 ( .A1(n7418), .A2(n6498), .ZN(n9272) );
  NAND3_X1 U9644 ( .A1(n7785), .A2(n9064), .A3(n7401), .ZN(n6809) );
  NAND2_X1 U9645 ( .A1(n12506), .A2(n6582), .ZN(n7135) );
  NAND2_X1 U9646 ( .A1(n7132), .A2(n7135), .ZN(n7136) );
  NAND2_X1 U9647 ( .A1(n12559), .A2(n6816), .ZN(n6813) );
  NAND3_X1 U9648 ( .A1(n6814), .A2(n6813), .A3(n7150), .ZN(n15214) );
  NAND3_X1 U9649 ( .A1(n12192), .A2(n6571), .A3(n9726), .ZN(n7534) );
  INV_X2 U9650 ( .A(n9590), .ZN(n13214) );
  NAND2_X1 U9651 ( .A1(n9587), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6827) );
  NAND3_X1 U9652 ( .A1(n11760), .A2(n11876), .A3(n10652), .ZN(n6828) );
  OAI21_X1 U9653 ( .B1(n10501), .B2(n6839), .A(n6460), .ZN(n6840) );
  INV_X2 U9654 ( .A(n9631), .ZN(n9848) );
  NAND2_X2 U9655 ( .A1(n9632), .A2(n10817), .ZN(n9631) );
  XNOR2_X2 U9656 ( .A(n9605), .B(n9604), .ZN(n15436) );
  XNOR2_X2 U9657 ( .A(n9602), .B(n9601), .ZN(n9986) );
  NAND2_X1 U9658 ( .A1(n6841), .A2(n7389), .ZN(n10589) );
  NAND3_X1 U9659 ( .A1(n6843), .A2(n7391), .A3(n6842), .ZN(n6841) );
  OAI211_X1 U9660 ( .C1(n10580), .C2(n7379), .A(n7376), .B(n7377), .ZN(n6842)
         );
  NAND2_X1 U9661 ( .A1(n6844), .A2(n10583), .ZN(n6843) );
  NAND2_X1 U9662 ( .A1(n7374), .A2(n7375), .ZN(n6844) );
  NAND2_X1 U9663 ( .A1(n11316), .A2(n6845), .ZN(n15520) );
  NAND2_X1 U9664 ( .A1(n11315), .A2(n11314), .ZN(n6845) );
  OAI21_X1 U9665 ( .B1(n12421), .B2(n6850), .A(n6474), .ZN(n12555) );
  NAND2_X1 U9666 ( .A1(n6848), .A2(n6846), .ZN(n7717) );
  NAND2_X1 U9667 ( .A1(n12421), .A2(n6474), .ZN(n6848) );
  AOI21_X1 U9668 ( .B1(n6858), .B2(n6856), .A(n6491), .ZN(n6851) );
  NAND2_X1 U9669 ( .A1(n6857), .A2(n6858), .ZN(n6852) );
  NAND2_X1 U9670 ( .A1(n6855), .A2(n6858), .ZN(n15144) );
  NAND2_X1 U9671 ( .A1(n15178), .A2(n7277), .ZN(n6855) );
  INV_X1 U9672 ( .A(n7277), .ZN(n6856) );
  INV_X1 U9673 ( .A(n15178), .ZN(n6857) );
  AOI21_X2 U9674 ( .B1(n7277), .B2(n6441), .A(n15139), .ZN(n6858) );
  NAND2_X1 U9675 ( .A1(n7581), .A2(n7579), .ZN(n6865) );
  NAND2_X1 U9676 ( .A1(n11932), .A2(n6870), .ZN(n6868) );
  NAND3_X1 U9677 ( .A1(n6443), .A2(n10416), .A3(n7788), .ZN(n14246) );
  NAND3_X1 U9678 ( .A1(n6443), .A2(n10416), .A3(n6876), .ZN(n6875) );
  OAI21_X1 U9679 ( .B1(n10422), .B2(n7567), .A(n7564), .ZN(n10426) );
  XNOR2_X1 U9680 ( .A(n6881), .B(n14102), .ZN(n14094) );
  NAND2_X1 U9681 ( .A1(n6886), .A2(n6883), .ZN(n10995) );
  NAND2_X1 U9682 ( .A1(n10994), .A2(n10993), .ZN(n11303) );
  NAND2_X1 U9683 ( .A1(n10770), .A2(n14856), .ZN(n6896) );
  NAND2_X1 U9684 ( .A1(n11707), .A2(n6899), .ZN(n6898) );
  NAND2_X1 U9685 ( .A1(n10349), .A2(n6908), .ZN(n6907) );
  AND2_X1 U9686 ( .A1(n9364), .A2(n11710), .ZN(n7797) );
  XNOR2_X1 U9687 ( .A(n13978), .B(n13827), .ZN(n11710) );
  NAND2_X1 U9688 ( .A1(n7794), .A2(n11297), .ZN(n11296) );
  NAND2_X1 U9689 ( .A1(n11144), .A2(n10092), .ZN(n11297) );
  INV_X1 U9690 ( .A(n11147), .ZN(n6923) );
  NAND2_X1 U9691 ( .A1(n10100), .A2(n10099), .ZN(n10101) );
  INV_X1 U9692 ( .A(n10100), .ZN(n6925) );
  OAI21_X2 U9693 ( .B1(n11816), .B2(n6935), .A(n6933), .ZN(n12214) );
  INV_X1 U9694 ( .A(n12214), .ZN(n10156) );
  NAND2_X1 U9695 ( .A1(n14721), .A2(n6941), .ZN(n6940) );
  NAND2_X1 U9696 ( .A1(n8732), .A2(n7792), .ZN(n6947) );
  OAI21_X1 U9697 ( .B1(n8732), .B2(n6950), .A(n6948), .ZN(n8756) );
  NAND2_X1 U9698 ( .A1(n8732), .A2(n6948), .ZN(n6946) );
  OAI22_X2 U9699 ( .A1(n7088), .A2(n6540), .B1(n6952), .B2(n6951), .ZN(n9455)
         );
  INV_X1 U9700 ( .A(n9446), .ZN(n7074) );
  NAND2_X2 U9701 ( .A1(n12893), .A2(n13194), .ZN(n8153) );
  XNOR2_X2 U9702 ( .A(n6958), .B(n12945), .ZN(n13194) );
  AOI21_X2 U9703 ( .B1(n12784), .B2(n12783), .A(n12782), .ZN(n12897) );
  OAI21_X2 U9704 ( .B1(n12342), .B2(n6444), .A(n6550), .ZN(n12531) );
  INV_X1 U9705 ( .A(n13732), .ZN(n6959) );
  NAND3_X1 U9706 ( .A1(n6962), .A2(n6439), .A3(n6959), .ZN(n13064) );
  NAND2_X2 U9707 ( .A1(n6439), .A2(n6962), .ZN(n11181) );
  NAND3_X1 U9708 ( .A1(n6439), .A2(n6962), .A3(n13732), .ZN(n11442) );
  NAND3_X1 U9709 ( .A1(n11442), .A2(n11289), .A3(n6430), .ZN(n6961) );
  AND2_X1 U9710 ( .A1(n7822), .A2(n7823), .ZN(n6965) );
  NAND3_X1 U9711 ( .A1(n7822), .A2(n7823), .A3(n7914), .ZN(n6967) );
  NAND3_X1 U9712 ( .A1(n11553), .A2(n11777), .A3(n11552), .ZN(n6969) );
  XNOR2_X1 U9713 ( .A(n13307), .B(n13308), .ZN(n13309) );
  OAI21_X1 U9714 ( .B1(n6971), .B2(n13351), .A(n13315), .ZN(P3_U3169) );
  XNOR2_X1 U9715 ( .A(n6972), .B(n13311), .ZN(n6971) );
  OAI21_X2 U9716 ( .B1(n13226), .B2(n7433), .A(n7431), .ZN(n13291) );
  NAND2_X1 U9717 ( .A1(n13567), .A2(n13150), .ZN(n13558) );
  INV_X2 U9718 ( .A(n13721), .ZN(n6974) );
  NAND2_X2 U9719 ( .A1(n7966), .A2(n7929), .ZN(n8471) );
  NAND2_X1 U9720 ( .A1(n13007), .A2(n11437), .ZN(n11439) );
  NAND2_X1 U9721 ( .A1(n13716), .A2(n13063), .ZN(n11288) );
  NAND3_X1 U9722 ( .A1(n11379), .A2(n13720), .A3(n7041), .ZN(n11378) );
  NAND2_X1 U9723 ( .A1(n11777), .A2(n11586), .ZN(n11587) );
  INV_X4 U9724 ( .A(n8110), .ZN(n12983) );
  OAI211_X1 U9725 ( .C1(n10329), .C2(n10328), .A(n6975), .B(n10327), .ZN(
        P1_U3220) );
  NAND2_X1 U9726 ( .A1(n10329), .A2(n10326), .ZN(n6975) );
  INV_X1 U9727 ( .A(n11537), .ZN(n10113) );
  NAND2_X1 U9728 ( .A1(n13301), .A2(n13300), .ZN(n13299) );
  NAND3_X1 U9729 ( .A1(n9448), .A2(n6593), .A3(n9449), .ZN(n7088) );
  OAI21_X1 U9730 ( .B1(n8895), .B2(n7582), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8542) );
  NAND2_X1 U9731 ( .A1(n7378), .A2(n10579), .ZN(n7377) );
  INV_X1 U9732 ( .A(n8633), .ZN(n8634) );
  NOR2_X1 U9733 ( .A1(n10606), .A2(n10605), .ZN(n10608) );
  NAND2_X1 U9734 ( .A1(n8656), .A2(n8655), .ZN(n7123) );
  NAND2_X1 U9735 ( .A1(n7015), .A2(n7124), .ZN(n8656) );
  NAND2_X1 U9736 ( .A1(n9599), .A2(n8552), .ZN(n8560) );
  NAND2_X1 U9737 ( .A1(n10426), .A2(n10425), .ZN(n10428) );
  NAND2_X1 U9738 ( .A1(n10539), .A2(n10556), .ZN(n7019) );
  XNOR2_X1 U9739 ( .A(n10457), .B(n10456), .ZN(n7545) );
  NAND2_X1 U9740 ( .A1(n6976), .A2(n15670), .ZN(n7259) );
  NOR2_X1 U9741 ( .A1(n15598), .A2(n15599), .ZN(n15596) );
  MUX2_X2 U9742 ( .A(n15390), .B(n15389), .S(n15550), .Z(n15391) );
  NOR2_X2 U9743 ( .A1(n15110), .A2(n15111), .ZN(n15109) );
  NAND2_X1 U9744 ( .A1(n8811), .A2(n8810), .ZN(n8817) );
  NAND2_X1 U9745 ( .A1(n6980), .A2(n6521), .ZN(n9501) );
  XNOR2_X1 U9746 ( .A(n8864), .B(n8863), .ZN(n10639) );
  INV_X1 U9747 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10808) );
  INV_X1 U9748 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7068) );
  INV_X1 U9749 ( .A(n9500), .ZN(n6980) );
  OAI21_X1 U9750 ( .B1(n7464), .B2(n7460), .A(n7458), .ZN(n8864) );
  NAND2_X1 U9751 ( .A1(n6996), .A2(n8610), .ZN(n8616) );
  INV_X1 U9752 ( .A(n8847), .ZN(n7464) );
  NOR2_X1 U9753 ( .A1(n9487), .A2(n6519), .ZN(n9488) );
  NAND2_X1 U9754 ( .A1(n12087), .A2(n8478), .ZN(n6999) );
  NAND2_X1 U9755 ( .A1(n6999), .A2(n6574), .ZN(n6998) );
  NAND3_X1 U9756 ( .A1(n7009), .A2(n6983), .A3(n10491), .ZN(n7354) );
  OAI21_X1 U9757 ( .B1(n7368), .B2(n7367), .A(n7369), .ZN(n10501) );
  NOR2_X1 U9758 ( .A1(n10494), .A2(n10492), .ZN(n7353) );
  NAND2_X1 U9759 ( .A1(n10481), .A2(n10480), .ZN(n6983) );
  NAND2_X1 U9760 ( .A1(n12725), .A2(n10345), .ZN(n14319) );
  INV_X1 U9761 ( .A(n9513), .ZN(n11484) );
  NAND2_X1 U9762 ( .A1(n10594), .A2(n10593), .ZN(n10596) );
  NAND2_X1 U9763 ( .A1(n7011), .A2(n7010), .ZN(n10511) );
  NAND2_X1 U9764 ( .A1(n7255), .A2(n7253), .ZN(n10447) );
  NAND2_X1 U9765 ( .A1(n10755), .A2(n10754), .ZN(n10753) );
  NAND2_X1 U9766 ( .A1(n8839), .A2(n7454), .ZN(n8843) );
  NAND2_X1 U9767 ( .A1(n15305), .A2(n6606), .ZN(P1_U3553) );
  NAND2_X1 U9768 ( .A1(n6986), .A2(n7797), .ZN(n7097) );
  AOI21_X1 U9769 ( .B1(n9531), .B2(n9489), .A(n9488), .ZN(n9496) );
  INV_X1 U9770 ( .A(n11255), .ZN(n11250) );
  NAND2_X1 U9771 ( .A1(n7102), .A2(n7101), .ZN(n7100) );
  NAND2_X1 U9772 ( .A1(n7275), .A2(n10011), .ZN(n15211) );
  NOR2_X1 U9773 ( .A1(n6602), .A2(n6992), .ZN(n6991) );
  NOR3_X2 U9774 ( .A1(n15109), .A2(n10023), .A3(n15092), .ZN(n15087) );
  NAND2_X1 U9775 ( .A1(n7648), .A2(n7647), .ZN(n13603) );
  NAND2_X2 U9776 ( .A1(n13064), .A2(n13063), .ZN(n11375) );
  INV_X1 U9777 ( .A(n8316), .ZN(n7047) );
  NAND2_X1 U9778 ( .A1(n12614), .A2(n8304), .ZN(n12796) );
  NAND2_X1 U9779 ( .A1(n8166), .A2(n8165), .ZN(n11740) );
  NAND2_X1 U9780 ( .A1(n7210), .A2(n7208), .ZN(n12393) );
  NAND2_X1 U9781 ( .A1(n10156), .A2(n10155), .ZN(n12212) );
  NAND2_X1 U9782 ( .A1(n7246), .A2(n7245), .ZN(n7242) );
  NAND2_X1 U9783 ( .A1(n14740), .A2(n7691), .ZN(n14649) );
  NAND2_X1 U9784 ( .A1(n10051), .A2(n10050), .ZN(n6989) );
  OR2_X2 U9785 ( .A1(n12109), .A2(n6989), .ZN(n10084) );
  OAI21_X1 U9786 ( .B1(n14354), .B2(n15664), .A(n7544), .ZN(P2_U3496) );
  NAND2_X1 U9787 ( .A1(n13299), .A2(n12905), .ZN(n13337) );
  NAND2_X1 U9788 ( .A1(n11378), .A2(n7084), .ZN(n11290) );
  AOI21_X2 U9789 ( .B1(n12897), .B2(n12896), .A(n12895), .ZN(n13226) );
  NAND2_X1 U9790 ( .A1(n11288), .A2(n12935), .ZN(n7041) );
  NAND2_X1 U9791 ( .A1(n7928), .A2(n11107), .ZN(n11332) );
  XNOR2_X2 U9792 ( .A(n7961), .B(n6599), .ZN(n13508) );
  NAND3_X1 U9793 ( .A1(n7005), .A2(n7089), .A3(n8004), .ZN(P3_U3201) );
  NAND2_X1 U9794 ( .A1(n7110), .A2(n7107), .ZN(n12318) );
  OAI21_X1 U9795 ( .B1(n12499), .B2(n6446), .A(n12828), .ZN(n7299) );
  NAND3_X1 U9796 ( .A1(n8607), .A2(n8606), .A3(n6997), .ZN(n6996) );
  INV_X1 U9797 ( .A(n9400), .ZN(n7382) );
  NAND2_X1 U9798 ( .A1(n7109), .A2(n7108), .ZN(n7107) );
  NAND2_X1 U9799 ( .A1(n7296), .A2(n7295), .ZN(n7120) );
  OAI21_X1 U9800 ( .B1(n12318), .B2(n12317), .A(n12316), .ZN(n12320) );
  NOR2_X1 U9801 ( .A1(n7668), .A2(n13041), .ZN(n7667) );
  NAND2_X1 U9802 ( .A1(n13670), .A2(n6605), .ZN(P3_U3487) );
  NAND2_X1 U9803 ( .A1(n13740), .A2(n6615), .ZN(P3_U3455) );
  NAND2_X1 U9804 ( .A1(n7673), .A2(n13167), .ZN(n7104) );
  NAND2_X1 U9805 ( .A1(n9861), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U9806 ( .A1(n15035), .A2(n15034), .ZN(n7072) );
  OAI21_X1 U9807 ( .B1(n9455), .B2(n9454), .A(n9453), .ZN(n9457) );
  NAND4_X2 U9808 ( .A1(n9025), .A2(n9024), .A3(n9023), .A4(n9022), .ZN(n13975)
         );
  NAND2_X1 U9809 ( .A1(n11201), .A2(n7865), .ZN(n7871) );
  INV_X1 U9810 ( .A(n7046), .ZN(n7045) );
  NAND2_X1 U9811 ( .A1(n7483), .A2(n7045), .ZN(n13492) );
  NAND2_X1 U9812 ( .A1(n7241), .A2(n6596), .ZN(n14682) );
  NAND2_X1 U9813 ( .A1(n7692), .A2(n7696), .ZN(n7695) );
  NOR2_X1 U9814 ( .A1(n14943), .A2(n14944), .ZN(n14954) );
  NOR2_X1 U9815 ( .A1(n10708), .A2(n7004), .ZN(n7994) );
  NAND2_X1 U9816 ( .A1(n14877), .A2(n14876), .ZN(n14875) );
  INV_X1 U9817 ( .A(n13455), .ZN(n7343) );
  NAND4_X1 U9818 ( .A1(n10489), .A2(n10490), .A3(n11321), .A4(n11255), .ZN(
        n7009) );
  INV_X1 U9819 ( .A(n10510), .ZN(n7011) );
  OAI21_X1 U9820 ( .B1(n10496), .B2(n10497), .A(n6586), .ZN(n7367) );
  NAND2_X1 U9821 ( .A1(n11759), .A2(n9998), .ZN(n7012) );
  NAND2_X1 U9822 ( .A1(n15309), .A2(n6607), .ZN(P1_U3552) );
  NAND2_X1 U9823 ( .A1(n7731), .A2(n7732), .ZN(n12421) );
  OAI21_X2 U9824 ( .B1(n15087), .B2(n15067), .A(n15066), .ZN(n15069) );
  NAND2_X2 U9825 ( .A1(n8087), .A2(n8086), .ZN(n8138) );
  NAND2_X1 U9826 ( .A1(n8711), .A2(n8666), .ZN(n7262) );
  NAND2_X1 U9827 ( .A1(n10540), .A2(n10550), .ZN(n7018) );
  INV_X4 U9828 ( .A(n10786), .ZN(n8812) );
  XNOR2_X1 U9829 ( .A(n9633), .B(n9634), .ZN(n14863) );
  NOR2_X1 U9830 ( .A1(n10958), .A2(n10957), .ZN(n10960) );
  NAND2_X1 U9831 ( .A1(n7464), .A2(n8848), .ZN(n7463) );
  NOR2_X1 U9832 ( .A1(n7611), .A2(n14081), .ZN(n7610) );
  INV_X1 U9833 ( .A(n7024), .ZN(n14350) );
  AOI21_X1 U9834 ( .B1(n14583), .B2(n15670), .A(n7025), .ZN(n7024) );
  INV_X1 U9835 ( .A(n7026), .ZN(n14584) );
  AOI21_X1 U9836 ( .B1(n14583), .B2(n15666), .A(n7027), .ZN(n7026) );
  INV_X1 U9837 ( .A(n8582), .ZN(n8601) );
  NAND2_X1 U9838 ( .A1(n8650), .A2(n10806), .ZN(n7028) );
  AND2_X1 U9839 ( .A1(n7030), .A2(n14079), .ZN(n14348) );
  NAND2_X1 U9840 ( .A1(n7608), .A2(n7607), .ZN(n14079) );
  AOI21_X1 U9841 ( .B1(n14080), .B2(n14081), .A(n14320), .ZN(n7030) );
  NAND2_X1 U9842 ( .A1(n13187), .A2(n7167), .ZN(n7031) );
  OAI21_X1 U9843 ( .B1(n9385), .B2(n9384), .A(n9388), .ZN(n9390) );
  NAND2_X2 U9844 ( .A1(n10015), .A2(n10014), .ZN(n15178) );
  INV_X1 U9845 ( .A(n7125), .ZN(n7124) );
  NAND2_X1 U9846 ( .A1(n13414), .A2(n13413), .ZN(n7347) );
  NAND2_X1 U9847 ( .A1(n7259), .A2(n6618), .ZN(P2_U3528) );
  NAND2_X1 U9848 ( .A1(n7373), .A2(n7372), .ZN(n10518) );
  NAND3_X1 U9849 ( .A1(n7040), .A2(n7044), .A3(n8473), .ZN(n13530) );
  NAND2_X1 U9850 ( .A1(n13534), .A2(n13718), .ZN(n7040) );
  NAND2_X1 U9851 ( .A1(n7136), .A2(n7407), .ZN(n13926) );
  NAND2_X1 U9852 ( .A1(n13898), .A2(n13897), .ZN(n13896) );
  INV_X1 U9853 ( .A(n7440), .ZN(n7439) );
  OAI21_X1 U9854 ( .B1(n8838), .B2(n14412), .A(n8837), .ZN(n7454) );
  NAND3_X1 U9855 ( .A1(n9475), .A2(n9531), .A3(n7042), .ZN(n9490) );
  NAND2_X1 U9856 ( .A1(n12616), .A2(n12615), .ZN(n12614) );
  AOI21_X2 U9857 ( .B1(n13421), .B2(n10714), .A(n10715), .ZN(n10713) );
  OAI21_X1 U9858 ( .B1(n13494), .B2(P3_REG1_REG_17__SCAN_IN), .A(n13493), .ZN(
        n7046) );
  NAND2_X1 U9859 ( .A1(n12276), .A2(n7665), .ZN(n7210) );
  NOR2_X1 U9860 ( .A1(n7490), .A2(n7489), .ZN(n7095) );
  NAND2_X2 U9861 ( .A1(n7049), .A2(n7048), .ZN(n11317) );
  INV_X2 U9862 ( .A(n11259), .ZN(n7048) );
  NOR2_X2 U9863 ( .A1(n15054), .A2(n15053), .ZN(n15041) );
  NAND2_X1 U9864 ( .A1(n7475), .A2(n8779), .ZN(n8792) );
  NAND2_X1 U9865 ( .A1(n7074), .A2(n7073), .ZN(n9449) );
  NAND2_X1 U9866 ( .A1(n7981), .A2(n11202), .ZN(n11206) );
  NAND2_X1 U9867 ( .A1(n7994), .A2(n7993), .ZN(n7345) );
  NAND3_X1 U9868 ( .A1(n6442), .A2(n8000), .A3(n7318), .ZN(n7317) );
  NAND3_X1 U9869 ( .A1(n7496), .A2(P3_REG1_REG_3__SCAN_IN), .A3(n11198), .ZN(
        n11328) );
  NAND2_X1 U9870 ( .A1(n11104), .A2(n7860), .ZN(n7498) );
  NAND2_X1 U9871 ( .A1(n11818), .A2(n11817), .ZN(n11816) );
  NAND2_X1 U9872 ( .A1(n7503), .A2(n7502), .ZN(n7877) );
  NOR2_X2 U9873 ( .A1(n13508), .A2(n13507), .ZN(n13511) );
  OR2_X1 U9874 ( .A1(n11585), .A2(n11782), .ZN(n11586) );
  INV_X1 U9875 ( .A(n7818), .ZN(n7804) );
  AND2_X1 U9876 ( .A1(n7424), .A2(n11582), .ZN(n7083) );
  NAND2_X1 U9877 ( .A1(n7064), .A2(n13116), .ZN(n13120) );
  NAND3_X1 U9878 ( .A1(n13115), .A2(n13113), .A3(n13114), .ZN(n7064) );
  INV_X1 U9879 ( .A(n10492), .ZN(n7352) );
  NAND2_X1 U9880 ( .A1(n13166), .A2(n7224), .ZN(n13173) );
  AOI21_X1 U9881 ( .B1(n10561), .B2(n7086), .A(n7149), .ZN(n10578) );
  AOI21_X2 U9882 ( .B1(n9503), .B2(n9502), .A(n9501), .ZN(n9535) );
  NAND3_X1 U9883 ( .A1(n10039), .A2(n10038), .A3(n7728), .ZN(n10076) );
  OAI21_X2 U9884 ( .B1(n8650), .B2(P2_DATAO_REG_4__SCAN_IN), .A(n7069), .ZN(
        n8604) );
  NAND2_X1 U9885 ( .A1(n8650), .A2(n10808), .ZN(n7069) );
  NAND2_X1 U9886 ( .A1(n7470), .A2(n7468), .ZN(n8811) );
  NAND2_X1 U9887 ( .A1(n15462), .A2(n15463), .ZN(n7115) );
  NAND2_X1 U9888 ( .A1(n10773), .A2(n10772), .ZN(n7106) );
  NAND2_X1 U9889 ( .A1(n13481), .A2(n13480), .ZN(n13479) );
  NAND2_X1 U9890 ( .A1(n9475), .A2(n9531), .ZN(n9487) );
  NAND2_X1 U9891 ( .A1(n9481), .A2(n9482), .ZN(n9475) );
  NAND2_X1 U9892 ( .A1(n8847), .A2(n8846), .ZN(n8849) );
  NAND2_X1 U9893 ( .A1(n14634), .A2(n8834), .ZN(n8852) );
  OAI21_X1 U9894 ( .B1(n9426), .B2(n7359), .A(n7075), .ZN(n9430) );
  INV_X4 U9895 ( .A(n9476), .ZN(n9478) );
  AND2_X2 U9896 ( .A1(n7077), .A2(n9586), .ZN(n9600) );
  OR2_X1 U9897 ( .A1(n9614), .A2(n11501), .ZN(n9606) );
  NAND2_X1 U9898 ( .A1(n8475), .A2(n13073), .ZN(n11694) );
  NAND2_X1 U9899 ( .A1(n7274), .A2(n10029), .ZN(n15031) );
  NAND2_X1 U9900 ( .A1(n7717), .A2(n7276), .ZN(n7275) );
  NAND2_X1 U9901 ( .A1(n11250), .A2(n11251), .ZN(n7702) );
  NOR2_X1 U9902 ( .A1(n13530), .A2(n7800), .ZN(n13742) );
  NAND2_X1 U9903 ( .A1(n7457), .A2(n7456), .ZN(n7122) );
  NOR2_X1 U9904 ( .A1(n7087), .A2(n10552), .ZN(n7086) );
  NAND3_X1 U9905 ( .A1(n8539), .A2(n8538), .A3(n8742), .ZN(n8895) );
  AOI21_X1 U9906 ( .B1(n9383), .B2(n9382), .A(n9381), .ZN(n9384) );
  NAND2_X1 U9907 ( .A1(n8765), .A2(n8764), .ZN(n8869) );
  XNOR2_X1 U9908 ( .A(n8767), .B(n8766), .ZN(n8934) );
  NAND3_X1 U9909 ( .A1(n10512), .A2(n10511), .A3(n6592), .ZN(n7373) );
  NAND2_X1 U9910 ( .A1(n7426), .A2(n7425), .ZN(n13318) );
  NAND2_X1 U9911 ( .A1(n14981), .A2(n14983), .ZN(n7091) );
  OR2_X1 U9912 ( .A1(n9370), .A2(n9369), .ZN(n7096) );
  OAI21_X1 U9913 ( .B1(n7479), .B2(n7252), .A(n8649), .ZN(n7125) );
  NAND2_X1 U9914 ( .A1(n10764), .A2(n10763), .ZN(n10773) );
  NAND2_X1 U9915 ( .A1(n7106), .A2(n10768), .ZN(n10769) );
  NAND2_X1 U9916 ( .A1(n7106), .A2(n6575), .ZN(n10770) );
  INV_X1 U9917 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7105) );
  NAND2_X1 U9918 ( .A1(n11790), .A2(n11789), .ZN(n7114) );
  NAND2_X1 U9919 ( .A1(n11794), .A2(n7113), .ZN(n7109) );
  AND2_X2 U9920 ( .A1(n7116), .A2(n7115), .ZN(n15471) );
  NAND2_X1 U9921 ( .A1(n7120), .A2(n7121), .ZN(n10799) );
  NAND3_X1 U9922 ( .A1(n7120), .A2(n7121), .A3(n15496), .ZN(n7119) );
  NAND2_X1 U9923 ( .A1(n7122), .A2(n8708), .ZN(n8703) );
  NAND2_X1 U9924 ( .A1(n7122), .A2(n8684), .ZN(n8677) );
  NAND2_X1 U9925 ( .A1(n7131), .A2(n9300), .ZN(P2_U3186) );
  NAND3_X1 U9926 ( .A1(n13854), .A2(n9273), .A3(n13915), .ZN(n7131) );
  NAND2_X2 U9927 ( .A1(n9590), .A2(n15428), .ZN(n9614) );
  NAND2_X1 U9928 ( .A1(n11760), .A2(n10652), .ZN(n7142) );
  NAND2_X1 U9929 ( .A1(n7144), .A2(n7143), .ZN(n9901) );
  AOI21_X1 U9930 ( .B1(n6572), .B2(n15193), .A(n7145), .ZN(n7144) );
  NAND3_X1 U9931 ( .A1(n13185), .A2(n7171), .A3(n15674), .ZN(n7165) );
  NAND2_X1 U9932 ( .A1(n8266), .A2(n7176), .ZN(n7175) );
  NAND2_X1 U9933 ( .A1(n8016), .A2(n7184), .ZN(n7183) );
  NAND2_X1 U9934 ( .A1(n8053), .A2(n7190), .ZN(n7187) );
  NAND2_X1 U9935 ( .A1(n7187), .A2(n7188), .ZN(n8056) );
  NAND2_X1 U9936 ( .A1(n8053), .A2(n7193), .ZN(n7189) );
  NAND2_X1 U9937 ( .A1(n8053), .A2(n8052), .ZN(n8393) );
  NAND2_X1 U9938 ( .A1(n8331), .A2(n6603), .ZN(n7197) );
  NAND2_X1 U9939 ( .A1(n8331), .A2(n8330), .ZN(n8329) );
  INV_X1 U9940 ( .A(n13557), .ZN(n7213) );
  OAI21_X1 U9941 ( .B1(n7672), .B2(n7222), .A(n7219), .ZN(n9325) );
  NAND2_X1 U9942 ( .A1(n8066), .A2(n6579), .ZN(n8241) );
  NAND2_X1 U9943 ( .A1(n8074), .A2(n8073), .ZN(n8396) );
  NAND3_X1 U9944 ( .A1(n8064), .A2(n11732), .A3(n8063), .ZN(n8180) );
  NAND2_X1 U9945 ( .A1(n10096), .A2(n10292), .ZN(n10094) );
  NAND2_X1 U9946 ( .A1(n6459), .A2(n12968), .ZN(n11539) );
  NAND2_X2 U9947 ( .A1(n12969), .A2(n12970), .ZN(n12968) );
  NAND2_X1 U9948 ( .A1(n14649), .A2(n10207), .ZN(n10212) );
  NAND3_X1 U9949 ( .A1(n14782), .A2(n6597), .A3(n7242), .ZN(n7241) );
  NAND2_X1 U9950 ( .A1(n14649), .A2(n7243), .ZN(n7246) );
  INV_X1 U9951 ( .A(n7246), .ZN(n14784) );
  AND2_X2 U9952 ( .A1(n9579), .A2(n9791), .ZN(n9586) );
  NAND2_X1 U9953 ( .A1(n9976), .A2(n6501), .ZN(n10044) );
  NAND2_X1 U9954 ( .A1(n9976), .A2(n7247), .ZN(n7249) );
  NAND2_X1 U9955 ( .A1(n7251), .A2(n7479), .ZN(n8646) );
  INV_X1 U9956 ( .A(n8645), .ZN(n7252) );
  INV_X1 U9957 ( .A(n7743), .ZN(n7742) );
  INV_X1 U9958 ( .A(n7269), .ZN(n7741) );
  NAND2_X1 U9959 ( .A1(n15059), .A2(n15058), .ZN(n7274) );
  NAND2_X1 U9960 ( .A1(n7457), .A2(n7285), .ZN(n7282) );
  NAND2_X1 U9961 ( .A1(n7282), .A2(n7283), .ZN(n8678) );
  NAND2_X2 U9962 ( .A1(n7288), .A2(n9772), .ZN(n12720) );
  NOR2_X1 U9963 ( .A1(n15448), .A2(n15449), .ZN(n15452) );
  NAND2_X1 U9964 ( .A1(n15449), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n7292) );
  INV_X1 U9965 ( .A(n15449), .ZN(n7294) );
  INV_X1 U9966 ( .A(n10771), .ZN(n7296) );
  NAND2_X1 U9967 ( .A1(n12495), .A2(n7300), .ZN(n7297) );
  NAND2_X1 U9968 ( .A1(n7298), .A2(n7297), .ZN(n12838) );
  NAND2_X1 U9969 ( .A1(n7310), .A2(n7311), .ZN(n11359) );
  MUX2_X1 U9970 ( .A(n7922), .B(n11410), .S(n11365), .Z(n7923) );
  MUX2_X1 U9971 ( .A(n15725), .B(n7980), .S(n11365), .Z(n7934) );
  OAI211_X1 U9972 ( .C1(n6442), .C2(n8000), .A(n7317), .B(n7316), .ZN(n8003)
         );
  NAND2_X1 U9973 ( .A1(n7343), .A2(n7342), .ZN(n7339) );
  NAND2_X1 U9974 ( .A1(n6556), .A2(n12659), .ZN(n7349) );
  NAND4_X1 U9975 ( .A1(n7351), .A2(n7350), .A3(n8530), .A4(n8529), .ZN(n8669)
         );
  AOI21_X1 U9976 ( .B1(n9426), .B2(n7358), .A(n7356), .ZN(n7355) );
  NAND2_X1 U9977 ( .A1(n9390), .A2(n7363), .ZN(n7360) );
  NAND2_X1 U9978 ( .A1(n10580), .A2(n7377), .ZN(n7374) );
  AOI21_X1 U9979 ( .B1(n7379), .B2(n7377), .A(n7376), .ZN(n7375) );
  AOI21_X1 U9980 ( .B1(n7383), .B2(n9403), .A(n7382), .ZN(n7381) );
  NAND4_X1 U9981 ( .A1(n8742), .A2(n8539), .A3(n8538), .A4(n6496), .ZN(n8901)
         );
  NAND2_X1 U9982 ( .A1(n7395), .A2(n11574), .ZN(n7394) );
  NAND3_X1 U9983 ( .A1(n7394), .A2(n7393), .A3(n12003), .ZN(n12002) );
  INV_X1 U9984 ( .A(n7785), .ZN(n7403) );
  XNOR2_X1 U9985 ( .A(n7406), .B(n11979), .ZN(n8982) );
  XNOR2_X1 U9986 ( .A(n15657), .B(n7406), .ZN(n9001) );
  XNOR2_X1 U9987 ( .A(n11914), .B(n7406), .ZN(n9014) );
  XNOR2_X1 U9988 ( .A(n12064), .B(n7406), .ZN(n9026) );
  XNOR2_X1 U9989 ( .A(n12445), .B(n7406), .ZN(n9045) );
  XNOR2_X1 U9990 ( .A(n12409), .B(n7406), .ZN(n9059) );
  XNOR2_X1 U9991 ( .A(n12735), .B(n7406), .ZN(n9085) );
  XNOR2_X1 U9992 ( .A(n14571), .B(n7406), .ZN(n9079) );
  XNOR2_X1 U9993 ( .A(n12609), .B(n7406), .ZN(n9100) );
  XNOR2_X1 U9994 ( .A(n14562), .B(n7406), .ZN(n9124) );
  XNOR2_X1 U9995 ( .A(n12678), .B(n7406), .ZN(n9110) );
  XNOR2_X1 U9996 ( .A(n14546), .B(n7406), .ZN(n9147) );
  XNOR2_X1 U9997 ( .A(n14275), .B(n7406), .ZN(n9159) );
  XNOR2_X1 U9998 ( .A(n14537), .B(n7406), .ZN(n9172) );
  XNOR2_X1 U9999 ( .A(n14196), .B(n7406), .ZN(n9200) );
  XNOR2_X1 U10000 ( .A(n14149), .B(n7406), .ZN(n9228) );
  XNOR2_X1 U10001 ( .A(n14135), .B(n7406), .ZN(n9238) );
  XNOR2_X1 U10002 ( .A(n14356), .B(n7406), .ZN(n9267) );
  INV_X1 U10003 ( .A(n7418), .ZN(n13934) );
  NOR2_X2 U10004 ( .A1(n8669), .A2(n7420), .ZN(n8742) );
  NAND4_X1 U10005 ( .A1(n8531), .A2(n8532), .A3(n8533), .A4(n7421), .ZN(n7420)
         );
  AND2_X1 U10006 ( .A1(n8743), .A2(n6598), .ZN(n7422) );
  NAND2_X1 U10007 ( .A1(n8744), .A2(n7422), .ZN(n7423) );
  INV_X1 U10008 ( .A(n7423), .ZN(n8881) );
  INV_X1 U10009 ( .A(n11587), .ZN(n7424) );
  NAND2_X1 U10010 ( .A1(n13337), .A2(n7427), .ZN(n7426) );
  NAND3_X2 U10011 ( .A1(n8511), .A2(n8512), .A3(n7172), .ZN(n11287) );
  NAND2_X1 U10012 ( .A1(n7449), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U10013 ( .A1(n7899), .A2(n7449), .ZN(n13485) );
  NAND2_X1 U10014 ( .A1(n8460), .A2(n7451), .ZN(n7450) );
  NAND2_X1 U10015 ( .A1(n7450), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7808) );
  NAND2_X1 U10016 ( .A1(n12507), .A2(n12508), .ZN(n12506) );
  NAND2_X2 U10017 ( .A1(n8957), .A2(n10377), .ZN(n8969) );
  NAND2_X1 U10018 ( .A1(n8773), .A2(n7471), .ZN(n7470) );
  NAND2_X1 U10019 ( .A1(n8773), .A2(n7476), .ZN(n7475) );
  NAND2_X1 U10020 ( .A1(n8772), .A2(n8777), .ZN(n7477) );
  OAI21_X2 U10021 ( .B1(n8815), .B2(n7478), .A(n8818), .ZN(n8826) );
  INV_X1 U10022 ( .A(n13477), .ZN(n7485) );
  NAND2_X1 U10023 ( .A1(n7901), .A2(n13477), .ZN(n7483) );
  NOR2_X1 U10024 ( .A1(n7484), .A2(n13493), .ZN(n13496) );
  INV_X1 U10025 ( .A(n7881), .ZN(n7487) );
  INV_X1 U10026 ( .A(n7494), .ZN(n7489) );
  INV_X1 U10027 ( .A(n11344), .ZN(n7497) );
  INV_X1 U10028 ( .A(n10738), .ZN(n7509) );
  NAND2_X1 U10029 ( .A1(n7513), .A2(n7515), .ZN(n7514) );
  INV_X1 U10030 ( .A(n13459), .ZN(n7513) );
  OR2_X1 U10031 ( .A1(n11017), .A2(n13713), .ZN(n7518) );
  NAND2_X2 U10032 ( .A1(n7519), .A2(n9645), .ZN(n11830) );
  AOI21_X2 U10033 ( .B1(n7522), .B2(n12710), .A(n7521), .ZN(n7520) );
  OAI21_X1 U10034 ( .B1(n15030), .B2(n7528), .A(n7525), .ZN(n7529) );
  NAND2_X1 U10035 ( .A1(n12023), .A2(n12028), .ZN(n7542) );
  NOR2_X2 U10036 ( .A1(n9974), .A2(n9584), .ZN(n9585) );
  INV_X1 U10037 ( .A(n8895), .ZN(n7581) );
  NAND2_X1 U10038 ( .A1(n8160), .A2(n7586), .ZN(n7585) );
  NAND2_X1 U10039 ( .A1(n8211), .A2(n7592), .ZN(n7591) );
  NAND2_X1 U10040 ( .A1(n8444), .A2(n7603), .ZN(n7600) );
  INV_X1 U10041 ( .A(n14096), .ZN(n7607) );
  XNOR2_X1 U10042 ( .A(n14079), .B(n9474), .ZN(n8884) );
  NAND2_X1 U10043 ( .A1(n8056), .A2(n12111), .ZN(n7623) );
  NAND2_X1 U10044 ( .A1(n7623), .A2(n12110), .ZN(n7622) );
  NAND2_X1 U10045 ( .A1(n7624), .A2(n7623), .ZN(n8418) );
  NAND2_X1 U10046 ( .A1(n7624), .A2(n7622), .ZN(n8431) );
  XNOR2_X1 U10047 ( .A(n12981), .B(n13028), .ZN(n9566) );
  NAND2_X1 U10048 ( .A1(n13121), .A2(n7637), .ZN(n7635) );
  OAI22_X1 U10049 ( .A1(n8429), .A2(n7644), .B1(n8488), .B2(n13582), .ZN(n7642) );
  NAND2_X1 U10050 ( .A1(n13634), .A2(n6437), .ZN(n7647) );
  INV_X1 U10051 ( .A(n13611), .ZN(n7656) );
  OAI21_X1 U10052 ( .B1(n13592), .B2(n13147), .A(n13145), .ZN(n13581) );
  NAND2_X1 U10053 ( .A1(n7673), .A2(n6573), .ZN(n9347) );
  AOI21_X1 U10054 ( .B1(n14707), .B2(n14708), .A(n7782), .ZN(n14714) );
  INV_X1 U10055 ( .A(n7782), .ZN(n7679) );
  NAND2_X1 U10056 ( .A1(n8602), .A2(n7682), .ZN(n8606) );
  NAND3_X1 U10057 ( .A1(n8599), .A2(n7682), .A3(n8600), .ZN(n8607) );
  NAND2_X1 U10058 ( .A1(n8590), .A2(n7682), .ZN(n8591) );
  NAND2_X1 U10059 ( .A1(n8589), .A2(SI_4_), .ZN(n7682) );
  NAND2_X1 U10060 ( .A1(n12212), .A2(n7693), .ZN(n7692) );
  NAND2_X1 U10061 ( .A1(n7695), .A2(n7694), .ZN(n12626) );
  NAND2_X1 U10062 ( .A1(n10904), .A2(n9902), .ZN(n7697) );
  OAI21_X1 U10063 ( .B1(n7701), .B2(n15354), .A(n12031), .ZN(n12032) );
  NAND2_X1 U10064 ( .A1(n7702), .A2(n9994), .ZN(n11315) );
  OAI21_X1 U10065 ( .B1(n11250), .B2(n11251), .A(n7702), .ZN(n11680) );
  NAND2_X1 U10066 ( .A1(n15127), .A2(n7713), .ZN(n7712) );
  OAI21_X1 U10067 ( .B1(n15127), .B2(n7716), .A(n7713), .ZN(n15068) );
  OAI21_X1 U10068 ( .B1(n12555), .B2(n12714), .A(n7718), .ZN(n12763) );
  NAND2_X1 U10069 ( .A1(n15014), .A2(n6578), .ZN(n7722) );
  NAND3_X1 U10070 ( .A1(n7721), .A2(n7720), .A3(n7722), .ZN(n7728) );
  NAND3_X1 U10071 ( .A1(n7722), .A2(n7724), .A3(n7721), .ZN(n13198) );
  NAND2_X1 U10072 ( .A1(n12188), .A2(n7733), .ZN(n7731) );
  NAND2_X1 U10073 ( .A1(n9586), .A2(n9585), .ZN(n9603) );
  NAND2_X1 U10074 ( .A1(n10369), .A2(n10368), .ZN(n14112) );
  NAND2_X1 U10075 ( .A1(n7755), .A2(n7753), .ZN(n10349) );
  NOR3_X2 U10076 ( .A1(n15054), .A2(n10626), .A3(n7757), .ZN(n14998) );
  AND2_X2 U10077 ( .A1(n15041), .A2(n7759), .ZN(n15020) );
  AND3_X2 U10078 ( .A1(n7763), .A2(n7760), .A3(n12565), .ZN(n15269) );
  NAND3_X1 U10079 ( .A1(n7763), .A2(n12565), .A3(n7762), .ZN(n7764) );
  INV_X1 U10080 ( .A(n7764), .ZN(n15268) );
  NAND2_X1 U10081 ( .A1(n11508), .A2(n11564), .ZN(n7765) );
  NAND4_X1 U10082 ( .A1(n11770), .A2(n11508), .A3(n11564), .A4(n7768), .ZN(
        n12020) );
  NOR2_X2 U10083 ( .A1(n7766), .A2(n7765), .ZN(n12021) );
  NAND3_X1 U10084 ( .A1(n11770), .A2(n7768), .A3(n7767), .ZN(n7766) );
  NAND2_X1 U10085 ( .A1(n15328), .A2(n15183), .ZN(n15167) );
  INV_X1 U10086 ( .A(n7772), .ZN(n15219) );
  AOI21_X1 U10087 ( .B1(n10604), .B2(n10603), .A(n10602), .ZN(n10606) );
  NOR2_X1 U10088 ( .A1(n10604), .A2(n10603), .ZN(n10605) );
  XNOR2_X1 U10089 ( .A(n8831), .B(n8827), .ZN(n12543) );
  NAND2_X1 U10090 ( .A1(n9355), .A2(n9354), .ZN(n9513) );
  NAND2_X1 U10091 ( .A1(n11375), .A2(n13720), .ZN(n11441) );
  AOI21_X1 U10092 ( .B1(n13668), .B2(n13676), .A(n13667), .ZN(n13738) );
  NAND2_X1 U10093 ( .A1(n13524), .A2(n13523), .ZN(n13667) );
  NAND2_X1 U10094 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), 
        .ZN(n7855) );
  OAI21_X1 U10095 ( .B1(n10478), .B2(n7048), .A(n10474), .ZN(n10477) );
  MUX2_X2 U10096 ( .A(n15277), .B(n15373), .S(n15554), .Z(n15278) );
  MUX2_X2 U10097 ( .A(n15374), .B(n15373), .S(n15550), .Z(n15375) );
  INV_X1 U10098 ( .A(n15012), .ZN(n15380) );
  CLKBUF_X1 U10099 ( .A(n11440), .Z(n11725) );
  AOI21_X1 U10100 ( .B1(n11154), .B2(n10292), .A(n10090), .ZN(n11147) );
  XNOR2_X1 U10101 ( .A(n9346), .B(n13165), .ZN(n13534) );
  NAND2_X1 U10102 ( .A1(n9516), .A2(n10385), .ZN(n10331) );
  OAI22_X1 U10103 ( .A1(n10105), .A2(n11159), .B1(n7048), .B2(n10299), .ZN(
        n10106) );
  NAND2_X1 U10104 ( .A1(n10096), .A2(n11498), .ZN(n10488) );
  INV_X1 U10105 ( .A(n8950), .ZN(n8891) );
  OR2_X1 U10106 ( .A1(n13412), .A2(n8273), .ZN(n7773) );
  OR2_X1 U10107 ( .A1(n13412), .A2(n12284), .ZN(n7774) );
  INV_X1 U10108 ( .A(n10252), .ZN(n10117) );
  OR2_X1 U10109 ( .A1(n14355), .A2(n14346), .ZN(n7775) );
  AND2_X1 U10110 ( .A1(n12916), .A2(n13239), .ZN(n7776) );
  AND2_X1 U10111 ( .A1(n15151), .A2(n14756), .ZN(n7777) );
  OR2_X1 U10112 ( .A1(n8789), .A2(SI_21_), .ZN(n7778) );
  AND3_X1 U10113 ( .A1(n8741), .A2(n8740), .A3(n8739), .ZN(n7779) );
  AND2_X1 U10114 ( .A1(n7609), .A2(n14093), .ZN(n7780) );
  OR2_X1 U10115 ( .A1(n7609), .A2(n14627), .ZN(n7781) );
  AND2_X1 U10116 ( .A1(n10218), .A2(n10217), .ZN(n7782) );
  AND3_X1 U10117 ( .A1(n13849), .A2(n13848), .A3(n13915), .ZN(n7783) );
  NOR2_X1 U10118 ( .A1(n12482), .A2(n9091), .ZN(n7785) );
  AND2_X1 U10119 ( .A1(n12160), .A2(n12165), .ZN(n7787) );
  AND2_X1 U10120 ( .A1(n14247), .A2(n14245), .ZN(n7788) );
  INV_X1 U10121 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14630) );
  AND2_X1 U10122 ( .A1(n12983), .A2(SI_30_), .ZN(n7789) );
  NAND2_X1 U10123 ( .A1(n9226), .A2(n9225), .ZN(n14160) );
  INV_X1 U10124 ( .A(n13724), .ZN(n13641) );
  INV_X1 U10125 ( .A(n14582), .ZN(n8939) );
  INV_X1 U10126 ( .A(n14797), .ZN(n14754) );
  INV_X1 U10127 ( .A(n9523), .ZN(n14289) );
  AND2_X1 U10128 ( .A1(n10638), .A2(n7784), .ZN(n7790) );
  INV_X1 U10129 ( .A(n12046), .ZN(n10695) );
  XOR2_X1 U10130 ( .A(P1_IR_REG_19__SCAN_IN), .B(P1_IR_REG_31__SCAN_IN), .Z(
        n7791) );
  AND2_X1 U10131 ( .A1(n8733), .A2(n8725), .ZN(n7792) );
  INV_X1 U10132 ( .A(n13180), .ZN(n12998) );
  XOR2_X1 U10133 ( .A(n9532), .B(n11455), .Z(n7793) );
  INV_X1 U10134 ( .A(n9474), .ZN(n14077) );
  OR2_X1 U10135 ( .A1(n12855), .A2(n13275), .ZN(n7795) );
  INV_X1 U10136 ( .A(n12189), .ZN(n9725) );
  XNOR2_X1 U10137 ( .A(n12735), .B(n14329), .ZN(n12724) );
  INV_X1 U10138 ( .A(n12724), .ZN(n10344) );
  INV_X1 U10139 ( .A(n15236), .ZN(n9812) );
  OR2_X1 U10140 ( .A1(n8787), .A2(SI_20_), .ZN(n7796) );
  INV_X1 U10141 ( .A(n15213), .ZN(n9825) );
  NOR2_X1 U10142 ( .A1(n12487), .A2(n12486), .ZN(n7798) );
  AND2_X1 U10143 ( .A1(n10558), .A2(n10557), .ZN(n7799) );
  AND2_X1 U10144 ( .A1(n13534), .A2(n15720), .ZN(n7800) );
  INV_X1 U10145 ( .A(n10475), .ZN(n10476) );
  NAND2_X1 U10146 ( .A1(n9355), .A2(n6514), .ZN(n9361) );
  INV_X1 U10147 ( .A(n9411), .ZN(n9412) );
  AOI21_X1 U10148 ( .B1(n9414), .B2(n9413), .A(n9412), .ZN(n9423) );
  AND2_X1 U10149 ( .A1(n10575), .A2(n10574), .ZN(n10576) );
  INV_X1 U10150 ( .A(n13007), .ZN(n13060) );
  INV_X1 U10151 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8740) );
  INV_X1 U10152 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9581) );
  OR2_X1 U10153 ( .A1(n7978), .A2(n11344), .ZN(n7979) );
  AND2_X1 U10154 ( .A1(n13009), .A2(n11724), .ZN(n8150) );
  INV_X1 U10155 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7801) );
  INV_X1 U10156 ( .A(n8577), .ZN(n8539) );
  NAND2_X1 U10157 ( .A1(n10017), .A2(n15159), .ZN(n9879) );
  INV_X1 U10158 ( .A(n13018), .ZN(n8279) );
  INV_X1 U10159 ( .A(n11146), .ZN(n10091) );
  INV_X1 U10160 ( .A(n15085), .ZN(n10023) );
  NAND2_X1 U10161 ( .A1(n8838), .A2(n14412), .ZN(n8839) );
  NAND2_X1 U10162 ( .A1(n8817), .A2(SI_24_), .ZN(n8818) );
  INV_X1 U10163 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9727) );
  INV_X1 U10164 ( .A(n11580), .ZN(n11581) );
  INV_X1 U10165 ( .A(n13194), .ZN(n8086) );
  OR2_X1 U10166 ( .A1(n11017), .A2(n7995), .ZN(n7996) );
  XNOR2_X1 U10167 ( .A(n12994), .B(n13522), .ZN(n13028) );
  INV_X1 U10168 ( .A(n13537), .ZN(n13539) );
  INV_X1 U10169 ( .A(n12076), .ZN(n8479) );
  NAND2_X1 U10170 ( .A1(n10808), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8011) );
  AND2_X1 U10171 ( .A1(n9151), .A2(n13876), .ZN(n9152) );
  INV_X1 U10172 ( .A(n11639), .ZN(n9006) );
  INV_X1 U10173 ( .A(n9213), .ZN(n9204) );
  NAND2_X1 U10174 ( .A1(n9254), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9280) );
  INV_X1 U10175 ( .A(n14143), .ZN(n10365) );
  INV_X1 U10176 ( .A(n11485), .ZN(n9354) );
  AND2_X1 U10177 ( .A1(n12403), .A2(n12402), .ZN(n14330) );
  OR2_X1 U10178 ( .A1(n10255), .A2(n10254), .ZN(n10256) );
  NAND2_X1 U10179 ( .A1(n10690), .A2(n10689), .ZN(n10691) );
  INV_X1 U10180 ( .A(n10662), .ZN(n15058) );
  NOR2_X1 U10181 ( .A1(n10023), .A2(n10022), .ZN(n10024) );
  INV_X1 U10182 ( .A(n15139), .ZN(n10020) );
  OR2_X1 U10183 ( .A1(n9691), .A2(n9588), .ZN(n9595) );
  CLKBUF_X3 U10184 ( .A(n9654), .Z(n9902) );
  INV_X1 U10185 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9570) );
  NAND2_X1 U10186 ( .A1(n8704), .A2(n10973), .ZN(n8722) );
  INV_X1 U10187 ( .A(n12924), .ZN(n12925) );
  INV_X1 U10188 ( .A(n13613), .ZN(n13320) );
  INV_X1 U10189 ( .A(n13357), .ZN(n13331) );
  OR2_X1 U10190 ( .A1(n11282), .A2(n11281), .ZN(n13359) );
  CLKBUF_X3 U10191 ( .A(n8126), .Z(n9327) );
  INV_X1 U10192 ( .A(n13722), .ZN(n13643) );
  AND2_X1 U10193 ( .A1(n8025), .A2(n8024), .ZN(n8234) );
  AND2_X1 U10194 ( .A1(n8550), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8122) );
  INV_X1 U10195 ( .A(n9270), .ZN(n9271) );
  AND2_X1 U10196 ( .A1(n9280), .A2(n9257), .ZN(n14097) );
  INV_X1 U10197 ( .A(n14378), .ZN(n14168) );
  XNOR2_X1 U10198 ( .A(n14180), .B(n14191), .ZN(n14177) );
  INV_X1 U10199 ( .A(n13967), .ZN(n12675) );
  INV_X1 U10200 ( .A(n9522), .ZN(n12573) );
  INV_X1 U10201 ( .A(n9619), .ZN(n9654) );
  NAND2_X1 U10202 ( .A1(n14742), .A2(n14741), .ZN(n14740) );
  INV_X1 U10203 ( .A(n14766), .ZN(n14778) );
  INV_X1 U10204 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14823) );
  XNOR2_X1 U10205 ( .A(n15049), .B(n15058), .ZN(n15050) );
  XNOR2_X1 U10206 ( .A(n15113), .B(n15089), .ZN(n15111) );
  NOR2_X1 U10207 ( .A1(n12763), .A2(n12764), .ZN(n15250) );
  AND2_X1 U10208 ( .A1(n10869), .A2(n14839), .ZN(n15257) );
  OR2_X1 U10209 ( .A1(n15533), .A2(n11497), .ZN(n15234) );
  INV_X1 U10210 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n10067) );
  AND2_X1 U10211 ( .A1(n8755), .A2(n8736), .ZN(n8749) );
  INV_X1 U10212 ( .A(n8204), .ZN(n12168) );
  INV_X1 U10213 ( .A(n13570), .ZN(n13541) );
  AND2_X1 U10214 ( .A1(n8002), .A2(n13188), .ZN(n13495) );
  INV_X1 U10215 ( .A(n11412), .ZN(n13645) );
  NAND2_X1 U10216 ( .A1(n15731), .A2(n9322), .ZN(n9544) );
  AND4_X1 U10217 ( .A1(n9549), .A2(n8521), .A3(n11171), .A4(n8520), .ZN(n8522)
         );
  INV_X1 U10218 ( .A(n13790), .ZN(n13774) );
  OR2_X1 U10219 ( .A1(n11047), .A2(n11046), .ZN(n11064) );
  INV_X1 U10220 ( .A(n14159), .ZN(n14191) );
  AND2_X1 U10221 ( .A1(n9277), .A2(n9269), .ZN(n13915) );
  OR2_X1 U10222 ( .A1(n13845), .A2(n9464), .ZN(n9286) );
  NOR2_X1 U10223 ( .A1(n11077), .A2(n11078), .ZN(n11418) );
  INV_X1 U10224 ( .A(n15591), .ZN(n15613) );
  AND2_X1 U10225 ( .A1(n9288), .A2(n8885), .ZN(n14286) );
  INV_X1 U10226 ( .A(n14341), .ZN(n15622) );
  NAND2_X1 U10227 ( .A1(n15645), .A2(n9275), .ZN(n15619) );
  INV_X1 U10228 ( .A(n14627), .ZN(n10703) );
  AND2_X1 U10229 ( .A1(n8931), .A2(n8912), .ZN(n15634) );
  AND2_X1 U10230 ( .A1(n10316), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14776) );
  AND2_X1 U10231 ( .A1(n10315), .A2(n11496), .ZN(n14771) );
  AND2_X1 U10232 ( .A1(n14771), .A2(n15547), .ZN(n14795) );
  OR2_X1 U10233 ( .A1(n9691), .A2(n9613), .ZN(n9616) );
  NOR2_X1 U10234 ( .A1(n11266), .A2(n11265), .ZN(n11606) );
  INV_X1 U10235 ( .A(n14989), .ZN(n15513) );
  NAND2_X1 U10236 ( .A1(n14998), .A2(n15380), .ZN(n15008) );
  AND2_X1 U10237 ( .A1(n10562), .A2(n10564), .ZN(n15192) );
  NAND2_X1 U10238 ( .A1(n10471), .A2(n9984), .ZN(n15260) );
  INV_X1 U10239 ( .A(n15174), .ZN(n15522) );
  OR2_X1 U10240 ( .A1(n12033), .A2(n12032), .ZN(n15545) );
  INV_X1 U10241 ( .A(n15354), .ZN(n15370) );
  AND2_X1 U10242 ( .A1(n10084), .A2(n10856), .ZN(n11496) );
  AND2_X1 U10243 ( .A1(n7969), .A2(n7968), .ZN(n15671) );
  AND2_X1 U10244 ( .A1(n11187), .A2(n11186), .ZN(n13351) );
  INV_X1 U10245 ( .A(n13569), .ZN(n13595) );
  INV_X1 U10246 ( .A(n13293), .ZN(n13374) );
  OR2_X1 U10247 ( .A1(n15691), .A2(n9348), .ZN(n13663) );
  INV_X1 U10248 ( .A(n15734), .ZN(n15731) );
  OR2_X1 U10249 ( .A1(n15721), .A2(n9564), .ZN(n13793) );
  INV_X1 U10250 ( .A(n8087), .ZN(n12893) );
  INV_X1 U10251 ( .A(n9299), .ZN(n9300) );
  INV_X1 U10252 ( .A(n13915), .ZN(n13956) );
  OR2_X1 U10253 ( .A1(n9541), .A2(n9540), .ZN(n9542) );
  NAND2_X1 U10254 ( .A1(n9236), .A2(n9235), .ZN(n13962) );
  INV_X1 U10255 ( .A(n15622), .ZN(n14312) );
  AND2_X1 U10256 ( .A1(n10452), .A2(n15619), .ZN(n14341) );
  AOI21_X1 U10257 ( .B1(n9474), .B2(n8939), .A(n8938), .ZN(n8940) );
  OR2_X1 U10258 ( .A1(n10440), .A2(n8936), .ZN(n15668) );
  INV_X1 U10259 ( .A(n14232), .ZN(n14608) );
  INV_X1 U10260 ( .A(n12735), .ZN(n14628) );
  OR2_X1 U10261 ( .A1(n10448), .A2(n10440), .ZN(n15664) );
  INV_X1 U10262 ( .A(n15639), .ZN(n15637) );
  AND2_X1 U10263 ( .A1(n9293), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15645) );
  INV_X1 U10265 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10905) );
  INV_X1 U10266 ( .A(n15171), .ZN(n15328) );
  INV_X1 U10267 ( .A(n12964), .ZN(n15038) );
  OR2_X1 U10268 ( .A1(n15533), .A2(n14993), .ZN(n15174) );
  AND2_X1 U10269 ( .A1(n13202), .A2(n15217), .ZN(n15533) );
  NAND2_X1 U10270 ( .A1(n10626), .A2(n12686), .ZN(n10081) );
  OR2_X1 U10271 ( .A1(n10075), .A2(n11489), .ZN(n15552) );
  INV_X1 U10272 ( .A(n15271), .ZN(n15414) );
  OR2_X1 U10273 ( .A1(n10075), .A2(n10066), .ZN(n15549) );
  AND2_X1 U10274 ( .A1(n10868), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10856) );
  INV_X1 U10275 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11022) );
  INV_X1 U10276 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10906) );
  AND2_X1 U10277 ( .A1(n12838), .A2(n12837), .ZN(n12863) );
  NAND2_X1 U10278 ( .A1(n7775), .A2(n10470), .ZN(P2_U3236) );
  NOR2_X1 U10279 ( .A1(n7819), .A2(n7817), .ZN(n7803) );
  AND2_X2 U10280 ( .A1(n7803), .A2(n7846), .ZN(n7833) );
  NAND2_X1 U10281 ( .A1(n7804), .A2(n7813), .ZN(n7834) );
  NOR2_X2 U10282 ( .A1(n7834), .A2(n7814), .ZN(n7805) );
  INV_X1 U10283 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8462) );
  INV_X1 U10284 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7806) );
  INV_X1 U10285 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7807) );
  XNOR2_X1 U10286 ( .A(n7808), .B(n7809), .ZN(n8510) );
  NOR2_X1 U10287 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_22__SCAN_IN), 
        .ZN(n7811) );
  NAND2_X1 U10288 ( .A1(n7826), .A2(n7816), .ZN(n7829) );
  NAND2_X1 U10289 ( .A1(n7829), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7812) );
  INV_X1 U10290 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7815) );
  INV_X1 U10291 ( .A(n7826), .ZN(n7827) );
  NAND2_X1 U10292 ( .A1(n7827), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7828) );
  MUX2_X1 U10293 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7828), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n7830) );
  NAND2_X1 U10294 ( .A1(n7830), .A2(n7829), .ZN(n13809) );
  OR3_X1 U10295 ( .A1(n8510), .A2(n12959), .A3(n13809), .ZN(n11170) );
  INV_X1 U10296 ( .A(n11170), .ZN(n7832) );
  NAND2_X1 U10297 ( .A1(n7909), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7831) );
  XNOR2_X1 U10298 ( .A(n7831), .B(n7452), .ZN(n11169) );
  AND2_X2 U10299 ( .A1(n7832), .A2(n13797), .ZN(P3_U3897) );
  INV_X1 U10300 ( .A(n7833), .ZN(n7843) );
  INV_X1 U10301 ( .A(n7882), .ZN(n7838) );
  INV_X1 U10302 ( .A(n7834), .ZN(n7835) );
  NAND2_X1 U10303 ( .A1(n7838), .A2(n7835), .ZN(n7897) );
  NAND2_X1 U10304 ( .A1(n7897), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7836) );
  INV_X1 U10305 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13713) );
  NAND2_X1 U10306 ( .A1(n7838), .A2(n7837), .ZN(n7888) );
  OR2_X1 U10307 ( .A1(n7888), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n7890) );
  INV_X1 U10308 ( .A(n7890), .ZN(n7839) );
  INV_X1 U10309 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7891) );
  NAND2_X1 U10310 ( .A1(n7839), .A2(n7891), .ZN(n7841) );
  NAND2_X1 U10311 ( .A1(n7841), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7840) );
  MUX2_X1 U10312 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7840), .S(
        P3_IR_REG_14__SCAN_IN), .Z(n7842) );
  OR2_X1 U10313 ( .A1(n7841), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n7894) );
  NAND2_X1 U10314 ( .A1(n7842), .A2(n7894), .ZN(n10977) );
  NAND2_X1 U10315 ( .A1(n7843), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7844) );
  MUX2_X1 U10316 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7844), .S(
        P3_IR_REG_10__SCAN_IN), .Z(n7845) );
  NAND2_X1 U10317 ( .A1(n7845), .A2(n7882), .ZN(n10845) );
  INV_X1 U10318 ( .A(n7863), .ZN(n7848) );
  NOR2_X1 U10319 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .ZN(
        n7847) );
  NAND2_X1 U10320 ( .A1(n7848), .A2(n7847), .ZN(n7851) );
  NAND2_X1 U10321 ( .A1(n7849), .A2(n7874), .ZN(n7878) );
  NAND2_X1 U10322 ( .A1(n7878), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7850) );
  INV_X1 U10323 ( .A(n11529), .ZN(n10824) );
  NAND2_X1 U10324 ( .A1(n7851), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7852) );
  XNOR2_X1 U10325 ( .A(n7852), .B(P3_IR_REG_6__SCAN_IN), .ZN(n8188) );
  INV_X1 U10326 ( .A(n8188), .ZN(n10820) );
  INV_X1 U10327 ( .A(n7975), .ZN(n7853) );
  INV_X1 U10328 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n11451) );
  XNOR2_X1 U10329 ( .A(n7973), .B(n11451), .ZN(n11106) );
  NAND2_X1 U10330 ( .A1(n7802), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7856) );
  NAND2_X1 U10331 ( .A1(n8113), .A2(n7856), .ZN(n7858) );
  INV_X1 U10332 ( .A(n7856), .ZN(n11369) );
  INV_X1 U10333 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7857) );
  NAND2_X1 U10334 ( .A1(n11369), .A2(n7857), .ZN(n7859) );
  NAND2_X1 U10335 ( .A1(n7858), .A2(n7859), .ZN(n11402) );
  INV_X1 U10336 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n11401) );
  NAND2_X1 U10337 ( .A1(n11404), .A2(n7859), .ZN(n11105) );
  NAND2_X1 U10338 ( .A1(n11106), .A2(n11105), .ZN(n11104) );
  NAND2_X1 U10339 ( .A1(n11122), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7860) );
  NAND2_X1 U10340 ( .A1(n7861), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7862) );
  NAND2_X1 U10341 ( .A1(n11328), .A2(n11198), .ZN(n7864) );
  NAND2_X1 U10342 ( .A1(n7863), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7867) );
  INV_X1 U10343 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15725) );
  XNOR2_X1 U10344 ( .A(n11219), .B(n15725), .ZN(n11197) );
  NAND2_X1 U10345 ( .A1(n7864), .A2(n11197), .ZN(n11201) );
  NAND2_X1 U10346 ( .A1(n11219), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7865) );
  NAND2_X1 U10347 ( .A1(n7867), .A2(n7866), .ZN(n7868) );
  NAND2_X1 U10348 ( .A1(n7868), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7870) );
  XNOR2_X1 U10349 ( .A(n7869), .B(n7870), .ZN(n11041) );
  NAND2_X1 U10350 ( .A1(n7871), .A2(n11041), .ZN(n10737) );
  AND2_X2 U10351 ( .A1(n7872), .A2(n10737), .ZN(n11027) );
  INV_X1 U10352 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15729) );
  XNOR2_X1 U10353 ( .A(n8188), .B(n15729), .ZN(n10738) );
  NAND2_X1 U10354 ( .A1(n7873), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7875) );
  XNOR2_X1 U10355 ( .A(n7875), .B(n7874), .ZN(n11352) );
  INV_X1 U10356 ( .A(n11352), .ZN(n7986) );
  AOI21_X1 U10357 ( .B1(n7876), .B2(n7986), .A(n7877), .ZN(n11345) );
  NAND2_X1 U10358 ( .A1(n11345), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n11346) );
  INV_X1 U10359 ( .A(n7877), .ZN(n11530) );
  INV_X1 U10360 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n12184) );
  XNOR2_X1 U10361 ( .A(n11529), .B(n12184), .ZN(n11531) );
  OAI21_X1 U10362 ( .B1(n7878), .B2(P3_IR_REG_8__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7880) );
  XNOR2_X1 U10363 ( .A(n7880), .B(n7879), .ZN(n11849) );
  XNOR2_X1 U10364 ( .A(n10845), .B(P3_REG1_REG_10__SCAN_IN), .ZN(n13394) );
  INV_X1 U10365 ( .A(n7885), .ZN(n7887) );
  NAND2_X1 U10366 ( .A1(n7882), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7883) );
  MUX2_X1 U10367 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7883), .S(
        P3_IR_REG_11__SCAN_IN), .Z(n7884) );
  NAND2_X1 U10368 ( .A1(n7884), .A2(n7888), .ZN(n10850) );
  INV_X1 U10369 ( .A(n10850), .ZN(n12659) );
  INV_X1 U10370 ( .A(n7511), .ZN(n7886) );
  INV_X1 U10371 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n12656) );
  NAND2_X1 U10372 ( .A1(n7888), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7889) );
  XNOR2_X1 U10373 ( .A(n7889), .B(P3_IR_REG_12__SCAN_IN), .ZN(n13412) );
  XNOR2_X1 U10374 ( .A(n13412), .B(P3_REG1_REG_12__SCAN_IN), .ZN(n13416) );
  INV_X1 U10375 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n8273) );
  NAND2_X1 U10376 ( .A1(n7890), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7892) );
  OAI21_X1 U10377 ( .B1(n7893), .B2(n13430), .A(n10714), .ZN(n13423) );
  INV_X1 U10378 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n13424) );
  OR2_X2 U10379 ( .A1(n13423), .A2(n13424), .ZN(n13421) );
  XNOR2_X1 U10380 ( .A(n10977), .B(P3_REG1_REG_14__SCAN_IN), .ZN(n10715) );
  NAND2_X1 U10381 ( .A1(n7894), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7895) );
  XNOR2_X1 U10382 ( .A(n7895), .B(n6752), .ZN(n13449) );
  INV_X1 U10383 ( .A(n13449), .ZN(n7993) );
  XNOR2_X1 U10384 ( .A(n11017), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n13458) );
  OAI21_X1 U10385 ( .B1(n7897), .B2(P3_IR_REG_16__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7898) );
  MUX2_X1 U10386 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7898), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n7899) );
  NAND2_X1 U10387 ( .A1(n7900), .A2(n13485), .ZN(n7901) );
  OAI21_X1 U10388 ( .B1(n7900), .B2(n13485), .A(n7901), .ZN(n13477) );
  INV_X1 U10389 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13705) );
  INV_X1 U10390 ( .A(n7901), .ZN(n13494) );
  MUX2_X1 U10391 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7902), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n7903) );
  INV_X1 U10392 ( .A(n6599), .ZN(n11222) );
  NAND2_X1 U10393 ( .A1(n11222), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n7905) );
  INV_X1 U10394 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13703) );
  NAND2_X1 U10395 ( .A1(n6599), .A2(n13703), .ZN(n7904) );
  AND2_X1 U10396 ( .A1(n7905), .A2(n7904), .ZN(n13493) );
  NAND2_X1 U10397 ( .A1(n13492), .A2(n7905), .ZN(n7907) );
  XNOR2_X2 U10398 ( .A(n7906), .B(P3_IR_REG_19__SCAN_IN), .ZN(n11284) );
  XNOR2_X1 U10399 ( .A(n11284), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n7962) );
  NAND2_X1 U10400 ( .A1(n11170), .A2(n13797), .ZN(n9557) );
  OR2_X1 U10401 ( .A1(n11169), .A2(P3_U3151), .ZN(n13193) );
  NAND2_X1 U10402 ( .A1(n9557), .A2(n13193), .ZN(n7969) );
  NAND2_X1 U10403 ( .A1(n6473), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7908) );
  MUX2_X1 U10404 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7908), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n7910) );
  NAND2_X1 U10405 ( .A1(n6547), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7911) );
  NAND2_X1 U10406 ( .A1(n13168), .A2(n11169), .ZN(n7917) );
  INV_X1 U10407 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7914) );
  XNOR2_X2 U10408 ( .A(n7916), .B(n7913), .ZN(n7929) );
  NAND2_X1 U10409 ( .A1(n7917), .A2(n8471), .ZN(n7968) );
  INV_X1 U10410 ( .A(n7968), .ZN(n7918) );
  INV_X2 U10411 ( .A(n7929), .ZN(n11365) );
  MUX2_X1 U10412 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13188), .Z(n7960) );
  MUX2_X1 U10413 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n13188), .Z(n7958) );
  INV_X1 U10414 ( .A(n7958), .ZN(n7959) );
  MUX2_X1 U10415 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n13188), .Z(n7956) );
  MUX2_X1 U10416 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13188), .Z(n7955) );
  MUX2_X1 U10417 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13188), .Z(n7954) );
  INV_X1 U10418 ( .A(n13412), .ZN(n10874) );
  INV_X1 U10419 ( .A(n10845), .ZN(n13393) );
  MUX2_X1 U10420 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13188), .Z(n7951) );
  INV_X1 U10421 ( .A(n7951), .ZN(n7952) );
  MUX2_X1 U10422 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13188), .Z(n7947) );
  INV_X1 U10423 ( .A(n7947), .ZN(n7948) );
  INV_X1 U10424 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15689) );
  NAND2_X1 U10425 ( .A1(n7919), .A2(n8113), .ZN(n11108) );
  INV_X1 U10426 ( .A(n7919), .ZN(n7920) );
  INV_X1 U10427 ( .A(n8113), .ZN(n11409) );
  NAND2_X1 U10428 ( .A1(n7920), .A2(n11409), .ZN(n7921) );
  INV_X1 U10429 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11410) );
  INV_X1 U10430 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n7922) );
  NAND2_X1 U10431 ( .A1(n7923), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11394) );
  NAND2_X1 U10432 ( .A1(n11396), .A2(n11108), .ZN(n7928) );
  INV_X1 U10433 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15680) );
  MUX2_X1 U10434 ( .A(n15680), .B(n11451), .S(n7929), .Z(n7925) );
  INV_X1 U10435 ( .A(n11122), .ZN(n7924) );
  NAND2_X1 U10436 ( .A1(n7925), .A2(n7924), .ZN(n11331) );
  INV_X1 U10437 ( .A(n7925), .ZN(n7926) );
  NAND2_X1 U10438 ( .A1(n7926), .A2(n11122), .ZN(n7927) );
  AND2_X1 U10439 ( .A1(n11331), .A2(n7927), .ZN(n11107) );
  INV_X1 U10440 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11730) );
  INV_X1 U10441 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15723) );
  MUX2_X1 U10442 ( .A(n11730), .B(n15723), .S(n7929), .Z(n7930) );
  NAND2_X1 U10443 ( .A1(n7930), .A2(n7497), .ZN(n7933) );
  INV_X1 U10444 ( .A(n7930), .ZN(n7931) );
  NAND2_X1 U10445 ( .A1(n7931), .A2(n11344), .ZN(n7932) );
  NAND2_X1 U10446 ( .A1(n7933), .A2(n7932), .ZN(n11330) );
  INV_X1 U10447 ( .A(n7933), .ZN(n11212) );
  INV_X1 U10448 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n7980) );
  INV_X1 U10449 ( .A(n11219), .ZN(n10865) );
  NAND2_X1 U10450 ( .A1(n7934), .A2(n10865), .ZN(n11036) );
  INV_X1 U10451 ( .A(n7934), .ZN(n7935) );
  NAND2_X1 U10452 ( .A1(n7935), .A2(n11219), .ZN(n7936) );
  AND2_X1 U10453 ( .A1(n11036), .A2(n7936), .ZN(n11211) );
  INV_X1 U10454 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n14433) );
  INV_X1 U10455 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15727) );
  MUX2_X1 U10456 ( .A(n14433), .B(n15727), .S(n13188), .Z(n7937) );
  NAND2_X1 U10457 ( .A1(n7937), .A2(n7054), .ZN(n7940) );
  INV_X1 U10458 ( .A(n7937), .ZN(n7938) );
  NAND2_X1 U10459 ( .A1(n7938), .A2(n11041), .ZN(n7939) );
  NAND2_X1 U10460 ( .A1(n7940), .A2(n7939), .ZN(n11035) );
  INV_X1 U10461 ( .A(n7940), .ZN(n10741) );
  INV_X1 U10462 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n7985) );
  MUX2_X1 U10463 ( .A(n7985), .B(n15729), .S(n13188), .Z(n7941) );
  INV_X1 U10464 ( .A(n7941), .ZN(n7942) );
  INV_X1 U10465 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n12094) );
  INV_X1 U10466 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15732) );
  MUX2_X1 U10467 ( .A(n12094), .B(n15732), .S(n13188), .Z(n7943) );
  NAND2_X1 U10468 ( .A1(n7943), .A2(n7986), .ZN(n7946) );
  INV_X1 U10469 ( .A(n7943), .ZN(n7944) );
  NAND2_X1 U10470 ( .A1(n7944), .A2(n11352), .ZN(n7945) );
  NAND2_X1 U10471 ( .A1(n7946), .A2(n7945), .ZN(n11355) );
  XOR2_X1 U10472 ( .A(n11529), .B(n7947), .Z(n11521) );
  INV_X1 U10473 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n12225) );
  INV_X1 U10474 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n12297) );
  MUX2_X1 U10475 ( .A(n12225), .B(n12297), .S(n13188), .Z(n7949) );
  NOR2_X1 U10476 ( .A1(n7492), .A2(n7949), .ZN(n11844) );
  INV_X1 U10477 ( .A(n7949), .ZN(n7950) );
  NOR2_X1 U10478 ( .A1(n11849), .A2(n7950), .ZN(n11845) );
  XNOR2_X1 U10479 ( .A(n7951), .B(n10845), .ZN(n13388) );
  MUX2_X1 U10480 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13188), .Z(n7953) );
  XNOR2_X1 U10481 ( .A(n7953), .B(n10850), .ZN(n12657) );
  OAI22_X1 U10482 ( .A1(n12658), .A2(n12657), .B1(n7953), .B2(n10850), .ZN(
        n13408) );
  XOR2_X1 U10483 ( .A(n13412), .B(n7954), .Z(n13409) );
  XOR2_X1 U10484 ( .A(n7955), .B(n13430), .Z(n13426) );
  XNOR2_X1 U10485 ( .A(n10977), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n10710) );
  MUX2_X1 U10486 ( .A(n10715), .B(n10710), .S(n11365), .Z(n10720) );
  XNOR2_X1 U10487 ( .A(n7957), .B(n13449), .ZN(n13445) );
  MUX2_X1 U10488 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n13188), .Z(n13444) );
  XNOR2_X1 U10489 ( .A(n7958), .B(n11017), .ZN(n13465) );
  XOR2_X1 U10490 ( .A(n7960), .B(n13485), .Z(n13480) );
  MUX2_X1 U10491 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13188), .Z(n13507) );
  INV_X1 U10492 ( .A(n7962), .ZN(n7963) );
  INV_X1 U10493 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13625) );
  XNOR2_X1 U10494 ( .A(n11284), .B(n13625), .ZN(n8000) );
  MUX2_X1 U10495 ( .A(n7963), .B(n8000), .S(n11365), .Z(n7964) );
  XNOR2_X1 U10496 ( .A(n7965), .B(n7964), .ZN(n7972) );
  AND2_X1 U10497 ( .A1(n7966), .A2(P3_U3897), .ZN(n13509) );
  INV_X1 U10498 ( .A(n8002), .ZN(n7967) );
  INV_X1 U10499 ( .A(n7966), .ZN(n13800) );
  MUX2_X1 U10500 ( .A(n7967), .B(n13372), .S(n13800), .Z(n13486) );
  INV_X1 U10501 ( .A(n11284), .ZN(n13031) );
  NAND2_X1 U10502 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13250)
         );
  NAND2_X1 U10503 ( .A1(n15671), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7970) );
  OAI211_X1 U10504 ( .C1(n13486), .C2(n13031), .A(n13250), .B(n7970), .ZN(
        n7971) );
  NAND2_X1 U10505 ( .A1(n7802), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7974) );
  NAND2_X1 U10506 ( .A1(n7975), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7976) );
  NAND2_X1 U10507 ( .A1(n11393), .A2(n7976), .ZN(n11113) );
  NAND2_X1 U10508 ( .A1(n11122), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7977) );
  NAND2_X1 U10509 ( .A1(n11112), .A2(n7977), .ZN(n7978) );
  NAND2_X1 U10510 ( .A1(n7978), .A2(n11344), .ZN(n11203) );
  NAND2_X1 U10511 ( .A1(n11335), .A2(n11203), .ZN(n7981) );
  XNOR2_X1 U10512 ( .A(n11219), .B(n7980), .ZN(n11202) );
  NAND2_X1 U10513 ( .A1(n11219), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7982) );
  XNOR2_X1 U10514 ( .A(n8188), .B(n7985), .ZN(n10735) );
  AOI21_X1 U10515 ( .B1(n7987), .B2(n7986), .A(n7988), .ZN(n11349) );
  INV_X1 U10516 ( .A(n7988), .ZN(n11524) );
  INV_X1 U10517 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n12116) );
  XNOR2_X1 U10518 ( .A(n11529), .B(n12116), .ZN(n11525) );
  INV_X1 U10519 ( .A(n7989), .ZN(n13398) );
  XNOR2_X1 U10520 ( .A(n10845), .B(P3_REG2_REG_10__SCAN_IN), .ZN(n13399) );
  INV_X1 U10521 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12662) );
  XNOR2_X1 U10522 ( .A(n13412), .B(P3_REG2_REG_12__SCAN_IN), .ZN(n13413) );
  INV_X1 U10523 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12284) );
  INV_X1 U10524 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13431) );
  AOI21_X1 U10525 ( .B1(n13434), .B2(n10709), .A(n10710), .ZN(n10708) );
  XNOR2_X1 U10526 ( .A(n11017), .B(P3_REG2_REG_16__SCAN_IN), .ZN(n13454) );
  INV_X1 U10527 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n7995) );
  INV_X1 U10528 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13657) );
  NAND2_X1 U10529 ( .A1(n11222), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7999) );
  INV_X1 U10530 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13647) );
  NAND2_X1 U10531 ( .A1(n6599), .A2(n13647), .ZN(n7998) );
  NAND2_X1 U10532 ( .A1(n7999), .A2(n7998), .ZN(n13502) );
  NAND2_X1 U10533 ( .A1(n13800), .A2(n11365), .ZN(n8470) );
  INV_X1 U10534 ( .A(n8470), .ZN(n8001) );
  NAND2_X1 U10535 ( .A1(n8003), .A2(n13504), .ZN(n8004) );
  NAND2_X1 U10536 ( .A1(n8122), .A2(n8112), .ZN(n8111) );
  NAND2_X1 U10537 ( .A1(n8111), .A2(n8005), .ZN(n8133) );
  AND2_X1 U10538 ( .A1(n8007), .A2(n8006), .ZN(n8132) );
  NAND2_X1 U10539 ( .A1(n8133), .A2(n8132), .ZN(n8131) );
  NAND2_X1 U10540 ( .A1(n10790), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8008) );
  NAND2_X1 U10541 ( .A1(n10795), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8010) );
  NAND2_X1 U10542 ( .A1(n10810), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8013) );
  INV_X1 U10543 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10788) );
  NAND2_X1 U10544 ( .A1(n10788), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8012) );
  AND2_X1 U10545 ( .A1(n8013), .A2(n8012), .ZN(n8173) );
  NAND2_X1 U10546 ( .A1(n10792), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U10547 ( .A1(n8187), .A2(n8014), .ZN(n8016) );
  NAND2_X1 U10548 ( .A1(n10814), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8015) );
  NAND2_X1 U10549 ( .A1(n10828), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8017) );
  NAND2_X1 U10550 ( .A1(n10862), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8021) );
  INV_X1 U10551 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10861) );
  NAND2_X1 U10552 ( .A1(n10861), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8020) );
  NAND2_X1 U10553 ( .A1(n10878), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8023) );
  NAND2_X1 U10554 ( .A1(n10880), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8022) );
  INV_X1 U10555 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10901) );
  NAND2_X1 U10556 ( .A1(n10901), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8025) );
  INV_X1 U10557 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10899) );
  NAND2_X1 U10558 ( .A1(n10899), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8024) );
  NAND2_X1 U10559 ( .A1(n10906), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8027) );
  NAND2_X1 U10560 ( .A1(n10905), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8026) );
  AND2_X1 U10561 ( .A1(n8027), .A2(n8026), .ZN(n8253) );
  INV_X1 U10562 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10999) );
  NAND2_X1 U10563 ( .A1(n10999), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8029) );
  INV_X1 U10564 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10983) );
  NAND2_X1 U10565 ( .A1(n10983), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8028) );
  AND2_X1 U10566 ( .A1(n8029), .A2(n8028), .ZN(n8265) );
  AND2_X1 U10567 ( .A1(n11103), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U10568 ( .A1(n11022), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8033) );
  NAND2_X1 U10569 ( .A1(n11021), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8030) );
  NAND2_X1 U10570 ( .A1(n8033), .A2(n8030), .ZN(n8294) );
  AND2_X1 U10571 ( .A1(n11025), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n8031) );
  INV_X1 U10572 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10979) );
  NAND2_X1 U10573 ( .A1(n10979), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8035) );
  INV_X1 U10574 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10980) );
  NAND2_X1 U10575 ( .A1(n10980), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8034) );
  AND2_X1 U10576 ( .A1(n8035), .A2(n8034), .ZN(n8305) );
  NAND2_X1 U10577 ( .A1(n8306), .A2(n8305), .ZN(n8036) );
  NAND2_X1 U10578 ( .A1(n8036), .A2(n8035), .ZN(n8318) );
  INV_X1 U10579 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11124) );
  NAND2_X1 U10580 ( .A1(n11124), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8039) );
  INV_X1 U10581 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11069) );
  NAND2_X1 U10582 ( .A1(n11069), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8037) );
  NAND2_X1 U10583 ( .A1(n8039), .A2(n8037), .ZN(n8317) );
  INV_X1 U10584 ( .A(n8317), .ZN(n8038) );
  NAND2_X1 U10585 ( .A1(n8318), .A2(n8038), .ZN(n8040) );
  NAND2_X1 U10586 ( .A1(n8040), .A2(n8039), .ZN(n8331) );
  INV_X1 U10587 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11249) );
  NAND2_X1 U10588 ( .A1(n11249), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8042) );
  INV_X1 U10589 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11196) );
  NAND2_X1 U10590 ( .A1(n11196), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8041) );
  AND2_X1 U10591 ( .A1(n8042), .A2(n8041), .ZN(n8330) );
  INV_X1 U10592 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11482) );
  NAND2_X1 U10593 ( .A1(n11482), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8044) );
  INV_X1 U10594 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11434) );
  NAND2_X1 U10595 ( .A1(n11434), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8043) );
  AND2_X1 U10596 ( .A1(n8044), .A2(n8043), .ZN(n8343) );
  INV_X1 U10597 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11456) );
  NAND2_X1 U10598 ( .A1(n11456), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8046) );
  INV_X1 U10599 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11454) );
  NAND2_X1 U10600 ( .A1(n11454), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8045) );
  AND2_X1 U10601 ( .A1(n8046), .A2(n8045), .ZN(n8358) );
  INV_X1 U10602 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11824) );
  NAND2_X1 U10603 ( .A1(n11824), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8052) );
  INV_X1 U10604 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12979) );
  NAND2_X1 U10605 ( .A1(n12979), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8050) );
  NAND2_X1 U10606 ( .A1(n8052), .A2(n8050), .ZN(n8381) );
  INV_X1 U10607 ( .A(n8381), .ZN(n8051) );
  INV_X1 U10608 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11926) );
  XNOR2_X1 U10609 ( .A(n11926), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8392) );
  NAND2_X1 U10610 ( .A1(n11926), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8054) );
  XNOR2_X1 U10611 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8404) );
  INV_X1 U10612 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n12043) );
  INV_X1 U10613 ( .A(n8056), .ZN(n8055) );
  INV_X1 U10614 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12111) );
  INV_X1 U10615 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12244) );
  NAND2_X1 U10616 ( .A1(n12244), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8057) );
  INV_X1 U10617 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12242) );
  NAND2_X1 U10618 ( .A1(n12242), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8058) );
  INV_X1 U10619 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12547) );
  INV_X1 U10620 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n12544) );
  NAND2_X1 U10621 ( .A1(n12544), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8060) );
  NAND3_X1 U10622 ( .A1(n14072), .A2(n8061), .A3(P3_ADDR_REG_19__SCAN_IN), 
        .ZN(n8062) );
  XNOR2_X1 U10623 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8523) );
  INV_X1 U10624 ( .A(n8523), .ZN(n8097) );
  NAND2_X1 U10625 ( .A1(n12988), .A2(n8097), .ZN(n8095) );
  INV_X4 U10626 ( .A(n10786), .ZN(n8650) );
  NAND2_X1 U10627 ( .A1(n12983), .A2(SI_27_), .ZN(n8524) );
  NAND2_X1 U10628 ( .A1(n8524), .A2(n8523), .ZN(n8094) );
  INV_X1 U10629 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n8068) );
  INV_X1 U10630 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8070) );
  INV_X1 U10631 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n14485) );
  INV_X1 U10632 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8073) );
  INV_X1 U10633 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8075) );
  INV_X1 U10634 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8077) );
  INV_X1 U10635 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8079) );
  NAND2_X1 U10636 ( .A1(n8449), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8080) );
  INV_X1 U10637 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8082) );
  NAND2_X1 U10638 ( .A1(n8084), .A2(n8082), .ZN(n12944) );
  INV_X1 U10639 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12945) );
  INV_X1 U10640 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8083) );
  INV_X1 U10641 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n8090) );
  NAND2_X1 U10642 ( .A1(n12875), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U10643 ( .A1(n9327), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8088) );
  OAI211_X1 U10644 ( .C1(n12880), .C2(n8090), .A(n8089), .B(n8088), .ZN(n8091)
         );
  INV_X1 U10645 ( .A(n8091), .ZN(n8092) );
  MUX2_X1 U10646 ( .A(n8095), .B(n8094), .S(n13542), .Z(n8096) );
  NAND2_X1 U10647 ( .A1(n12988), .A2(n8523), .ZN(n8099) );
  NAND3_X1 U10648 ( .A1(n13542), .A2(n8097), .A3(n8524), .ZN(n8098) );
  OAI21_X1 U10649 ( .B1(n13542), .B2(n8099), .A(n8098), .ZN(n8100) );
  NAND2_X1 U10650 ( .A1(n9304), .A2(n8100), .ZN(n8104) );
  INV_X1 U10651 ( .A(n8524), .ZN(n8102) );
  OAI21_X1 U10652 ( .B1(n12988), .B2(n8102), .A(n13542), .ZN(n8101) );
  OAI21_X1 U10653 ( .B1(n8102), .B2(n13542), .A(n8101), .ZN(n8103) );
  INV_X1 U10654 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11400) );
  OR2_X1 U10655 ( .A1(n8138), .A2(n11400), .ZN(n8109) );
  NAND2_X1 U10656 ( .A1(n9328), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8108) );
  INV_X1 U10657 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8105) );
  OAI21_X1 U10658 ( .B1(n8112), .B2(n8122), .A(n8111), .ZN(n10841) );
  NAND2_X1 U10659 ( .A1(n12988), .A2(n10841), .ZN(n8115) );
  INV_X4 U10660 ( .A(n8471), .ZN(n8361) );
  NAND2_X1 U10661 ( .A1(n8361), .A2(n8113), .ZN(n8114) );
  NAND2_X1 U10662 ( .A1(n11181), .A2(n13732), .ZN(n13063) );
  NAND2_X1 U10663 ( .A1(n9328), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8121) );
  INV_X1 U10664 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11366) );
  INV_X1 U10665 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n8117) );
  OR2_X1 U10666 ( .A1(n8137), .A2(n11410), .ZN(n8118) );
  INV_X1 U10667 ( .A(n8122), .ZN(n8124) );
  INV_X1 U10668 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U10669 ( .A1(n9596), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U10670 ( .A1(n8124), .A2(n8123), .ZN(n8125) );
  MUX2_X1 U10671 ( .A(n8125), .B(SI_0_), .S(n10817), .Z(n13810) );
  MUX2_X1 U10672 ( .A(P3_IR_REG_0__SCAN_IN), .B(n13810), .S(n8471), .Z(n11413)
         );
  NAND2_X1 U10673 ( .A1(n6432), .A2(n11413), .ZN(n13720) );
  NAND2_X1 U10674 ( .A1(n11441), .A2(n11442), .ZN(n8136) );
  NAND2_X1 U10675 ( .A1(n8126), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8130) );
  INV_X1 U10676 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n11295) );
  OR2_X1 U10677 ( .A1(n8137), .A2(n15680), .ZN(n8128) );
  OR2_X1 U10678 ( .A1(n9321), .A2(n11451), .ZN(n8127) );
  NAND4_X2 U10679 ( .A1(n8127), .A2(n8128), .A3(n8129), .A4(n8130), .ZN(n13721) );
  OAI21_X1 U10680 ( .B1(n8133), .B2(n8132), .A(n8131), .ZN(n10838) );
  INV_X1 U10681 ( .A(SI_2_), .ZN(n10839) );
  NAND2_X1 U10682 ( .A1(n12983), .A2(n10839), .ZN(n8135) );
  NAND2_X1 U10683 ( .A1(n8361), .A2(n11122), .ZN(n8134) );
  NAND2_X1 U10684 ( .A1(n13721), .A2(n11448), .ZN(n13066) );
  NAND2_X1 U10685 ( .A1(n8136), .A2(n13060), .ZN(n11440) );
  NAND2_X1 U10686 ( .A1(n8179), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8143) );
  OR2_X1 U10687 ( .A1(n8138), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8142) );
  INV_X1 U10688 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8139) );
  OR2_X1 U10689 ( .A1(n8153), .A2(n8139), .ZN(n8141) );
  OR2_X1 U10690 ( .A1(n9321), .A2(n15723), .ZN(n8140) );
  NAND4_X2 U10691 ( .A1(n8143), .A2(n8142), .A3(n8141), .A4(n8140), .ZN(n13385) );
  OR2_X1 U10692 ( .A1(n8145), .A2(n8144), .ZN(n8146) );
  AND2_X1 U10693 ( .A1(n8147), .A2(n8146), .ZN(n10836) );
  NAND2_X1 U10694 ( .A1(n12988), .A2(n10836), .ZN(n8149) );
  NAND2_X1 U10695 ( .A1(n8361), .A2(n11344), .ZN(n8148) );
  OAI211_X1 U10696 ( .C1(n8110), .C2(SI_3_), .A(n8149), .B(n8148), .ZN(n11731)
         );
  NAND2_X1 U10697 ( .A1(n13385), .A2(n11731), .ZN(n13072) );
  NAND2_X1 U10698 ( .A1(n13073), .A2(n13072), .ZN(n13009) );
  NAND2_X1 U10699 ( .A1(n6974), .A2(n11448), .ZN(n11724) );
  NAND2_X1 U10700 ( .A1(n11440), .A2(n8150), .ZN(n11723) );
  INV_X1 U10701 ( .A(n11731), .ZN(n11548) );
  NAND2_X1 U10702 ( .A1(n13385), .A2(n11548), .ZN(n8151) );
  NAND2_X1 U10703 ( .A1(n11723), .A2(n8151), .ZN(n11698) );
  NAND2_X1 U10704 ( .A1(n8179), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8158) );
  OR2_X1 U10705 ( .A1(n9321), .A2(n15725), .ZN(n8157) );
  NAND2_X1 U10706 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8152) );
  AND2_X1 U10707 ( .A1(n8167), .A2(n8152), .ZN(n11696) );
  INV_X1 U10708 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8154) );
  OR2_X1 U10709 ( .A1(n8160), .A2(n8159), .ZN(n8161) );
  NAND2_X1 U10710 ( .A1(n8162), .A2(n8161), .ZN(n10866) );
  INV_X1 U10711 ( .A(SI_4_), .ZN(n8603) );
  NAND2_X1 U10712 ( .A1(n12983), .A2(n8603), .ZN(n8164) );
  NAND2_X1 U10713 ( .A1(n8361), .A2(n11219), .ZN(n8163) );
  OR2_X1 U10714 ( .A1(n11554), .A2(n15699), .ZN(n13077) );
  NAND2_X1 U10715 ( .A1(n11554), .A2(n15699), .ZN(n13076) );
  NAND2_X1 U10716 ( .A1(n11698), .A2(n11697), .ZN(n8166) );
  NAND2_X1 U10717 ( .A1(n11554), .A2(n11584), .ZN(n8165) );
  NAND2_X1 U10718 ( .A1(n9327), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8172) );
  OR2_X1 U10719 ( .A1(n9321), .A2(n15727), .ZN(n8171) );
  NAND2_X1 U10720 ( .A1(n8167), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8168) );
  AND2_X1 U10721 ( .A1(n8180), .A2(n8168), .ZN(n11744) );
  OR2_X1 U10722 ( .A1(n8138), .A2(n11744), .ZN(n8170) );
  OR2_X1 U10723 ( .A1(n12880), .A2(n14433), .ZN(n8169) );
  AND4_X2 U10724 ( .A1(n8172), .A2(n8171), .A3(n8170), .A4(n8169), .ZN(n12165)
         );
  INV_X2 U10725 ( .A(n12165), .ZN(n13384) );
  OR2_X1 U10726 ( .A1(n8174), .A2(n8173), .ZN(n8175) );
  AND2_X1 U10727 ( .A1(n8176), .A2(n8175), .ZN(n10834) );
  NAND2_X1 U10728 ( .A1(n12988), .A2(n10834), .ZN(n8178) );
  NAND2_X1 U10729 ( .A1(n8361), .A2(n11041), .ZN(n8177) );
  OAI211_X1 U10730 ( .C1(n8110), .C2(SI_5_), .A(n8178), .B(n8177), .ZN(n11779)
         );
  NAND2_X1 U10731 ( .A1(n13384), .A2(n11779), .ZN(n13083) );
  NAND2_X1 U10732 ( .A1(n13082), .A2(n13083), .ZN(n8476) );
  NAND2_X1 U10733 ( .A1(n8179), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8185) );
  OR2_X1 U10734 ( .A1(n9321), .A2(n15729), .ZN(n8184) );
  NAND2_X1 U10735 ( .A1(n8180), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8181) );
  AND2_X1 U10736 ( .A1(n8197), .A2(n8181), .ZN(n12171) );
  OR2_X1 U10737 ( .A1(n8138), .A2(n12171), .ZN(n8183) );
  OR2_X1 U10738 ( .A1(n8153), .A2(n15714), .ZN(n8182) );
  NAND4_X1 U10739 ( .A1(n8185), .A2(n8184), .A3(n8183), .A4(n8182), .ZN(n13383) );
  XNOR2_X1 U10740 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .ZN(n8186) );
  XNOR2_X1 U10741 ( .A(n8187), .B(n8186), .ZN(n10819) );
  NAND2_X1 U10742 ( .A1(n10819), .A2(n12988), .ZN(n8190) );
  AOI22_X1 U10743 ( .A1(n12983), .A2(SI_6_), .B1(n8361), .B2(n8188), .ZN(n8189) );
  NAND2_X1 U10744 ( .A1(n13383), .A2(n12168), .ZN(n12083) );
  NAND2_X1 U10745 ( .A1(n8476), .A2(n12083), .ZN(n8206) );
  NAND2_X1 U10746 ( .A1(n8192), .A2(n8191), .ZN(n8193) );
  NAND2_X1 U10747 ( .A1(n8194), .A2(n8193), .ZN(n10837) );
  NAND2_X1 U10748 ( .A1(n10837), .A2(n12988), .ZN(n8196) );
  INV_X1 U10749 ( .A(SI_7_), .ZN(n14401) );
  AOI22_X1 U10750 ( .A1(n12983), .A2(n14401), .B1(n8361), .B2(n11352), .ZN(
        n8195) );
  NAND2_X1 U10751 ( .A1(n8196), .A2(n8195), .ZN(n15716) );
  NAND2_X1 U10752 ( .A1(n8179), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8203) );
  OR2_X1 U10753 ( .A1(n9321), .A2(n15732), .ZN(n8202) );
  NAND2_X1 U10754 ( .A1(n8197), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8198) );
  AND2_X1 U10755 ( .A1(n8226), .A2(n8198), .ZN(n12363) );
  OR2_X1 U10756 ( .A1(n8138), .A2(n12363), .ZN(n8201) );
  INV_X1 U10757 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n8199) );
  OR2_X1 U10758 ( .A1(n8153), .A2(n8199), .ZN(n8200) );
  NAND4_X1 U10759 ( .A1(n8203), .A2(n8202), .A3(n8201), .A4(n8200), .ZN(n13382) );
  XNOR2_X1 U10760 ( .A(n15716), .B(n13382), .ZN(n12085) );
  NAND2_X1 U10761 ( .A1(n13383), .A2(n8204), .ZN(n13089) );
  NAND2_X1 U10762 ( .A1(n13090), .A2(n13089), .ZN(n11990) );
  NAND2_X1 U10763 ( .A1(n12165), .A2(n11779), .ZN(n11991) );
  NAND2_X1 U10764 ( .A1(n11990), .A2(n11991), .ZN(n11992) );
  NAND2_X1 U10765 ( .A1(n11992), .A2(n12083), .ZN(n8205) );
  OAI211_X1 U10766 ( .C1(n11740), .C2(n8206), .A(n12085), .B(n8205), .ZN(n8208) );
  INV_X1 U10767 ( .A(n15716), .ZN(n12360) );
  NAND2_X1 U10768 ( .A1(n12360), .A2(n13382), .ZN(n8207) );
  NAND2_X1 U10769 ( .A1(n8208), .A2(n8207), .ZN(n12013) );
  OR2_X1 U10770 ( .A1(n8211), .A2(n8210), .ZN(n8212) );
  NAND2_X1 U10771 ( .A1(n8209), .A2(n8212), .ZN(n10847) );
  NAND2_X1 U10772 ( .A1(n10847), .A2(n12985), .ZN(n8214) );
  INV_X1 U10773 ( .A(SI_9_), .ZN(n10846) );
  AOI22_X1 U10774 ( .A1(n11849), .A2(n8361), .B1(n12983), .B2(n10846), .ZN(
        n8213) );
  NAND2_X1 U10775 ( .A1(n8214), .A2(n8213), .ZN(n12534) );
  NAND2_X1 U10776 ( .A1(n8179), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8220) );
  OR2_X1 U10777 ( .A1(n9321), .A2(n12297), .ZN(n8219) );
  NAND2_X1 U10778 ( .A1(n6490), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8215) );
  AND2_X1 U10779 ( .A1(n8241), .A2(n8215), .ZN(n12226) );
  OR2_X1 U10780 ( .A1(n8138), .A2(n12226), .ZN(n8218) );
  INV_X1 U10781 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n8216) );
  OR2_X1 U10782 ( .A1(n8153), .A2(n8216), .ZN(n8217) );
  NAND4_X1 U10783 ( .A1(n8220), .A2(n8219), .A3(n8218), .A4(n8217), .ZN(n13380) );
  OR2_X1 U10784 ( .A1(n12534), .A2(n12702), .ZN(n12075) );
  INV_X1 U10785 ( .A(n8221), .ZN(n8222) );
  XNOR2_X1 U10786 ( .A(n8223), .B(n8222), .ZN(n10823) );
  NAND2_X1 U10787 ( .A1(n10823), .A2(n12985), .ZN(n8225) );
  AOI22_X1 U10788 ( .A1(n12983), .A2(SI_8_), .B1(n11529), .B2(n8361), .ZN(
        n8224) );
  NAND2_X1 U10789 ( .A1(n8225), .A2(n8224), .ZN(n12351) );
  NAND2_X1 U10790 ( .A1(n12875), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8232) );
  OR2_X1 U10791 ( .A1(n12880), .A2(n12116), .ZN(n8231) );
  NAND2_X1 U10792 ( .A1(n8226), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8227) );
  AND2_X1 U10793 ( .A1(n6490), .A2(n8227), .ZN(n12349) );
  OR2_X1 U10794 ( .A1(n8138), .A2(n12349), .ZN(n8230) );
  INV_X1 U10795 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8228) );
  OR2_X1 U10796 ( .A1(n8153), .A2(n8228), .ZN(n8229) );
  NAND4_X1 U10797 ( .A1(n8232), .A2(n8231), .A3(n8230), .A4(n8229), .ZN(n13381) );
  OR2_X1 U10798 ( .A1(n12351), .A2(n12537), .ZN(n13099) );
  NAND2_X1 U10799 ( .A1(n12351), .A2(n12537), .ZN(n13100) );
  NAND2_X1 U10800 ( .A1(n12075), .A2(n13015), .ZN(n8249) );
  OR2_X1 U10801 ( .A1(n12534), .A2(n13380), .ZN(n13104) );
  NAND2_X1 U10802 ( .A1(n12534), .A2(n13380), .ZN(n13105) );
  NAND2_X1 U10803 ( .A1(n13104), .A2(n13105), .ZN(n13013) );
  OR2_X1 U10804 ( .A1(n12351), .A2(n13381), .ZN(n12073) );
  NAND2_X1 U10805 ( .A1(n13013), .A2(n12073), .ZN(n8233) );
  NAND2_X1 U10806 ( .A1(n8233), .A2(n12075), .ZN(n8247) );
  OR2_X1 U10807 ( .A1(n8235), .A2(n8234), .ZN(n8236) );
  NAND2_X1 U10808 ( .A1(n8237), .A2(n8236), .ZN(n10844) );
  NAND2_X1 U10809 ( .A1(n10844), .A2(n12985), .ZN(n8239) );
  INV_X1 U10810 ( .A(SI_10_), .ZN(n14402) );
  AOI22_X1 U10811 ( .A1(n12983), .A2(n14402), .B1(n8361), .B2(n10845), .ZN(
        n8238) );
  NAND2_X1 U10812 ( .A1(n8179), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8246) );
  INV_X1 U10813 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n8240) );
  OR2_X1 U10814 ( .A1(n9321), .A2(n8240), .ZN(n8245) );
  NAND2_X1 U10815 ( .A1(n8241), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8242) );
  AND2_X1 U10816 ( .A1(n8258), .A2(n8242), .ZN(n12703) );
  OR2_X1 U10817 ( .A1(n8138), .A2(n12703), .ZN(n8244) );
  INV_X1 U10818 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n14469) );
  OR2_X1 U10819 ( .A1(n8153), .A2(n14469), .ZN(n8243) );
  NAND4_X1 U10820 ( .A1(n8246), .A2(n8245), .A3(n8244), .A4(n8243), .ZN(n13379) );
  XNOR2_X1 U10821 ( .A(n13110), .B(n13379), .ZN(n12076) );
  INV_X1 U10822 ( .A(n13379), .ZN(n13109) );
  OR2_X1 U10823 ( .A1(n13110), .A2(n13109), .ZN(n8250) );
  NAND2_X1 U10824 ( .A1(n8251), .A2(n8250), .ZN(n12276) );
  OR2_X1 U10825 ( .A1(n8254), .A2(n8253), .ZN(n8255) );
  NAND2_X1 U10826 ( .A1(n8252), .A2(n8255), .ZN(n10849) );
  NAND2_X1 U10827 ( .A1(n10849), .A2(n12985), .ZN(n8257) );
  INV_X1 U10828 ( .A(SI_11_), .ZN(n10848) );
  AOI22_X1 U10829 ( .A1(n12983), .A2(n10848), .B1(n8361), .B2(n10850), .ZN(
        n8256) );
  NAND2_X1 U10830 ( .A1(n8257), .A2(n8256), .ZN(n12855) );
  NAND2_X1 U10831 ( .A1(n8258), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U10832 ( .A1(n8271), .A2(n8259), .ZN(n12860) );
  NAND2_X1 U10833 ( .A1(n9318), .A2(n12860), .ZN(n8263) );
  OR2_X1 U10834 ( .A1(n12880), .A2(n12662), .ZN(n8262) );
  OR2_X1 U10835 ( .A1(n9321), .A2(n12656), .ZN(n8261) );
  INV_X1 U10836 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n12291) );
  OR2_X1 U10837 ( .A1(n8153), .A2(n12291), .ZN(n8260) );
  NAND2_X1 U10838 ( .A1(n12855), .A2(n13275), .ZN(n8264) );
  OR2_X1 U10839 ( .A1(n8266), .A2(n8265), .ZN(n8267) );
  NAND2_X1 U10840 ( .A1(n8268), .A2(n8267), .ZN(n10873) );
  AOI22_X1 U10841 ( .A1(n12983), .A2(SI_12_), .B1(n8361), .B2(n13412), .ZN(
        n8269) );
  NAND2_X1 U10842 ( .A1(n8271), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8272) );
  NAND2_X1 U10843 ( .A1(n8286), .A2(n8272), .ZN(n13277) );
  NAND2_X1 U10844 ( .A1(n9318), .A2(n13277), .ZN(n8278) );
  OR2_X1 U10845 ( .A1(n12880), .A2(n12284), .ZN(n8277) );
  OR2_X1 U10846 ( .A1(n9321), .A2(n8273), .ZN(n8276) );
  INV_X1 U10847 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n8274) );
  OR2_X1 U10848 ( .A1(n8153), .A2(n8274), .ZN(n8275) );
  NAND2_X1 U10849 ( .A1(n13278), .A2(n13270), .ZN(n13118) );
  INV_X1 U10850 ( .A(n13270), .ZN(n13377) );
  NAND2_X1 U10851 ( .A1(n8280), .A2(n11103), .ZN(n8293) );
  OR2_X1 U10852 ( .A1(n8280), .A2(n11103), .ZN(n8281) );
  NAND2_X1 U10853 ( .A1(n8293), .A2(n8281), .ZN(n8282) );
  NAND2_X1 U10854 ( .A1(n8282), .A2(n11025), .ZN(n8283) );
  NAND2_X1 U10855 ( .A1(n8295), .A2(n8283), .ZN(n10910) );
  NAND2_X1 U10856 ( .A1(n10910), .A2(n12985), .ZN(n8285) );
  INV_X1 U10857 ( .A(SI_13_), .ZN(n10909) );
  AOI22_X1 U10858 ( .A1(n12983), .A2(n10909), .B1(n13430), .B2(n8361), .ZN(
        n8284) );
  NAND2_X1 U10859 ( .A1(n8286), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8287) );
  NAND2_X1 U10860 ( .A1(n8300), .A2(n8287), .ZN(n12793) );
  NAND2_X1 U10861 ( .A1(n12793), .A2(n9318), .ZN(n8291) );
  NAND2_X1 U10862 ( .A1(n8179), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U10863 ( .A1(n12875), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8289) );
  NAND2_X1 U10864 ( .A1(n9327), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8288) );
  NAND4_X1 U10865 ( .A1(n8291), .A2(n8290), .A3(n8289), .A4(n8288), .ZN(n13376) );
  NAND2_X1 U10866 ( .A1(n12790), .A2(n13376), .ZN(n13122) );
  NAND2_X1 U10867 ( .A1(n13121), .A2(n13122), .ZN(n13126) );
  NAND2_X1 U10868 ( .A1(n12393), .A2(n13126), .ZN(n12392) );
  INV_X1 U10869 ( .A(n13376), .ZN(n13231) );
  OR2_X1 U10870 ( .A1(n12790), .A2(n13231), .ZN(n8292) );
  NAND2_X1 U10871 ( .A1(n12392), .A2(n8292), .ZN(n12616) );
  NAND3_X1 U10872 ( .A1(n8295), .A2(n8294), .A3(n8293), .ZN(n8297) );
  NAND2_X1 U10873 ( .A1(n8297), .A2(n8296), .ZN(n10976) );
  NAND2_X1 U10874 ( .A1(n10976), .A2(n12985), .ZN(n8299) );
  INV_X1 U10875 ( .A(SI_14_), .ZN(n10975) );
  AOI22_X1 U10876 ( .A1(n10977), .A2(n8361), .B1(n12983), .B2(n10975), .ZN(
        n8298) );
  INV_X1 U10877 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12620) );
  NAND2_X1 U10878 ( .A1(n8300), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U10879 ( .A1(n8309), .A2(n8301), .ZN(n13233) );
  NAND2_X1 U10880 ( .A1(n13233), .A2(n9318), .ZN(n8303) );
  AOI22_X1 U10881 ( .A1(n8179), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n12875), 
        .B2(P3_REG1_REG_14__SCAN_IN), .ZN(n8302) );
  OAI211_X1 U10882 ( .C1(n8153), .C2(n12620), .A(n8303), .B(n8302), .ZN(n13375) );
  OR2_X1 U10883 ( .A1(n13236), .A2(n13375), .ZN(n13127) );
  NAND2_X1 U10884 ( .A1(n13236), .A2(n13375), .ZN(n13128) );
  NAND2_X1 U10885 ( .A1(n13127), .A2(n13128), .ZN(n12615) );
  INV_X1 U10886 ( .A(n13375), .ZN(n13360) );
  OR2_X1 U10887 ( .A1(n13236), .A2(n13360), .ZN(n8304) );
  XNOR2_X1 U10888 ( .A(n8306), .B(n8305), .ZN(n10974) );
  NAND2_X1 U10889 ( .A1(n10974), .A2(n12985), .ZN(n8308) );
  INV_X1 U10890 ( .A(SI_15_), .ZN(n10973) );
  AOI22_X1 U10891 ( .A1(n13449), .A2(n8361), .B1(n12983), .B2(n10973), .ZN(
        n8307) );
  NAND2_X1 U10892 ( .A1(n8309), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8310) );
  NAND2_X1 U10893 ( .A1(n8321), .A2(n8310), .ZN(n13363) );
  NAND2_X1 U10894 ( .A1(n13363), .A2(n9318), .ZN(n8313) );
  AOI22_X1 U10895 ( .A1(n12875), .A2(P3_REG1_REG_15__SCAN_IN), .B1(n9327), 
        .B2(P3_REG0_REG_15__SCAN_IN), .ZN(n8312) );
  NAND2_X1 U10896 ( .A1(n8179), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8311) );
  NAND2_X1 U10897 ( .A1(n13366), .A2(n13293), .ZN(n8314) );
  NAND2_X1 U10898 ( .A1(n12796), .A2(n8314), .ZN(n8316) );
  OR2_X1 U10899 ( .A1(n13366), .A2(n13293), .ZN(n8315) );
  XNOR2_X1 U10900 ( .A(n8318), .B(n8317), .ZN(n11016) );
  NAND2_X1 U10901 ( .A1(n11016), .A2(n12985), .ZN(n8320) );
  AOI22_X1 U10902 ( .A1(n12983), .A2(SI_16_), .B1(n8361), .B2(n11017), .ZN(
        n8319) );
  NAND2_X1 U10903 ( .A1(n8321), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U10904 ( .A1(n8335), .A2(n8322), .ZN(n13295) );
  NAND2_X1 U10905 ( .A1(n13295), .A2(n9318), .ZN(n8327) );
  INV_X1 U10906 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n14482) );
  NAND2_X1 U10907 ( .A1(n12875), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8324) );
  NAND2_X1 U10908 ( .A1(n8179), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8323) );
  OAI211_X1 U10909 ( .C1(n8153), .C2(n14482), .A(n8324), .B(n8323), .ZN(n8325)
         );
  INV_X1 U10910 ( .A(n8325), .ZN(n8326) );
  OR2_X1 U10911 ( .A1(n13712), .A2(n13654), .ZN(n8328) );
  OR2_X1 U10912 ( .A1(n8331), .A2(n8330), .ZN(n8332) );
  NAND2_X1 U10913 ( .A1(n8329), .A2(n8332), .ZN(n11101) );
  NAND2_X1 U10914 ( .A1(n11101), .A2(n12985), .ZN(n8334) );
  INV_X1 U10915 ( .A(SI_17_), .ZN(n14461) );
  AOI22_X1 U10916 ( .A1(n12983), .A2(n14461), .B1(n13485), .B2(n8361), .ZN(
        n8333) );
  NAND2_X1 U10917 ( .A1(n8335), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8336) );
  NAND2_X1 U10918 ( .A1(n8349), .A2(n8336), .ZN(n13658) );
  NAND2_X1 U10919 ( .A1(n13658), .A2(n9318), .ZN(n8341) );
  NAND2_X1 U10920 ( .A1(n9327), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8338) );
  NAND2_X1 U10921 ( .A1(n12875), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8337) );
  OAI211_X1 U10922 ( .C1(n12880), .C2(n13657), .A(n8338), .B(n8337), .ZN(n8339) );
  INV_X1 U10923 ( .A(n8339), .ZN(n8340) );
  NAND2_X1 U10924 ( .A1(n8341), .A2(n8340), .ZN(n13373) );
  NAND2_X1 U10925 ( .A1(n13789), .A2(n13373), .ZN(n13040) );
  INV_X1 U10926 ( .A(n13373), .ZN(n13640) );
  OR2_X1 U10927 ( .A1(n8344), .A2(n8343), .ZN(n8345) );
  NAND2_X1 U10928 ( .A1(n8342), .A2(n8345), .ZN(n11221) );
  AOI22_X1 U10929 ( .A1(n12983), .A2(SI_18_), .B1(n8361), .B2(n6599), .ZN(
        n8347) );
  NAND2_X1 U10930 ( .A1(n8349), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8350) );
  NAND2_X1 U10931 ( .A1(n8364), .A2(n8350), .ZN(n13644) );
  NAND2_X1 U10932 ( .A1(n13644), .A2(n9318), .ZN(n8355) );
  NAND2_X1 U10933 ( .A1(n9327), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8352) );
  NAND2_X1 U10934 ( .A1(n12875), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8351) );
  OAI211_X1 U10935 ( .C1(n12880), .C2(n13647), .A(n8352), .B(n8351), .ZN(n8353) );
  INV_X1 U10936 ( .A(n8353), .ZN(n8354) );
  NAND2_X1 U10937 ( .A1(n13702), .A2(n13249), .ZN(n13042) );
  OR2_X1 U10938 ( .A1(n13702), .A2(n13655), .ZN(n8356) );
  OR2_X1 U10939 ( .A1(n8359), .A2(n8358), .ZN(n8360) );
  NAND2_X1 U10940 ( .A1(n8357), .A2(n8360), .ZN(n11435) );
  AOI22_X1 U10941 ( .A1(n12983), .A2(SI_19_), .B1(n11284), .B2(n8361), .ZN(
        n8362) );
  NAND2_X1 U10942 ( .A1(n8364), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8365) );
  NAND2_X1 U10943 ( .A1(n8374), .A2(n8365), .ZN(n13626) );
  NAND2_X1 U10944 ( .A1(n13626), .A2(n9318), .ZN(n8370) );
  NAND2_X1 U10945 ( .A1(n9327), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8367) );
  NAND2_X1 U10946 ( .A1(n12875), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8366) );
  OAI211_X1 U10947 ( .C1(n12880), .C2(n13625), .A(n8367), .B(n8366), .ZN(n8368) );
  INV_X1 U10948 ( .A(n8368), .ZN(n8369) );
  NAND2_X1 U10949 ( .A1(n8370), .A2(n8369), .ZN(n13615) );
  NOR2_X1 U10950 ( .A1(n13775), .A2(n13615), .ZN(n13006) );
  NAND2_X1 U10951 ( .A1(n13775), .A2(n13615), .ZN(n13004) );
  INV_X1 U10952 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11776) );
  XNOR2_X1 U10953 ( .A(n8371), .B(n11776), .ZN(n11803) );
  NAND2_X1 U10954 ( .A1(n11803), .A2(n12985), .ZN(n8373) );
  NAND2_X1 U10955 ( .A1(n12983), .A2(SI_20_), .ZN(n8372) );
  NAND2_X1 U10956 ( .A1(n8374), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8375) );
  NAND2_X1 U10957 ( .A1(n8385), .A2(n8375), .ZN(n13617) );
  NAND2_X1 U10958 ( .A1(n13617), .A2(n9318), .ZN(n8380) );
  INV_X1 U10959 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13616) );
  NAND2_X1 U10960 ( .A1(n9327), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8377) );
  NAND2_X1 U10961 ( .A1(n12875), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8376) );
  OAI211_X1 U10962 ( .C1(n12880), .C2(n13616), .A(n8377), .B(n8376), .ZN(n8378) );
  INV_X1 U10963 ( .A(n8378), .ZN(n8379) );
  NAND2_X1 U10964 ( .A1(n13768), .A2(n13251), .ZN(n13035) );
  XNOR2_X1 U10965 ( .A(n8382), .B(n8381), .ZN(n11897) );
  NAND2_X1 U10966 ( .A1(n11897), .A2(n12985), .ZN(n8384) );
  NAND2_X1 U10967 ( .A1(n12983), .A2(SI_21_), .ZN(n8383) );
  NAND2_X1 U10968 ( .A1(n8385), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U10969 ( .A1(n8396), .A2(n8386), .ZN(n13607) );
  NAND2_X1 U10970 ( .A1(n13607), .A2(n9318), .ZN(n8391) );
  INV_X1 U10971 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13606) );
  NAND2_X1 U10972 ( .A1(n12875), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U10973 ( .A1(n9327), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8387) );
  OAI211_X1 U10974 ( .C1(n13606), .C2(n12880), .A(n8388), .B(n8387), .ZN(n8389) );
  INV_X1 U10975 ( .A(n8389), .ZN(n8390) );
  NAND2_X1 U10976 ( .A1(n8391), .A2(n8390), .ZN(n13613) );
  AND2_X1 U10977 ( .A1(n13762), .A2(n13613), .ZN(n13003) );
  OR2_X1 U10978 ( .A1(n13762), .A2(n13613), .ZN(n13002) );
  XNOR2_X1 U10979 ( .A(n8393), .B(n8392), .ZN(n11966) );
  NAND2_X1 U10980 ( .A1(n11966), .A2(n12985), .ZN(n8395) );
  NAND2_X1 U10981 ( .A1(n12983), .A2(SI_22_), .ZN(n8394) );
  NAND2_X1 U10982 ( .A1(n8396), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U10983 ( .A1(n8408), .A2(n8397), .ZN(n13598) );
  NAND2_X1 U10984 ( .A1(n13598), .A2(n9318), .ZN(n8402) );
  INV_X1 U10985 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n14453) );
  NAND2_X1 U10986 ( .A1(n12875), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8399) );
  NAND2_X1 U10987 ( .A1(n8179), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8398) );
  OAI211_X1 U10988 ( .C1(n14453), .C2(n8153), .A(n8399), .B(n8398), .ZN(n8400)
         );
  INV_X1 U10989 ( .A(n8400), .ZN(n8401) );
  NOR2_X1 U10990 ( .A1(n13756), .A2(n13604), .ZN(n8403) );
  XNOR2_X1 U10991 ( .A(n8405), .B(n8404), .ZN(n12270) );
  NAND2_X1 U10992 ( .A1(n12270), .A2(n12985), .ZN(n8407) );
  NAND2_X1 U10993 ( .A1(n12983), .A2(SI_23_), .ZN(n8406) );
  NAND2_X1 U10994 ( .A1(n8408), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U10995 ( .A1(n8421), .A2(n8409), .ZN(n13586) );
  NAND2_X1 U10996 ( .A1(n13586), .A2(n9318), .ZN(n8415) );
  INV_X1 U10997 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n8412) );
  NAND2_X1 U10998 ( .A1(n12875), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8411) );
  NAND2_X1 U10999 ( .A1(n9327), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8410) );
  OAI211_X1 U11000 ( .C1(n12880), .C2(n8412), .A(n8411), .B(n8410), .ZN(n8413)
         );
  INV_X1 U11001 ( .A(n8413), .ZN(n8414) );
  NAND2_X1 U11002 ( .A1(n13243), .A2(n13569), .ZN(n8416) );
  NAND2_X1 U11003 ( .A1(n13243), .A2(n13595), .ZN(n8417) );
  INV_X1 U11004 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12110) );
  XNOR2_X1 U11005 ( .A(n8418), .B(n12110), .ZN(n12976) );
  NAND2_X1 U11006 ( .A1(n12976), .A2(n12985), .ZN(n8420) );
  NAND2_X1 U11007 ( .A1(n12983), .A2(SI_24_), .ZN(n8419) );
  NAND2_X1 U11008 ( .A1(n8421), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8422) );
  NAND2_X1 U11009 ( .A1(n8434), .A2(n8422), .ZN(n13574) );
  NAND2_X1 U11010 ( .A1(n13574), .A2(n9318), .ZN(n8428) );
  INV_X1 U11011 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U11012 ( .A1(n9327), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8424) );
  NAND2_X1 U11013 ( .A1(n12875), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8423) );
  OAI211_X1 U11014 ( .C1(n12880), .C2(n8425), .A(n8424), .B(n8423), .ZN(n8426)
         );
  INV_X1 U11015 ( .A(n8426), .ZN(n8427) );
  AND2_X1 U11016 ( .A1(n8488), .A2(n13582), .ZN(n8429) );
  XNOR2_X1 U11017 ( .A(n12244), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8430) );
  XNOR2_X1 U11018 ( .A(n8431), .B(n8430), .ZN(n13804) );
  NAND2_X1 U11019 ( .A1(n13804), .A2(n12985), .ZN(n8433) );
  NAND2_X1 U11020 ( .A1(n12983), .A2(SI_25_), .ZN(n8432) );
  NAND2_X1 U11021 ( .A1(n8434), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8435) );
  NAND2_X1 U11022 ( .A1(n8447), .A2(n8435), .ZN(n13559) );
  NAND2_X1 U11023 ( .A1(n13559), .A2(n9318), .ZN(n8441) );
  INV_X1 U11024 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n8438) );
  NAND2_X1 U11025 ( .A1(n9327), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8437) );
  NAND2_X1 U11026 ( .A1(n12875), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8436) );
  OAI211_X1 U11027 ( .C1(n12880), .C2(n8438), .A(n8437), .B(n8436), .ZN(n8439)
         );
  INV_X1 U11028 ( .A(n8439), .ZN(n8440) );
  NAND2_X1 U11029 ( .A1(n13675), .A2(n13570), .ZN(n13160) );
  NAND2_X1 U11030 ( .A1(n13675), .A2(n13541), .ZN(n8442) );
  XNOR2_X1 U11031 ( .A(n12547), .B(P1_DATAO_REG_26__SCAN_IN), .ZN(n8443) );
  XNOR2_X1 U11032 ( .A(n8444), .B(n8443), .ZN(n12956) );
  NAND2_X1 U11033 ( .A1(n12956), .A2(n12985), .ZN(n8446) );
  NAND2_X1 U11034 ( .A1(n12983), .A2(SI_26_), .ZN(n8445) );
  NAND2_X1 U11035 ( .A1(n8447), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8448) );
  NAND2_X1 U11036 ( .A1(n8449), .A2(n8448), .ZN(n13546) );
  NAND2_X1 U11037 ( .A1(n13546), .A2(n9318), .ZN(n8455) );
  INV_X1 U11038 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U11039 ( .A1(n12875), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8451) );
  NAND2_X1 U11040 ( .A1(n9327), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8450) );
  OAI211_X1 U11041 ( .C1(n8452), .C2(n12880), .A(n8451), .B(n8450), .ZN(n8453)
         );
  INV_X1 U11042 ( .A(n8453), .ZN(n8454) );
  OR2_X1 U11043 ( .A1(n13671), .A2(n13371), .ZN(n8456) );
  NAND2_X1 U11044 ( .A1(n13671), .A2(n13371), .ZN(n8457) );
  INV_X1 U11045 ( .A(n9302), .ZN(n8458) );
  AOI21_X1 U11046 ( .B1(n13165), .B2(n8459), .A(n8458), .ZN(n8474) );
  NAND2_X1 U11047 ( .A1(n13191), .A2(n11284), .ZN(n9551) );
  INV_X1 U11048 ( .A(n8460), .ZN(n8461) );
  NAND2_X1 U11049 ( .A1(n8461), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8463) );
  NAND2_X1 U11050 ( .A1(n13054), .A2(n9552), .ZN(n13000) );
  INV_X1 U11051 ( .A(n13728), .ZN(n13638) );
  NAND2_X1 U11052 ( .A1(n8464), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8465) );
  INV_X1 U11053 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n8468) );
  NAND2_X1 U11054 ( .A1(n12875), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U11055 ( .A1(n9327), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8466) );
  OAI211_X1 U11056 ( .C1(n8468), .C2(n12880), .A(n8467), .B(n8466), .ZN(n8469)
         );
  INV_X1 U11057 ( .A(n9308), .ZN(n13370) );
  NAND2_X1 U11058 ( .A1(n8471), .A2(n8470), .ZN(n11281) );
  INV_X1 U11059 ( .A(n11281), .ZN(n8472) );
  AOI22_X1 U11060 ( .A1(n13370), .A2(n13722), .B1(n13724), .B2(n13371), .ZN(
        n8473) );
  INV_X1 U11061 ( .A(n11413), .ZN(n11390) );
  NAND2_X1 U11062 ( .A1(n11288), .A2(n13064), .ZN(n11437) );
  NAND2_X1 U11063 ( .A1(n11439), .A2(n13065), .ZN(n11721) );
  INV_X1 U11064 ( .A(n13009), .ZN(n11722) );
  NAND2_X1 U11065 ( .A1(n11721), .A2(n11722), .ZN(n8475) );
  NAND2_X1 U11066 ( .A1(n11737), .A2(n13079), .ZN(n11739) );
  INV_X1 U11067 ( .A(n11990), .ZN(n13011) );
  NAND2_X1 U11068 ( .A1(n8477), .A2(n13090), .ZN(n12088) );
  INV_X1 U11069 ( .A(n12085), .ZN(n13092) );
  NAND2_X1 U11070 ( .A1(n12088), .A2(n13092), .ZN(n12087) );
  OR2_X1 U11071 ( .A1(n13382), .A2(n15716), .ZN(n13094) );
  AND2_X1 U11072 ( .A1(n13100), .A2(n13094), .ZN(n8478) );
  INV_X1 U11073 ( .A(n12070), .ZN(n8480) );
  INV_X1 U11074 ( .A(n13275), .ZN(n13378) );
  NAND2_X1 U11075 ( .A1(n12855), .A2(n13378), .ZN(n13051) );
  NAND2_X1 U11076 ( .A1(n13110), .A2(n13379), .ZN(n12201) );
  INV_X1 U11077 ( .A(n12855), .ZN(n12280) );
  INV_X1 U11078 ( .A(n13118), .ZN(n8481) );
  AOI21_X1 U11079 ( .B1(n13018), .B2(n13049), .A(n8481), .ZN(n8482) );
  INV_X1 U11080 ( .A(n13128), .ZN(n8483) );
  NAND2_X1 U11081 ( .A1(n13366), .A2(n13374), .ZN(n13131) );
  XNOR2_X1 U11082 ( .A(n13712), .B(n13654), .ZN(n13021) );
  INV_X1 U11083 ( .A(n13654), .ZN(n13303) );
  AND2_X1 U11084 ( .A1(n13712), .A2(n13303), .ZN(n13134) );
  NAND2_X1 U11085 ( .A1(n13040), .A2(n13134), .ZN(n8484) );
  NAND2_X1 U11086 ( .A1(n8484), .A2(n13037), .ZN(n8485) );
  NOR2_X1 U11087 ( .A1(n7207), .A2(n8485), .ZN(n8486) );
  INV_X1 U11088 ( .A(n13615), .ZN(n13642) );
  NOR2_X1 U11089 ( .A1(n13775), .A2(n13642), .ZN(n13046) );
  NAND2_X1 U11090 ( .A1(n13775), .A2(n13642), .ZN(n13038) );
  NAND2_X1 U11091 ( .A1(n13762), .A2(n13320), .ZN(n13033) );
  OR2_X1 U11092 ( .A1(n8488), .A2(n13551), .ZN(n13152) );
  NAND2_X1 U11093 ( .A1(n8488), .A2(n13551), .ZN(n13150) );
  NAND2_X1 U11094 ( .A1(n13152), .A2(n13150), .ZN(n13565) );
  NAND2_X1 U11095 ( .A1(n13568), .A2(n8489), .ZN(n13567) );
  NAND2_X1 U11096 ( .A1(n13558), .A2(n13557), .ZN(n13556) );
  OAI21_X1 U11097 ( .B1(n11964), .B2(n9552), .A(n11284), .ZN(n8490) );
  NAND2_X1 U11098 ( .A1(n8490), .A2(n13059), .ZN(n8492) );
  OAI21_X1 U11099 ( .B1(n13054), .B2(n9552), .A(n11964), .ZN(n8491) );
  NAND2_X1 U11100 ( .A1(n8492), .A2(n8491), .ZN(n11182) );
  NAND2_X1 U11101 ( .A1(n11804), .A2(n13031), .ZN(n13183) );
  INV_X1 U11102 ( .A(n13183), .ZN(n9550) );
  NAND2_X1 U11103 ( .A1(n11964), .A2(n13059), .ZN(n15715) );
  NAND3_X1 U11104 ( .A1(n11182), .A2(n9550), .A3(n15715), .ZN(n8494) );
  NOR2_X1 U11105 ( .A1(n11804), .A2(n11284), .ZN(n8493) );
  NAND2_X1 U11106 ( .A1(n13191), .A2(n8493), .ZN(n8519) );
  NAND2_X1 U11107 ( .A1(n8494), .A2(n8519), .ZN(n13718) );
  NAND2_X1 U11108 ( .A1(n11804), .A2(n11284), .ZN(n15683) );
  INV_X1 U11109 ( .A(n15683), .ZN(n15674) );
  AND2_X1 U11110 ( .A1(n11964), .A2(n15674), .ZN(n15720) );
  INV_X1 U11111 ( .A(n12959), .ZN(n8498) );
  XNOR2_X1 U11112 ( .A(P3_IR_REG_23__SCAN_IN), .B(P3_IR_REG_24__SCAN_IN), .ZN(
        n8495) );
  XNOR2_X1 U11113 ( .A(n8495), .B(P3_B_REG_SCAN_IN), .ZN(n8496) );
  NAND2_X1 U11114 ( .A1(n13809), .A2(n8496), .ZN(n8497) );
  NAND2_X1 U11115 ( .A1(n8498), .A2(n8497), .ZN(n10859) );
  NOR2_X1 U11116 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n8502) );
  NOR4_X1 U11117 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8501) );
  NOR4_X1 U11118 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8500) );
  NOR4_X1 U11119 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8499) );
  NAND4_X1 U11120 ( .A1(n8502), .A2(n8501), .A3(n8500), .A4(n8499), .ZN(n8508)
         );
  NOR4_X1 U11121 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8506) );
  NOR4_X1 U11122 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8505) );
  NOR4_X1 U11123 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8504) );
  NOR4_X1 U11124 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8503) );
  NAND4_X1 U11125 ( .A1(n8506), .A2(n8505), .A3(n8504), .A4(n8503), .ZN(n8507)
         );
  NOR2_X1 U11126 ( .A1(n8508), .A2(n8507), .ZN(n8509) );
  NOR2_X1 U11127 ( .A1(n10859), .A2(n8509), .ZN(n9555) );
  NOR2_X1 U11128 ( .A1(n9557), .A2(n9555), .ZN(n8515) );
  NAND2_X1 U11129 ( .A1(n8510), .A2(n12959), .ZN(n8512) );
  OR2_X2 U11130 ( .A1(n10859), .A2(P3_D_REG_0__SCAN_IN), .ZN(n8511) );
  OR2_X1 U11131 ( .A1(n10859), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8514) );
  NAND2_X1 U11132 ( .A1(n12959), .A2(n13809), .ZN(n8513) );
  NAND2_X1 U11133 ( .A1(n8514), .A2(n8513), .ZN(n9338) );
  NAND2_X1 U11134 ( .A1(n13796), .A2(n9338), .ZN(n9556) );
  AND2_X1 U11135 ( .A1(n8515), .A2(n9556), .ZN(n9344) );
  OR2_X1 U11136 ( .A1(n13796), .A2(n9338), .ZN(n9549) );
  OAI22_X1 U11137 ( .A1(n15715), .A2(n9552), .B1(n11284), .B2(n11964), .ZN(
        n8516) );
  NAND2_X1 U11138 ( .A1(n8516), .A2(n13183), .ZN(n8517) );
  NAND2_X1 U11139 ( .A1(n8517), .A2(n13172), .ZN(n8518) );
  NAND2_X1 U11140 ( .A1(n8518), .A2(n9338), .ZN(n8521) );
  AND2_X1 U11141 ( .A1(n13168), .A2(n13183), .ZN(n9340) );
  INV_X1 U11142 ( .A(n9340), .ZN(n11171) );
  INV_X1 U11143 ( .A(n9338), .ZN(n13795) );
  AND2_X1 U11144 ( .A1(n13172), .A2(n8519), .ZN(n9337) );
  NAND2_X1 U11145 ( .A1(n13795), .A2(n9337), .ZN(n8520) );
  AND2_X2 U11146 ( .A1(n9344), .A2(n8522), .ZN(n15734) );
  XNOR2_X1 U11147 ( .A(n9304), .B(n8523), .ZN(n12954) );
  NAND2_X1 U11148 ( .A1(n12954), .A2(n12988), .ZN(n8525) );
  INV_X1 U11149 ( .A(n15715), .ZN(n15703) );
  NAND2_X1 U11150 ( .A1(n15734), .A2(n15703), .ZN(n13709) );
  INV_X1 U11151 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n8526) );
  INV_X1 U11152 ( .A(n8527), .ZN(n8528) );
  NOR2_X1 U11153 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), 
        .ZN(n8535) );
  INV_X1 U11154 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8534) );
  NAND4_X1 U11155 ( .A1(n8535), .A2(n8740), .A3(n8741), .A4(n8534), .ZN(n8537)
         );
  NAND4_X1 U11156 ( .A1(n8882), .A2(n8764), .A3(n8873), .A4(n8766), .ZN(n8536)
         );
  NOR2_X1 U11157 ( .A1(n8537), .A2(n8536), .ZN(n8538) );
  INV_X1 U11158 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8540) );
  INV_X1 U11159 ( .A(n8544), .ZN(n8554) );
  AND2_X1 U11160 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8545) );
  AND2_X1 U11161 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U11162 ( .A1(n10818), .A2(n8546), .ZN(n8552) );
  INV_X1 U11163 ( .A(SI_1_), .ZN(n10842) );
  XNOR2_X1 U11164 ( .A(n8560), .B(n10842), .ZN(n8548) );
  OR2_X1 U11165 ( .A1(n8566), .A2(n10875), .ZN(n8549) );
  NAND2_X1 U11166 ( .A1(n10817), .A2(SI_0_), .ZN(n8551) );
  NAND2_X1 U11167 ( .A1(n8551), .A2(n8550), .ZN(n8553) );
  AND2_X1 U11168 ( .A1(n8553), .A2(n8552), .ZN(n14648) );
  NAND2_X1 U11169 ( .A1(n8554), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8555) );
  MUX2_X1 U11170 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8555), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n8557) );
  INV_X1 U11171 ( .A(n8556), .ZN(n8572) );
  INV_X1 U11172 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10798) );
  NAND2_X1 U11173 ( .A1(n10818), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8558) );
  OAI211_X1 U11174 ( .C1(n10798), .C2(n10818), .A(n8558), .B(n10842), .ZN(
        n8559) );
  NAND2_X1 U11175 ( .A1(n8560), .A2(n8559), .ZN(n8563) );
  NAND2_X1 U11176 ( .A1(n10818), .A2(n10876), .ZN(n8561) );
  OAI211_X1 U11177 ( .C1(P2_DATAO_REG_1__SCAN_IN), .C2(n10818), .A(n8561), .B(
        SI_1_), .ZN(n8562) );
  INV_X1 U11178 ( .A(n9620), .ZN(n10813) );
  OR2_X1 U11179 ( .A1(n10813), .A2(n8566), .ZN(n8565) );
  OAI211_X2 U11180 ( .C1(n11042), .C2(n11071), .A(n8565), .B(n8564), .ZN(
        n11979) );
  INV_X1 U11181 ( .A(n8567), .ZN(n8568) );
  XNOR2_X1 U11182 ( .A(n8582), .B(SI_3_), .ZN(n8580) );
  XNOR2_X1 U11183 ( .A(n8600), .B(n8580), .ZN(n10789) );
  NAND2_X1 U11184 ( .A1(n8592), .A2(n10789), .ZN(n8576) );
  NAND2_X1 U11185 ( .A1(n8572), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8574) );
  XNOR2_X1 U11186 ( .A(n8574), .B(n8573), .ZN(n15560) );
  OR2_X1 U11187 ( .A1(n11042), .A2(n15560), .ZN(n8575) );
  INV_X1 U11188 ( .A(n13827), .ZN(n12264) );
  NAND2_X1 U11189 ( .A1(n11972), .A2(n12264), .ZN(n11937) );
  NAND2_X1 U11190 ( .A1(n8577), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8578) );
  MUX2_X1 U11191 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8578), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8579) );
  NOR2_X2 U11192 ( .A1(n8577), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8743) );
  INV_X1 U11193 ( .A(n8743), .ZN(n8594) );
  NAND2_X1 U11194 ( .A1(n8579), .A2(n8594), .ZN(n14005) );
  INV_X1 U11195 ( .A(n14005), .ZN(n14000) );
  INV_X1 U11196 ( .A(n8600), .ZN(n8581) );
  NAND2_X1 U11197 ( .A1(n8581), .A2(n8580), .ZN(n8583) );
  NAND2_X1 U11198 ( .A1(n8583), .A2(n8599), .ZN(n8588) );
  XNOR2_X1 U11199 ( .A(n8604), .B(SI_4_), .ZN(n8587) );
  INV_X1 U11200 ( .A(n8587), .ZN(n8584) );
  XNOR2_X1 U11201 ( .A(n8588), .B(n8584), .ZN(n10794) );
  NAND2_X1 U11202 ( .A1(n10794), .A2(n8834), .ZN(n8585) );
  MUX2_X1 U11203 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n10818), .Z(n8609) );
  XNOR2_X1 U11204 ( .A(n8609), .B(SI_5_), .ZN(n8598) );
  NAND2_X1 U11205 ( .A1(n8588), .A2(n8587), .ZN(n8590) );
  INV_X1 U11206 ( .A(n8604), .ZN(n8589) );
  XNOR2_X1 U11207 ( .A(n8598), .B(n8591), .ZN(n10787) );
  CLKBUF_X3 U11208 ( .A(n8592), .Z(n8834) );
  NAND2_X1 U11209 ( .A1(n10787), .A2(n8834), .ZN(n8597) );
  NAND2_X1 U11210 ( .A1(n8594), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8593) );
  MUX2_X1 U11211 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8593), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8595) );
  AND2_X1 U11212 ( .A1(n8595), .A2(n8619), .ZN(n11087) );
  AOI22_X1 U11213 ( .A1(n8769), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8768), .B2(
        n11087), .ZN(n8596) );
  NOR2_X1 U11214 ( .A1(n8601), .A2(SI_3_), .ZN(n8602) );
  NAND2_X1 U11215 ( .A1(n8604), .A2(n8603), .ZN(n8605) );
  NAND2_X1 U11216 ( .A1(n8609), .A2(SI_5_), .ZN(n8610) );
  MUX2_X1 U11217 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n8650), .Z(n8617) );
  XNOR2_X1 U11218 ( .A(n8616), .B(n8614), .ZN(n10791) );
  NAND2_X1 U11219 ( .A1(n10791), .A2(n8834), .ZN(n8613) );
  NAND2_X1 U11220 ( .A1(n8619), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8611) );
  XNOR2_X1 U11221 ( .A(n8611), .B(P2_IR_REG_6__SCAN_IN), .ZN(n14023) );
  AOI22_X1 U11222 ( .A1(n8769), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8768), .B2(
        n14023), .ZN(n8612) );
  NAND2_X1 U11223 ( .A1(n8617), .A2(SI_6_), .ZN(n8618) );
  MUX2_X1 U11224 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10818), .Z(n8625) );
  INV_X1 U11225 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8620) );
  NAND2_X1 U11226 ( .A1(n8726), .A2(n8620), .ZN(n8627) );
  NAND2_X1 U11227 ( .A1(n8627), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8621) );
  XNOR2_X1 U11228 ( .A(n8621), .B(P2_IR_REG_7__SCAN_IN), .ZN(n11228) );
  AOI22_X1 U11229 ( .A1(n8769), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8768), .B2(
        n11228), .ZN(n8622) );
  NAND2_X1 U11230 ( .A1(n12252), .A2(n12375), .ZN(n12251) );
  NAND2_X1 U11231 ( .A1(n8625), .A2(SI_7_), .ZN(n8626) );
  XNOR2_X1 U11232 ( .A(n8633), .B(n8635), .ZN(n10860) );
  NAND2_X1 U11233 ( .A1(n10860), .A2(n8834), .ZN(n8632) );
  NAND2_X1 U11234 ( .A1(n8629), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8628) );
  MUX2_X1 U11235 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8628), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8630) );
  NAND2_X1 U11236 ( .A1(n8630), .A2(n8638), .ZN(n11243) );
  INV_X1 U11237 ( .A(n11243), .ZN(n11093) );
  AOI22_X1 U11238 ( .A1(n8769), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8768), .B2(
        n11093), .ZN(n8631) );
  MUX2_X1 U11239 ( .A(n10878), .B(n10880), .S(n8650), .Z(n8647) );
  XNOR2_X1 U11240 ( .A(n8646), .B(n7252), .ZN(n10877) );
  NAND2_X1 U11241 ( .A1(n10877), .A2(n8834), .ZN(n8644) );
  NAND2_X1 U11242 ( .A1(n8638), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8637) );
  MUX2_X1 U11243 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8637), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n8641) );
  INV_X1 U11244 ( .A(n8638), .ZN(n8640) );
  INV_X1 U11245 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8639) );
  NAND2_X1 U11246 ( .A1(n8640), .A2(n8639), .ZN(n8662) );
  NAND2_X1 U11247 ( .A1(n8641), .A2(n8662), .ZN(n11422) );
  OAI22_X1 U11248 ( .A1(n10880), .A2(n8866), .B1(n11422), .B2(n11042), .ZN(
        n8642) );
  INV_X1 U11249 ( .A(n8642), .ZN(n8643) );
  INV_X1 U11250 ( .A(n8647), .ZN(n8648) );
  NAND2_X1 U11251 ( .A1(n8648), .A2(SI_9_), .ZN(n8649) );
  MUX2_X1 U11252 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n8650), .Z(n8657) );
  XNOR2_X1 U11253 ( .A(n8656), .B(n8654), .ZN(n10898) );
  NAND2_X1 U11254 ( .A1(n10898), .A2(n8834), .ZN(n8653) );
  NAND2_X1 U11255 ( .A1(n8662), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8651) );
  AOI22_X1 U11256 ( .A1(n11462), .A2(n8768), .B1(P1_DATAO_REG_10__SCAN_IN), 
        .B2(n8769), .ZN(n8652) );
  NAND2_X1 U11257 ( .A1(n8657), .A2(SI_10_), .ZN(n8658) );
  MUX2_X1 U11258 ( .A(n10906), .B(n10905), .S(n8812), .Z(n8659) );
  INV_X1 U11259 ( .A(n8659), .ZN(n8660) );
  NAND2_X1 U11260 ( .A1(n8660), .A2(SI_11_), .ZN(n8661) );
  NAND2_X1 U11261 ( .A1(n10904), .A2(n8834), .ZN(n8665) );
  OAI21_X1 U11262 ( .B1(n8662), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8663) );
  XNOR2_X1 U11263 ( .A(n8663), .B(P2_IR_REG_11__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U11264 ( .A1(n12453), .A2(n8768), .B1(P1_DATAO_REG_11__SCAN_IN), 
        .B2(n8769), .ZN(n8664) );
  INV_X1 U11265 ( .A(n14571), .ZN(n14327) );
  MUX2_X1 U11266 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n8812), .Z(n8667) );
  NAND2_X1 U11267 ( .A1(n8667), .A2(SI_12_), .ZN(n8685) );
  INV_X1 U11268 ( .A(n8667), .ZN(n8668) );
  INV_X1 U11269 ( .A(SI_12_), .ZN(n10872) );
  AND2_X1 U11270 ( .A1(n8685), .A2(n8687), .ZN(n8676) );
  NAND2_X1 U11271 ( .A1(n10982), .A2(n8834), .ZN(n8675) );
  INV_X1 U11272 ( .A(n8669), .ZN(n8670) );
  NAND2_X1 U11273 ( .A1(n8726), .A2(n8670), .ZN(n8672) );
  NAND2_X1 U11274 ( .A1(n8672), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8671) );
  MUX2_X1 U11275 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8671), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8673) );
  AOI22_X1 U11276 ( .A1(n8769), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8768), 
        .B2(n15580), .ZN(n8674) );
  MUX2_X1 U11277 ( .A(n11103), .B(n11025), .S(n8812), .Z(n8689) );
  NAND2_X1 U11278 ( .A1(n11024), .A2(n8834), .ZN(n8683) );
  NAND2_X1 U11279 ( .A1(n8680), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8679) );
  MUX2_X1 U11280 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8679), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8681) );
  NAND2_X1 U11281 ( .A1(n8681), .A2(n8718), .ZN(n12457) );
  AOI22_X1 U11282 ( .A1(n8769), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8768), 
        .B2(n15586), .ZN(n8682) );
  INV_X1 U11283 ( .A(n8685), .ZN(n8702) );
  NAND2_X1 U11284 ( .A1(n6431), .A2(n8685), .ZN(n8686) );
  INV_X1 U11285 ( .A(n8689), .ZN(n8690) );
  NAND2_X1 U11286 ( .A1(n8690), .A2(SI_13_), .ZN(n8700) );
  NAND2_X1 U11287 ( .A1(n8691), .A2(n8700), .ZN(n8695) );
  INV_X1 U11288 ( .A(n8692), .ZN(n8693) );
  NAND2_X1 U11289 ( .A1(n8693), .A2(SI_14_), .ZN(n8694) );
  XNOR2_X2 U11290 ( .A(n8699), .B(n8695), .ZN(n11020) );
  NAND2_X1 U11291 ( .A1(n11020), .A2(n8834), .ZN(n8698) );
  NAND2_X1 U11292 ( .A1(n8718), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8696) );
  XNOR2_X1 U11293 ( .A(n8696), .B(P2_IR_REG_14__SCAN_IN), .ZN(n12466) );
  AOI22_X1 U11294 ( .A1(n8769), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n12466), 
        .B2(n8768), .ZN(n8697) );
  NAND2_X1 U11295 ( .A1(n8703), .A2(n8712), .ZN(n8707) );
  MUX2_X1 U11296 ( .A(n10979), .B(n10980), .S(n8812), .Z(n8704) );
  INV_X1 U11297 ( .A(n8704), .ZN(n8705) );
  NAND2_X1 U11298 ( .A1(n8705), .A2(SI_15_), .ZN(n8706) );
  NAND3_X1 U11299 ( .A1(n8707), .A2(n8714), .A3(n8713), .ZN(n8717) );
  INV_X1 U11300 ( .A(n8714), .ZN(n8709) );
  NAND2_X1 U11301 ( .A1(n10978), .A2(n8834), .ZN(n8721) );
  OAI21_X1 U11302 ( .B1(n8718), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8719) );
  XNOR2_X1 U11303 ( .A(n8719), .B(P2_IR_REG_15__SCAN_IN), .ZN(n12640) );
  AOI22_X1 U11304 ( .A1(n8768), .A2(n12640), .B1(n8769), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n8720) );
  NAND2_X1 U11305 ( .A1(n14311), .A2(n14617), .ZN(n14297) );
  MUX2_X1 U11306 ( .A(n11124), .B(n11069), .S(n8812), .Z(n8723) );
  INV_X1 U11307 ( .A(SI_16_), .ZN(n11019) );
  NAND2_X1 U11308 ( .A1(n8723), .A2(n11019), .ZN(n8733) );
  INV_X1 U11309 ( .A(n8723), .ZN(n8724) );
  NAND2_X1 U11310 ( .A1(n8724), .A2(SI_16_), .ZN(n8725) );
  XNOR2_X1 U11311 ( .A(n8732), .B(n7792), .ZN(n11068) );
  NAND2_X1 U11312 ( .A1(n11068), .A2(n8834), .ZN(n8731) );
  NAND2_X1 U11313 ( .A1(n8726), .A2(n8742), .ZN(n8728) );
  NAND2_X1 U11314 ( .A1(n8728), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8727) );
  MUX2_X1 U11315 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8727), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8729) );
  OR2_X1 U11316 ( .A1(n8728), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n8737) );
  AND2_X1 U11317 ( .A1(n8729), .A2(n8737), .ZN(n12645) );
  AOI22_X1 U11318 ( .A1(n8769), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8768), 
        .B2(n12645), .ZN(n8730) );
  MUX2_X1 U11319 ( .A(n11249), .B(n11196), .S(n8812), .Z(n8734) );
  INV_X1 U11320 ( .A(n8734), .ZN(n8735) );
  NAND2_X1 U11321 ( .A1(n8735), .A2(SI_17_), .ZN(n8736) );
  NAND2_X1 U11322 ( .A1(n11195), .A2(n8834), .ZN(n8747) );
  NAND2_X1 U11323 ( .A1(n8737), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8738) );
  MUX2_X1 U11324 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8738), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8745) );
  INV_X1 U11325 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8739) );
  INV_X1 U11326 ( .A(n8765), .ZN(n8751) );
  NAND2_X1 U11327 ( .A1(n8745), .A2(n8751), .ZN(n12648) );
  INV_X1 U11328 ( .A(n12648), .ZN(n14050) );
  AOI22_X1 U11329 ( .A1(n8769), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8768), 
        .B2(n14050), .ZN(n8746) );
  MUX2_X1 U11330 ( .A(n11482), .B(n11434), .S(n8812), .Z(n8757) );
  XNOR2_X1 U11331 ( .A(n8757), .B(SI_18_), .ZN(n8750) );
  XNOR2_X1 U11332 ( .A(n8773), .B(n8750), .ZN(n11433) );
  NAND2_X1 U11333 ( .A1(n11433), .A2(n8592), .ZN(n8754) );
  NAND2_X1 U11334 ( .A1(n8751), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8752) );
  XNOR2_X1 U11335 ( .A(n8752), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14062) );
  AOI22_X1 U11336 ( .A1(n8769), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8768), 
        .B2(n14062), .ZN(n8753) );
  INV_X1 U11337 ( .A(n14537), .ZN(n14257) );
  INV_X1 U11338 ( .A(SI_18_), .ZN(n11220) );
  NAND2_X1 U11339 ( .A1(n8757), .A2(n11220), .ZN(n8774) );
  NAND3_X1 U11340 ( .A1(n8756), .A2(n8755), .A3(n8774), .ZN(n8759) );
  INV_X1 U11341 ( .A(n8757), .ZN(n8758) );
  NAND2_X1 U11342 ( .A1(n8758), .A2(SI_18_), .ZN(n8772) );
  NAND2_X1 U11343 ( .A1(n8759), .A2(n8772), .ZN(n8763) );
  MUX2_X1 U11344 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n8812), .Z(n8760) );
  NAND2_X1 U11345 ( .A1(n8760), .A2(SI_19_), .ZN(n8777) );
  INV_X1 U11346 ( .A(n8760), .ZN(n8761) );
  INV_X1 U11347 ( .A(SI_19_), .ZN(n11436) );
  NAND2_X1 U11348 ( .A1(n8761), .A2(n11436), .ZN(n8775) );
  NAND2_X1 U11349 ( .A1(n8777), .A2(n8775), .ZN(n8762) );
  NAND2_X1 U11350 ( .A1(n11453), .A2(n8834), .ZN(n8771) );
  NAND2_X1 U11351 ( .A1(n8869), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8767) );
  INV_X1 U11352 ( .A(n8934), .ZN(n14070) );
  AOI22_X1 U11353 ( .A1(n8769), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n14070), 
        .B2(n8768), .ZN(n8770) );
  INV_X1 U11354 ( .A(n8774), .ZN(n8778) );
  INV_X1 U11355 ( .A(n8775), .ZN(n8776) );
  AOI21_X1 U11356 ( .B1(n8778), .B2(n8777), .A(n8776), .ZN(n8779) );
  INV_X1 U11357 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11814) );
  MUX2_X1 U11358 ( .A(n11776), .B(n11814), .S(n8812), .Z(n8788) );
  OR2_X1 U11359 ( .A1(n8866), .A2(n11814), .ZN(n8780) );
  NAND2_X1 U11360 ( .A1(n8781), .A2(n8787), .ZN(n8783) );
  INV_X1 U11361 ( .A(SI_20_), .ZN(n11806) );
  OR2_X1 U11362 ( .A1(n8792), .A2(n11806), .ZN(n8782) );
  MUX2_X1 U11363 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n8812), .Z(n8789) );
  XNOR2_X1 U11364 ( .A(n8789), .B(SI_21_), .ZN(n8784) );
  NAND2_X1 U11365 ( .A1(n11823), .A2(n8834), .ZN(n8786) );
  OR2_X1 U11366 ( .A1(n8866), .A2(n12979), .ZN(n8785) );
  NOR2_X1 U11367 ( .A1(n8788), .A2(n11806), .ZN(n8790) );
  AOI22_X1 U11368 ( .A1(n8790), .A2(n7778), .B1(SI_21_), .B2(n8789), .ZN(n8791) );
  INV_X1 U11369 ( .A(SI_22_), .ZN(n8804) );
  MUX2_X1 U11370 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n8812), .Z(n8807) );
  XNOR2_X1 U11371 ( .A(n9882), .B(n8805), .ZN(n11923) );
  NAND2_X1 U11372 ( .A1(n11923), .A2(n8834), .ZN(n8794) );
  OR2_X1 U11373 ( .A1(n8866), .A2(n11926), .ZN(n8793) );
  AND2_X2 U11374 ( .A1(n14195), .A2(n14599), .ZN(n14178) );
  NAND2_X1 U11375 ( .A1(n9882), .A2(n8807), .ZN(n8796) );
  NAND2_X1 U11376 ( .A1(n8803), .A2(SI_22_), .ZN(n8795) );
  MUX2_X1 U11377 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n8812), .Z(n8808) );
  XNOR2_X1 U11378 ( .A(n8808), .B(SI_23_), .ZN(n8797) );
  OR2_X1 U11379 ( .A1(n8866), .A2(n12043), .ZN(n8799) );
  INV_X1 U11380 ( .A(n8808), .ZN(n8801) );
  INV_X1 U11381 ( .A(SI_23_), .ZN(n12272) );
  AOI22_X1 U11382 ( .A1(n8804), .A2(n8805), .B1(n8801), .B2(n12272), .ZN(n8802) );
  OAI21_X1 U11383 ( .B1(n8805), .B2(n8804), .A(n12272), .ZN(n8809) );
  AND2_X1 U11384 ( .A1(SI_23_), .A2(SI_22_), .ZN(n8806) );
  AOI22_X1 U11385 ( .A1(n8809), .A2(n8808), .B1(n8807), .B2(n8806), .ZN(n8810)
         );
  MUX2_X1 U11386 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n8812), .Z(n8816) );
  NAND2_X1 U11387 ( .A1(n12108), .A2(n8834), .ZN(n8814) );
  OR2_X1 U11388 ( .A1(n8866), .A2(n12111), .ZN(n8813) );
  MUX2_X1 U11389 ( .A(n12242), .B(n12244), .S(n10817), .Z(n8819) );
  INV_X1 U11390 ( .A(SI_25_), .ZN(n13806) );
  NAND2_X1 U11391 ( .A1(n8819), .A2(n13806), .ZN(n8824) );
  INV_X1 U11392 ( .A(n8819), .ZN(n8820) );
  NAND2_X1 U11393 ( .A1(n8820), .A2(SI_25_), .ZN(n8821) );
  NAND2_X1 U11394 ( .A1(n8824), .A2(n8821), .ZN(n8825) );
  OR2_X1 U11395 ( .A1(n8866), .A2(n12244), .ZN(n8822) );
  MUX2_X1 U11396 ( .A(n12547), .B(n12544), .S(n10817), .Z(n8830) );
  XNOR2_X1 U11397 ( .A(n8830), .B(SI_26_), .ZN(n8827) );
  OR2_X1 U11398 ( .A1(n8866), .A2(n12544), .ZN(n8828) );
  INV_X1 U11399 ( .A(SI_26_), .ZN(n12957) );
  NAND2_X1 U11400 ( .A1(n8831), .A2(n12957), .ZN(n8832) );
  INV_X1 U11401 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15434) );
  INV_X1 U11402 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14645) );
  MUX2_X1 U11403 ( .A(n15434), .B(n14645), .S(n10817), .Z(n8837) );
  XNOR2_X1 U11404 ( .A(n8837), .B(SI_27_), .ZN(n8833) );
  OR2_X1 U11405 ( .A1(n8866), .A2(n14645), .ZN(n8835) );
  INV_X1 U11406 ( .A(SI_27_), .ZN(n14412) );
  INV_X1 U11407 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12891) );
  INV_X1 U11408 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9312) );
  MUX2_X1 U11409 ( .A(n12891), .B(n9312), .S(n10817), .Z(n8845) );
  XNOR2_X1 U11410 ( .A(n8845), .B(SI_28_), .ZN(n8842) );
  OR2_X1 U11411 ( .A1(n8866), .A2(n9312), .ZN(n8840) );
  NAND2_X1 U11412 ( .A1(n8843), .A2(n8842), .ZN(n8847) );
  INV_X1 U11413 ( .A(SI_28_), .ZN(n8844) );
  NAND2_X1 U11414 ( .A1(n8845), .A2(n8844), .ZN(n8846) );
  INV_X1 U11415 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15431) );
  INV_X1 U11416 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14638) );
  MUX2_X1 U11417 ( .A(n15431), .B(n14638), .S(n10817), .Z(n8854) );
  XNOR2_X1 U11418 ( .A(n8854), .B(SI_29_), .ZN(n8848) );
  OR2_X1 U11419 ( .A1(n8866), .A2(n14638), .ZN(n8851) );
  INV_X1 U11420 ( .A(n14352), .ZN(n8853) );
  INV_X1 U11421 ( .A(SI_29_), .ZN(n14491) );
  MUX2_X1 U11422 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10817), .Z(n8859) );
  XNOR2_X1 U11423 ( .A(n8859), .B(SI_30_), .ZN(n8860) );
  INV_X1 U11424 ( .A(n8860), .ZN(n8856) );
  NAND2_X1 U11425 ( .A1(n13212), .A2(n8592), .ZN(n8858) );
  INV_X1 U11426 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13217) );
  OR2_X1 U11427 ( .A1(n8866), .A2(n13217), .ZN(n8857) );
  MUX2_X1 U11428 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10817), .Z(n8862) );
  XNOR2_X1 U11429 ( .A(n8862), .B(SI_31_), .ZN(n8863) );
  NAND2_X1 U11430 ( .A1(n10639), .A2(n8834), .ZN(n8868) );
  INV_X1 U11431 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8865) );
  OR2_X1 U11432 ( .A1(n8866), .A2(n8865), .ZN(n8867) );
  NAND2_X2 U11433 ( .A1(n8868), .A2(n8867), .ZN(n9474) );
  NAND2_X1 U11434 ( .A1(n8870), .A2(n8873), .ZN(n8871) );
  INV_X1 U11435 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8876) );
  NAND2_X1 U11436 ( .A1(n8873), .A2(n8876), .ZN(n8879) );
  NAND3_X1 U11437 ( .A1(n8880), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_22__SCAN_IN), .ZN(n8878) );
  NAND2_X1 U11438 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n8874) );
  NAND2_X1 U11439 ( .A1(n8874), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8875) );
  OAI21_X1 U11440 ( .B1(n8876), .B2(P2_IR_REG_31__SCAN_IN), .A(n8875), .ZN(
        n8877) );
  XNOR2_X1 U11441 ( .A(n8883), .B(n8882), .ZN(n8926) );
  BUF_X4 U11442 ( .A(n8989), .Z(n14320) );
  NAND2_X1 U11443 ( .A1(n10453), .A2(n10430), .ZN(n11044) );
  INV_X1 U11444 ( .A(P2_B_REG_SCAN_IN), .ZN(n8910) );
  OR2_X1 U11445 ( .A1(n14647), .A2(n8910), .ZN(n8886) );
  AND2_X1 U11446 ( .A1(n14286), .A2(n8886), .ZN(n10458) );
  INV_X1 U11447 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8889) );
  XNOR2_X1 U11448 ( .A(n8890), .B(n8889), .ZN(n13216) );
  INV_X1 U11449 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8888) );
  INV_X1 U11450 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8937) );
  AND2_X2 U11451 ( .A1(n8891), .A2(n14635), .ZN(n8996) );
  INV_X2 U11452 ( .A(n9262), .ZN(n9245) );
  NAND2_X1 U11453 ( .A1(n9245), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8894) );
  INV_X1 U11454 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8892) );
  OR2_X1 U11455 ( .A1(n8984), .A2(n8892), .ZN(n8893) );
  OAI211_X1 U11456 ( .C1(n9469), .C2(n8937), .A(n8894), .B(n8893), .ZN(n13958)
         );
  AND2_X1 U11457 ( .A1(n10458), .A2(n13958), .ZN(n14347) );
  NOR2_X1 U11458 ( .A1(n14073), .A2(n14347), .ZN(n10701) );
  OR2_X1 U11459 ( .A1(n8895), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n8906) );
  INV_X1 U11460 ( .A(n8906), .ZN(n8897) );
  NAND2_X1 U11461 ( .A1(n8897), .A2(n8896), .ZN(n8908) );
  INV_X1 U11462 ( .A(n8908), .ZN(n8899) );
  NAND2_X1 U11463 ( .A1(n8899), .A2(n8898), .ZN(n8904) );
  NAND2_X1 U11464 ( .A1(n8904), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8900) );
  MUX2_X1 U11465 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8900), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8902) );
  AND2_X1 U11466 ( .A1(n8902), .A2(n8901), .ZN(n8931) );
  NAND2_X1 U11467 ( .A1(n8908), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8903) );
  MUX2_X1 U11468 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8903), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8905) );
  NAND2_X1 U11469 ( .A1(n8905), .A2(n8904), .ZN(n12246) );
  NAND2_X1 U11470 ( .A1(n8906), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8907) );
  MUX2_X1 U11471 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8907), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8909) );
  NAND2_X1 U11472 ( .A1(n8909), .A2(n8908), .ZN(n12113) );
  XOR2_X1 U11473 ( .A(n8910), .B(n12113), .Z(n8911) );
  NAND2_X1 U11474 ( .A1(n12246), .A2(n8911), .ZN(n8912) );
  NOR2_X1 U11475 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .ZN(
        n8916) );
  NOR4_X1 U11476 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n8915) );
  NOR4_X1 U11477 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8914) );
  NOR4_X1 U11478 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n8913) );
  AND4_X1 U11479 ( .A1(n8916), .A2(n8915), .A3(n8914), .A4(n8913), .ZN(n8922)
         );
  NOR4_X1 U11480 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8920) );
  NOR4_X1 U11481 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8919) );
  NOR4_X1 U11482 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8918) );
  NOR4_X1 U11483 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8917) );
  AND4_X1 U11484 ( .A1(n8920), .A2(n8919), .A3(n8918), .A4(n8917), .ZN(n8921)
         );
  NAND2_X1 U11485 ( .A1(n8922), .A2(n8921), .ZN(n8923) );
  AND2_X1 U11486 ( .A1(n15634), .A2(n8923), .ZN(n9268) );
  INV_X1 U11487 ( .A(n9268), .ZN(n8927) );
  INV_X1 U11488 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15643) );
  NAND2_X1 U11489 ( .A1(n15634), .A2(n15643), .ZN(n8925) );
  INV_X1 U11490 ( .A(n8931), .ZN(n12545) );
  NAND2_X1 U11491 ( .A1(n12545), .A2(n12246), .ZN(n8924) );
  NAND2_X1 U11492 ( .A1(n8925), .A2(n8924), .ZN(n15644) );
  AND2_X2 U11493 ( .A1(n8926), .A2(n14070), .ZN(n11596) );
  AND2_X2 U11494 ( .A1(n11596), .A2(n11924), .ZN(n15653) );
  NAND2_X1 U11495 ( .A1(n15653), .A2(n9533), .ZN(n9290) );
  NAND3_X1 U11496 ( .A1(n8927), .A2(n15644), .A3(n9290), .ZN(n10440) );
  INV_X1 U11497 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15640) );
  NAND2_X1 U11498 ( .A1(n15634), .A2(n15640), .ZN(n8929) );
  NAND2_X1 U11499 ( .A1(n12545), .A2(n12113), .ZN(n8928) );
  NAND2_X1 U11500 ( .A1(n8929), .A2(n8928), .ZN(n15641) );
  INV_X1 U11501 ( .A(n15641), .ZN(n8935) );
  NOR2_X1 U11502 ( .A1(n12246), .A2(n12113), .ZN(n8930) );
  NAND2_X1 U11503 ( .A1(n8931), .A2(n8930), .ZN(n10707) );
  NAND2_X1 U11504 ( .A1(n8895), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8933) );
  XNOR2_X1 U11505 ( .A(n8933), .B(n8932), .ZN(n10706) );
  NAND2_X1 U11506 ( .A1(n11815), .A2(n11455), .ZN(n9539) );
  NAND2_X1 U11507 ( .A1(n9288), .A2(n9539), .ZN(n10439) );
  NAND3_X1 U11508 ( .A1(n8935), .A2(n15645), .A3(n10439), .ZN(n8936) );
  INV_X2 U11509 ( .A(n15668), .ZN(n15670) );
  NAND2_X1 U11510 ( .A1(n9274), .A2(n9539), .ZN(n15648) );
  NAND2_X1 U11511 ( .A1(n15670), .A2(n15656), .ZN(n14582) );
  NOR2_X1 U11512 ( .A1(n15670), .A2(n8937), .ZN(n8938) );
  OAI21_X1 U11513 ( .B1(n10701), .B2(n15668), .A(n8940), .ZN(P2_U3530) );
  INV_X1 U11514 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11460) );
  INV_X1 U11515 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U11516 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n8944) );
  INV_X1 U11517 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9130) );
  INV_X1 U11518 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9173) );
  INV_X1 U11519 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13920) );
  INV_X1 U11520 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13817) );
  NAND2_X1 U11521 ( .A1(n9207), .A2(n13817), .ZN(n8948) );
  NAND2_X1 U11522 ( .A1(n9220), .A2(n8948), .ZN(n14162) );
  OR2_X1 U11523 ( .A1(n14162), .A2(n9464), .ZN(n8956) );
  INV_X1 U11524 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8953) );
  NAND2_X1 U11525 ( .A1(n9465), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8952) );
  NAND2_X1 U11526 ( .A1(n9245), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8951) );
  OAI211_X1 U11527 ( .C1(n9469), .C2(n8953), .A(n8952), .B(n8951), .ZN(n8954)
         );
  INV_X1 U11528 ( .A(n8954), .ZN(n8955) );
  NAND2_X1 U11529 ( .A1(n8956), .A2(n8955), .ZN(n13963) );
  NAND2_X1 U11530 ( .A1(n10430), .A2(n11455), .ZN(n8957) );
  NAND2_X1 U11531 ( .A1(n8996), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8961) );
  INV_X1 U11532 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11599) );
  INV_X1 U11533 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n11049) );
  NAND2_X1 U11534 ( .A1(n14310), .A2(n11485), .ZN(n8962) );
  NAND2_X1 U11535 ( .A1(n10747), .A2(n8962), .ZN(n11483) );
  AND2_X1 U11536 ( .A1(n9354), .A2(n8969), .ZN(n8963) );
  OR2_X1 U11537 ( .A1(n8984), .A2(n13984), .ZN(n8968) );
  NAND2_X1 U11538 ( .A1(n8996), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8967) );
  INV_X1 U11539 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n13980) );
  INV_X1 U11540 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n8964) );
  OR2_X1 U11541 ( .A1(n8983), .A2(n8964), .ZN(n8965) );
  AND4_X2 U11542 ( .A1(n8968), .A2(n8967), .A3(n8966), .A4(n8965), .ZN(n10330)
         );
  NAND2_X1 U11543 ( .A1(n9353), .A2(n8989), .ZN(n8979) );
  XNOR2_X1 U11544 ( .A(n13859), .B(n8969), .ZN(n8978) );
  XNOR2_X1 U11545 ( .A(n8979), .B(n8978), .ZN(n13862) );
  INV_X1 U11546 ( .A(n8982), .ZN(n8977) );
  NAND2_X1 U11547 ( .A1(n8996), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8975) );
  NAND2_X1 U11548 ( .A1(n8970), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8974) );
  INV_X1 U11549 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11975) );
  INV_X1 U11550 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n8971) );
  OR2_X1 U11551 ( .A1(n8983), .A2(n8971), .ZN(n8972) );
  NAND4_X4 U11552 ( .A1(n8975), .A2(n8974), .A3(n8973), .A4(n8972), .ZN(n9514)
         );
  NAND2_X1 U11553 ( .A1(n9514), .A2(n8989), .ZN(n8981) );
  INV_X1 U11554 ( .A(n8981), .ZN(n8976) );
  INV_X1 U11555 ( .A(n11473), .ZN(n8991) );
  INV_X1 U11556 ( .A(n8978), .ZN(n8980) );
  AND2_X1 U11557 ( .A1(n8980), .A2(n8979), .ZN(n11471) );
  XNOR2_X1 U11558 ( .A(n13827), .B(n8969), .ZN(n8993) );
  NAND2_X1 U11559 ( .A1(n8996), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8988) );
  NAND2_X1 U11560 ( .A1(n9259), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8987) );
  OR2_X1 U11561 ( .A1(n9464), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8986) );
  INV_X1 U11562 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n12262) );
  OR2_X1 U11563 ( .A1(n8984), .A2(n12262), .ZN(n8985) );
  NAND2_X1 U11564 ( .A1(n13978), .A2(n8989), .ZN(n8992) );
  XNOR2_X1 U11565 ( .A(n8993), .B(n8992), .ZN(n13825) );
  INV_X1 U11566 ( .A(n8992), .ZN(n8994) );
  NAND2_X1 U11567 ( .A1(n8994), .A2(n8993), .ZN(n8995) );
  NAND2_X1 U11568 ( .A1(n9259), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9000) );
  NAND2_X1 U11569 ( .A1(n9245), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8999) );
  OAI21_X1 U11570 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n9008), .ZN(n11940) );
  OR2_X1 U11571 ( .A1(n9464), .A2(n11940), .ZN(n8998) );
  INV_X1 U11572 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11083) );
  OR2_X1 U11573 ( .A1(n8984), .A2(n11083), .ZN(n8997) );
  NAND2_X1 U11574 ( .A1(n13977), .A2(n8989), .ZN(n9002) );
  NAND2_X1 U11575 ( .A1(n9001), .A2(n9002), .ZN(n9007) );
  INV_X1 U11576 ( .A(n9001), .ZN(n9004) );
  INV_X1 U11577 ( .A(n9002), .ZN(n9003) );
  NAND2_X1 U11578 ( .A1(n9004), .A2(n9003), .ZN(n9005) );
  NAND2_X1 U11579 ( .A1(n9007), .A2(n9005), .ZN(n11639) );
  NAND2_X1 U11580 ( .A1(n11637), .A2(n9007), .ZN(n11575) );
  NAND2_X1 U11581 ( .A1(n9259), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9013) );
  NAND2_X1 U11582 ( .A1(n8996), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9012) );
  NAND2_X1 U11583 ( .A1(n9008), .A2(n6691), .ZN(n9009) );
  NAND2_X1 U11584 ( .A1(n9020), .A2(n9009), .ZN(n11958) );
  OR2_X1 U11585 ( .A1(n9464), .A2(n11958), .ZN(n9011) );
  INV_X1 U11586 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11957) );
  OR2_X1 U11587 ( .A1(n8984), .A2(n11957), .ZN(n9010) );
  NAND4_X1 U11588 ( .A1(n9013), .A2(n9012), .A3(n9011), .A4(n9010), .ZN(n13976) );
  NAND2_X1 U11589 ( .A1(n13976), .A2(n8989), .ZN(n9015) );
  NAND2_X1 U11590 ( .A1(n9014), .A2(n9015), .ZN(n9019) );
  INV_X1 U11591 ( .A(n9014), .ZN(n9017) );
  INV_X1 U11592 ( .A(n9015), .ZN(n9016) );
  NAND2_X1 U11593 ( .A1(n9017), .A2(n9016), .ZN(n9018) );
  AND2_X1 U11594 ( .A1(n9019), .A2(n9018), .ZN(n11576) );
  NAND2_X1 U11595 ( .A1(n9245), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9025) );
  NAND2_X1 U11596 ( .A1(n9465), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9024) );
  NAND2_X1 U11597 ( .A1(n9020), .A2(n6692), .ZN(n9021) );
  NAND2_X1 U11598 ( .A1(n9032), .A2(n9021), .ZN(n12065) );
  OR2_X1 U11599 ( .A1(n9464), .A2(n12065), .ZN(n9023) );
  INV_X1 U11600 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n11075) );
  OR2_X1 U11601 ( .A1(n9469), .A2(n11075), .ZN(n9022) );
  NAND2_X1 U11602 ( .A1(n13975), .A2(n8989), .ZN(n9027) );
  XNOR2_X1 U11603 ( .A(n9026), .B(n9027), .ZN(n11627) );
  INV_X1 U11604 ( .A(n9026), .ZN(n9029) );
  INV_X1 U11605 ( .A(n9027), .ZN(n9028) );
  NAND2_X1 U11606 ( .A1(n9029), .A2(n9028), .ZN(n9030) );
  XNOR2_X1 U11607 ( .A(n15624), .B(n8969), .ZN(n9040) );
  NAND2_X1 U11608 ( .A1(n9259), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9037) );
  NAND2_X1 U11609 ( .A1(n9245), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9036) );
  INV_X1 U11610 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9031) );
  NAND2_X1 U11611 ( .A1(n9032), .A2(n9031), .ZN(n9033) );
  NAND2_X1 U11612 ( .A1(n9053), .A2(n9033), .ZN(n15620) );
  OR2_X1 U11613 ( .A1(n9464), .A2(n15620), .ZN(n9035) );
  INV_X1 U11614 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n15621) );
  OR2_X1 U11615 ( .A1(n8984), .A2(n15621), .ZN(n9034) );
  NAND4_X1 U11616 ( .A1(n9037), .A2(n9036), .A3(n9035), .A4(n9034), .ZN(n13974) );
  NAND2_X1 U11617 ( .A1(n13974), .A2(n14320), .ZN(n9038) );
  INV_X1 U11618 ( .A(n9038), .ZN(n9039) );
  NAND2_X1 U11619 ( .A1(n9259), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9044) );
  NAND2_X1 U11620 ( .A1(n9245), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9043) );
  INV_X1 U11621 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9052) );
  XNOR2_X1 U11622 ( .A(n9053), .B(n9052), .ZN(n12384) );
  OR2_X1 U11623 ( .A1(n9464), .A2(n12384), .ZN(n9042) );
  INV_X1 U11624 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n12382) );
  OR2_X1 U11625 ( .A1(n8984), .A2(n12382), .ZN(n9041) );
  NAND4_X1 U11626 ( .A1(n9044), .A2(n9043), .A3(n9042), .A4(n9041), .ZN(n13973) );
  NAND2_X1 U11627 ( .A1(n13973), .A2(n14320), .ZN(n9046) );
  NAND2_X1 U11628 ( .A1(n9045), .A2(n9046), .ZN(n9050) );
  INV_X1 U11629 ( .A(n9045), .ZN(n9048) );
  INV_X1 U11630 ( .A(n9046), .ZN(n9047) );
  NAND2_X1 U11631 ( .A1(n9048), .A2(n9047), .ZN(n9049) );
  AND2_X1 U11632 ( .A1(n9050), .A2(n9049), .ZN(n12003) );
  NAND2_X1 U11633 ( .A1(n9245), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9058) );
  NAND2_X1 U11634 ( .A1(n9465), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9057) );
  INV_X1 U11635 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11070) );
  OR2_X1 U11636 ( .A1(n9469), .A2(n11070), .ZN(n9056) );
  INV_X1 U11637 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9051) );
  OAI21_X1 U11638 ( .B1(n9053), .B2(n9052), .A(n9051), .ZN(n9054) );
  NAND2_X1 U11639 ( .A1(n9054), .A2(n9066), .ZN(n12595) );
  OR2_X1 U11640 ( .A1(n9464), .A2(n12595), .ZN(n9055) );
  NAND4_X1 U11641 ( .A1(n9058), .A2(n9057), .A3(n9056), .A4(n9055), .ZN(n13971) );
  NAND2_X1 U11642 ( .A1(n13971), .A2(n14320), .ZN(n9060) );
  NAND2_X1 U11643 ( .A1(n9059), .A2(n9060), .ZN(n9064) );
  INV_X1 U11644 ( .A(n9059), .ZN(n9062) );
  INV_X1 U11645 ( .A(n9060), .ZN(n9061) );
  NAND2_X1 U11646 ( .A1(n9062), .A2(n9061), .ZN(n9063) );
  AND2_X1 U11647 ( .A1(n9064), .A2(n9063), .ZN(n12136) );
  NAND2_X1 U11648 ( .A1(n9259), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9071) );
  NAND2_X1 U11649 ( .A1(n9465), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9070) );
  INV_X1 U11650 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14625) );
  OR2_X1 U11651 ( .A1(n9262), .A2(n14625), .ZN(n9069) );
  INV_X1 U11652 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9065) );
  NAND2_X1 U11653 ( .A1(n9066), .A2(n9065), .ZN(n9067) );
  NAND2_X1 U11654 ( .A1(n9072), .A2(n9067), .ZN(n12736) );
  OR2_X1 U11655 ( .A1(n9464), .A2(n12736), .ZN(n9068) );
  NAND4_X1 U11656 ( .A1(n9071), .A2(n9070), .A3(n9069), .A4(n9068), .ZN(n14329) );
  NAND2_X1 U11657 ( .A1(n14329), .A2(n14320), .ZN(n9086) );
  XNOR2_X1 U11658 ( .A(n9085), .B(n9086), .ZN(n12482) );
  NAND2_X1 U11659 ( .A1(n9259), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9078) );
  NAND2_X1 U11660 ( .A1(n9245), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n9077) );
  NAND2_X1 U11661 ( .A1(n9072), .A2(n11460), .ZN(n9073) );
  NAND2_X1 U11662 ( .A1(n9094), .A2(n9073), .ZN(n14322) );
  OR2_X1 U11663 ( .A1(n9464), .A2(n14322), .ZN(n9076) );
  INV_X1 U11664 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9074) );
  OR2_X1 U11665 ( .A1(n8984), .A2(n9074), .ZN(n9075) );
  NAND4_X1 U11666 ( .A1(n9078), .A2(n9077), .A3(n9076), .A4(n9075), .ZN(n13970) );
  NAND2_X1 U11667 ( .A1(n13970), .A2(n14320), .ZN(n9080) );
  NAND2_X1 U11668 ( .A1(n9079), .A2(n9080), .ZN(n9084) );
  INV_X1 U11669 ( .A(n9084), .ZN(n9091) );
  INV_X1 U11670 ( .A(n9079), .ZN(n9082) );
  INV_X1 U11671 ( .A(n9080), .ZN(n9081) );
  NAND2_X1 U11672 ( .A1(n9082), .A2(n9081), .ZN(n9083) );
  NAND2_X1 U11673 ( .A1(n9084), .A2(n9083), .ZN(n12486) );
  INV_X1 U11674 ( .A(n12486), .ZN(n9089) );
  INV_X1 U11675 ( .A(n9085), .ZN(n9088) );
  INV_X1 U11676 ( .A(n9086), .ZN(n9087) );
  NAND2_X1 U11677 ( .A1(n9088), .A2(n9087), .ZN(n12484) );
  AND2_X1 U11678 ( .A1(n9089), .A2(n12484), .ZN(n9090) );
  INV_X1 U11679 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9092) );
  OR2_X1 U11680 ( .A1(n9469), .A2(n9092), .ZN(n9099) );
  NAND2_X1 U11681 ( .A1(n9245), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9098) );
  NAND2_X1 U11682 ( .A1(n9094), .A2(n9093), .ZN(n9095) );
  NAND2_X1 U11683 ( .A1(n9117), .A2(n9095), .ZN(n12604) );
  OR2_X1 U11684 ( .A1(n9464), .A2(n12604), .ZN(n9097) );
  INV_X1 U11685 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n12605) );
  OR2_X1 U11686 ( .A1(n8984), .A2(n12605), .ZN(n9096) );
  NAND4_X1 U11687 ( .A1(n9099), .A2(n9098), .A3(n9097), .A4(n9096), .ZN(n13969) );
  NAND2_X1 U11688 ( .A1(n13969), .A2(n14320), .ZN(n9101) );
  NAND2_X1 U11689 ( .A1(n9100), .A2(n9101), .ZN(n9105) );
  INV_X1 U11690 ( .A(n9100), .ZN(n9103) );
  INV_X1 U11691 ( .A(n9101), .ZN(n9102) );
  NAND2_X1 U11692 ( .A1(n9103), .A2(n9102), .ZN(n9104) );
  NAND2_X1 U11693 ( .A1(n9259), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U11694 ( .A1(n9245), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9108) );
  INV_X1 U11695 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9116) );
  XNOR2_X1 U11696 ( .A(n9117), .B(n9116), .ZN(n12679) );
  OR2_X1 U11697 ( .A1(n9464), .A2(n12679), .ZN(n9107) );
  INV_X1 U11698 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n12680) );
  OR2_X1 U11699 ( .A1(n8984), .A2(n12680), .ZN(n9106) );
  NAND4_X1 U11700 ( .A1(n9109), .A2(n9108), .A3(n9107), .A4(n9106), .ZN(n13968) );
  NAND2_X1 U11701 ( .A1(n13968), .A2(n14320), .ZN(n9111) );
  XNOR2_X1 U11702 ( .A(n9110), .B(n9111), .ZN(n12549) );
  INV_X1 U11703 ( .A(n12549), .ZN(n9114) );
  INV_X1 U11704 ( .A(n9110), .ZN(n9113) );
  INV_X1 U11705 ( .A(n9111), .ZN(n9112) );
  NAND2_X1 U11706 ( .A1(n9259), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9123) );
  NAND2_X1 U11707 ( .A1(n9245), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n9122) );
  INV_X1 U11708 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9115) );
  OAI21_X1 U11709 ( .B1(n9117), .B2(n9116), .A(n9115), .ZN(n9118) );
  NAND2_X1 U11710 ( .A1(n9137), .A2(n9118), .ZN(n12807) );
  OR2_X1 U11711 ( .A1(n9464), .A2(n12807), .ZN(n9121) );
  INV_X1 U11712 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9119) );
  OR2_X1 U11713 ( .A1(n8984), .A2(n9119), .ZN(n9120) );
  NAND4_X1 U11714 ( .A1(n9123), .A2(n9122), .A3(n9121), .A4(n9120), .ZN(n13967) );
  NAND2_X1 U11715 ( .A1(n13967), .A2(n14320), .ZN(n9125) );
  NAND2_X1 U11716 ( .A1(n9124), .A2(n9125), .ZN(n9129) );
  INV_X1 U11717 ( .A(n9124), .ZN(n9127) );
  INV_X1 U11718 ( .A(n9125), .ZN(n9126) );
  NAND2_X1 U11719 ( .A1(n9127), .A2(n9126), .ZN(n9128) );
  NAND2_X1 U11720 ( .A1(n9139), .A2(n9130), .ZN(n9131) );
  NAND2_X1 U11721 ( .A1(n9155), .A2(n9131), .ZN(n14283) );
  NAND2_X1 U11722 ( .A1(n9465), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9132) );
  OAI21_X1 U11723 ( .B1(n14283), .B2(n9464), .A(n9132), .ZN(n9135) );
  INV_X1 U11724 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n12637) );
  NAND2_X1 U11725 ( .A1(n9245), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n9133) );
  OAI21_X1 U11726 ( .B1(n12637), .B2(n9469), .A(n9133), .ZN(n9134) );
  NAND2_X1 U11727 ( .A1(n13966), .A2(n14320), .ZN(n9148) );
  NAND2_X1 U11728 ( .A1(n9147), .A2(n9148), .ZN(n13877) );
  XNOR2_X1 U11729 ( .A(n14313), .B(n8969), .ZN(n9145) );
  INV_X1 U11730 ( .A(n9145), .ZN(n13879) );
  NAND2_X1 U11731 ( .A1(n9245), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n9143) );
  NAND2_X1 U11732 ( .A1(n9465), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n9142) );
  INV_X1 U11733 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14558) );
  OR2_X1 U11734 ( .A1(n9469), .A2(n14558), .ZN(n9141) );
  INV_X1 U11735 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9136) );
  NAND2_X1 U11736 ( .A1(n9137), .A2(n9136), .ZN(n9138) );
  NAND2_X1 U11737 ( .A1(n9139), .A2(n9138), .ZN(n14309) );
  OR2_X1 U11738 ( .A1(n9464), .A2(n14309), .ZN(n9140) );
  NAND4_X1 U11739 ( .A1(n9143), .A2(n9142), .A3(n9141), .A4(n9140), .ZN(n14284) );
  AND2_X1 U11740 ( .A1(n14284), .A2(n14320), .ZN(n9146) );
  INV_X1 U11741 ( .A(n9146), .ZN(n13945) );
  NAND2_X1 U11742 ( .A1(n13879), .A2(n13945), .ZN(n9144) );
  NAND2_X1 U11743 ( .A1(n13877), .A2(n9144), .ZN(n9153) );
  NAND3_X1 U11744 ( .A1(n13877), .A2(n9146), .A3(n9145), .ZN(n9151) );
  INV_X1 U11745 ( .A(n9147), .ZN(n9150) );
  INV_X1 U11746 ( .A(n9148), .ZN(n9149) );
  NAND2_X1 U11747 ( .A1(n9150), .A2(n9149), .ZN(n13876) );
  INV_X1 U11748 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n14277) );
  INV_X1 U11749 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9154) );
  NAND2_X1 U11750 ( .A1(n9155), .A2(n9154), .ZN(n9156) );
  NAND2_X1 U11751 ( .A1(n9166), .A2(n9156), .ZN(n14276) );
  OR2_X1 U11752 ( .A1(n14276), .A2(n9464), .ZN(n9158) );
  AOI22_X1 U11753 ( .A1(n9259), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n9245), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n9157) );
  OAI211_X1 U11754 ( .C1(n8984), .C2(n14277), .A(n9158), .B(n9157), .ZN(n14287) );
  NAND2_X1 U11755 ( .A1(n14287), .A2(n14320), .ZN(n9160) );
  NAND2_X1 U11756 ( .A1(n9159), .A2(n9160), .ZN(n9164) );
  INV_X1 U11757 ( .A(n9159), .ZN(n9162) );
  INV_X1 U11758 ( .A(n9160), .ZN(n9161) );
  NAND2_X1 U11759 ( .A1(n9162), .A2(n9161), .ZN(n9163) );
  NAND2_X1 U11760 ( .A1(n9164), .A2(n9163), .ZN(n13888) );
  INV_X1 U11761 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9170) );
  INV_X1 U11762 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9165) );
  NAND2_X1 U11763 ( .A1(n9166), .A2(n9165), .ZN(n9167) );
  NAND2_X1 U11764 ( .A1(n9174), .A2(n9167), .ZN(n14254) );
  OR2_X1 U11765 ( .A1(n14254), .A2(n9464), .ZN(n9169) );
  AOI22_X1 U11766 ( .A1(n9259), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n9245), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n9168) );
  OAI211_X1 U11767 ( .C1(n8984), .C2(n9170), .A(n9169), .B(n9168), .ZN(n13965)
         );
  NAND2_X1 U11768 ( .A1(n13965), .A2(n14320), .ZN(n9171) );
  XNOR2_X1 U11769 ( .A(n9172), .B(n9171), .ZN(n13927) );
  XNOR2_X1 U11770 ( .A(n14232), .B(n8969), .ZN(n9178) );
  NAND2_X1 U11771 ( .A1(n9174), .A2(n9173), .ZN(n9175) );
  NAND2_X1 U11772 ( .A1(n9192), .A2(n9175), .ZN(n14233) );
  AOI22_X1 U11773 ( .A1(n9259), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n9245), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n9177) );
  NAND2_X1 U11774 ( .A1(n9465), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n9176) );
  OAI211_X1 U11775 ( .C1(n14233), .C2(n9464), .A(n9177), .B(n9176), .ZN(n14207) );
  AND2_X1 U11776 ( .A1(n14207), .A2(n14320), .ZN(n9179) );
  INV_X1 U11777 ( .A(n9178), .ZN(n9181) );
  INV_X1 U11778 ( .A(n9179), .ZN(n9180) );
  NAND2_X1 U11779 ( .A1(n9181), .A2(n9180), .ZN(n13832) );
  XNOR2_X1 U11780 ( .A(n14393), .B(n8969), .ZN(n9188) );
  XNOR2_X1 U11781 ( .A(n9192), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n14210) );
  NAND2_X1 U11782 ( .A1(n14210), .A2(n9258), .ZN(n9187) );
  INV_X1 U11783 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9184) );
  NAND2_X1 U11784 ( .A1(n9465), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9183) );
  NAND2_X1 U11785 ( .A1(n9245), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9182) );
  OAI211_X1 U11786 ( .C1(n9469), .C2(n9184), .A(n9183), .B(n9182), .ZN(n9185)
         );
  INV_X1 U11787 ( .A(n9185), .ZN(n9186) );
  NAND2_X1 U11788 ( .A1(n9187), .A2(n9186), .ZN(n13964) );
  NAND2_X1 U11789 ( .A1(n13964), .A2(n14320), .ZN(n9189) );
  XNOR2_X1 U11790 ( .A(n9188), .B(n9189), .ZN(n13905) );
  INV_X1 U11791 ( .A(n9188), .ZN(n9190) );
  NAND2_X1 U11792 ( .A1(n9190), .A2(n9189), .ZN(n9191) );
  INV_X1 U11793 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13907) );
  INV_X1 U11794 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n14435) );
  OAI21_X1 U11795 ( .B1(n9192), .B2(n13907), .A(n14435), .ZN(n9193) );
  NAND2_X1 U11796 ( .A1(n9205), .A2(n9193), .ZN(n14197) );
  OR2_X1 U11797 ( .A1(n14197), .A2(n9464), .ZN(n9198) );
  INV_X1 U11798 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14390) );
  NAND2_X1 U11799 ( .A1(n9465), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9195) );
  NAND2_X1 U11800 ( .A1(n9245), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9194) );
  OAI211_X1 U11801 ( .C1(n9469), .C2(n14390), .A(n9195), .B(n9194), .ZN(n9196)
         );
  INV_X1 U11802 ( .A(n9196), .ZN(n9197) );
  NAND2_X1 U11803 ( .A1(n9198), .A2(n9197), .ZN(n14206) );
  NAND2_X1 U11804 ( .A1(n14206), .A2(n14320), .ZN(n9201) );
  XNOR2_X1 U11805 ( .A(n9200), .B(n9201), .ZN(n10728) );
  INV_X1 U11806 ( .A(n10728), .ZN(n9199) );
  INV_X1 U11807 ( .A(n9200), .ZN(n9203) );
  INV_X1 U11808 ( .A(n9201), .ZN(n9202) );
  XNOR2_X1 U11809 ( .A(n14180), .B(n8969), .ZN(n9213) );
  NAND2_X1 U11810 ( .A1(n9205), .A2(n13920), .ZN(n9206) );
  AND2_X1 U11811 ( .A1(n9207), .A2(n9206), .ZN(n14181) );
  NAND2_X1 U11812 ( .A1(n14181), .A2(n9258), .ZN(n9212) );
  INV_X1 U11813 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14385) );
  NAND2_X1 U11814 ( .A1(n9465), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9209) );
  NAND2_X1 U11815 ( .A1(n9245), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9208) );
  OAI211_X1 U11816 ( .C1(n9469), .C2(n14385), .A(n9209), .B(n9208), .ZN(n9210)
         );
  INV_X1 U11817 ( .A(n9210), .ZN(n9211) );
  NAND2_X1 U11818 ( .A1(n9212), .A2(n9211), .ZN(n14159) );
  AND2_X1 U11819 ( .A1(n14159), .A2(n14320), .ZN(n13917) );
  OAI211_X1 U11820 ( .C1(n13963), .C2(n13814), .A(n13811), .B(n13917), .ZN(
        n9219) );
  AND2_X1 U11821 ( .A1(n13963), .A2(n14320), .ZN(n13813) );
  OAI21_X1 U11822 ( .B1(n13813), .B2(n13814), .A(n13812), .ZN(n9217) );
  INV_X1 U11823 ( .A(n13814), .ZN(n9216) );
  INV_X1 U11824 ( .A(n13813), .ZN(n9215) );
  AND2_X1 U11825 ( .A1(n9217), .A2(n7786), .ZN(n9218) );
  NAND2_X1 U11826 ( .A1(n9219), .A2(n9218), .ZN(n13898) );
  INV_X1 U11827 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13900) );
  NAND2_X1 U11828 ( .A1(n9220), .A2(n13900), .ZN(n9221) );
  NAND2_X1 U11829 ( .A1(n9243), .A2(n9221), .ZN(n14150) );
  INV_X1 U11830 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n14375) );
  NAND2_X1 U11831 ( .A1(n8996), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9223) );
  NAND2_X1 U11832 ( .A1(n9465), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9222) );
  OAI211_X1 U11833 ( .C1(n14375), .C2(n9469), .A(n9223), .B(n9222), .ZN(n9224)
         );
  INV_X1 U11834 ( .A(n9224), .ZN(n9225) );
  NAND2_X1 U11835 ( .A1(n14160), .A2(n14320), .ZN(n9227) );
  AOI21_X1 U11836 ( .B1(n9228), .B2(n9227), .A(n9229), .ZN(n13897) );
  INV_X1 U11837 ( .A(n9229), .ZN(n9230) );
  XNOR2_X1 U11838 ( .A(n9243), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n14134) );
  NAND2_X1 U11839 ( .A1(n14134), .A2(n9258), .ZN(n9236) );
  INV_X1 U11840 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9233) );
  NAND2_X1 U11841 ( .A1(n9465), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9232) );
  NAND2_X1 U11842 ( .A1(n8996), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9231) );
  OAI211_X1 U11843 ( .C1(n9469), .C2(n9233), .A(n9232), .B(n9231), .ZN(n9234)
         );
  INV_X1 U11844 ( .A(n9234), .ZN(n9235) );
  NAND2_X1 U11845 ( .A1(n13962), .A2(n14320), .ZN(n9237) );
  AOI21_X1 U11846 ( .B1(n9238), .B2(n9237), .A(n9239), .ZN(n13868) );
  INV_X1 U11847 ( .A(n9239), .ZN(n9240) );
  NAND2_X1 U11848 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n9241) );
  INV_X1 U11849 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13870) );
  INV_X1 U11850 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9242) );
  OAI21_X1 U11851 ( .B1(n9243), .B2(n13870), .A(n9242), .ZN(n9244) );
  INV_X1 U11852 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9248) );
  NAND2_X1 U11853 ( .A1(n9245), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9247) );
  NAND2_X1 U11854 ( .A1(n9259), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9246) );
  OAI211_X1 U11855 ( .C1(n8984), .C2(n9248), .A(n9247), .B(n9246), .ZN(n9249)
         );
  INV_X1 U11856 ( .A(n9249), .ZN(n9250) );
  NAND2_X1 U11857 ( .A1(n14125), .A2(n14320), .ZN(n9252) );
  XOR2_X1 U11858 ( .A(n9252), .B(n9251), .Z(n13936) );
  INV_X1 U11859 ( .A(n9251), .ZN(n9253) );
  INV_X1 U11860 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9255) );
  NAND2_X1 U11861 ( .A1(n9256), .A2(n9255), .ZN(n9257) );
  NAND2_X1 U11862 ( .A1(n14097), .A2(n9258), .ZN(n9265) );
  INV_X1 U11863 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n14444) );
  NAND2_X1 U11864 ( .A1(n9259), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9261) );
  NAND2_X1 U11865 ( .A1(n9465), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9260) );
  OAI211_X1 U11866 ( .C1(n9262), .C2(n14444), .A(n9261), .B(n9260), .ZN(n9263)
         );
  INV_X1 U11867 ( .A(n9263), .ZN(n9264) );
  NAND2_X1 U11868 ( .A1(n13961), .A2(n14320), .ZN(n9266) );
  NOR2_X1 U11869 ( .A1(n9267), .A2(n9266), .ZN(n13844) );
  AOI21_X1 U11870 ( .B1(n9267), .B2(n9266), .A(n13844), .ZN(n9270) );
  OR2_X1 U11871 ( .A1(n9268), .A2(n15644), .ZN(n10449) );
  NOR2_X1 U11872 ( .A1(n10449), .A2(n15641), .ZN(n9289) );
  AND2_X1 U11873 ( .A1(n9289), .A2(n15645), .ZN(n9277) );
  AND2_X1 U11874 ( .A1(n15648), .A2(n11044), .ZN(n9269) );
  NAND2_X1 U11875 ( .A1(n9272), .A2(n9271), .ZN(n9273) );
  INV_X1 U11876 ( .A(n9274), .ZN(n11595) );
  NOR2_X1 U11877 ( .A1(n11595), .A2(n11815), .ZN(n10462) );
  NAND2_X1 U11878 ( .A1(n9277), .A2(n10462), .ZN(n9276) );
  INV_X1 U11879 ( .A(n9290), .ZN(n9275) );
  NAND2_X1 U11880 ( .A1(n9276), .A2(n15619), .ZN(n13954) );
  INV_X1 U11881 ( .A(n13954), .ZN(n13925) );
  INV_X1 U11882 ( .A(n9539), .ZN(n9507) );
  NAND2_X1 U11883 ( .A1(n9277), .A2(n9507), .ZN(n13891) );
  OR2_X1 U11884 ( .A1(n13891), .A2(n14192), .ZN(n13908) );
  INV_X1 U11885 ( .A(n13908), .ZN(n13937) );
  INV_X1 U11886 ( .A(n9280), .ZN(n9278) );
  NAND2_X1 U11887 ( .A1(n9278), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n10464) );
  INV_X1 U11888 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9279) );
  NAND2_X1 U11889 ( .A1(n9280), .A2(n9279), .ZN(n9281) );
  NAND2_X1 U11890 ( .A1(n10464), .A2(n9281), .ZN(n13845) );
  INV_X1 U11891 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10438) );
  NAND2_X1 U11892 ( .A1(n8996), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9283) );
  NAND2_X1 U11893 ( .A1(n9465), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9282) );
  OAI211_X1 U11894 ( .C1(n10438), .C2(n9469), .A(n9283), .B(n9282), .ZN(n9284)
         );
  INV_X1 U11895 ( .A(n9284), .ZN(n9285) );
  INV_X1 U11896 ( .A(n14125), .ZN(n13871) );
  INV_X1 U11897 ( .A(n13891), .ZN(n13949) );
  INV_X1 U11898 ( .A(n8885), .ZN(n9287) );
  NAND2_X1 U11899 ( .A1(n13949), .A2(n14285), .ZN(n13941) );
  INV_X1 U11900 ( .A(n9289), .ZN(n9291) );
  NAND2_X1 U11901 ( .A1(n9291), .A2(n9290), .ZN(n9292) );
  NAND2_X1 U11902 ( .A1(n9292), .A2(n10439), .ZN(n11477) );
  INV_X1 U11903 ( .A(n9293), .ZN(n9294) );
  OR2_X1 U11904 ( .A1(n11477), .A2(n9294), .ZN(n9295) );
  AOI22_X1 U11905 ( .A1(n14097), .A2(n13938), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9296) );
  OAI21_X1 U11906 ( .B1(n13871), .B2(n13941), .A(n9296), .ZN(n9297) );
  AOI21_X1 U11907 ( .B1(n13937), .B2(n14093), .A(n9297), .ZN(n9298) );
  OR2_X1 U11908 ( .A1(n12933), .A2(n13542), .ZN(n9301) );
  AND2_X1 U11909 ( .A1(n14645), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9303) );
  XNOR2_X1 U11910 ( .A(n12891), .B(P1_DATAO_REG_28__SCAN_IN), .ZN(n9305) );
  NAND2_X1 U11911 ( .A1(n12983), .A2(SI_28_), .ZN(n9306) );
  NAND2_X1 U11912 ( .A1(n9309), .A2(n9308), .ZN(n13169) );
  AND2_X1 U11913 ( .A1(n12891), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9310) );
  NAND2_X1 U11914 ( .A1(n9312), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9313) );
  XNOR2_X1 U11915 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .ZN(n12871) );
  XNOR2_X1 U11916 ( .A(n12874), .B(n12871), .ZN(n12892) );
  NAND2_X1 U11917 ( .A1(n12892), .A2(n12988), .ZN(n9316) );
  NAND2_X1 U11918 ( .A1(n12983), .A2(SI_29_), .ZN(n9315) );
  INV_X1 U11919 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9322) );
  NAND2_X1 U11920 ( .A1(n8179), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9320) );
  NAND2_X1 U11921 ( .A1(n9327), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9319) );
  OAI211_X1 U11922 ( .C1(n9322), .C2(n9321), .A(n9320), .B(n9319), .ZN(n9323)
         );
  INV_X1 U11923 ( .A(n9323), .ZN(n9324) );
  XNOR2_X1 U11924 ( .A(n9325), .B(n13028), .ZN(n9326) );
  NAND2_X1 U11925 ( .A1(n9326), .A2(n13728), .ZN(n9336) );
  INV_X1 U11926 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n9331) );
  NAND2_X1 U11927 ( .A1(n9327), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9330) );
  NAND2_X1 U11928 ( .A1(n12875), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9329) );
  OAI211_X1 U11929 ( .C1(n12880), .C2(n9331), .A(n9330), .B(n9329), .ZN(n9332)
         );
  INV_X1 U11930 ( .A(n9332), .ZN(n9333) );
  NAND2_X1 U11931 ( .A1(n12883), .A2(n9333), .ZN(n13369) );
  NAND2_X1 U11932 ( .A1(n13800), .A2(P3_B_REG_SCAN_IN), .ZN(n9334) );
  AND2_X1 U11933 ( .A1(n13722), .A2(n9334), .ZN(n12884) );
  AOI22_X1 U11934 ( .A1(n13724), .A2(n13370), .B1(n13369), .B2(n12884), .ZN(
        n9335) );
  NAND2_X1 U11935 ( .A1(n9336), .A2(n9335), .ZN(n9560) );
  OR2_X1 U11936 ( .A1(n9557), .A2(n15715), .ZN(n11190) );
  NOR2_X1 U11937 ( .A1(n11190), .A2(n15683), .ZN(n11412) );
  NAND2_X1 U11938 ( .A1(n13796), .A2(n9337), .ZN(n9342) );
  INV_X1 U11939 ( .A(n9337), .ZN(n9339) );
  NAND2_X1 U11940 ( .A1(n9339), .A2(n9338), .ZN(n9341) );
  AOI21_X1 U11941 ( .B1(n9342), .B2(n9341), .A(n9340), .ZN(n9343) );
  NAND2_X1 U11942 ( .A1(n9344), .A2(n9343), .ZN(n9349) );
  AND2_X2 U11943 ( .A1(n13645), .A2(n9349), .ZN(n15691) );
  AOI21_X1 U11944 ( .B1(n9560), .B2(n9345), .A(n6617), .ZN(n9352) );
  INV_X1 U11945 ( .A(n13542), .ZN(n12939) );
  NAND2_X1 U11946 ( .A1(n12933), .A2(n12939), .ZN(n13167) );
  NAND2_X1 U11947 ( .A1(n9347), .A2(n13171), .ZN(n12981) );
  NOR2_X1 U11948 ( .A1(n13059), .A2(n15683), .ZN(n11695) );
  NOR2_X1 U11949 ( .A1(n13718), .A2(n11695), .ZN(n9348) );
  INV_X1 U11950 ( .A(n13663), .ZN(n13563) );
  INV_X1 U11951 ( .A(n12994), .ZN(n9565) );
  OR2_X1 U11952 ( .A1(n9349), .A2(n15674), .ZN(n11989) );
  NAND2_X1 U11953 ( .A1(n9350), .A2(n15685), .ZN(n12887) );
  OAI21_X1 U11954 ( .B1(n9565), .B2(n13588), .A(n12887), .ZN(n9351) );
  INV_X1 U11955 ( .A(n9401), .ZN(n9476) );
  MUX2_X1 U11956 ( .A(n13977), .B(n15657), .S(n9497), .Z(n9372) );
  INV_X1 U11957 ( .A(n13978), .ZN(n11982) );
  AOI21_X1 U11958 ( .B1(n13978), .B2(n9473), .A(n13827), .ZN(n9369) );
  NOR2_X1 U11959 ( .A1(n9513), .A2(n9478), .ZN(n9356) );
  INV_X1 U11960 ( .A(n10377), .ZN(n9357) );
  OR2_X1 U11961 ( .A1(n9357), .A2(n11485), .ZN(n9358) );
  NAND2_X1 U11962 ( .A1(n9358), .A2(n9401), .ZN(n9360) );
  INV_X1 U11963 ( .A(n9360), .ZN(n9359) );
  NOR2_X1 U11964 ( .A1(n9353), .A2(n9360), .ZN(n9362) );
  XNOR2_X1 U11965 ( .A(n9514), .B(n11979), .ZN(n9364) );
  INV_X1 U11966 ( .A(n9514), .ZN(n9515) );
  NAND3_X1 U11967 ( .A1(n9515), .A2(n9478), .A3(n11979), .ZN(n9366) );
  NAND3_X1 U11968 ( .A1(n9514), .A2(n15649), .A3(n9476), .ZN(n9365) );
  NAND2_X1 U11969 ( .A1(n9366), .A2(n9365), .ZN(n9367) );
  MUX2_X1 U11970 ( .A(n15657), .B(n13977), .S(n9497), .Z(n9371) );
  AND2_X1 U11971 ( .A1(n13976), .A2(n9473), .ZN(n9374) );
  OAI21_X1 U11972 ( .B1(n13976), .B2(n9476), .A(n11914), .ZN(n9373) );
  OAI21_X1 U11973 ( .B1(n9374), .B2(n11914), .A(n9373), .ZN(n9375) );
  XNOR2_X1 U11974 ( .A(n13975), .B(n12064), .ZN(n10390) );
  OAI21_X1 U11975 ( .B1(n13975), .B2(n9478), .A(n12064), .ZN(n9379) );
  NAND2_X1 U11976 ( .A1(n13975), .A2(n9478), .ZN(n9377) );
  NAND2_X1 U11977 ( .A1(n12104), .A2(n9377), .ZN(n9378) );
  NAND2_X1 U11978 ( .A1(n9379), .A2(n9378), .ZN(n9380) );
  MUX2_X1 U11979 ( .A(n13974), .B(n15624), .S(n9473), .Z(n9382) );
  XNOR2_X1 U11980 ( .A(n12445), .B(n13973), .ZN(n12371) );
  OAI21_X1 U11981 ( .B1(n9383), .B2(n9382), .A(n12371), .ZN(n9385) );
  MUX2_X1 U11982 ( .A(n12372), .B(n12375), .S(n9497), .Z(n9381) );
  AND2_X1 U11983 ( .A1(n13973), .A2(n9478), .ZN(n9387) );
  OAI21_X1 U11984 ( .B1(n9478), .B2(n13973), .A(n12445), .ZN(n9386) );
  OAI21_X1 U11985 ( .B1(n9387), .B2(n12445), .A(n9386), .ZN(n9388) );
  MUX2_X1 U11986 ( .A(n13971), .B(n12409), .S(n9473), .Z(n9391) );
  MUX2_X1 U11987 ( .A(n13971), .B(n12409), .S(n9497), .Z(n9389) );
  INV_X1 U11988 ( .A(n9391), .ZN(n9392) );
  AND2_X1 U11989 ( .A1(n14329), .A2(n9478), .ZN(n9394) );
  OAI21_X1 U11990 ( .B1(n9478), .B2(n14329), .A(n12735), .ZN(n9393) );
  OAI21_X1 U11991 ( .B1(n9394), .B2(n12735), .A(n9393), .ZN(n9395) );
  MUX2_X1 U11992 ( .A(n13970), .B(n14571), .S(n9473), .Z(n9397) );
  XNOR2_X1 U11993 ( .A(n12609), .B(n13969), .ZN(n9522) );
  INV_X1 U11994 ( .A(n13970), .ZN(n10398) );
  MUX2_X1 U11995 ( .A(n10398), .B(n14327), .S(n9497), .Z(n9396) );
  AND2_X1 U11996 ( .A1(n13969), .A2(n9497), .ZN(n9399) );
  OAI21_X1 U11997 ( .B1(n9478), .B2(n13969), .A(n12609), .ZN(n9398) );
  OAI21_X1 U11998 ( .B1(n9399), .B2(n12609), .A(n9398), .ZN(n9400) );
  MUX2_X1 U11999 ( .A(n13968), .B(n12678), .S(n9473), .Z(n9403) );
  MUX2_X1 U12000 ( .A(n13968), .B(n12678), .S(n9497), .Z(n9402) );
  MUX2_X1 U12001 ( .A(n13967), .B(n14562), .S(n9497), .Z(n9413) );
  MUX2_X1 U12002 ( .A(n14287), .B(n14275), .S(n9473), .Z(n9418) );
  NAND2_X1 U12003 ( .A1(n14275), .A2(n14287), .ZN(n9404) );
  NAND2_X1 U12004 ( .A1(n9418), .A2(n9404), .ZN(n9408) );
  AND2_X1 U12005 ( .A1(n13966), .A2(n9497), .ZN(n9406) );
  OAI21_X1 U12006 ( .B1(n9478), .B2(n13966), .A(n14546), .ZN(n9405) );
  OAI21_X1 U12007 ( .B1(n9406), .B2(n14546), .A(n9405), .ZN(n9407) );
  NAND2_X1 U12008 ( .A1(n9408), .A2(n9407), .ZN(n9415) );
  INV_X1 U12009 ( .A(n14284), .ZN(n13882) );
  MUX2_X1 U12010 ( .A(n13882), .B(n14617), .S(n9497), .Z(n9417) );
  MUX2_X1 U12011 ( .A(n14284), .B(n14313), .S(n9473), .Z(n9416) );
  AND2_X1 U12012 ( .A1(n9417), .A2(n9416), .ZN(n9409) );
  NOR2_X1 U12013 ( .A1(n9415), .A2(n9409), .ZN(n9410) );
  OAI21_X1 U12014 ( .B1(n9414), .B2(n9413), .A(n9410), .ZN(n9424) );
  MUX2_X1 U12015 ( .A(n13967), .B(n14562), .S(n9473), .Z(n9411) );
  INV_X1 U12016 ( .A(n9415), .ZN(n9421) );
  XNOR2_X1 U12017 ( .A(n14546), .B(n13966), .ZN(n9523) );
  OAI21_X1 U12018 ( .B1(n9417), .B2(n9416), .A(n9523), .ZN(n9420) );
  NOR2_X1 U12019 ( .A1(n14275), .A2(n14287), .ZN(n14261) );
  NOR2_X1 U12020 ( .A1(n9418), .A2(n14261), .ZN(n9419) );
  AOI21_X1 U12021 ( .B1(n9421), .B2(n9420), .A(n9419), .ZN(n9422) );
  MUX2_X1 U12022 ( .A(n13965), .B(n14537), .S(n9497), .Z(n9427) );
  MUX2_X1 U12023 ( .A(n13965), .B(n14537), .S(n9473), .Z(n9425) );
  MUX2_X1 U12024 ( .A(n14207), .B(n14232), .S(n9473), .Z(n9429) );
  MUX2_X1 U12025 ( .A(n14207), .B(n14232), .S(n9497), .Z(n9428) );
  MUX2_X1 U12026 ( .A(n13964), .B(n14393), .S(n9497), .Z(n9432) );
  MUX2_X1 U12027 ( .A(n13964), .B(n14393), .S(n9473), .Z(n9431) );
  MUX2_X1 U12028 ( .A(n14206), .B(n14196), .S(n9473), .Z(n9436) );
  MUX2_X1 U12029 ( .A(n14206), .B(n14196), .S(n9478), .Z(n9433) );
  NAND2_X1 U12030 ( .A1(n9434), .A2(n9433), .ZN(n9440) );
  INV_X1 U12031 ( .A(n9435), .ZN(n9438) );
  INV_X1 U12032 ( .A(n9436), .ZN(n9437) );
  NAND2_X1 U12033 ( .A1(n9438), .A2(n9437), .ZN(n9439) );
  MUX2_X1 U12034 ( .A(n14159), .B(n14180), .S(n9478), .Z(n9442) );
  MUX2_X1 U12035 ( .A(n14159), .B(n14180), .S(n9473), .Z(n9441) );
  INV_X1 U12036 ( .A(n9442), .ZN(n9443) );
  MUX2_X1 U12037 ( .A(n13963), .B(n14378), .S(n9473), .Z(n9445) );
  MUX2_X1 U12038 ( .A(n13963), .B(n14378), .S(n9478), .Z(n9444) );
  MUX2_X1 U12039 ( .A(n14160), .B(n14149), .S(n9478), .Z(n9450) );
  MUX2_X1 U12040 ( .A(n14160), .B(n14149), .S(n9473), .Z(n9447) );
  MUX2_X1 U12041 ( .A(n13962), .B(n14135), .S(n9473), .Z(n9452) );
  MUX2_X1 U12042 ( .A(n13962), .B(n14135), .S(n9478), .Z(n9451) );
  MUX2_X1 U12043 ( .A(n13871), .B(n7629), .S(n9478), .Z(n9454) );
  MUX2_X1 U12044 ( .A(n14113), .B(n14125), .S(n9478), .Z(n9453) );
  NAND2_X1 U12045 ( .A1(n9455), .A2(n9454), .ZN(n9456) );
  NAND2_X1 U12046 ( .A1(n9457), .A2(n9456), .ZN(n9503) );
  MUX2_X1 U12047 ( .A(n13961), .B(n14356), .S(n9473), .Z(n9491) );
  INV_X1 U12048 ( .A(n9491), .ZN(n9480) );
  INV_X1 U12049 ( .A(n13961), .ZN(n14110) );
  MUX2_X1 U12050 ( .A(n14110), .B(n14099), .S(n9478), .Z(n9492) );
  INV_X1 U12051 ( .A(n9492), .ZN(n9479) );
  INV_X1 U12052 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14349) );
  NAND2_X1 U12053 ( .A1(n8996), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9460) );
  INV_X1 U12054 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n9458) );
  OR2_X1 U12055 ( .A1(n8984), .A2(n9458), .ZN(n9459) );
  OAI211_X1 U12056 ( .C1(n9469), .C2(n14349), .A(n9460), .B(n9459), .ZN(n13959) );
  MUX2_X1 U12057 ( .A(n13959), .B(n14081), .S(n9478), .Z(n9484) );
  NAND2_X1 U12058 ( .A1(n13958), .A2(n9478), .ZN(n9461) );
  NAND2_X1 U12059 ( .A1(n10430), .A2(n11596), .ZN(n9504) );
  NAND4_X1 U12060 ( .A1(n9461), .A2(n10453), .A3(n9539), .A4(n9504), .ZN(n9462) );
  AND2_X1 U12061 ( .A1(n9462), .A2(n13959), .ZN(n9463) );
  AOI21_X1 U12062 ( .B1(n14081), .B2(n9476), .A(n9463), .ZN(n9483) );
  OR2_X1 U12063 ( .A1(n10464), .A2(n9464), .ZN(n9472) );
  INV_X1 U12064 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9468) );
  NAND2_X1 U12065 ( .A1(n9465), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9467) );
  NAND2_X1 U12066 ( .A1(n8996), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9466) );
  OAI211_X1 U12067 ( .C1(n9469), .C2(n9468), .A(n9467), .B(n9466), .ZN(n9470)
         );
  INV_X1 U12068 ( .A(n9470), .ZN(n9471) );
  NAND2_X1 U12069 ( .A1(n9472), .A2(n9471), .ZN(n13960) );
  INV_X1 U12070 ( .A(n14093), .ZN(n9477) );
  MUX2_X1 U12071 ( .A(n9477), .B(n7609), .S(n9476), .Z(n9486) );
  MUX2_X1 U12072 ( .A(n14093), .B(n14087), .S(n9478), .Z(n9485) );
  OAI22_X1 U12073 ( .A1(n9484), .A2(n9483), .B1(n9482), .B2(n9481), .ZN(n9489)
         );
  INV_X1 U12074 ( .A(n9490), .ZN(n9493) );
  NAND3_X1 U12075 ( .A1(n9493), .A2(n9492), .A3(n9491), .ZN(n9495) );
  AOI21_X1 U12076 ( .B1(n9496), .B2(n9495), .A(n9494), .ZN(n9500) );
  AND2_X1 U12077 ( .A1(n14077), .A2(n13958), .ZN(n9499) );
  NOR2_X1 U12078 ( .A1(n14077), .A2(n13958), .ZN(n9498) );
  NAND2_X1 U12079 ( .A1(n10453), .A2(n14070), .ZN(n9505) );
  OAI21_X1 U12080 ( .B1(n9505), .B2(n11815), .A(n9504), .ZN(n9506) );
  INV_X1 U12081 ( .A(n9506), .ZN(n9511) );
  AOI21_X1 U12082 ( .B1(n10453), .B2(n11455), .A(n9507), .ZN(n9508) );
  OAI21_X1 U12083 ( .B1(n10430), .B2(n10377), .A(n9508), .ZN(n9509) );
  NAND2_X1 U12084 ( .A1(n9535), .A2(n9509), .ZN(n9510) );
  OAI21_X1 U12085 ( .B1(n9535), .B2(n9511), .A(n9510), .ZN(n9538) );
  NAND2_X1 U12086 ( .A1(n14087), .A2(n14093), .ZN(n10444) );
  INV_X1 U12087 ( .A(n14111), .ZN(n14106) );
  XNOR2_X1 U12088 ( .A(n14135), .B(n13962), .ZN(n14130) );
  INV_X1 U12089 ( .A(n14206), .ZN(n13918) );
  OR2_X1 U12090 ( .A1(n14196), .A2(n13918), .ZN(n10420) );
  NAND2_X1 U12091 ( .A1(n14196), .A2(n13918), .ZN(n10421) );
  NAND2_X1 U12092 ( .A1(n10420), .A2(n10421), .ZN(n14193) );
  INV_X1 U12093 ( .A(n13964), .ZN(n14189) );
  XNOR2_X1 U12094 ( .A(n14393), .B(n14189), .ZN(n14217) );
  INV_X1 U12095 ( .A(n11911), .ZN(n11908) );
  NAND2_X1 U12096 ( .A1(n9513), .A2(n10747), .ZN(n11622) );
  NAND2_X1 U12097 ( .A1(n9514), .A2(n15649), .ZN(n9516) );
  NAND2_X1 U12098 ( .A1(n9515), .A2(n11979), .ZN(n10385) );
  NOR4_X1 U12099 ( .A1(n11622), .A2(n11815), .A3(n10331), .A4(n10755), .ZN(
        n9517) );
  XNOR2_X1 U12100 ( .A(n13977), .B(n15657), .ZN(n11931) );
  NAND4_X1 U12101 ( .A1(n9517), .A2(n11710), .A3(n10390), .A4(n11931), .ZN(
        n9518) );
  INV_X1 U12102 ( .A(n12371), .ZN(n12377) );
  XNOR2_X1 U12103 ( .A(n15624), .B(n12372), .ZN(n12248) );
  NOR4_X1 U12104 ( .A1(n11908), .A2(n9518), .A3(n12377), .A4(n12248), .ZN(
        n9519) );
  XNOR2_X1 U12105 ( .A(n14571), .B(n13970), .ZN(n14336) );
  XNOR2_X1 U12106 ( .A(n12409), .B(n13971), .ZN(n12402) );
  AND4_X1 U12107 ( .A1(n9519), .A2(n12724), .A3(n14336), .A4(n12402), .ZN(
        n9521) );
  INV_X1 U12108 ( .A(n13968), .ZN(n12816) );
  NAND2_X1 U12109 ( .A1(n12678), .A2(n12816), .ZN(n10409) );
  OR2_X1 U12110 ( .A1(n12678), .A2(n12816), .ZN(n9520) );
  NAND2_X1 U12111 ( .A1(n10409), .A2(n9520), .ZN(n12672) );
  INV_X1 U12112 ( .A(n12672), .ZN(n12669) );
  XNOR2_X1 U12113 ( .A(n14313), .B(n14284), .ZN(n14305) );
  NAND3_X1 U12114 ( .A1(n9521), .A2(n12669), .A3(n14305), .ZN(n9524) );
  XNOR2_X1 U12115 ( .A(n14562), .B(n12675), .ZN(n12813) );
  NOR4_X1 U12116 ( .A1(n9524), .A2(n12573), .A3(n12813), .A4(n14289), .ZN(
        n9525) );
  INV_X1 U12117 ( .A(n14207), .ZN(n13929) );
  XNOR2_X1 U12118 ( .A(n14232), .B(n13929), .ZN(n14224) );
  INV_X1 U12119 ( .A(n14224), .ZN(n14229) );
  INV_X1 U12120 ( .A(n13965), .ZN(n13836) );
  XNOR2_X1 U12121 ( .A(n14537), .B(n13836), .ZN(n14260) );
  INV_X1 U12122 ( .A(n14260), .ZN(n14247) );
  XNOR2_X1 U12123 ( .A(n14275), .B(n14287), .ZN(n10413) );
  NAND4_X1 U12124 ( .A1(n9525), .A2(n14229), .A3(n14247), .A4(n10413), .ZN(
        n9526) );
  NOR4_X1 U12125 ( .A1(n14177), .A2(n14193), .A3(n14217), .A4(n9526), .ZN(
        n9527) );
  INV_X1 U12126 ( .A(n13963), .ZN(n13919) );
  XNOR2_X1 U12127 ( .A(n14378), .B(n13919), .ZN(n14157) );
  NAND4_X1 U12128 ( .A1(n14130), .A2(n9527), .A3(n14143), .A4(n7571), .ZN(
        n9528) );
  NOR4_X1 U12129 ( .A1(n10375), .A2(n10373), .A3(n14106), .A4(n9528), .ZN(
        n9530) );
  XOR2_X1 U12130 ( .A(n13959), .B(n14585), .Z(n9529) );
  NAND4_X1 U12131 ( .A1(n9531), .A2(n9530), .A3(n9529), .A4(n10456), .ZN(n9532) );
  AOI21_X1 U12132 ( .B1(n9535), .B2(n11596), .A(n9534), .ZN(n9537) );
  OR2_X1 U12133 ( .A1(n10706), .A2(P2_U3088), .ZN(n12041) );
  INV_X1 U12134 ( .A(n12041), .ZN(n9536) );
  OAI21_X1 U12135 ( .B1(n9538), .B2(n9537), .A(n9536), .ZN(n9543) );
  INV_X1 U12136 ( .A(n15645), .ZN(n15642) );
  INV_X1 U12137 ( .A(n14285), .ZN(n14190) );
  NOR4_X1 U12138 ( .A1(n15642), .A2(n14190), .A3(n9539), .A4(n14647), .ZN(
        n9541) );
  OAI21_X1 U12139 ( .B1(n10430), .B2(n12041), .A(P2_B_REG_SCAN_IN), .ZN(n9540)
         );
  NAND2_X1 U12140 ( .A1(n9543), .A2(n9542), .ZN(P2_U3328) );
  OR2_X1 U12141 ( .A1(n9560), .A2(n15731), .ZN(n9545) );
  NAND2_X1 U12142 ( .A1(n9545), .A2(n9544), .ZN(n9548) );
  NOR2_X1 U12143 ( .A1(n13718), .A2(n15720), .ZN(n9564) );
  INV_X1 U12144 ( .A(n9564), .ZN(n13676) );
  NAND2_X1 U12145 ( .A1(n15734), .A2(n13676), .ZN(n13715) );
  OAI22_X1 U12146 ( .A1(n9566), .A2(n13715), .B1(n9565), .B2(n13709), .ZN(
        n9546) );
  INV_X1 U12147 ( .A(n9546), .ZN(n9547) );
  NAND2_X1 U12148 ( .A1(n9548), .A2(n9547), .ZN(P3_U3488) );
  NOR2_X1 U12149 ( .A1(n9549), .A2(n9555), .ZN(n11189) );
  NAND2_X1 U12150 ( .A1(n13168), .A2(n9550), .ZN(n11384) );
  NOR2_X1 U12151 ( .A1(n9557), .A2(n11384), .ZN(n13189) );
  INV_X1 U12152 ( .A(n9551), .ZN(n9553) );
  NAND2_X1 U12153 ( .A1(n13059), .A2(n9552), .ZN(n13186) );
  NAND2_X1 U12154 ( .A1(n9553), .A2(n7172), .ZN(n11172) );
  NOR2_X1 U12155 ( .A1(n9557), .A2(n11172), .ZN(n11184) );
  OR2_X1 U12156 ( .A1(n13189), .A2(n11184), .ZN(n9554) );
  NAND2_X1 U12157 ( .A1(n11189), .A2(n9554), .ZN(n9559) );
  NOR2_X1 U12158 ( .A1(n9556), .A2(n9555), .ZN(n11185) );
  INV_X1 U12159 ( .A(n9557), .ZN(n11183) );
  NAND3_X1 U12160 ( .A1(n11185), .A2(n11183), .A3(n11182), .ZN(n9558) );
  AND2_X2 U12161 ( .A1(n9559), .A2(n9558), .ZN(n15721) );
  OR2_X1 U12162 ( .A1(n9560), .A2(n15721), .ZN(n9563) );
  INV_X1 U12163 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9561) );
  NAND2_X1 U12164 ( .A1(n15721), .A2(n9561), .ZN(n9562) );
  NAND2_X1 U12165 ( .A1(n9563), .A2(n9562), .ZN(n9569) );
  OAI22_X1 U12166 ( .A1(n9566), .A2(n13793), .B1(n9565), .B2(n13790), .ZN(
        n9567) );
  INV_X1 U12167 ( .A(n9567), .ZN(n9568) );
  NAND2_X1 U12168 ( .A1(n9569), .A2(n9568), .ZN(P3_U3456) );
  NAND4_X1 U12169 ( .A1(n9571), .A2(n9841), .A3(n9839), .A4(n9570), .ZN(n9844)
         );
  NAND2_X1 U12170 ( .A1(n9980), .A2(n9572), .ZN(n9573) );
  NOR2_X1 U12171 ( .A1(n9844), .A2(n9573), .ZN(n9579) );
  NOR2_X1 U12172 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .ZN(n9576) );
  NAND4_X1 U12173 ( .A1(n9576), .A2(n9575), .A3(n9574), .A4(n9769), .ZN(n9578)
         );
  NAND4_X1 U12174 ( .A1(n9727), .A2(n9766), .A3(n9699), .A4(n9656), .ZN(n9577)
         );
  NOR2_X2 U12175 ( .A1(n9578), .A2(n9577), .ZN(n9791) );
  INV_X2 U12176 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n15490) );
  NOR2_X1 U12177 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n9583) );
  NOR2_X1 U12178 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n9582) );
  NAND3_X1 U12179 ( .A1(n9583), .A2(n9582), .A3(n9581), .ZN(n9584) );
  INV_X1 U12180 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9588) );
  INV_X1 U12181 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11891) );
  OR2_X1 U12182 ( .A1(n6429), .A2(n11891), .ZN(n9594) );
  AND2_X2 U12183 ( .A1(n13214), .A2(n9589), .ZN(n9660) );
  INV_X1 U12184 ( .A(n9660), .ZN(n9646) );
  INV_X1 U12185 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10087) );
  OR2_X1 U12186 ( .A1(n9646), .A2(n10087), .ZN(n9593) );
  INV_X1 U12187 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9591) );
  OR2_X1 U12188 ( .A1(n9614), .A2(n9591), .ZN(n9592) );
  INV_X1 U12189 ( .A(SI_0_), .ZN(n9597) );
  OAI21_X1 U12190 ( .B1(n10817), .B2(n9597), .A(n9596), .ZN(n9598) );
  AND2_X1 U12191 ( .A1(n9599), .A2(n9598), .ZN(n15439) );
  INV_X1 U12192 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9604) );
  MUX2_X1 U12193 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15439), .S(n9632), .Z(n11128)
         );
  NAND2_X1 U12194 ( .A1(n11156), .A2(n11128), .ZN(n10483) );
  INV_X1 U12195 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14822) );
  NAND2_X1 U12196 ( .A1(n9660), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9607) );
  INV_X1 U12197 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11501) );
  INV_X1 U12198 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9609) );
  NAND2_X1 U12199 ( .A1(n9632), .A2(n6978), .ZN(n9619) );
  INV_X1 U12200 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9611) );
  INV_X1 U12201 ( .A(n11498), .ZN(n11166) );
  NAND2_X1 U12202 ( .A1(n9991), .A2(n11166), .ZN(n10487) );
  BUF_X4 U12203 ( .A(n9660), .Z(n10612) );
  INV_X1 U12204 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11675) );
  OR2_X1 U12205 ( .A1(n6429), .A2(n11675), .ZN(n9617) );
  INV_X1 U12206 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9613) );
  INV_X1 U12207 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10936) );
  NAND4_X4 U12208 ( .A1(n9618), .A2(n9617), .A3(n9616), .A4(n9615), .ZN(n14820) );
  NAND2_X1 U12209 ( .A1(n9654), .A2(n9620), .ZN(n9627) );
  NAND2_X1 U12210 ( .A1(n9622), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9621) );
  MUX2_X1 U12211 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9621), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n9625) );
  INV_X1 U12212 ( .A(n9622), .ZN(n9624) );
  INV_X1 U12213 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9623) );
  NAND2_X1 U12214 ( .A1(n9624), .A2(n9623), .ZN(n9643) );
  NAND2_X1 U12215 ( .A1(n9625), .A2(n9643), .ZN(n14843) );
  OR2_X1 U12216 ( .A1(n9632), .A2(n14843), .ZN(n9626) );
  XNOR2_X2 U12217 ( .A(n14820), .B(n11259), .ZN(n11255) );
  NAND2_X1 U12218 ( .A1(n11254), .A2(n11255), .ZN(n9630) );
  INV_X1 U12219 ( .A(n14820), .ZN(n11159) );
  NAND2_X1 U12220 ( .A1(n11159), .A2(n11259), .ZN(n9629) );
  NAND2_X1 U12221 ( .A1(n9630), .A2(n9629), .ZN(n11320) );
  NAND2_X1 U12222 ( .A1(n10789), .A2(n9654), .ZN(n9637) );
  OR2_X1 U12223 ( .A1(n9631), .A2(n10790), .ZN(n9636) );
  NAND2_X1 U12224 ( .A1(n9643), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9634) );
  OR2_X1 U12225 ( .A1(n9632), .A2(n14863), .ZN(n9635) );
  NAND2_X1 U12226 ( .A1(n9929), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9641) );
  INV_X1 U12227 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10917) );
  OR2_X1 U12228 ( .A1(n9646), .A2(n10917), .ZN(n9640) );
  INV_X1 U12229 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10939) );
  OR2_X1 U12230 ( .A1(n9614), .A2(n10939), .ZN(n9639) );
  OR2_X1 U12231 ( .A1(n6429), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9638) );
  NAND2_X1 U12232 ( .A1(n11320), .A2(n11321), .ZN(n9642) );
  NAND2_X1 U12233 ( .A1(n9995), .A2(n15523), .ZN(n10475) );
  NAND2_X1 U12234 ( .A1(n9642), .A2(n10475), .ZN(n11511) );
  NAND2_X1 U12235 ( .A1(n10794), .A2(n9902), .ZN(n9645) );
  OAI21_X1 U12236 ( .B1(n9643), .B2(P1_IR_REG_3__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9644) );
  NAND2_X1 U12237 ( .A1(n9929), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9650) );
  INV_X1 U12238 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10918) );
  OR2_X1 U12239 ( .A1(n9646), .A2(n10918), .ZN(n9649) );
  XNOR2_X1 U12240 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n11834) );
  OR2_X1 U12241 ( .A1(n6429), .A2(n11834), .ZN(n9648) );
  INV_X1 U12242 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11563) );
  OR2_X1 U12243 ( .A1(n9614), .A2(n11563), .ZN(n9647) );
  INV_X1 U12244 ( .A(n14818), .ZN(n11865) );
  NAND2_X1 U12245 ( .A1(n11830), .A2(n14818), .ZN(n9651) );
  NAND2_X1 U12246 ( .A1(n11761), .A2(n9651), .ZN(n10651) );
  NAND2_X1 U12247 ( .A1(n11511), .A2(n10651), .ZN(n9653) );
  NAND2_X1 U12248 ( .A1(n11865), .A2(n11830), .ZN(n9652) );
  NAND2_X1 U12249 ( .A1(n9653), .A2(n9652), .ZN(n11760) );
  NAND2_X1 U12250 ( .A1(n10787), .A2(n9902), .ZN(n9659) );
  NAND2_X1 U12251 ( .A1(n9974), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9655) );
  MUX2_X1 U12252 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9655), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n9657) );
  NAND2_X1 U12253 ( .A1(n9792), .A2(n9656), .ZN(n9684) );
  NAND2_X1 U12254 ( .A1(n9657), .A2(n9684), .ZN(n14879) );
  INV_X1 U12255 ( .A(n14879), .ZN(n14874) );
  AOI22_X1 U12256 ( .A1(n9848), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9847), .B2(
        n14874), .ZN(n9658) );
  NAND2_X1 U12257 ( .A1(n9959), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9668) );
  INV_X1 U12258 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9661) );
  OR2_X1 U12259 ( .A1(n9896), .A2(n9661), .ZN(n9667) );
  INV_X1 U12260 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n11863) );
  NAND2_X1 U12261 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9662) );
  NAND2_X1 U12262 ( .A1(n11863), .A2(n9662), .ZN(n9663) );
  NAND2_X1 U12263 ( .A1(n9673), .A2(n9663), .ZN(n11864) );
  OR2_X1 U12264 ( .A1(n6429), .A2(n11864), .ZN(n9666) );
  INV_X1 U12265 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9664) );
  OR2_X1 U12266 ( .A1(n9691), .A2(n9664), .ZN(n9665) );
  NAND4_X1 U12267 ( .A1(n9668), .A2(n9667), .A3(n9666), .A4(n9665), .ZN(n14817) );
  OR2_X1 U12268 ( .A1(n11868), .A2(n14817), .ZN(n11879) );
  NAND2_X1 U12269 ( .A1(n11868), .A2(n14817), .ZN(n9669) );
  INV_X1 U12270 ( .A(n14817), .ZN(n11819) );
  NAND2_X1 U12271 ( .A1(n11868), .A2(n11819), .ZN(n9670) );
  NAND2_X1 U12272 ( .A1(n9959), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9679) );
  INV_X1 U12273 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14895) );
  OR2_X1 U12274 ( .A1(n9896), .A2(n14895), .ZN(n9678) );
  INV_X1 U12275 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9672) );
  NAND2_X1 U12276 ( .A1(n9673), .A2(n9672), .ZN(n9674) );
  OR2_X1 U12277 ( .A1(n6429), .A2(n11886), .ZN(n9677) );
  INV_X1 U12278 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9675) );
  OR2_X1 U12279 ( .A1(n9691), .A2(n9675), .ZN(n9676) );
  NAND4_X1 U12280 ( .A1(n9679), .A2(n9678), .A3(n9677), .A4(n9676), .ZN(n14816) );
  NAND2_X1 U12281 ( .A1(n10791), .A2(n9902), .ZN(n9682) );
  NAND2_X1 U12282 ( .A1(n9684), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9680) );
  XNOR2_X1 U12283 ( .A(n9680), .B(P1_IR_REG_6__SCAN_IN), .ZN(n14894) );
  AOI22_X1 U12284 ( .A1(n9848), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9847), .B2(
        n14894), .ZN(n9681) );
  OR2_X1 U12285 ( .A1(n14816), .A2(n15543), .ZN(n12024) );
  NAND2_X1 U12286 ( .A1(n15543), .A2(n14816), .ZN(n9683) );
  NAND2_X1 U12287 ( .A1(n12024), .A2(n9683), .ZN(n11876) );
  INV_X1 U12288 ( .A(n14816), .ZN(n11903) );
  NAND2_X1 U12289 ( .A1(n10827), .A2(n9902), .ZN(n9687) );
  NAND2_X1 U12290 ( .A1(n9698), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9685) );
  XNOR2_X1 U12291 ( .A(n9685), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14911) );
  AOI22_X1 U12292 ( .A1(n9848), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9847), .B2(
        n14911), .ZN(n9686) );
  NAND2_X1 U12293 ( .A1(n9959), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9696) );
  INV_X1 U12294 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10923) );
  OR2_X1 U12295 ( .A1(n9896), .A2(n10923), .ZN(n9695) );
  INV_X1 U12296 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9689) );
  NAND2_X1 U12297 ( .A1(n9705), .A2(n9690), .ZN(n12036) );
  OR2_X1 U12298 ( .A1(n6429), .A2(n12036), .ZN(n9694) );
  INV_X1 U12299 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9692) );
  OR2_X1 U12300 ( .A1(n10615), .A2(n9692), .ZN(n9693) );
  INV_X1 U12301 ( .A(n14815), .ZN(n12154) );
  NAND2_X1 U12302 ( .A1(n15548), .A2(n12154), .ZN(n9697) );
  NAND2_X1 U12303 ( .A1(n10860), .A2(n9902), .ZN(n9703) );
  INV_X1 U12304 ( .A(n9698), .ZN(n9700) );
  NAND2_X1 U12305 ( .A1(n9700), .A2(n9699), .ZN(n9714) );
  NAND2_X1 U12306 ( .A1(n9714), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9701) );
  XNOR2_X1 U12307 ( .A(n9701), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10963) );
  AOI22_X1 U12308 ( .A1(n9848), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9847), .B2(
        n10963), .ZN(n9702) );
  NAND2_X1 U12309 ( .A1(n9959), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9711) );
  INV_X1 U12310 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9704) );
  OR2_X1 U12311 ( .A1(n9896), .A2(n9704), .ZN(n9710) );
  NAND2_X1 U12312 ( .A1(n9705), .A2(n6672), .ZN(n9706) );
  NAND2_X1 U12313 ( .A1(n9718), .A2(n9706), .ZN(n12303) );
  OR2_X1 U12314 ( .A1(n6429), .A2(n12303), .ZN(n9709) );
  INV_X1 U12315 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9707) );
  OR2_X1 U12316 ( .A1(n10615), .A2(n9707), .ZN(n9708) );
  NAND4_X1 U12317 ( .A1(n9711), .A2(n9710), .A3(n9709), .A4(n9708), .ZN(n14814) );
  OR2_X1 U12318 ( .A1(n12220), .A2(n14814), .ZN(n10004) );
  NAND2_X1 U12319 ( .A1(n12220), .A2(n14814), .ZN(n9712) );
  INV_X1 U12320 ( .A(n14814), .ZN(n12522) );
  OR2_X1 U12321 ( .A1(n12220), .A2(n12522), .ZN(n9713) );
  NAND2_X1 U12322 ( .A1(n10877), .A2(n9902), .ZN(n9716) );
  NAND2_X1 U12323 ( .A1(n9741), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9728) );
  XNOR2_X1 U12324 ( .A(n9728), .B(P1_IR_REG_9__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U12325 ( .A1(n9848), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9847), .B2(
        n11005), .ZN(n9715) );
  NAND2_X1 U12326 ( .A1(n9959), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9724) );
  INV_X1 U12327 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9717) );
  OR2_X1 U12328 ( .A1(n9896), .A2(n9717), .ZN(n9723) );
  NAND2_X1 U12329 ( .A1(n9718), .A2(n6674), .ZN(n9719) );
  NAND2_X1 U12330 ( .A1(n9735), .A2(n9719), .ZN(n12521) );
  OR2_X1 U12331 ( .A1(n6429), .A2(n12521), .ZN(n9722) );
  INV_X1 U12332 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9720) );
  OR2_X1 U12333 ( .A1(n10615), .A2(n9720), .ZN(n9721) );
  NAND4_X1 U12334 ( .A1(n9724), .A2(n9723), .A3(n9722), .A4(n9721), .ZN(n14813) );
  INV_X1 U12335 ( .A(n14813), .ZN(n12153) );
  XNOR2_X1 U12336 ( .A(n12516), .B(n12153), .ZN(n12189) );
  NAND2_X1 U12337 ( .A1(n12516), .A2(n12153), .ZN(n9726) );
  NAND2_X1 U12338 ( .A1(n10898), .A2(n9902), .ZN(n9732) );
  NAND2_X1 U12339 ( .A1(n9728), .A2(n9727), .ZN(n9729) );
  NAND2_X1 U12340 ( .A1(n9729), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9730) );
  XNOR2_X1 U12341 ( .A(n9730), .B(P1_IR_REG_10__SCAN_IN), .ZN(n14924) );
  AOI22_X1 U12342 ( .A1(n9848), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n14924), 
        .B2(n9847), .ZN(n9731) );
  NAND2_X1 U12343 ( .A1(n9959), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9740) );
  INV_X1 U12344 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9733) );
  OR2_X1 U12345 ( .A1(n9896), .A2(n9733), .ZN(n9739) );
  NAND2_X1 U12346 ( .A1(n9735), .A2(n9734), .ZN(n9736) );
  NAND2_X1 U12347 ( .A1(n9747), .A2(n9736), .ZN(n12336) );
  OR2_X1 U12348 ( .A1(n6429), .A2(n12336), .ZN(n9738) );
  INV_X1 U12349 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14432) );
  OR2_X1 U12350 ( .A1(n10615), .A2(n14432), .ZN(n9737) );
  NAND4_X1 U12351 ( .A1(n9740), .A2(n9739), .A3(n9738), .A4(n9737), .ZN(n14812) );
  XNOR2_X1 U12352 ( .A(n14674), .B(n12590), .ZN(n12332) );
  INV_X1 U12353 ( .A(n9741), .ZN(n9743) );
  NOR2_X1 U12354 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n9742) );
  NAND2_X1 U12355 ( .A1(n9743), .A2(n9742), .ZN(n9755) );
  NAND2_X1 U12356 ( .A1(n9755), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9744) );
  XNOR2_X1 U12357 ( .A(n9744), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U12358 ( .A1(n9848), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n11269), 
        .B2(n9847), .ZN(n9745) );
  NAND2_X1 U12359 ( .A1(n9959), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9752) );
  INV_X1 U12360 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14437) );
  OR2_X1 U12361 ( .A1(n9896), .A2(n14437), .ZN(n9751) );
  INV_X1 U12362 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9746) );
  NAND2_X1 U12363 ( .A1(n9747), .A2(n9746), .ZN(n9748) );
  NAND2_X1 U12364 ( .A1(n9759), .A2(n9748), .ZN(n12589) );
  OR2_X1 U12365 ( .A1(n6429), .A2(n12589), .ZN(n9750) );
  INV_X1 U12366 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n12692) );
  OR2_X1 U12367 ( .A1(n10615), .A2(n12692), .ZN(n9749) );
  NAND4_X1 U12368 ( .A1(n9752), .A2(n9751), .A3(n9750), .A4(n9749), .ZN(n14811) );
  OR2_X1 U12369 ( .A1(n12423), .A2(n14811), .ZN(n10006) );
  NAND2_X1 U12370 ( .A1(n12423), .A2(n14811), .ZN(n9753) );
  NAND2_X1 U12371 ( .A1(n10006), .A2(n9753), .ZN(n12430) );
  OR2_X1 U12372 ( .A1(n14674), .A2(n12590), .ZN(n12427) );
  INV_X1 U12373 ( .A(n14811), .ZN(n12629) );
  OR2_X1 U12374 ( .A1(n12423), .A2(n12629), .ZN(n9754) );
  NAND2_X1 U12375 ( .A1(n9756), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9767) );
  XNOR2_X1 U12376 ( .A(n9767), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U12377 ( .A1(n9847), .A2(n11609), .B1(n9848), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n9757) );
  NAND2_X1 U12378 ( .A1(n9959), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9764) );
  INV_X1 U12379 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n12750) );
  OR2_X1 U12380 ( .A1(n9896), .A2(n12750), .ZN(n9763) );
  INV_X1 U12381 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9758) );
  NAND2_X1 U12382 ( .A1(n9759), .A2(n9758), .ZN(n9760) );
  NAND2_X1 U12383 ( .A1(n9774), .A2(n9760), .ZN(n12628) );
  OR2_X1 U12384 ( .A1(n6429), .A2(n12628), .ZN(n9762) );
  INV_X1 U12385 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n12753) );
  OR2_X1 U12386 ( .A1(n10615), .A2(n12753), .ZN(n9761) );
  NAND4_X1 U12387 ( .A1(n9764), .A2(n9763), .A3(n9762), .A4(n9761), .ZN(n14810) );
  XNOR2_X1 U12388 ( .A(n12567), .B(n14810), .ZN(n12560) );
  NAND2_X1 U12389 ( .A1(n12561), .A2(n12560), .ZN(n12559) );
  INV_X1 U12390 ( .A(n14810), .ZN(n14745) );
  OR2_X1 U12391 ( .A1(n12567), .A2(n14745), .ZN(n9765) );
  NAND2_X1 U12392 ( .A1(n9767), .A2(n9766), .ZN(n9768) );
  NAND2_X1 U12393 ( .A1(n9768), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9770) );
  OR2_X1 U12394 ( .A1(n9770), .A2(n9769), .ZN(n9771) );
  NAND2_X1 U12395 ( .A1(n9770), .A2(n9769), .ZN(n9780) );
  AOI22_X1 U12396 ( .A1(n11663), .A2(n9847), .B1(P2_DATAO_REG_13__SCAN_IN), 
        .B2(n9848), .ZN(n9772) );
  NAND2_X1 U12397 ( .A1(n10612), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9779) );
  INV_X1 U12398 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n12717) );
  OR2_X1 U12399 ( .A1(n9614), .A2(n12717), .ZN(n9778) );
  INV_X1 U12400 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9773) );
  NAND2_X1 U12401 ( .A1(n9774), .A2(n9773), .ZN(n9775) );
  NAND2_X1 U12402 ( .A1(n9785), .A2(n9775), .ZN(n14744) );
  OR2_X1 U12403 ( .A1(n6429), .A2(n14744), .ZN(n9777) );
  INV_X1 U12404 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n15419) );
  OR2_X1 U12405 ( .A1(n10615), .A2(n15419), .ZN(n9776) );
  NAND4_X1 U12406 ( .A1(n9779), .A2(n9778), .A3(n9777), .A4(n9776), .ZN(n14809) );
  OR2_X1 U12407 ( .A1(n12720), .A2(n7287), .ZN(n12765) );
  NAND2_X1 U12408 ( .A1(n11020), .A2(n9902), .ZN(n9783) );
  NAND2_X1 U12409 ( .A1(n9780), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9781) );
  XNOR2_X1 U12410 ( .A(n9781), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12124) );
  AOI22_X1 U12411 ( .A1(n12124), .A2(n9847), .B1(P2_DATAO_REG_14__SCAN_IN), 
        .B2(n9848), .ZN(n9782) );
  INV_X1 U12412 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9784) );
  NAND2_X1 U12413 ( .A1(n9785), .A2(n9784), .ZN(n9786) );
  NAND2_X1 U12414 ( .A1(n9798), .A2(n9786), .ZN(n12771) );
  NAND2_X1 U12415 ( .A1(n9929), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9787) );
  OAI21_X1 U12416 ( .B1(n12771), .B2(n6429), .A(n9787), .ZN(n9790) );
  INV_X1 U12417 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n15363) );
  NAND2_X1 U12418 ( .A1(n9959), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9788) );
  OAI21_X1 U12419 ( .B1(n9896), .B2(n15363), .A(n9788), .ZN(n9789) );
  NAND2_X1 U12420 ( .A1(n12770), .A2(n14788), .ZN(n10534) );
  AND2_X2 U12421 ( .A1(n10531), .A2(n10534), .ZN(n12764) );
  NAND2_X1 U12422 ( .A1(n10978), .A2(n9902), .ZN(n9795) );
  NAND2_X1 U12423 ( .A1(n9791), .A2(n9792), .ZN(n9845) );
  NAND2_X1 U12424 ( .A1(n9845), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9793) );
  XNOR2_X1 U12425 ( .A(n9793), .B(P1_IR_REG_15__SCAN_IN), .ZN(n14940) );
  AOI22_X1 U12426 ( .A1(n9848), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9847), 
        .B2(n14940), .ZN(n9794) );
  INV_X1 U12427 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n15412) );
  INV_X1 U12428 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9797) );
  NAND2_X1 U12429 ( .A1(n9798), .A2(n9797), .ZN(n9799) );
  NAND2_X1 U12430 ( .A1(n9808), .A2(n9799), .ZN(n15249) );
  OR2_X1 U12431 ( .A1(n15249), .A2(n6429), .ZN(n9801) );
  AOI22_X1 U12432 ( .A1(n9959), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n10612), 
        .B2(P1_REG1_REG_15__SCAN_IN), .ZN(n9800) );
  OAI211_X1 U12433 ( .C1(n10615), .C2(n15412), .A(n9801), .B(n9800), .ZN(
        n14808) );
  INV_X1 U12434 ( .A(n14808), .ZN(n15240) );
  NAND2_X1 U12435 ( .A1(n11068), .A2(n9902), .ZN(n9806) );
  NAND2_X1 U12436 ( .A1(n9843), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9802) );
  MUX2_X1 U12437 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9802), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9804) );
  INV_X1 U12438 ( .A(n9843), .ZN(n9803) );
  INV_X1 U12439 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9840) );
  NAND2_X1 U12440 ( .A1(n9803), .A2(n9840), .ZN(n9826) );
  NAND2_X1 U12441 ( .A1(n9804), .A2(n9826), .ZN(n14951) );
  INV_X1 U12442 ( .A(n14951), .ZN(n14955) );
  AOI22_X1 U12443 ( .A1(n9848), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9847), 
        .B2(n14955), .ZN(n9805) );
  INV_X1 U12444 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9807) );
  NAND2_X1 U12445 ( .A1(n9808), .A2(n9807), .ZN(n9809) );
  NAND2_X1 U12446 ( .A1(n9817), .A2(n9809), .ZN(n14709) );
  AOI22_X1 U12447 ( .A1(n9959), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n10612), 
        .B2(P1_REG1_REG_16__SCAN_IN), .ZN(n9811) );
  NAND2_X1 U12448 ( .A1(n9929), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9810) );
  OAI211_X1 U12449 ( .C1(n14709), .C2(n6429), .A(n9811), .B(n9810), .ZN(n15259) );
  INV_X1 U12450 ( .A(n15259), .ZN(n14791) );
  XNOR2_X1 U12451 ( .A(n15351), .B(n14791), .ZN(n15236) );
  NAND2_X1 U12452 ( .A1(n11195), .A2(n9902), .ZN(n9815) );
  NAND2_X1 U12453 ( .A1(n9826), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9813) );
  XNOR2_X1 U12454 ( .A(n9813), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14965) );
  AOI22_X1 U12455 ( .A1(n9848), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9847), 
        .B2(n14965), .ZN(n9814) );
  INV_X1 U12456 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9816) );
  NAND2_X1 U12457 ( .A1(n9817), .A2(n9816), .ZN(n9818) );
  NAND2_X1 U12458 ( .A1(n9831), .A2(n9818), .ZN(n15216) );
  OR2_X1 U12459 ( .A1(n15216), .A2(n6429), .ZN(n9824) );
  INV_X1 U12460 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9821) );
  NAND2_X1 U12461 ( .A1(n9959), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9820) );
  NAND2_X1 U12462 ( .A1(n10612), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9819) );
  OAI211_X1 U12463 ( .C1(n9821), .C2(n10615), .A(n9820), .B(n9819), .ZN(n9822)
         );
  INV_X1 U12464 ( .A(n9822), .ZN(n9823) );
  NAND2_X1 U12465 ( .A1(n9824), .A2(n9823), .ZN(n14807) );
  INV_X1 U12466 ( .A(n14807), .ZN(n15242) );
  NAND2_X1 U12467 ( .A1(n15345), .A2(n15242), .ZN(n10547) );
  NAND2_X1 U12468 ( .A1(n10546), .A2(n10547), .ZN(n15213) );
  NAND2_X1 U12469 ( .A1(n15214), .A2(n10546), .ZN(n15193) );
  NAND2_X1 U12470 ( .A1(n11433), .A2(n9902), .ZN(n9829) );
  OAI21_X1 U12471 ( .B1(n9826), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9827) );
  XNOR2_X1 U12472 ( .A(n9827), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14983) );
  AOI22_X1 U12473 ( .A1(n9848), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9847), 
        .B2(n14983), .ZN(n9828) );
  INV_X1 U12474 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9830) );
  NAND2_X1 U12475 ( .A1(n9831), .A2(n9830), .ZN(n9832) );
  AND2_X1 U12476 ( .A1(n9852), .A2(n9832), .ZN(n15200) );
  INV_X1 U12477 ( .A(n6429), .ZN(n9944) );
  NAND2_X1 U12478 ( .A1(n15200), .A2(n9944), .ZN(n9838) );
  INV_X1 U12479 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9835) );
  NAND2_X1 U12480 ( .A1(n9959), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9834) );
  NAND2_X1 U12481 ( .A1(n10612), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9833) );
  OAI211_X1 U12482 ( .C1(n9835), .C2(n10615), .A(n9834), .B(n9833), .ZN(n9836)
         );
  INV_X1 U12483 ( .A(n9836), .ZN(n9837) );
  NAND2_X1 U12484 ( .A1(n9838), .A2(n9837), .ZN(n14806) );
  INV_X1 U12485 ( .A(n14806), .ZN(n10225) );
  NAND2_X1 U12486 ( .A1(n15199), .A2(n10225), .ZN(n10564) );
  NAND2_X1 U12487 ( .A1(n11453), .A2(n9902), .ZN(n9850) );
  NAND3_X1 U12488 ( .A1(n9841), .A2(n9840), .A3(n9839), .ZN(n9842) );
  AOI22_X1 U12489 ( .A1(n9848), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14993), 
        .B2(n9847), .ZN(n9849) );
  INV_X1 U12490 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9851) );
  NAND2_X1 U12491 ( .A1(n9852), .A2(n9851), .ZN(n9853) );
  NAND2_X1 U12492 ( .A1(n9870), .A2(n9853), .ZN(n15181) );
  OR2_X1 U12493 ( .A1(n15181), .A2(n6429), .ZN(n9859) );
  INV_X1 U12494 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14475) );
  NAND2_X1 U12495 ( .A1(n9959), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9856) );
  NAND2_X1 U12496 ( .A1(n9929), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9855) );
  OAI211_X1 U12497 ( .C1(n9896), .C2(n14475), .A(n9856), .B(n9855), .ZN(n9857)
         );
  INV_X1 U12498 ( .A(n9857), .ZN(n9858) );
  NAND2_X1 U12499 ( .A1(n9859), .A2(n9858), .ZN(n14805) );
  INV_X1 U12500 ( .A(n14805), .ZN(n14735) );
  OR2_X1 U12501 ( .A1(n15332), .A2(n14735), .ZN(n10570) );
  NAND2_X1 U12502 ( .A1(n15332), .A2(n14735), .ZN(n15159) );
  NAND2_X1 U12503 ( .A1(n10570), .A2(n15159), .ZN(n15177) );
  OR2_X1 U12504 ( .A1(n9631), .A2(n11824), .ZN(n9860) );
  INV_X1 U12505 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14694) );
  NAND2_X1 U12506 ( .A1(n9872), .A2(n14694), .ZN(n9862) );
  NAND2_X1 U12507 ( .A1(n9884), .A2(n9862), .ZN(n15149) );
  INV_X1 U12508 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n14409) );
  NAND2_X1 U12509 ( .A1(n10612), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9864) );
  NAND2_X1 U12510 ( .A1(n9959), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9863) );
  OAI211_X1 U12511 ( .C1(n14409), .C2(n10615), .A(n9864), .B(n9863), .ZN(n9865) );
  INV_X1 U12512 ( .A(n9865), .ZN(n9866) );
  INV_X1 U12513 ( .A(n15122), .ZN(n14756) );
  NAND2_X1 U12514 ( .A1(n11774), .A2(n9902), .ZN(n9869) );
  OR2_X1 U12515 ( .A1(n9631), .A2(n11776), .ZN(n9868) );
  NAND2_X2 U12516 ( .A1(n9869), .A2(n9868), .ZN(n15171) );
  INV_X1 U12517 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14736) );
  NAND2_X1 U12518 ( .A1(n9870), .A2(n14736), .ZN(n9871) );
  NAND2_X1 U12519 ( .A1(n9872), .A2(n9871), .ZN(n15169) );
  INV_X1 U12520 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9875) );
  NAND2_X1 U12521 ( .A1(n9959), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9874) );
  NAND2_X1 U12522 ( .A1(n10612), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n9873) );
  OAI211_X1 U12523 ( .C1(n9875), .C2(n10615), .A(n9874), .B(n9873), .ZN(n9876)
         );
  INV_X1 U12524 ( .A(n9876), .ZN(n9877) );
  INV_X1 U12525 ( .A(n14804), .ZN(n10567) );
  NAND2_X1 U12526 ( .A1(n15171), .A2(n10567), .ZN(n10017) );
  INV_X1 U12527 ( .A(n15151), .ZN(n15148) );
  INV_X1 U12528 ( .A(n15138), .ZN(n15121) );
  NAND2_X1 U12529 ( .A1(n15121), .A2(n14756), .ZN(n9881) );
  AOI22_X1 U12530 ( .A1(n15148), .A2(n9881), .B1(n15138), .B2(n15122), .ZN(
        n9889) );
  NAND2_X1 U12531 ( .A1(n9882), .A2(n6978), .ZN(n9883) );
  INV_X1 U12532 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14758) );
  NAND2_X1 U12533 ( .A1(n9884), .A2(n14758), .ZN(n9885) );
  INV_X1 U12534 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n15402) );
  NAND2_X1 U12535 ( .A1(n9959), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9887) );
  NAND2_X1 U12536 ( .A1(n10612), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9886) );
  OAI211_X1 U12537 ( .C1(n15402), .C2(n10615), .A(n9887), .B(n9886), .ZN(n9888) );
  XNOR2_X1 U12538 ( .A(n15404), .B(n14691), .ZN(n15124) );
  AND2_X1 U12539 ( .A1(n9889), .A2(n15124), .ZN(n9890) );
  INV_X1 U12540 ( .A(n14691), .ZN(n14803) );
  INV_X1 U12541 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12048) );
  OR2_X1 U12542 ( .A1(n9631), .A2(n12048), .ZN(n9892) );
  XNOR2_X1 U12543 ( .A(n9907), .B(P1_REG3_REG_23__SCAN_IN), .ZN(n15114) );
  NAND2_X1 U12544 ( .A1(n15114), .A2(n9944), .ZN(n9899) );
  INV_X1 U12545 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n15313) );
  NAND2_X1 U12546 ( .A1(n9959), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9895) );
  NAND2_X1 U12547 ( .A1(n9929), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9894) );
  OAI211_X1 U12548 ( .C1(n9896), .C2(n15313), .A(n9895), .B(n9894), .ZN(n9897)
         );
  INV_X1 U12549 ( .A(n9897), .ZN(n9898) );
  INV_X1 U12550 ( .A(n15089), .ZN(n14757) );
  NAND2_X1 U12551 ( .A1(n15113), .A2(n14757), .ZN(n9900) );
  NAND2_X1 U12552 ( .A1(n9901), .A2(n9900), .ZN(n15047) );
  OR2_X1 U12553 ( .A1(n9631), .A2(n12110), .ZN(n9903) );
  AND2_X1 U12554 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n9905) );
  INV_X1 U12555 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9906) );
  INV_X1 U12556 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14723) );
  OAI21_X1 U12557 ( .B1(n9907), .B2(n9906), .A(n14723), .ZN(n9908) );
  NAND2_X1 U12558 ( .A1(n9917), .A2(n9908), .ZN(n15100) );
  INV_X1 U12559 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n15394) );
  NAND2_X1 U12560 ( .A1(n9959), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9910) );
  NAND2_X1 U12561 ( .A1(n10612), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9909) );
  OAI211_X1 U12562 ( .C1(n15394), .C2(n10615), .A(n9910), .B(n9909), .ZN(n9911) );
  INV_X1 U12563 ( .A(n9911), .ZN(n9912) );
  OR2_X1 U12564 ( .A1(n9631), .A2(n12242), .ZN(n9914) );
  INV_X1 U12565 ( .A(n9917), .ZN(n9916) );
  INV_X1 U12566 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14702) );
  NAND2_X1 U12567 ( .A1(n9917), .A2(n14702), .ZN(n9918) );
  NAND2_X1 U12568 ( .A1(n9927), .A2(n9918), .ZN(n15078) );
  INV_X1 U12569 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n15390) );
  NAND2_X1 U12570 ( .A1(n9959), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9920) );
  NAND2_X1 U12571 ( .A1(n10612), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9919) );
  OAI211_X1 U12572 ( .C1(n15390), .C2(n10615), .A(n9920), .B(n9919), .ZN(n9921) );
  INV_X1 U12573 ( .A(n9921), .ZN(n9922) );
  INV_X1 U12574 ( .A(n15090), .ZN(n14724) );
  OAI21_X1 U12575 ( .B1(n15396), .B2(n14802), .A(n15048), .ZN(n9938) );
  OR2_X1 U12576 ( .A1(n9631), .A2(n12547), .ZN(n9924) );
  INV_X1 U12577 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U12578 ( .A1(n9927), .A2(n9926), .ZN(n9928) );
  NAND2_X1 U12579 ( .A1(n15052), .A2(n9944), .ZN(n9934) );
  INV_X1 U12580 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n15057) );
  NAND2_X1 U12581 ( .A1(n10612), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9931) );
  NAND2_X1 U12582 ( .A1(n9929), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9930) );
  OAI211_X1 U12583 ( .C1(n9614), .C2(n15057), .A(n9931), .B(n9930), .ZN(n9932)
         );
  INV_X1 U12584 ( .A(n9932), .ZN(n9933) );
  OR2_X1 U12585 ( .A1(n15298), .A2(n14724), .ZN(n10025) );
  INV_X1 U12586 ( .A(n14802), .ZN(n9935) );
  NAND2_X1 U12587 ( .A1(n10025), .A2(n15070), .ZN(n9936) );
  NAND2_X1 U12588 ( .A1(n9936), .A2(n15048), .ZN(n9937) );
  OAI211_X1 U12589 ( .C1(n15047), .C2(n9938), .A(n10662), .B(n9937), .ZN(n9941) );
  INV_X1 U12590 ( .A(n15037), .ZN(n9939) );
  NAND2_X1 U12591 ( .A1(n15053), .A2(n9939), .ZN(n9940) );
  OR2_X1 U12592 ( .A1(n9631), .A2(n15434), .ZN(n9942) );
  XNOR2_X1 U12593 ( .A(n9957), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n15043) );
  NAND2_X1 U12594 ( .A1(n15043), .A2(n9944), .ZN(n9949) );
  INV_X1 U12595 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n15385) );
  NAND2_X1 U12596 ( .A1(n9959), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9946) );
  NAND2_X1 U12597 ( .A1(n10612), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9945) );
  OAI211_X1 U12598 ( .C1(n15385), .C2(n10615), .A(n9946), .B(n9945), .ZN(n9947) );
  INV_X1 U12599 ( .A(n9947), .ZN(n9948) );
  INV_X1 U12600 ( .A(n14801), .ZN(n9950) );
  OR2_X1 U12601 ( .A1(n9631), .A2(n12891), .ZN(n9951) );
  INV_X1 U12602 ( .A(n9957), .ZN(n9954) );
  AND2_X1 U12603 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n9953) );
  NAND2_X1 U12604 ( .A1(n9954), .A2(n9953), .ZN(n13201) );
  INV_X1 U12605 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9956) );
  INV_X1 U12606 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9955) );
  OAI21_X1 U12607 ( .B1(n9957), .B2(n9956), .A(n9955), .ZN(n9958) );
  NAND2_X1 U12608 ( .A1(n13201), .A2(n9958), .ZN(n10313) );
  INV_X1 U12609 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n15382) );
  NAND2_X1 U12610 ( .A1(n9959), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9961) );
  NAND2_X1 U12611 ( .A1(n10612), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9960) );
  OAI211_X1 U12612 ( .C1(n15382), .C2(n10615), .A(n9961), .B(n9960), .ZN(n9962) );
  INV_X1 U12613 ( .A(n9962), .ZN(n9963) );
  AND2_X1 U12614 ( .A1(n15023), .A2(n12964), .ZN(n9965) );
  NAND2_X1 U12615 ( .A1(n14634), .A2(n9902), .ZN(n9967) );
  OR2_X1 U12616 ( .A1(n9631), .A2(n15431), .ZN(n9966) );
  NAND2_X2 U12617 ( .A1(n9967), .A2(n9966), .ZN(n10626) );
  OR2_X1 U12618 ( .A1(n13201), .A2(n6429), .ZN(n9972) );
  NAND2_X1 U12619 ( .A1(n10612), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9969) );
  INV_X1 U12620 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n13204) );
  OR2_X1 U12621 ( .A1(n9614), .A2(n13204), .ZN(n9968) );
  OAI211_X1 U12622 ( .C1(n10067), .C2(n10615), .A(n9969), .B(n9968), .ZN(n9970) );
  INV_X1 U12623 ( .A(n9970), .ZN(n9971) );
  NAND2_X1 U12624 ( .A1(n9972), .A2(n9971), .ZN(n14800) );
  INV_X1 U12625 ( .A(n14800), .ZN(n10625) );
  INV_X2 U12626 ( .A(n9982), .ZN(n9976) );
  AND2_X2 U12627 ( .A1(n9978), .A2(n9977), .ZN(n10031) );
  INV_X1 U12628 ( .A(n11775), .ZN(n11890) );
  NAND2_X1 U12629 ( .A1(n10031), .A2(n11890), .ZN(n10471) );
  INV_X1 U12630 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n14416) );
  XNOR2_X1 U12631 ( .A(n9983), .B(n14416), .ZN(n11127) );
  OR2_X1 U12632 ( .A1(n11127), .A2(n11458), .ZN(n9984) );
  NAND2_X1 U12633 ( .A1(n9985), .A2(n15260), .ZN(n9988) );
  INV_X1 U12634 ( .A(n11127), .ZN(n15438) );
  AND2_X1 U12635 ( .A1(n10031), .A2(n15438), .ZN(n10869) );
  INV_X1 U12636 ( .A(n14836), .ZN(n14839) );
  NAND2_X1 U12637 ( .A1(n15038), .A2(n15257), .ZN(n9987) );
  NAND2_X1 U12638 ( .A1(n9988), .A2(n9987), .ZN(n13199) );
  INV_X1 U12639 ( .A(n13199), .ZN(n10039) );
  NAND2_X1 U12640 ( .A1(n10031), .A2(n11775), .ZN(n10083) );
  NAND2_X1 U12641 ( .A1(n15438), .A2(n11458), .ZN(n9989) );
  INV_X2 U12642 ( .A(n10297), .ZN(n10281) );
  NAND2_X1 U12643 ( .A1(n10645), .A2(n15438), .ZN(n9990) );
  NAND2_X1 U12644 ( .A1(n10281), .A2(n9990), .ZN(n15354) );
  XNOR2_X1 U12645 ( .A(n10096), .B(n11498), .ZN(n10484) );
  INV_X1 U12646 ( .A(n11128), .ZN(n11151) );
  NAND2_X1 U12647 ( .A1(n10484), .A2(n11150), .ZN(n9993) );
  NAND2_X1 U12648 ( .A1(n9991), .A2(n11498), .ZN(n9992) );
  NAND2_X1 U12649 ( .A1(n9993), .A2(n9992), .ZN(n11251) );
  NAND2_X1 U12650 ( .A1(n11159), .A2(n7048), .ZN(n9994) );
  INV_X1 U12651 ( .A(n11321), .ZN(n11314) );
  NAND2_X1 U12652 ( .A1(n9995), .A2(n11545), .ZN(n9996) );
  NAND2_X1 U12653 ( .A1(n11507), .A2(n11512), .ZN(n11506) );
  NAND2_X1 U12654 ( .A1(n11506), .A2(n11761), .ZN(n9997) );
  INV_X1 U12655 ( .A(n10652), .ZN(n11764) );
  NAND2_X1 U12656 ( .A1(n9997), .A2(n11764), .ZN(n11759) );
  AND2_X1 U12657 ( .A1(n11879), .A2(n9999), .ZN(n9998) );
  INV_X1 U12658 ( .A(n9999), .ZN(n10001) );
  INV_X1 U12659 ( .A(n11876), .ZN(n11880) );
  INV_X1 U12660 ( .A(n12028), .ZN(n10654) );
  OR2_X1 U12661 ( .A1(n15548), .A2(n14815), .ZN(n10003) );
  OR2_X1 U12662 ( .A1(n12516), .A2(n14813), .ZN(n10005) );
  INV_X1 U12663 ( .A(n12430), .ZN(n12420) );
  INV_X1 U12664 ( .A(n12560), .ZN(n12557) );
  OR2_X1 U12665 ( .A1(n12567), .A2(n14810), .ZN(n10007) );
  NAND2_X1 U12666 ( .A1(n12770), .A2(n15256), .ZN(n15252) );
  OR2_X1 U12667 ( .A1(n15271), .A2(n14808), .ZN(n15227) );
  NAND2_X1 U12668 ( .A1(n15226), .A2(n15227), .ZN(n10009) );
  NAND2_X1 U12669 ( .A1(n15351), .A2(n15259), .ZN(n10008) );
  AND2_X1 U12670 ( .A1(n7521), .A2(n15227), .ZN(n15206) );
  OR2_X1 U12671 ( .A1(n15351), .A2(n15259), .ZN(n15208) );
  OAI211_X1 U12672 ( .C1(n15206), .C2(n6554), .A(n15213), .B(n15208), .ZN(
        n10010) );
  INV_X1 U12673 ( .A(n10010), .ZN(n10011) );
  NAND2_X1 U12674 ( .A1(n15345), .A2(n14807), .ZN(n10012) );
  OR2_X1 U12675 ( .A1(n15199), .A2(n14806), .ZN(n10013) );
  NAND2_X1 U12676 ( .A1(n15190), .A2(n10013), .ZN(n10015) );
  NAND2_X1 U12677 ( .A1(n15199), .A2(n14806), .ZN(n10014) );
  OR2_X1 U12678 ( .A1(n15332), .A2(n14805), .ZN(n10016) );
  NAND2_X1 U12679 ( .A1(n15171), .A2(n14804), .ZN(n10019) );
  XNOR2_X1 U12680 ( .A(n15151), .B(n15122), .ZN(n15139) );
  INV_X1 U12681 ( .A(n15124), .ZN(n15128) );
  NAND2_X1 U12682 ( .A1(n15404), .A2(n14691), .ZN(n10021) );
  NAND2_X1 U12683 ( .A1(n15113), .A2(n15089), .ZN(n15085) );
  NAND2_X1 U12684 ( .A1(n15099), .A2(n14802), .ZN(n10026) );
  INV_X1 U12685 ( .A(n10026), .ZN(n10022) );
  OR2_X1 U12686 ( .A1(n15099), .A2(n14802), .ZN(n15065) );
  INV_X1 U12687 ( .A(n15113), .ZN(n15400) );
  NAND3_X1 U12688 ( .A1(n10026), .A2(n15400), .A3(n14757), .ZN(n10027) );
  AND3_X1 U12689 ( .A1(n15071), .A2(n15065), .A3(n10027), .ZN(n10028) );
  NAND2_X1 U12690 ( .A1(n15053), .A2(n15037), .ZN(n10029) );
  NAND2_X1 U12691 ( .A1(n15023), .A2(n15038), .ZN(n10030) );
  NOR2_X4 U12692 ( .A1(n11317), .A2(n15523), .ZN(n11508) );
  INV_X1 U12693 ( .A(n11868), .ZN(n11770) );
  INV_X1 U12694 ( .A(n12220), .ZN(n12304) );
  NAND2_X1 U12695 ( .A1(n12021), .A2(n12304), .ZN(n12147) );
  INV_X1 U12696 ( .A(n15351), .ZN(n15235) );
  NAND2_X2 U12697 ( .A1(n15269), .A2(n15235), .ZN(n15230) );
  INV_X1 U12698 ( .A(n15332), .ZN(n15186) );
  OR2_X2 U12699 ( .A1(n15079), .A2(n15298), .ZN(n15054) );
  AND2_X1 U12700 ( .A1(n11775), .A2(n11127), .ZN(n10642) );
  NAND2_X4 U12701 ( .A1(n10642), .A2(n11825), .ZN(n15270) );
  AOI21_X1 U12702 ( .B1(n10032), .B2(n10626), .A(n15270), .ZN(n10033) );
  INV_X1 U12703 ( .A(n14998), .ZN(n15006) );
  NAND2_X1 U12704 ( .A1(n10033), .A2(n15006), .ZN(n13200) );
  INV_X1 U12705 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n15378) );
  NAND2_X1 U12706 ( .A1(n10612), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n10035) );
  INV_X1 U12707 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n15009) );
  OR2_X1 U12708 ( .A1(n9614), .A2(n15009), .ZN(n10034) );
  OAI211_X1 U12709 ( .C1(n10615), .C2(n15378), .A(n10035), .B(n10034), .ZN(
        n14799) );
  NAND2_X1 U12710 ( .A1(n10869), .A2(n14836), .ZN(n15241) );
  INV_X1 U12711 ( .A(P1_B_REG_SCAN_IN), .ZN(n10036) );
  NOR2_X1 U12712 ( .A1(n15436), .A2(n10036), .ZN(n10037) );
  NOR2_X1 U12713 ( .A1(n15241), .A2(n10037), .ZN(n15001) );
  NAND2_X1 U12714 ( .A1(n14799), .A2(n15001), .ZN(n13203) );
  INV_X1 U12715 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10047) );
  INV_X1 U12716 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10040) );
  MUX2_X1 U12717 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10042), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n10043) );
  NAND2_X1 U12718 ( .A1(n10044), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10045) );
  XNOR2_X1 U12719 ( .A(n10045), .B(P1_IR_REG_25__SCAN_IN), .ZN(n10051) );
  NAND2_X1 U12720 ( .A1(n11775), .A2(n11458), .ZN(n10046) );
  NAND2_X1 U12721 ( .A1(n10869), .A2(n10046), .ZN(n11143) );
  NAND2_X1 U12722 ( .A1(n6612), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10048) );
  XNOR2_X1 U12723 ( .A(n10048), .B(n10047), .ZN(n10868) );
  AND2_X1 U12724 ( .A1(n11143), .A2(n10868), .ZN(n10049) );
  AND2_X1 U12725 ( .A1(n10084), .A2(n10049), .ZN(n10314) );
  INV_X1 U12726 ( .A(n10051), .ZN(n12243) );
  NAND3_X1 U12727 ( .A1(n12243), .A2(P1_B_REG_SCAN_IN), .A3(n12109), .ZN(
        n10052) );
  OAI211_X1 U12728 ( .C1(P1_B_REG_SCAN_IN), .C2(n12109), .A(n10050), .B(n10052), .ZN(n10851) );
  NOR2_X1 U12729 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .ZN(
        n14411) );
  NOR4_X1 U12730 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_30__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n10055) );
  NOR4_X1 U12731 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n10054) );
  NOR4_X1 U12732 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n10053) );
  NAND4_X1 U12733 ( .A1(n14411), .A2(n10055), .A3(n10054), .A4(n10053), .ZN(
        n10061) );
  NOR4_X1 U12734 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10059) );
  NOR4_X1 U12735 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n10058) );
  NOR4_X1 U12736 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n10057) );
  NOR4_X1 U12737 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n10056) );
  NAND4_X1 U12738 ( .A1(n10059), .A2(n10058), .A3(n10057), .A4(n10056), .ZN(
        n10060) );
  NOR2_X1 U12739 ( .A1(n10061), .A2(n10060), .ZN(n10062) );
  NOR2_X1 U12740 ( .A1(n10851), .A2(n10062), .ZN(n10303) );
  INV_X1 U12741 ( .A(n10303), .ZN(n10063) );
  OR2_X1 U12742 ( .A1(n15270), .A2(n11458), .ZN(n11494) );
  INV_X1 U12743 ( .A(n10050), .ZN(n12548) );
  NAND2_X1 U12744 ( .A1(n12548), .A2(n12243), .ZN(n10855) );
  OAI21_X1 U12745 ( .B1(n10851), .B2(P1_D_REG_1__SCAN_IN), .A(n10855), .ZN(
        n10304) );
  NAND4_X1 U12746 ( .A1(n11490), .A2(n10063), .A3(n11494), .A4(n10304), .ZN(
        n10075) );
  INV_X1 U12747 ( .A(n10851), .ZN(n10064) );
  INV_X1 U12748 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10854) );
  NAND2_X1 U12749 ( .A1(n10064), .A2(n10854), .ZN(n10065) );
  NAND2_X1 U12750 ( .A1(n12548), .A2(n12109), .ZN(n10852) );
  NAND2_X1 U12751 ( .A1(n10065), .A2(n10852), .ZN(n11489) );
  INV_X1 U12752 ( .A(n11489), .ZN(n10066) );
  INV_X2 U12753 ( .A(n15549), .ZN(n15550) );
  NAND2_X1 U12754 ( .A1(n15549), .A2(n10067), .ZN(n10068) );
  NAND2_X1 U12755 ( .A1(n10069), .A2(n10068), .ZN(n10074) );
  INV_X1 U12756 ( .A(n10626), .ZN(n10070) );
  AND2_X1 U12757 ( .A1(n11825), .A2(n11890), .ZN(n10670) );
  NAND2_X1 U12758 ( .A1(n10670), .A2(n11127), .ZN(n11497) );
  NAND3_X1 U12759 ( .A1(n11825), .A2(n14993), .A3(n11127), .ZN(n10071) );
  NAND2_X1 U12760 ( .A1(n11497), .A2(n10071), .ZN(n15547) );
  INV_X1 U12761 ( .A(n15547), .ZN(n15327) );
  NOR2_X1 U12762 ( .A1(n15549), .A2(n15327), .ZN(n12478) );
  INV_X1 U12763 ( .A(n12478), .ZN(n10072) );
  NAND2_X1 U12764 ( .A1(n10074), .A2(n10073), .ZN(P1_U3525) );
  INV_X2 U12765 ( .A(n15552), .ZN(n15554) );
  INV_X1 U12766 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n10077) );
  NAND2_X1 U12767 ( .A1(n15552), .A2(n10077), .ZN(n10078) );
  NAND2_X1 U12768 ( .A1(n10079), .A2(n10078), .ZN(n10082) );
  NOR2_X1 U12769 ( .A1(n15552), .A2(n15327), .ZN(n12686) );
  INV_X1 U12770 ( .A(n12686), .ZN(n10080) );
  NAND2_X1 U12771 ( .A1(n10082), .A2(n10081), .ZN(P1_U3557) );
  AND2_X4 U12772 ( .A1(n10117), .A2(n15270), .ZN(n10294) );
  INV_X1 U12773 ( .A(n10084), .ZN(n10085) );
  AOI22_X1 U12774 ( .A1(n10292), .A2(n11128), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n10085), .ZN(n10086) );
  INV_X1 U12775 ( .A(n11156), .ZN(n11154) );
  OR2_X1 U12776 ( .A1(n10252), .A2(n11151), .ZN(n10089) );
  OR2_X1 U12777 ( .A1(n10084), .A2(n10087), .ZN(n10088) );
  NAND2_X1 U12778 ( .A1(n10089), .A2(n10088), .ZN(n10090) );
  NAND2_X1 U12779 ( .A1(n11147), .A2(n10281), .ZN(n10092) );
  NAND2_X1 U12780 ( .A1(n10094), .A2(n10093), .ZN(n10095) );
  XNOR2_X1 U12781 ( .A(n10095), .B(n10297), .ZN(n10100) );
  NAND2_X1 U12782 ( .A1(n10294), .A2(n10096), .ZN(n10098) );
  OR2_X1 U12783 ( .A1(n10299), .A2(n11498), .ZN(n10097) );
  NAND2_X1 U12784 ( .A1(n11296), .A2(n10101), .ZN(n12969) );
  NAND2_X1 U12785 ( .A1(n10191), .A2(n14820), .ZN(n10103) );
  OR2_X1 U12786 ( .A1(n10252), .A2(n7048), .ZN(n10102) );
  NAND2_X1 U12787 ( .A1(n10103), .A2(n10102), .ZN(n10104) );
  XNOR2_X1 U12788 ( .A(n10104), .B(n10297), .ZN(n10107) );
  XNOR2_X1 U12789 ( .A(n10107), .B(n10106), .ZN(n12970) );
  INV_X1 U12790 ( .A(n10106), .ZN(n10108) );
  NAND2_X1 U12791 ( .A1(n10108), .A2(n10107), .ZN(n10109) );
  NAND2_X1 U12792 ( .A1(n10191), .A2(n14819), .ZN(n10111) );
  OR2_X1 U12793 ( .A1(n11545), .A2(n10252), .ZN(n10110) );
  NAND2_X1 U12794 ( .A1(n10111), .A2(n10110), .ZN(n10112) );
  XNOR2_X1 U12795 ( .A(n10112), .B(n10281), .ZN(n10115) );
  OAI22_X1 U12796 ( .A1(n10105), .A2(n9995), .B1(n11545), .B2(n10299), .ZN(
        n10114) );
  XNOR2_X1 U12797 ( .A(n10115), .B(n10114), .ZN(n11537) );
  NAND2_X1 U12798 ( .A1(n10115), .A2(n10114), .ZN(n10116) );
  NAND2_X1 U12799 ( .A1(n11539), .A2(n10116), .ZN(n11826) );
  NAND2_X1 U12800 ( .A1(n11868), .A2(n10287), .ZN(n10119) );
  NAND2_X1 U12801 ( .A1(n10191), .A2(n14817), .ZN(n10118) );
  NAND2_X1 U12802 ( .A1(n10119), .A2(n10118), .ZN(n10120) );
  XNOR2_X1 U12803 ( .A(n10120), .B(n10297), .ZN(n11860) );
  NAND2_X1 U12804 ( .A1(n10294), .A2(n14817), .ZN(n10122) );
  NAND2_X1 U12805 ( .A1(n11868), .A2(n10283), .ZN(n10121) );
  AND2_X1 U12806 ( .A1(n10122), .A2(n10121), .ZN(n11859) );
  NAND2_X1 U12807 ( .A1(n11860), .A2(n11859), .ZN(n11858) );
  NAND2_X1 U12808 ( .A1(n10287), .A2(n11830), .ZN(n10124) );
  NAND2_X1 U12809 ( .A1(n10191), .A2(n14818), .ZN(n10123) );
  NAND2_X1 U12810 ( .A1(n10124), .A2(n10123), .ZN(n10125) );
  XNOR2_X1 U12811 ( .A(n10125), .B(n10297), .ZN(n11829) );
  NAND2_X1 U12812 ( .A1(n10294), .A2(n14818), .ZN(n10127) );
  NAND2_X1 U12813 ( .A1(n10191), .A2(n11830), .ZN(n10126) );
  AND2_X1 U12814 ( .A1(n10127), .A2(n10126), .ZN(n11828) );
  NAND2_X1 U12815 ( .A1(n11829), .A2(n11828), .ZN(n10128) );
  AND2_X1 U12816 ( .A1(n11858), .A2(n10128), .ZN(n10129) );
  NAND2_X1 U12817 ( .A1(n11826), .A2(n10129), .ZN(n10136) );
  INV_X1 U12818 ( .A(n11829), .ZN(n11856) );
  INV_X1 U12819 ( .A(n11828), .ZN(n11855) );
  NAND2_X1 U12820 ( .A1(n11856), .A2(n11855), .ZN(n10130) );
  NAND2_X1 U12821 ( .A1(n10130), .A2(n11859), .ZN(n10134) );
  INV_X1 U12822 ( .A(n11860), .ZN(n10133) );
  INV_X1 U12823 ( .A(n11859), .ZN(n10131) );
  AND2_X1 U12824 ( .A1(n11855), .A2(n10131), .ZN(n10132) );
  AOI22_X1 U12825 ( .A1(n10134), .A2(n10133), .B1(n10132), .B2(n11856), .ZN(
        n10135) );
  NAND2_X1 U12826 ( .A1(n15543), .A2(n10287), .ZN(n10138) );
  NAND2_X1 U12827 ( .A1(n10191), .A2(n14816), .ZN(n10137) );
  NAND2_X1 U12828 ( .A1(n10138), .A2(n10137), .ZN(n10139) );
  XNOR2_X1 U12829 ( .A(n10139), .B(n10297), .ZN(n10141) );
  NAND2_X1 U12830 ( .A1(n15543), .A2(n10283), .ZN(n10140) );
  OAI21_X1 U12831 ( .B1(n10105), .B2(n11903), .A(n10140), .ZN(n10142) );
  XNOR2_X1 U12832 ( .A(n10141), .B(n10142), .ZN(n11817) );
  INV_X1 U12833 ( .A(n10141), .ZN(n10143) );
  NAND2_X1 U12834 ( .A1(n10143), .A2(n10142), .ZN(n10144) );
  NAND2_X1 U12835 ( .A1(n15548), .A2(n10287), .ZN(n10146) );
  NAND2_X1 U12836 ( .A1(n10191), .A2(n14815), .ZN(n10145) );
  NAND2_X1 U12837 ( .A1(n10146), .A2(n10145), .ZN(n10147) );
  XNOR2_X1 U12838 ( .A(n10147), .B(n10281), .ZN(n10148) );
  AOI22_X1 U12839 ( .A1(n15548), .A2(n10283), .B1(n10294), .B2(n14815), .ZN(
        n10149) );
  XNOR2_X1 U12840 ( .A(n10148), .B(n10149), .ZN(n11901) );
  INV_X1 U12841 ( .A(n10148), .ZN(n10150) );
  NAND2_X1 U12842 ( .A1(n12220), .A2(n10287), .ZN(n10152) );
  NAND2_X1 U12843 ( .A1(n10292), .A2(n14814), .ZN(n10151) );
  NAND2_X1 U12844 ( .A1(n10152), .A2(n10151), .ZN(n10153) );
  XNOR2_X1 U12845 ( .A(n10153), .B(n10297), .ZN(n10158) );
  NOR2_X1 U12846 ( .A1(n10105), .A2(n12522), .ZN(n10154) );
  AOI21_X1 U12847 ( .B1(n12220), .B2(n10283), .A(n10154), .ZN(n10157) );
  XNOR2_X1 U12848 ( .A(n10158), .B(n10157), .ZN(n12215) );
  INV_X1 U12849 ( .A(n12215), .ZN(n10155) );
  NAND2_X1 U12850 ( .A1(n10158), .A2(n10157), .ZN(n10159) );
  NAND2_X1 U12851 ( .A1(n14674), .A2(n10287), .ZN(n10161) );
  NAND2_X1 U12852 ( .A1(n10191), .A2(n14812), .ZN(n10160) );
  NAND2_X1 U12853 ( .A1(n10161), .A2(n10160), .ZN(n10162) );
  XNOR2_X1 U12854 ( .A(n10162), .B(n10281), .ZN(n14667) );
  NAND2_X1 U12855 ( .A1(n14674), .A2(n10283), .ZN(n10164) );
  NAND2_X1 U12856 ( .A1(n10294), .A2(n14812), .ZN(n10163) );
  NAND2_X1 U12857 ( .A1(n10164), .A2(n10163), .ZN(n14666) );
  NAND2_X1 U12858 ( .A1(n12516), .A2(n10287), .ZN(n10166) );
  NAND2_X1 U12859 ( .A1(n10292), .A2(n14813), .ZN(n10165) );
  NAND2_X1 U12860 ( .A1(n10166), .A2(n10165), .ZN(n10167) );
  XNOR2_X1 U12861 ( .A(n10167), .B(n10281), .ZN(n12519) );
  NAND2_X1 U12862 ( .A1(n12516), .A2(n10283), .ZN(n10169) );
  NAND2_X1 U12863 ( .A1(n10294), .A2(n14813), .ZN(n10168) );
  NAND2_X1 U12864 ( .A1(n10169), .A2(n10168), .ZN(n12518) );
  OAI22_X1 U12865 ( .A1(n14667), .A2(n14666), .B1(n12519), .B2(n12518), .ZN(
        n12581) );
  NAND2_X1 U12866 ( .A1(n10292), .A2(n14811), .ZN(n10170) );
  NAND2_X1 U12867 ( .A1(n10171), .A2(n10170), .ZN(n10172) );
  XNOR2_X1 U12868 ( .A(n10172), .B(n10281), .ZN(n10176) );
  INV_X1 U12869 ( .A(n10176), .ZN(n10174) );
  NOR2_X1 U12870 ( .A1(n10105), .A2(n12629), .ZN(n10173) );
  AOI21_X1 U12871 ( .B1(n12423), .B2(n10292), .A(n10173), .ZN(n10175) );
  AND2_X1 U12872 ( .A1(n10174), .A2(n10175), .ZN(n10181) );
  XNOR2_X1 U12873 ( .A(n10176), .B(n10175), .ZN(n12587) );
  INV_X1 U12874 ( .A(n12519), .ZN(n10178) );
  INV_X1 U12875 ( .A(n12518), .ZN(n14665) );
  INV_X1 U12876 ( .A(n14666), .ZN(n10177) );
  OAI21_X1 U12877 ( .B1(n10178), .B2(n14665), .A(n10177), .ZN(n10180) );
  AND2_X1 U12878 ( .A1(n14666), .A2(n12518), .ZN(n10179) );
  AOI22_X1 U12879 ( .A1(n10180), .A2(n14667), .B1(n10179), .B2(n12519), .ZN(
        n12582) );
  NAND2_X1 U12880 ( .A1(n12567), .A2(n10287), .ZN(n10183) );
  NAND2_X1 U12881 ( .A1(n10191), .A2(n14810), .ZN(n10182) );
  NAND2_X1 U12882 ( .A1(n10183), .A2(n10182), .ZN(n10184) );
  XNOR2_X1 U12883 ( .A(n10184), .B(n10297), .ZN(n10186) );
  NOR2_X1 U12884 ( .A1(n10105), .A2(n14745), .ZN(n10185) );
  AOI21_X1 U12885 ( .B1(n12567), .B2(n10283), .A(n10185), .ZN(n10187) );
  XNOR2_X1 U12886 ( .A(n10186), .B(n10187), .ZN(n12624) );
  INV_X1 U12887 ( .A(n10186), .ZN(n10189) );
  INV_X1 U12888 ( .A(n10187), .ZN(n10188) );
  NAND2_X1 U12889 ( .A1(n10189), .A2(n10188), .ZN(n10190) );
  NAND2_X1 U12890 ( .A1(n12626), .A2(n10190), .ZN(n14742) );
  NAND2_X1 U12891 ( .A1(n12720), .A2(n10287), .ZN(n10193) );
  NAND2_X1 U12892 ( .A1(n10191), .A2(n14809), .ZN(n10192) );
  NAND2_X1 U12893 ( .A1(n10193), .A2(n10192), .ZN(n10194) );
  XNOR2_X1 U12894 ( .A(n10194), .B(n10281), .ZN(n10198) );
  NOR2_X1 U12895 ( .A1(n10105), .A2(n7287), .ZN(n10195) );
  AOI21_X1 U12896 ( .B1(n12720), .B2(n10292), .A(n10195), .ZN(n10196) );
  XNOR2_X1 U12897 ( .A(n10198), .B(n10196), .ZN(n14741) );
  INV_X1 U12898 ( .A(n10196), .ZN(n10197) );
  NAND2_X1 U12899 ( .A1(n10198), .A2(n10197), .ZN(n10199) );
  NAND2_X1 U12900 ( .A1(n12770), .A2(n10287), .ZN(n10201) );
  NAND2_X1 U12901 ( .A1(n15256), .A2(n10283), .ZN(n10200) );
  NAND2_X1 U12902 ( .A1(n10201), .A2(n10200), .ZN(n10202) );
  XNOR2_X1 U12903 ( .A(n10202), .B(n10281), .ZN(n10204) );
  NOR2_X1 U12904 ( .A1(n14788), .A2(n10105), .ZN(n10203) );
  XNOR2_X1 U12905 ( .A(n10204), .B(n10205), .ZN(n14650) );
  INV_X1 U12906 ( .A(n10204), .ZN(n10206) );
  NAND2_X1 U12907 ( .A1(n10206), .A2(n10205), .ZN(n10207) );
  NAND2_X1 U12908 ( .A1(n15271), .A2(n10287), .ZN(n10209) );
  NAND2_X1 U12909 ( .A1(n14808), .A2(n10283), .ZN(n10208) );
  NAND2_X1 U12910 ( .A1(n10209), .A2(n10208), .ZN(n10210) );
  XNOR2_X1 U12911 ( .A(n10210), .B(n10297), .ZN(n10211) );
  OAI22_X1 U12912 ( .A1(n15414), .A2(n10299), .B1(n15240), .B2(n10105), .ZN(
        n14785) );
  NAND2_X1 U12913 ( .A1(n15351), .A2(n10287), .ZN(n10214) );
  NAND2_X1 U12914 ( .A1(n15259), .A2(n10283), .ZN(n10213) );
  NAND2_X1 U12915 ( .A1(n10214), .A2(n10213), .ZN(n10215) );
  XNOR2_X1 U12916 ( .A(n10215), .B(n10281), .ZN(n10216) );
  AOI22_X1 U12917 ( .A1(n15351), .A2(n10283), .B1(n10294), .B2(n15259), .ZN(
        n10217) );
  XNOR2_X1 U12918 ( .A(n10216), .B(n10217), .ZN(n14708) );
  INV_X1 U12919 ( .A(n10216), .ZN(n10218) );
  AOI22_X1 U12920 ( .A1(n15345), .A2(n10283), .B1(n10294), .B2(n14807), .ZN(
        n10222) );
  NAND2_X1 U12921 ( .A1(n15345), .A2(n10287), .ZN(n10220) );
  NAND2_X1 U12922 ( .A1(n14807), .A2(n10283), .ZN(n10219) );
  NAND2_X1 U12923 ( .A1(n10220), .A2(n10219), .ZN(n10221) );
  XNOR2_X1 U12924 ( .A(n10221), .B(n10281), .ZN(n10224) );
  XOR2_X1 U12925 ( .A(n10222), .B(n10224), .Z(n14715) );
  INV_X1 U12926 ( .A(n10222), .ZN(n10223) );
  INV_X1 U12927 ( .A(n15199), .ZN(n15202) );
  OAI22_X1 U12928 ( .A1(n15202), .A2(n10299), .B1(n10225), .B2(n10105), .ZN(
        n10230) );
  NAND2_X1 U12929 ( .A1(n15199), .A2(n10287), .ZN(n10227) );
  NAND2_X1 U12930 ( .A1(n14806), .A2(n10283), .ZN(n10226) );
  NAND2_X1 U12931 ( .A1(n10227), .A2(n10226), .ZN(n10228) );
  XNOR2_X1 U12932 ( .A(n10228), .B(n10281), .ZN(n10229) );
  XOR2_X1 U12933 ( .A(n10230), .B(n10229), .Z(n14765) );
  INV_X1 U12934 ( .A(n10229), .ZN(n10232) );
  INV_X1 U12935 ( .A(n10230), .ZN(n10231) );
  NAND2_X1 U12936 ( .A1(n15332), .A2(n10287), .ZN(n10234) );
  NAND2_X1 U12937 ( .A1(n14805), .A2(n10283), .ZN(n10233) );
  NAND2_X1 U12938 ( .A1(n10234), .A2(n10233), .ZN(n10235) );
  XNOR2_X1 U12939 ( .A(n10235), .B(n10281), .ZN(n10237) );
  AND2_X1 U12940 ( .A1(n14805), .A2(n10294), .ZN(n10236) );
  AOI21_X1 U12941 ( .B1(n15332), .B2(n10283), .A(n10236), .ZN(n10238) );
  XNOR2_X1 U12942 ( .A(n10237), .B(n10238), .ZN(n14681) );
  INV_X1 U12943 ( .A(n10238), .ZN(n10239) );
  NAND2_X1 U12944 ( .A1(n10237), .A2(n10239), .ZN(n10240) );
  NAND2_X1 U12945 ( .A1(n15171), .A2(n10287), .ZN(n10242) );
  NAND2_X1 U12946 ( .A1(n14804), .A2(n10283), .ZN(n10241) );
  NAND2_X1 U12947 ( .A1(n10242), .A2(n10241), .ZN(n10243) );
  XNOR2_X1 U12948 ( .A(n10243), .B(n10281), .ZN(n10246) );
  AOI22_X1 U12949 ( .A1(n15171), .A2(n10283), .B1(n10294), .B2(n14804), .ZN(
        n10244) );
  XNOR2_X1 U12950 ( .A(n10246), .B(n10244), .ZN(n14734) );
  INV_X1 U12951 ( .A(n10244), .ZN(n10245) );
  AND2_X1 U12952 ( .A1(n10246), .A2(n10245), .ZN(n10247) );
  AOI22_X1 U12953 ( .A1(n15151), .A2(n10283), .B1(n10294), .B2(n15122), .ZN(
        n10250) );
  AOI22_X1 U12954 ( .A1(n15151), .A2(n10287), .B1(n10283), .B2(n15122), .ZN(
        n10248) );
  XNOR2_X1 U12955 ( .A(n10248), .B(n10281), .ZN(n10249) );
  XOR2_X1 U12956 ( .A(n10250), .B(n10249), .Z(n14689) );
  NAND2_X1 U12957 ( .A1(n10249), .A2(n10250), .ZN(n10251) );
  OAI22_X1 U12958 ( .A1(n15404), .A2(n10299), .B1(n14691), .B2(n10105), .ZN(
        n10254) );
  OAI22_X1 U12959 ( .A1(n15404), .A2(n10252), .B1(n14691), .B2(n10299), .ZN(
        n10253) );
  XNOR2_X1 U12960 ( .A(n10253), .B(n10281), .ZN(n10255) );
  XOR2_X1 U12961 ( .A(n10254), .B(n10255), .Z(n14753) );
  NAND2_X1 U12962 ( .A1(n15113), .A2(n10287), .ZN(n10258) );
  NAND2_X1 U12963 ( .A1(n15089), .A2(n10283), .ZN(n10257) );
  NAND2_X1 U12964 ( .A1(n10258), .A2(n10257), .ZN(n10259) );
  XNOR2_X1 U12965 ( .A(n10259), .B(n10281), .ZN(n10262) );
  AOI22_X1 U12966 ( .A1(n15113), .A2(n10283), .B1(n10294), .B2(n15089), .ZN(
        n10260) );
  XNOR2_X1 U12967 ( .A(n10262), .B(n10260), .ZN(n14659) );
  INV_X1 U12968 ( .A(n10260), .ZN(n10261) );
  OR2_X1 U12969 ( .A1(n10262), .A2(n10261), .ZN(n10263) );
  NAND2_X1 U12970 ( .A1(n10264), .A2(n10263), .ZN(n14721) );
  NAND2_X1 U12971 ( .A1(n15099), .A2(n10287), .ZN(n10266) );
  NAND2_X1 U12972 ( .A1(n14802), .A2(n10283), .ZN(n10265) );
  NAND2_X1 U12973 ( .A1(n10266), .A2(n10265), .ZN(n10267) );
  XNOR2_X1 U12974 ( .A(n10267), .B(n10281), .ZN(n10270) );
  AOI22_X1 U12975 ( .A1(n15099), .A2(n10283), .B1(n10294), .B2(n14802), .ZN(
        n10268) );
  XNOR2_X1 U12976 ( .A(n10270), .B(n10268), .ZN(n14722) );
  INV_X1 U12977 ( .A(n10268), .ZN(n10269) );
  NAND2_X1 U12978 ( .A1(n15298), .A2(n10287), .ZN(n10273) );
  NAND2_X1 U12979 ( .A1(n15090), .A2(n10283), .ZN(n10272) );
  NAND2_X1 U12980 ( .A1(n10273), .A2(n10272), .ZN(n10274) );
  XNOR2_X1 U12981 ( .A(n10274), .B(n10281), .ZN(n10275) );
  AOI22_X1 U12982 ( .A1(n15298), .A2(n10283), .B1(n10294), .B2(n15090), .ZN(
        n10276) );
  XNOR2_X1 U12983 ( .A(n10275), .B(n10276), .ZN(n14700) );
  INV_X1 U12984 ( .A(n10275), .ZN(n10277) );
  NAND2_X1 U12985 ( .A1(n10277), .A2(n10276), .ZN(n10278) );
  NAND2_X1 U12986 ( .A1(n15053), .A2(n10287), .ZN(n10280) );
  NAND2_X1 U12987 ( .A1(n15037), .A2(n10283), .ZN(n10279) );
  NAND2_X1 U12988 ( .A1(n10280), .A2(n10279), .ZN(n10282) );
  XNOR2_X1 U12989 ( .A(n10282), .B(n10281), .ZN(n10284) );
  AOI22_X1 U12990 ( .A1(n15053), .A2(n10283), .B1(n10294), .B2(n15037), .ZN(
        n10285) );
  XNOR2_X1 U12991 ( .A(n10284), .B(n10285), .ZN(n14774) );
  INV_X1 U12992 ( .A(n10284), .ZN(n10286) );
  NAND2_X1 U12993 ( .A1(n15042), .A2(n10287), .ZN(n10289) );
  NAND2_X1 U12994 ( .A1(n14801), .A2(n10283), .ZN(n10288) );
  NAND2_X1 U12995 ( .A1(n10289), .A2(n10288), .ZN(n10290) );
  XNOR2_X1 U12996 ( .A(n10290), .B(n10297), .ZN(n10319) );
  AND2_X1 U12997 ( .A1(n14801), .A2(n10294), .ZN(n10291) );
  AOI21_X1 U12998 ( .B1(n15042), .B2(n10292), .A(n10291), .ZN(n10318) );
  XNOR2_X1 U12999 ( .A(n10319), .B(n10318), .ZN(n12960) );
  INV_X1 U13000 ( .A(n12960), .ZN(n10293) );
  NAND2_X1 U13001 ( .A1(n12961), .A2(n10293), .ZN(n10329) );
  NAND2_X1 U13002 ( .A1(n15023), .A2(n10283), .ZN(n10296) );
  NAND2_X1 U13003 ( .A1(n15038), .A2(n10294), .ZN(n10295) );
  NAND2_X1 U13004 ( .A1(n10296), .A2(n10295), .ZN(n10298) );
  XNOR2_X1 U13005 ( .A(n10298), .B(n10297), .ZN(n10302) );
  NOR2_X1 U13006 ( .A1(n12964), .A2(n10299), .ZN(n10300) );
  AOI21_X1 U13007 ( .B1(n15023), .B2(n10287), .A(n10300), .ZN(n10301) );
  XNOR2_X1 U13008 ( .A(n10302), .B(n10301), .ZN(n10325) );
  INV_X1 U13009 ( .A(n10325), .ZN(n10308) );
  OR2_X1 U13010 ( .A1(n10304), .A2(n10303), .ZN(n11491) );
  NOR2_X1 U13011 ( .A1(n11491), .A2(n11489), .ZN(n10312) );
  INV_X1 U13012 ( .A(n11496), .ZN(n10306) );
  INV_X1 U13013 ( .A(n10869), .ZN(n10644) );
  NAND2_X1 U13014 ( .A1(n15327), .A2(n10644), .ZN(n10305) );
  NOR2_X1 U13015 ( .A1(n10306), .A2(n10305), .ZN(n10307) );
  NAND2_X1 U13016 ( .A1(n10312), .A2(n10307), .ZN(n14797) );
  NAND2_X1 U13017 ( .A1(n10308), .A2(n14754), .ZN(n10328) );
  INV_X1 U13018 ( .A(n10312), .ZN(n10309) );
  NAND2_X1 U13019 ( .A1(n10309), .A2(n11494), .ZN(n10315) );
  NAND2_X1 U13020 ( .A1(n14801), .A2(n15257), .ZN(n10311) );
  NAND2_X1 U13021 ( .A1(n14800), .A2(n15258), .ZN(n10310) );
  AND2_X1 U13022 ( .A1(n10311), .A2(n10310), .ZN(n15018) );
  INV_X1 U13023 ( .A(n10313), .ZN(n15024) );
  NAND2_X1 U13024 ( .A1(n10315), .A2(n10314), .ZN(n10316) );
  AOI22_X1 U13025 ( .A1(n15024), .A2(n14776), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10317) );
  OAI21_X1 U13026 ( .B1(n15018), .B2(n14778), .A(n10317), .ZN(n10321) );
  NAND2_X1 U13027 ( .A1(n10319), .A2(n10318), .ZN(n10322) );
  NOR3_X1 U13028 ( .A1(n10325), .A2(n14797), .A3(n10322), .ZN(n10320) );
  AOI211_X1 U13029 ( .C1(n14795), .C2(n15023), .A(n10321), .B(n10320), .ZN(
        n10327) );
  INV_X1 U13030 ( .A(n10322), .ZN(n10323) );
  NOR2_X1 U13031 ( .A1(n10323), .A2(n14797), .ZN(n10324) );
  AND2_X1 U13032 ( .A1(n10325), .A2(n10324), .ZN(n10326) );
  NAND2_X1 U13033 ( .A1(n9515), .A2(n15649), .ZN(n11706) );
  NAND3_X1 U13034 ( .A1(n10753), .A2(n11705), .A3(n11706), .ZN(n10335) );
  INV_X1 U13035 ( .A(n10331), .ZN(n10332) );
  NAND2_X1 U13036 ( .A1(n10332), .A2(n11706), .ZN(n10334) );
  INV_X1 U13037 ( .A(n11710), .ZN(n10333) );
  NAND3_X1 U13038 ( .A1(n10335), .A2(n10334), .A3(n10333), .ZN(n11707) );
  NAND2_X1 U13039 ( .A1(n11982), .A2(n12264), .ZN(n10336) );
  INV_X1 U13040 ( .A(n13977), .ZN(n10387) );
  INV_X1 U13041 ( .A(n13976), .ZN(n10389) );
  NAND2_X1 U13042 ( .A1(n7628), .A2(n10389), .ZN(n10338) );
  NAND2_X1 U13043 ( .A1(n11907), .A2(n10338), .ZN(n12049) );
  INV_X1 U13044 ( .A(n10390), .ZN(n12053) );
  INV_X1 U13045 ( .A(n13975), .ZN(n11571) );
  NAND2_X1 U13046 ( .A1(n11571), .A2(n12104), .ZN(n10339) );
  AND2_X1 U13047 ( .A1(n12445), .A2(n13973), .ZN(n12398) );
  INV_X1 U13048 ( .A(n12402), .ZN(n10343) );
  INV_X1 U13049 ( .A(n12445), .ZN(n12442) );
  NOR2_X1 U13050 ( .A1(n15624), .A2(n13974), .ZN(n10340) );
  INV_X1 U13051 ( .A(n10340), .ZN(n12368) );
  NAND2_X1 U13052 ( .A1(n12368), .A2(n13973), .ZN(n10341) );
  INV_X1 U13053 ( .A(n13973), .ZN(n10392) );
  AOI22_X1 U13054 ( .A1(n12442), .A2(n10341), .B1(n10340), .B2(n10392), .ZN(
        n10342) );
  OR2_X1 U13055 ( .A1(n12735), .A2(n14329), .ZN(n10345) );
  NAND2_X1 U13056 ( .A1(n14571), .A2(n13970), .ZN(n10346) );
  OR2_X1 U13057 ( .A1(n14571), .A2(n13970), .ZN(n10347) );
  NAND2_X1 U13058 ( .A1(n12609), .A2(n13969), .ZN(n10348) );
  NAND2_X1 U13059 ( .A1(n12678), .A2(n13968), .ZN(n10350) );
  NAND2_X1 U13060 ( .A1(n14562), .A2(n13967), .ZN(n10351) );
  OR2_X1 U13061 ( .A1(n14313), .A2(n14284), .ZN(n10353) );
  NAND2_X1 U13062 ( .A1(n14546), .A2(n13966), .ZN(n10354) );
  INV_X1 U13063 ( .A(n14287), .ZN(n13928) );
  NAND2_X1 U13064 ( .A1(n10354), .A2(n13928), .ZN(n10355) );
  INV_X1 U13065 ( .A(n10354), .ZN(n14259) );
  AOI22_X1 U13066 ( .A1(n14275), .A2(n10355), .B1(n14259), .B2(n14287), .ZN(
        n10356) );
  AND2_X1 U13067 ( .A1(n14260), .A2(n10356), .ZN(n10357) );
  OR2_X1 U13068 ( .A1(n14537), .A2(n13965), .ZN(n14214) );
  OAI21_X1 U13069 ( .B1(n14232), .B2(n14207), .A(n14214), .ZN(n10358) );
  AND2_X1 U13070 ( .A1(n14232), .A2(n14207), .ZN(n14215) );
  AOI21_X1 U13071 ( .B1(n14393), .B2(n13964), .A(n14215), .ZN(n10360) );
  OR2_X1 U13072 ( .A1(n14196), .A2(n14206), .ZN(n10361) );
  NAND2_X1 U13073 ( .A1(n14180), .A2(n14159), .ZN(n10362) );
  AND2_X1 U13074 ( .A1(n14378), .A2(n13963), .ZN(n10363) );
  OR2_X1 U13075 ( .A1(n14378), .A2(n13963), .ZN(n10364) );
  NAND2_X1 U13076 ( .A1(n14149), .A2(n14160), .ZN(n10366) );
  OR2_X1 U13077 ( .A1(n14135), .A2(n13962), .ZN(n10367) );
  NAND2_X1 U13078 ( .A1(n14131), .A2(n10367), .ZN(n10369) );
  NAND2_X1 U13079 ( .A1(n14135), .A2(n13962), .ZN(n10368) );
  AND2_X1 U13080 ( .A1(n14113), .A2(n14125), .ZN(n10370) );
  OR2_X1 U13081 ( .A1(n14113), .A2(n14125), .ZN(n10371) );
  NAND2_X1 U13082 ( .A1(n14356), .A2(n13961), .ZN(n10374) );
  XNOR2_X1 U13083 ( .A(n10377), .B(n10430), .ZN(n10378) );
  NAND2_X1 U13084 ( .A1(n10378), .A2(n11455), .ZN(n11986) );
  INV_X1 U13085 ( .A(n15653), .ZN(n15660) );
  AOI21_X1 U13086 ( .B1(n14096), .B2(n14087), .A(n14320), .ZN(n10380) );
  NAND2_X1 U13087 ( .A1(n10380), .A2(n10461), .ZN(n14089) );
  INV_X1 U13088 ( .A(n10413), .ZN(n10381) );
  OR2_X1 U13089 ( .A1(n14289), .A2(n10381), .ZN(n14244) );
  NAND2_X1 U13090 ( .A1(n14313), .A2(n13882), .ZN(n14242) );
  INV_X1 U13091 ( .A(n14242), .ZN(n10382) );
  INV_X1 U13092 ( .A(n10411), .ZN(n10383) );
  NAND2_X1 U13093 ( .A1(n10749), .A2(n10384), .ZN(n11980) );
  NAND2_X1 U13094 ( .A1(n11980), .A2(n10332), .ZN(n11981) );
  NAND2_X1 U13095 ( .A1(n11981), .A2(n10385), .ZN(n11711) );
  NAND2_X1 U13096 ( .A1(n11711), .A2(n11710), .ZN(n11709) );
  NAND2_X1 U13097 ( .A1(n11982), .A2(n13827), .ZN(n10386) );
  NAND2_X1 U13098 ( .A1(n11709), .A2(n10386), .ZN(n11932) );
  NAND2_X1 U13099 ( .A1(n10387), .A2(n15657), .ZN(n10388) );
  NAND2_X1 U13100 ( .A1(n10389), .A2(n11914), .ZN(n12052) );
  NAND2_X1 U13101 ( .A1(n12445), .A2(n10392), .ZN(n10391) );
  OAI21_X1 U13102 ( .B1(n12375), .B2(n13974), .A(n10391), .ZN(n10397) );
  OAI21_X1 U13103 ( .B1(n15624), .B2(n12372), .A(n10392), .ZN(n10395) );
  NAND2_X1 U13104 ( .A1(n13974), .A2(n13973), .ZN(n10393) );
  NOR2_X1 U13105 ( .A1(n15624), .A2(n10393), .ZN(n10394) );
  AOI21_X1 U13106 ( .B1(n12442), .B2(n10395), .A(n10394), .ZN(n10396) );
  NAND2_X1 U13107 ( .A1(n14571), .A2(n10398), .ZN(n10404) );
  INV_X1 U13108 ( .A(n14329), .ZN(n10400) );
  NAND2_X1 U13109 ( .A1(n12735), .A2(n10400), .ZN(n14331) );
  NAND4_X1 U13110 ( .A1(n12403), .A2(n12402), .A3(n10404), .A4(n14331), .ZN(
        n10406) );
  INV_X1 U13111 ( .A(n13971), .ZN(n10399) );
  NOR2_X1 U13112 ( .A1(n12409), .A2(n10399), .ZN(n12727) );
  INV_X1 U13113 ( .A(n12727), .ZN(n10401) );
  NAND2_X1 U13114 ( .A1(n10401), .A2(n10400), .ZN(n10402) );
  AOI22_X1 U13115 ( .A1(n14628), .A2(n10402), .B1(n12727), .B2(n14329), .ZN(
        n10403) );
  NAND2_X1 U13116 ( .A1(n14336), .A2(n10403), .ZN(n14334) );
  NAND2_X1 U13117 ( .A1(n14334), .A2(n10404), .ZN(n10405) );
  NAND2_X1 U13118 ( .A1(n10406), .A2(n10405), .ZN(n12574) );
  INV_X1 U13119 ( .A(n13969), .ZN(n12674) );
  NAND2_X1 U13120 ( .A1(n12609), .A2(n12674), .ZN(n10407) );
  OR2_X1 U13121 ( .A1(n12609), .A2(n12674), .ZN(n10408) );
  OR2_X1 U13122 ( .A1(n14562), .A2(n12675), .ZN(n10410) );
  NAND2_X1 U13123 ( .A1(n12814), .A2(n10410), .ZN(n14241) );
  NAND2_X1 U13124 ( .A1(n14562), .A2(n12675), .ZN(n14240) );
  AND2_X1 U13125 ( .A1(n14240), .A2(n10411), .ZN(n10412) );
  NAND2_X1 U13126 ( .A1(n14241), .A2(n10412), .ZN(n10416) );
  INV_X1 U13127 ( .A(n13966), .ZN(n10414) );
  OR2_X1 U13128 ( .A1(n14546), .A2(n10414), .ZN(n14269) );
  OR2_X1 U13129 ( .A1(n10381), .A2(n14269), .ZN(n14267) );
  OR2_X1 U13130 ( .A1(n14275), .A2(n13928), .ZN(n10415) );
  AND2_X1 U13131 ( .A1(n14267), .A2(n10415), .ZN(n14245) );
  NAND2_X1 U13132 ( .A1(n14537), .A2(n13836), .ZN(n10417) );
  OR2_X1 U13133 ( .A1(n14232), .A2(n13929), .ZN(n10418) );
  NAND2_X1 U13134 ( .A1(n14393), .A2(n14189), .ZN(n10419) );
  OR2_X1 U13135 ( .A1(n14180), .A2(n14191), .ZN(n10423) );
  NAND2_X1 U13136 ( .A1(n14378), .A2(n13919), .ZN(n14121) );
  INV_X1 U13137 ( .A(n14160), .ZN(n14127) );
  NAND2_X1 U13138 ( .A1(n14149), .A2(n14127), .ZN(n14122) );
  NAND2_X1 U13139 ( .A1(n14594), .A2(n14160), .ZN(n10424) );
  INV_X1 U13140 ( .A(n13962), .ZN(n14109) );
  NAND2_X1 U13141 ( .A1(n14135), .A2(n14109), .ZN(n10427) );
  NAND2_X1 U13142 ( .A1(n14113), .A2(n13871), .ZN(n10429) );
  NAND2_X1 U13143 ( .A1(n10430), .A2(n14070), .ZN(n10431) );
  OAI21_X2 U13144 ( .B1(n9533), .B2(n11815), .A(n10431), .ZN(n14339) );
  OAI21_X1 U13145 ( .B1(n10433), .B2(n10432), .A(n14339), .ZN(n10434) );
  NAND2_X1 U13146 ( .A1(n13961), .A2(n14285), .ZN(n10436) );
  NAND2_X1 U13147 ( .A1(n13960), .A2(n14286), .ZN(n10435) );
  AND2_X1 U13148 ( .A1(n10436), .A2(n10435), .ZN(n13847) );
  INV_X1 U13149 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10442) );
  NAND3_X1 U13150 ( .A1(n15645), .A2(n15641), .A3(n10439), .ZN(n10448) );
  INV_X2 U13151 ( .A(n15664), .ZN(n15666) );
  MUX2_X1 U13152 ( .A(n10442), .B(n10441), .S(n15666), .Z(n10443) );
  NAND2_X1 U13153 ( .A1(n15666), .A2(n15656), .ZN(n14627) );
  NAND2_X1 U13154 ( .A1(n10443), .A2(n7781), .ZN(P2_U3495) );
  INV_X1 U13155 ( .A(n10448), .ZN(n10451) );
  INV_X1 U13156 ( .A(n10449), .ZN(n10450) );
  NAND2_X1 U13157 ( .A1(n10451), .A2(n10450), .ZN(n10452) );
  NAND2_X1 U13158 ( .A1(n10453), .A2(n11596), .ZN(n10759) );
  AND2_X1 U13159 ( .A1(n11986), .A2(n10759), .ZN(n10454) );
  NOR2_X1 U13160 ( .A1(n10455), .A2(n7780), .ZN(n10457) );
  NAND2_X1 U13161 ( .A1(n14093), .A2(n14285), .ZN(n10460) );
  NAND2_X1 U13162 ( .A1(n10458), .A2(n13959), .ZN(n10459) );
  AOI211_X1 U13163 ( .C1(n7611), .C2(n10461), .A(n14320), .B(n14078), .ZN(
        n14351) );
  INV_X1 U13164 ( .A(n10462), .ZN(n10463) );
  OR2_X2 U13165 ( .A1(n14341), .A2(n10463), .ZN(n14326) );
  INV_X1 U13166 ( .A(n10464), .ZN(n10465) );
  INV_X1 U13167 ( .A(n15619), .ZN(n14323) );
  AOI22_X1 U13168 ( .A1(n10465), .A2(n14323), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14312), .ZN(n10466) );
  OAI21_X1 U13169 ( .B1(n8853), .B2(n14326), .A(n10466), .ZN(n10467) );
  INV_X1 U13170 ( .A(n10527), .ZN(n10616) );
  NOR2_X1 U13171 ( .A1(n14820), .A2(n6435), .ZN(n10478) );
  NAND2_X1 U13172 ( .A1(n14820), .A2(n6433), .ZN(n10473) );
  NAND2_X1 U13173 ( .A1(n10473), .A2(n7048), .ZN(n10474) );
  OAI22_X1 U13174 ( .A1(n10477), .A2(n10476), .B1(n6435), .B2(n14819), .ZN(
        n10481) );
  NAND3_X1 U13175 ( .A1(n10478), .A2(n9995), .A3(n11259), .ZN(n10479) );
  NAND3_X1 U13176 ( .A1(n10479), .A2(n11545), .A3(n10527), .ZN(n10480) );
  NAND2_X1 U13177 ( .A1(n11156), .A2(n11151), .ZN(n10482) );
  NAND2_X1 U13178 ( .A1(n11150), .A2(n10482), .ZN(n11125) );
  NAND2_X1 U13179 ( .A1(n11125), .A2(n10645), .ZN(n10486) );
  XNOR2_X1 U13180 ( .A(n10483), .B(n10506), .ZN(n10485) );
  INV_X1 U13181 ( .A(n10484), .ZN(n11153) );
  NAND3_X1 U13182 ( .A1(n10486), .A2(n10485), .A3(n11153), .ZN(n10490) );
  NAND3_X1 U13183 ( .A1(n14819), .A2(n11545), .A3(n6434), .ZN(n10491) );
  MUX2_X1 U13184 ( .A(n14818), .B(n11830), .S(n10582), .Z(n10493) );
  MUX2_X1 U13185 ( .A(n14817), .B(n11868), .S(n6435), .Z(n10497) );
  MUX2_X1 U13186 ( .A(n14817), .B(n11868), .S(n10582), .Z(n10495) );
  MUX2_X1 U13187 ( .A(n14816), .B(n15543), .S(n10582), .Z(n10499) );
  MUX2_X1 U13188 ( .A(n14816), .B(n15543), .S(n6435), .Z(n10498) );
  MUX2_X1 U13189 ( .A(n14815), .B(n15548), .S(n6434), .Z(n10502) );
  MUX2_X1 U13190 ( .A(n14815), .B(n15548), .S(n10506), .Z(n10500) );
  MUX2_X1 U13191 ( .A(n14814), .B(n12220), .S(n10506), .Z(n10504) );
  MUX2_X1 U13192 ( .A(n14814), .B(n12220), .S(n6434), .Z(n10503) );
  INV_X1 U13193 ( .A(n10504), .ZN(n10505) );
  MUX2_X1 U13194 ( .A(n14813), .B(n12516), .S(n6434), .Z(n10509) );
  NAND2_X1 U13195 ( .A1(n10510), .A2(n10509), .ZN(n10508) );
  MUX2_X1 U13196 ( .A(n14813), .B(n12516), .S(n10506), .Z(n10507) );
  NAND2_X1 U13197 ( .A1(n10508), .A2(n10507), .ZN(n10512) );
  MUX2_X1 U13198 ( .A(n14812), .B(n14674), .S(n10582), .Z(n10514) );
  MUX2_X1 U13199 ( .A(n14812), .B(n14674), .S(n6434), .Z(n10513) );
  INV_X1 U13200 ( .A(n10514), .ZN(n10515) );
  MUX2_X1 U13201 ( .A(n14811), .B(n12423), .S(n6434), .Z(n10519) );
  NAND2_X1 U13202 ( .A1(n10518), .A2(n10519), .ZN(n10517) );
  MUX2_X1 U13203 ( .A(n14811), .B(n12423), .S(n10582), .Z(n10516) );
  NAND2_X1 U13204 ( .A1(n10517), .A2(n10516), .ZN(n10523) );
  INV_X1 U13205 ( .A(n10518), .ZN(n10521) );
  INV_X1 U13206 ( .A(n10519), .ZN(n10520) );
  NAND2_X1 U13207 ( .A1(n10521), .A2(n10520), .ZN(n10522) );
  NAND2_X1 U13208 ( .A1(n10523), .A2(n10522), .ZN(n10543) );
  MUX2_X1 U13209 ( .A(n14791), .B(n15235), .S(n6434), .Z(n10544) );
  NAND2_X1 U13210 ( .A1(n10544), .A2(n10547), .ZN(n10524) );
  NAND2_X1 U13211 ( .A1(n15351), .A2(n10582), .ZN(n10545) );
  NAND2_X1 U13212 ( .A1(n10524), .A2(n10545), .ZN(n10525) );
  NAND2_X1 U13213 ( .A1(n10525), .A2(n10546), .ZN(n10540) );
  AND2_X1 U13214 ( .A1(n15259), .A2(n6435), .ZN(n10526) );
  NAND2_X1 U13215 ( .A1(n10547), .A2(n10526), .ZN(n10550) );
  MUX2_X1 U13216 ( .A(n10533), .B(n10530), .S(n6435), .Z(n10556) );
  NAND2_X1 U13217 ( .A1(n14809), .A2(n6435), .ZN(n10529) );
  MUX2_X1 U13218 ( .A(n14809), .B(n12720), .S(n6435), .Z(n10555) );
  NAND2_X1 U13219 ( .A1(n12720), .A2(n10582), .ZN(n10528) );
  NAND4_X1 U13220 ( .A1(n12764), .A2(n10529), .A3(n10555), .A4(n10528), .ZN(
        n10538) );
  NAND2_X1 U13221 ( .A1(n10531), .A2(n10530), .ZN(n10532) );
  NAND2_X1 U13222 ( .A1(n10532), .A2(n10582), .ZN(n10537) );
  NAND2_X1 U13223 ( .A1(n10534), .A2(n10533), .ZN(n10535) );
  NAND2_X1 U13224 ( .A1(n10535), .A2(n6434), .ZN(n10536) );
  NAND3_X1 U13225 ( .A1(n10538), .A2(n10537), .A3(n10536), .ZN(n10539) );
  MUX2_X1 U13226 ( .A(n14745), .B(n12755), .S(n10582), .Z(n10558) );
  MUX2_X1 U13227 ( .A(n14810), .B(n12567), .S(n6434), .Z(n10557) );
  NAND2_X1 U13228 ( .A1(n10543), .A2(n10542), .ZN(n10561) );
  INV_X1 U13229 ( .A(n10544), .ZN(n10551) );
  OR3_X1 U13230 ( .A1(n15213), .A2(n10545), .A3(n10551), .ZN(n10549) );
  MUX2_X1 U13231 ( .A(n10547), .B(n10546), .S(n6434), .Z(n10548) );
  OAI211_X1 U13232 ( .C1(n10551), .C2(n10550), .A(n10549), .B(n10548), .ZN(
        n10552) );
  NAND2_X1 U13233 ( .A1(n7287), .A2(n6434), .ZN(n10553) );
  OAI21_X1 U13234 ( .B1(n12720), .B2(n6435), .A(n10553), .ZN(n10554) );
  OAI211_X1 U13235 ( .C1(n10558), .C2(n10557), .A(n12764), .B(n10556), .ZN(
        n10560) );
  XNOR2_X1 U13236 ( .A(n15171), .B(n14804), .ZN(n10566) );
  AND2_X1 U13237 ( .A1(n10570), .A2(n10562), .ZN(n10563) );
  MUX2_X1 U13238 ( .A(n10564), .B(n10563), .S(n6435), .Z(n10565) );
  NAND3_X1 U13239 ( .A1(n10566), .A2(n10565), .A3(n15159), .ZN(n10577) );
  AOI21_X1 U13240 ( .B1(n10570), .B2(n10567), .A(n6434), .ZN(n10572) );
  NAND2_X1 U13241 ( .A1(n14804), .A2(n10582), .ZN(n10569) );
  OR3_X1 U13242 ( .A1(n15159), .A2(n14804), .A3(n10582), .ZN(n10568) );
  OAI21_X1 U13243 ( .B1(n10570), .B2(n10569), .A(n10568), .ZN(n10571) );
  AOI21_X1 U13244 ( .B1(n15328), .B2(n10572), .A(n10571), .ZN(n10575) );
  AOI21_X1 U13245 ( .B1(n15159), .B2(n14804), .A(n10582), .ZN(n10573) );
  NAND2_X1 U13246 ( .A1(n15171), .A2(n10573), .ZN(n10574) );
  MUX2_X1 U13247 ( .A(n15122), .B(n15151), .S(n6433), .Z(n10581) );
  MUX2_X1 U13248 ( .A(n15122), .B(n15151), .S(n10582), .Z(n10579) );
  MUX2_X1 U13249 ( .A(n14803), .B(n15132), .S(n10582), .Z(n10584) );
  MUX2_X1 U13250 ( .A(n14803), .B(n15132), .S(n6434), .Z(n10583) );
  MUX2_X1 U13251 ( .A(n15089), .B(n15113), .S(n6434), .Z(n10586) );
  MUX2_X1 U13252 ( .A(n15089), .B(n15113), .S(n10582), .Z(n10585) );
  MUX2_X1 U13253 ( .A(n14802), .B(n15099), .S(n10506), .Z(n10590) );
  NAND2_X1 U13254 ( .A1(n10589), .A2(n10590), .ZN(n10588) );
  MUX2_X1 U13255 ( .A(n14802), .B(n15099), .S(n6435), .Z(n10587) );
  NAND2_X1 U13256 ( .A1(n10588), .A2(n10587), .ZN(n10594) );
  INV_X1 U13257 ( .A(n10589), .ZN(n10592) );
  INV_X1 U13258 ( .A(n10590), .ZN(n10591) );
  NAND2_X1 U13259 ( .A1(n10592), .A2(n10591), .ZN(n10593) );
  MUX2_X1 U13260 ( .A(n15090), .B(n15298), .S(n6433), .Z(n10597) );
  MUX2_X1 U13261 ( .A(n15090), .B(n15298), .S(n10582), .Z(n10595) );
  INV_X1 U13262 ( .A(n10597), .ZN(n10598) );
  MUX2_X1 U13263 ( .A(n15037), .B(n15053), .S(n10506), .Z(n10600) );
  MUX2_X1 U13264 ( .A(n15037), .B(n15053), .S(n6435), .Z(n10599) );
  MUX2_X1 U13265 ( .A(n14801), .B(n15042), .S(n6433), .Z(n10603) );
  MUX2_X1 U13266 ( .A(n14801), .B(n15042), .S(n10506), .Z(n10601) );
  INV_X1 U13267 ( .A(n10601), .ZN(n10602) );
  MUX2_X1 U13268 ( .A(n12964), .B(n15383), .S(n10582), .Z(n10609) );
  MUX2_X1 U13269 ( .A(n15023), .B(n15038), .S(n10506), .Z(n10607) );
  NAND2_X1 U13270 ( .A1(n13212), .A2(n9902), .ZN(n10611) );
  INV_X1 U13271 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13213) );
  OR2_X1 U13272 ( .A1(n9631), .A2(n13213), .ZN(n10610) );
  INV_X1 U13273 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n15374) );
  NAND2_X1 U13274 ( .A1(n10612), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n10614) );
  INV_X1 U13275 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n15000) );
  OR2_X1 U13276 ( .A1(n9614), .A2(n15000), .ZN(n10613) );
  OAI211_X1 U13277 ( .C1(n10615), .C2(n15374), .A(n10614), .B(n10613), .ZN(
        n15002) );
  NAND2_X1 U13278 ( .A1(n15002), .A2(n6434), .ZN(n10618) );
  NAND2_X1 U13279 ( .A1(n10618), .A2(n10617), .ZN(n10619) );
  AND2_X1 U13280 ( .A1(n10619), .A2(n14799), .ZN(n10620) );
  AOI21_X1 U13281 ( .B1(n15012), .B2(n10506), .A(n10620), .ZN(n10636) );
  INV_X1 U13282 ( .A(n10621), .ZN(n10622) );
  OAI21_X1 U13283 ( .B1(n15002), .B2(n10622), .A(n14799), .ZN(n10623) );
  INV_X1 U13284 ( .A(n10623), .ZN(n10624) );
  MUX2_X1 U13285 ( .A(n10624), .B(n15012), .S(n6434), .Z(n10632) );
  MUX2_X1 U13286 ( .A(n10625), .B(n10070), .S(n10582), .Z(n10629) );
  MUX2_X1 U13287 ( .A(n14800), .B(n10626), .S(n6434), .Z(n10628) );
  AOI22_X1 U13288 ( .A1(n10636), .A2(n10632), .B1(n10629), .B2(n10628), .ZN(
        n10627) );
  INV_X1 U13289 ( .A(n10628), .ZN(n10631) );
  INV_X1 U13290 ( .A(n10629), .ZN(n10630) );
  INV_X1 U13291 ( .A(n10636), .ZN(n10634) );
  INV_X1 U13292 ( .A(n10632), .ZN(n10633) );
  OAI21_X1 U13293 ( .B1(n10635), .B2(n10634), .A(n10633), .ZN(n10638) );
  INV_X1 U13294 ( .A(n10635), .ZN(n10637) );
  NAND2_X1 U13295 ( .A1(n10639), .A2(n9902), .ZN(n10641) );
  INV_X1 U13296 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14473) );
  OR2_X1 U13297 ( .A1(n9631), .A2(n14473), .ZN(n10640) );
  INV_X1 U13298 ( .A(n15376), .ZN(n15004) );
  XNOR2_X1 U13299 ( .A(n15004), .B(n15002), .ZN(n10668) );
  INV_X1 U13300 ( .A(n10668), .ZN(n10648) );
  INV_X1 U13301 ( .A(n10642), .ZN(n10643) );
  NAND2_X1 U13302 ( .A1(n10644), .A2(n10643), .ZN(n10647) );
  NAND2_X1 U13303 ( .A1(n10645), .A2(n14993), .ZN(n10646) );
  AND2_X1 U13304 ( .A1(n10647), .A2(n10646), .ZN(n10671) );
  INV_X1 U13305 ( .A(n10671), .ZN(n10677) );
  NOR2_X1 U13306 ( .A1(n10648), .A2(n10677), .ZN(n10649) );
  INV_X1 U13307 ( .A(n10650), .ZN(n15034) );
  AND4_X1 U13308 ( .A1(n10651), .A2(n11153), .A3(n11125), .A4(n11255), .ZN(
        n10653) );
  NAND4_X1 U13309 ( .A1(n10653), .A2(n11876), .A3(n10652), .A4(n11321), .ZN(
        n10655) );
  NOR3_X1 U13310 ( .A1(n12152), .A2(n10655), .A3(n10654), .ZN(n10656) );
  NAND3_X1 U13311 ( .A1(n12430), .A2(n10656), .A3(n9725), .ZN(n10657) );
  NOR4_X1 U13312 ( .A1(n7521), .A2(n15251), .A3(n12332), .A4(n10657), .ZN(
        n10658) );
  NAND2_X1 U13313 ( .A1(n10658), .A2(n12560), .ZN(n10659) );
  NOR4_X1 U13314 ( .A1(n10659), .A2(n12710), .A3(n15236), .A4(n15213), .ZN(
        n10660) );
  NAND4_X1 U13315 ( .A1(n15158), .A2(n7736), .A3(n15192), .A4(n10660), .ZN(
        n10661) );
  NOR4_X1 U13316 ( .A1(n15071), .A2(n15128), .A3(n10020), .A4(n10661), .ZN(
        n10663) );
  XNOR2_X1 U13317 ( .A(n15099), .B(n14802), .ZN(n15092) );
  NAND4_X1 U13318 ( .A1(n10663), .A2(n15111), .A3(n10662), .A4(n15092), .ZN(
        n10664) );
  NOR3_X1 U13319 ( .A1(n10665), .A2(n15034), .A3(n10664), .ZN(n10667) );
  XNOR2_X1 U13320 ( .A(n15012), .B(n14799), .ZN(n10666) );
  NAND4_X1 U13321 ( .A1(n10668), .A2(n10667), .A3(n15017), .A4(n10666), .ZN(
        n10669) );
  XNOR2_X1 U13322 ( .A(n10669), .B(n11458), .ZN(n10682) );
  INV_X1 U13323 ( .A(n10670), .ZN(n10681) );
  NOR2_X1 U13324 ( .A1(n10671), .A2(n10670), .ZN(n10686) );
  INV_X1 U13325 ( .A(n10686), .ZN(n10672) );
  NOR3_X1 U13326 ( .A1(n15376), .A2(n15002), .A3(n10672), .ZN(n10675) );
  NOR2_X1 U13327 ( .A1(n15376), .A2(n10506), .ZN(n10690) );
  INV_X1 U13328 ( .A(n10690), .ZN(n10674) );
  NOR3_X1 U13329 ( .A1(n10674), .A2(n15002), .A3(n10677), .ZN(n10673) );
  AOI21_X1 U13330 ( .B1(n10675), .B2(n10674), .A(n10673), .ZN(n10680) );
  NAND2_X1 U13331 ( .A1(n15376), .A2(n10582), .ZN(n10687) );
  INV_X1 U13332 ( .A(n10687), .ZN(n10676) );
  XOR2_X1 U13333 ( .A(n10677), .B(n10676), .Z(n10678) );
  NAND3_X1 U13334 ( .A1(n10678), .A2(n15376), .A3(n15002), .ZN(n10679) );
  OAI211_X1 U13335 ( .C1(n10682), .C2(n10681), .A(n10680), .B(n10679), .ZN(
        n10683) );
  NAND2_X1 U13336 ( .A1(n10685), .A2(n10684), .ZN(n10697) );
  INV_X1 U13337 ( .A(n15002), .ZN(n10689) );
  OAI21_X1 U13338 ( .B1(n10687), .B2(n10689), .A(n10686), .ZN(n10688) );
  INV_X1 U13339 ( .A(n10688), .ZN(n10692) );
  NAND2_X1 U13340 ( .A1(n10692), .A2(n10691), .ZN(n10693) );
  NOR2_X1 U13341 ( .A1(n10694), .A2(n10693), .ZN(n10696) );
  OR2_X1 U13342 ( .A1(n10868), .A2(P1_U3086), .ZN(n12046) );
  OAI21_X1 U13343 ( .B1(n10697), .B2(n10696), .A(n10695), .ZN(n10700) );
  INV_X1 U13344 ( .A(n15436), .ZN(n15489) );
  NAND3_X1 U13345 ( .A1(n11490), .A2(n15489), .A3(n15257), .ZN(n10698) );
  OAI211_X1 U13346 ( .C1(n15438), .C2(n12046), .A(n10698), .B(P1_B_REG_SCAN_IN), .ZN(n10699) );
  NAND2_X1 U13347 ( .A1(n10700), .A2(n10699), .ZN(P1_U3242) );
  INV_X1 U13348 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n10702) );
  MUX2_X1 U13349 ( .A(n10702), .B(n10701), .S(n15666), .Z(n10705) );
  NAND2_X1 U13350 ( .A1(n9474), .A2(n10703), .ZN(n10704) );
  NAND2_X1 U13351 ( .A1(n10705), .A2(n10704), .ZN(P2_U3498) );
  INV_X1 U13352 ( .A(n10706), .ZN(n11043) );
  NOR2_X1 U13353 ( .A1(n10707), .A2(n11043), .ZN(n11046) );
  AND2_X1 U13354 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11046), .ZN(P2_U3947) );
  INV_X1 U13355 ( .A(n10708), .ZN(n10712) );
  NAND3_X1 U13356 ( .A1(n13434), .A2(n10710), .A3(n10709), .ZN(n10711) );
  INV_X1 U13357 ( .A(n13504), .ZN(n13490) );
  AOI21_X1 U13358 ( .B1(n10712), .B2(n10711), .A(n13490), .ZN(n10725) );
  INV_X1 U13359 ( .A(n10713), .ZN(n10717) );
  NAND3_X1 U13360 ( .A1(n13421), .A2(n10715), .A3(n10714), .ZN(n10716) );
  INV_X1 U13361 ( .A(n13495), .ZN(n13461) );
  AOI21_X1 U13362 ( .B1(n10717), .B2(n10716), .A(n13461), .ZN(n10724) );
  INV_X1 U13363 ( .A(n13509), .ZN(n13407) );
  AOI211_X1 U13364 ( .C1(n10720), .C2(n10719), .A(n13407), .B(n10718), .ZN(
        n10723) );
  NAND2_X1 U13365 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n13229)
         );
  NAND2_X1 U13366 ( .A1(n15671), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n10721) );
  OAI211_X1 U13367 ( .C1(n13486), .C2(n10977), .A(n13229), .B(n10721), .ZN(
        n10722) );
  OR4_X1 U13368 ( .A1(n10725), .A2(n10724), .A3(n10723), .A4(n10722), .ZN(
        P3_U3196) );
  INV_X1 U13369 ( .A(n10856), .ZN(n10726) );
  OR2_X2 U13370 ( .A1(n10084), .A2(n10726), .ZN(n14821) );
  INV_X1 U13371 ( .A(n14821), .ZN(P1_U4016) );
  AOI211_X1 U13372 ( .C1(n10728), .C2(n10727), .A(n13956), .B(n6516), .ZN(
        n10732) );
  INV_X1 U13373 ( .A(n14196), .ZN(n14603) );
  NOR2_X1 U13374 ( .A1(n14603), .A2(n13925), .ZN(n10731) );
  OAI22_X1 U13375 ( .A1(n13941), .A2(n14189), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14435), .ZN(n10730) );
  OAI22_X1 U13376 ( .A1(n14191), .A2(n13908), .B1(n13952), .B2(n14197), .ZN(
        n10729) );
  OR4_X1 U13377 ( .A1(n10732), .A2(n10731), .A3(n10730), .A4(n10729), .ZN(
        P2_U3195) );
  AND2_X1 U13378 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n12167) );
  AOI21_X1 U13379 ( .B1(n15671), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n12167), .ZN(
        n10733) );
  OAI21_X1 U13380 ( .B1(n13486), .B2(n10820), .A(n10733), .ZN(n10746) );
  NAND3_X1 U13381 ( .A1(n11029), .A2(n10735), .A3(n10734), .ZN(n10736) );
  AOI21_X1 U13382 ( .B1(n6620), .B2(n10736), .A(n13490), .ZN(n10745) );
  NAND3_X1 U13383 ( .A1(n11026), .A2(n10738), .A3(n10737), .ZN(n10739) );
  AOI21_X1 U13384 ( .B1(n6621), .B2(n10739), .A(n13461), .ZN(n10744) );
  OR3_X1 U13385 ( .A1(n6994), .A2(n10741), .A3(n10740), .ZN(n10742) );
  AOI21_X1 U13386 ( .B1(n11357), .B2(n10742), .A(n13407), .ZN(n10743) );
  OR4_X1 U13387 ( .A1(n10746), .A2(n10745), .A3(n10744), .A4(n10743), .ZN(
        P3_U3188) );
  NAND2_X1 U13388 ( .A1(n10755), .A2(n10747), .ZN(n10748) );
  NAND2_X1 U13389 ( .A1(n10749), .A2(n10748), .ZN(n10752) );
  NAND2_X1 U13390 ( .A1(n9514), .A2(n14286), .ZN(n10750) );
  OAI21_X1 U13391 ( .B1(n13856), .B2(n14190), .A(n10750), .ZN(n10751) );
  AOI21_X1 U13392 ( .B1(n10752), .B2(n14339), .A(n10751), .ZN(n10757) );
  OAI21_X1 U13393 ( .B1(n10755), .B2(n10754), .A(n10753), .ZN(n10758) );
  INV_X1 U13394 ( .A(n11986), .ZN(n12060) );
  NAND2_X1 U13395 ( .A1(n10758), .A2(n12060), .ZN(n10756) );
  NAND2_X1 U13396 ( .A1(n10757), .A2(n10756), .ZN(n11683) );
  MUX2_X1 U13397 ( .A(n11683), .B(P2_REG2_REG_1__SCAN_IN), .S(n14341), .Z(
        n10762) );
  OAI22_X1 U13398 ( .A1(n14326), .A2(n11690), .B1(n15619), .B2(n13980), .ZN(
        n10761) );
  INV_X1 U13399 ( .A(n10758), .ZN(n11686) );
  OR2_X1 U13400 ( .A1(n14341), .A2(n10759), .ZN(n12069) );
  OAI211_X1 U13401 ( .C1(n11690), .C2(n9354), .A(n14310), .B(n11971), .ZN(
        n11684) );
  OAI22_X1 U13402 ( .A1(n11686), .A2(n12069), .B1(n15627), .B2(n11684), .ZN(
        n10760) );
  OR3_X1 U13403 ( .A1(n10762), .A2(n10761), .A3(n10760), .ZN(P2_U3264) );
  NAND2_X1 U13404 ( .A1(n10774), .A2(n10775), .ZN(n10764) );
  NAND2_X1 U13405 ( .A1(n14823), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10763) );
  NAND2_X1 U13406 ( .A1(n10765), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10768) );
  INV_X1 U13407 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10766) );
  NAND2_X1 U13408 ( .A1(n10766), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n10767) );
  INV_X1 U13409 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15496) );
  XNOR2_X1 U13410 ( .A(n10773), .B(n10772), .ZN(n15486) );
  NAND2_X1 U13411 ( .A1(n15486), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n10779) );
  XNOR2_X1 U13412 ( .A(n10774), .B(n10775), .ZN(n10778) );
  INV_X1 U13413 ( .A(n10775), .ZN(n10776) );
  OAI21_X1 U13414 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n10777), .A(n10776), .ZN(
        n15440) );
  NAND2_X1 U13415 ( .A1(n15440), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n15740) );
  XNOR2_X1 U13416 ( .A(n10778), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(n15739) );
  NOR2_X1 U13417 ( .A1(n15740), .A2(n15739), .ZN(n15738) );
  AOI21_X1 U13418 ( .B1(n10778), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n15738), .ZN(
        n15485) );
  NAND2_X1 U13419 ( .A1(n10779), .A2(n15485), .ZN(n10781) );
  OR2_X1 U13420 ( .A1(n15486), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n10780) );
  NAND2_X1 U13421 ( .A1(n10781), .A2(n10780), .ZN(n15735) );
  INV_X1 U13422 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10783) );
  INV_X1 U13423 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14856) );
  XNOR2_X1 U13424 ( .A(n10782), .B(n14856), .ZN(n15736) );
  OAI21_X1 U13425 ( .B1(n15735), .B2(n10783), .A(n15736), .ZN(n10785) );
  NAND2_X1 U13426 ( .A1(n15735), .A2(n10783), .ZN(n10784) );
  NAND2_X1 U13427 ( .A1(n10785), .A2(n10784), .ZN(n10801) );
  XNOR2_X1 U13428 ( .A(n10802), .B(n10801), .ZN(SUB_1596_U59) );
  NAND2_X1 U13429 ( .A1(n6978), .A2(P1_U3086), .ZN(n15433) );
  INV_X1 U13430 ( .A(n15433), .ZN(n12044) );
  INV_X1 U13431 ( .A(n12044), .ZN(n15426) );
  INV_X1 U13432 ( .A(n10787), .ZN(n10811) );
  AND2_X1 U13433 ( .A1(n10817), .A2(P1_U3086), .ZN(n15424) );
  INV_X2 U13434 ( .A(n15424), .ZN(n15435) );
  OAI222_X1 U13435 ( .A1(n14879), .A2(P1_U3086), .B1(n15426), .B2(n10811), 
        .C1(n10788), .C2(n15435), .ZN(P1_U3350) );
  INV_X1 U13436 ( .A(n10789), .ZN(n10807) );
  OAI222_X1 U13437 ( .A1(n14863), .A2(P1_U3086), .B1(n15426), .B2(n10807), 
        .C1(n10790), .C2(n15435), .ZN(P1_U3352) );
  INV_X1 U13438 ( .A(n14894), .ZN(n10793) );
  INV_X1 U13439 ( .A(n10791), .ZN(n10815) );
  OAI222_X1 U13440 ( .A1(n10793), .A2(P1_U3086), .B1(n15426), .B2(n10815), 
        .C1(n10792), .C2(n15435), .ZN(P1_U3349) );
  INV_X1 U13441 ( .A(n15507), .ZN(n10796) );
  INV_X1 U13442 ( .A(n10794), .ZN(n10809) );
  OAI222_X1 U13443 ( .A1(n10796), .A2(P1_U3086), .B1(n15426), .B2(n10809), 
        .C1(n10795), .C2(n15435), .ZN(P1_U3351) );
  OAI222_X1 U13444 ( .A1(n14843), .A2(P1_U3086), .B1(n15426), .B2(n10813), 
        .C1(n10797), .C2(n15435), .ZN(P1_U3353) );
  OAI222_X1 U13445 ( .A1(n14828), .A2(P1_U3086), .B1(n15426), .B2(n10875), 
        .C1(n10798), .C2(n15435), .ZN(P1_U3354) );
  INV_X1 U13446 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n10800) );
  INV_X1 U13447 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14872) );
  XNOR2_X1 U13448 ( .A(n10890), .B(n14872), .ZN(n10885) );
  NAND2_X1 U13449 ( .A1(n10802), .A2(n10801), .ZN(n10805) );
  INV_X1 U13450 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n13998) );
  NAND2_X1 U13451 ( .A1(n10803), .A2(n13998), .ZN(n10804) );
  INV_X1 U13452 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10883) );
  XNOR2_X1 U13453 ( .A(n10884), .B(n10883), .ZN(SUB_1596_U58) );
  NAND2_X1 U13454 ( .A1(n10817), .A2(P2_U3088), .ZN(n14644) );
  NOR2_X1 U13455 ( .A1(n8650), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14640) );
  OAI222_X1 U13456 ( .A1(n15560), .A2(P2_U3088), .B1(n14644), .B2(n10807), 
        .C1(n10806), .C2(n14646), .ZN(P2_U3324) );
  OAI222_X1 U13457 ( .A1(n14005), .A2(P2_U3088), .B1(n14644), .B2(n10809), 
        .C1(n10808), .C2(n14646), .ZN(P2_U3323) );
  INV_X1 U13458 ( .A(n11087), .ZN(n11142) );
  OAI222_X1 U13459 ( .A1(n11142), .A2(P2_U3088), .B1(n14644), .B2(n10811), 
        .C1(n10810), .C2(n14646), .ZN(P2_U3322) );
  OAI222_X1 U13460 ( .A1(n11071), .A2(P2_U3088), .B1(n14644), .B2(n10813), 
        .C1(n10812), .C2(n14646), .ZN(P2_U3325) );
  INV_X1 U13461 ( .A(n14023), .ZN(n10816) );
  OAI222_X1 U13462 ( .A1(n10816), .A2(P2_U3088), .B1(n14644), .B2(n10815), 
        .C1(n10814), .C2(n14646), .ZN(P2_U3321) );
  INV_X1 U13463 ( .A(SI_6_), .ZN(n10822) );
  NOR2_X1 U13464 ( .A1(n8650), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13801) );
  INV_X1 U13465 ( .A(n10819), .ZN(n10821) );
  OAI222_X1 U13466 ( .A1(n13805), .A2(n10822), .B1(n13808), .B2(n10821), .C1(
        P3_U3151), .C2(n10820), .ZN(P3_U3289) );
  INV_X1 U13467 ( .A(SI_8_), .ZN(n10826) );
  INV_X1 U13468 ( .A(n10823), .ZN(n10825) );
  OAI222_X1 U13469 ( .A1(n13805), .A2(n10826), .B1(n13808), .B2(n10825), .C1(
        P3_U3151), .C2(n10824), .ZN(P3_U3287) );
  INV_X1 U13470 ( .A(n11228), .ZN(n10829) );
  INV_X1 U13471 ( .A(n10827), .ZN(n10831) );
  OAI222_X1 U13472 ( .A1(n10829), .A2(P2_U3088), .B1(n14644), .B2(n10831), 
        .C1(n10828), .C2(n14646), .ZN(P2_U3320) );
  INV_X1 U13473 ( .A(n14911), .ZN(n10832) );
  OAI222_X1 U13474 ( .A1(n10832), .A2(P1_U3086), .B1(n15426), .B2(n10831), 
        .C1(n10830), .C2(n15435), .ZN(P1_U3348) );
  INV_X1 U13475 ( .A(SI_5_), .ZN(n10833) );
  INV_X1 U13476 ( .A(SI_3_), .ZN(n10835) );
  OAI222_X1 U13477 ( .A1(P3_U3151), .A2(n11344), .B1(n13808), .B2(n10836), 
        .C1(n10835), .C2(n13805), .ZN(P3_U3292) );
  OAI222_X1 U13478 ( .A1(n11352), .A2(P3_U3151), .B1(n13808), .B2(n10837), 
        .C1(n14401), .C2(n13805), .ZN(P3_U3288) );
  INV_X1 U13479 ( .A(n10838), .ZN(n10840) );
  OAI222_X1 U13480 ( .A1(P3_U3151), .A2(n11122), .B1(n13808), .B2(n10840), 
        .C1(n10839), .C2(n13805), .ZN(P3_U3293) );
  INV_X1 U13481 ( .A(n10841), .ZN(n10843) );
  OAI222_X1 U13482 ( .A1(n11409), .A2(P3_U3151), .B1(n13808), .B2(n10843), 
        .C1(n10842), .C2(n13805), .ZN(P3_U3294) );
  OAI222_X1 U13483 ( .A1(n10845), .A2(P3_U3151), .B1(n13808), .B2(n10844), 
        .C1(n14402), .C2(n13805), .ZN(P3_U3285) );
  OAI222_X1 U13484 ( .A1(n11849), .A2(P3_U3151), .B1(n13808), .B2(n10847), 
        .C1(n10846), .C2(n13805), .ZN(P3_U3286) );
  OAI222_X1 U13485 ( .A1(n10850), .A2(P3_U3151), .B1(n13808), .B2(n10849), 
        .C1(n10848), .C2(n13805), .ZN(P3_U3284) );
  NAND2_X1 U13486 ( .A1(n11496), .A2(n10851), .ZN(n15539) );
  INV_X1 U13487 ( .A(n10852), .ZN(n10853) );
  AOI22_X1 U13488 ( .A1(n15539), .A2(n10854), .B1(n10853), .B2(n10856), .ZN(
        P1_U3445) );
  INV_X1 U13489 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10858) );
  INV_X1 U13490 ( .A(n10855), .ZN(n10857) );
  AOI22_X1 U13491 ( .A1(n15539), .A2(n10858), .B1(n10857), .B2(n10856), .ZN(
        P1_U3446) );
  NAND2_X1 U13492 ( .A1(n13797), .A2(n10859), .ZN(n10908) );
  AND2_X1 U13493 ( .A1(n10908), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U13494 ( .A1(n10908), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U13495 ( .A1(n10908), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U13496 ( .A1(n10908), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U13497 ( .A1(n10908), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U13498 ( .A1(n10908), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U13499 ( .A1(n10908), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U13500 ( .A1(n10908), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U13501 ( .A1(n10908), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U13502 ( .A1(n10908), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U13503 ( .A1(n10908), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U13504 ( .A1(n10908), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U13505 ( .A1(n10908), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U13506 ( .A1(n10908), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U13507 ( .A1(n10908), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U13508 ( .A1(n10908), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  INV_X1 U13509 ( .A(n10860), .ZN(n10863) );
  OAI222_X1 U13510 ( .A1(n11243), .A2(P2_U3088), .B1(n14644), .B2(n10863), 
        .C1(n10861), .C2(n14646), .ZN(P2_U3319) );
  INV_X1 U13511 ( .A(n10963), .ZN(n10864) );
  OAI222_X1 U13512 ( .A1(n10864), .A2(P1_U3086), .B1(n15426), .B2(n10863), 
        .C1(n10862), .C2(n15435), .ZN(P1_U3347) );
  INV_X1 U13513 ( .A(n13805), .ZN(n13799) );
  AOI222_X1 U13514 ( .A1(n10866), .A2(n13801), .B1(n10865), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n13799), .ZN(n10867) );
  INV_X1 U13515 ( .A(n10867), .ZN(P3_U3291) );
  OR2_X1 U13516 ( .A1(n11496), .A2(n10695), .ZN(n10931) );
  NAND2_X1 U13517 ( .A1(n10869), .A2(n10868), .ZN(n10870) );
  AND2_X1 U13518 ( .A1(n10870), .A2(n9632), .ZN(n10930) );
  INV_X1 U13519 ( .A(n10930), .ZN(n10871) );
  AND2_X1 U13520 ( .A1(n10931), .A2(n10871), .ZN(n15492) );
  NOR2_X1 U13521 ( .A1(n15492), .A2(P1_U4016), .ZN(P1_U3085) );
  OAI222_X1 U13522 ( .A1(P3_U3151), .A2(n10874), .B1(n13808), .B2(n10873), 
        .C1(n10872), .C2(n13805), .ZN(P3_U3283) );
  INV_X1 U13523 ( .A(n14644), .ZN(n12040) );
  INV_X1 U13524 ( .A(n12040), .ZN(n14637) );
  OAI222_X1 U13525 ( .A1(n14646), .A2(n10876), .B1(n14637), .B2(n10875), .C1(
        P2_U3088), .C2(n13983), .ZN(P2_U3326) );
  INV_X1 U13526 ( .A(n11005), .ZN(n10879) );
  INV_X1 U13527 ( .A(n10877), .ZN(n10881) );
  OAI222_X1 U13528 ( .A1(n10879), .A2(P1_U3086), .B1(n15426), .B2(n10881), 
        .C1(n10878), .C2(n15435), .ZN(P1_U3346) );
  OAI222_X1 U13529 ( .A1(n11422), .A2(P2_U3088), .B1(n14644), .B2(n10881), 
        .C1(n10880), .C2(n14646), .ZN(P2_U3318) );
  INV_X1 U13530 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n14483) );
  NAND2_X1 U13531 ( .A1(P3_U3897), .A2(n11554), .ZN(n10882) );
  OAI21_X1 U13532 ( .B1(P3_U3897), .B2(n14483), .A(n10882), .ZN(P3_U3495) );
  NAND2_X1 U13533 ( .A1(n10884), .A2(n10883), .ZN(n10889) );
  INV_X1 U13534 ( .A(n10885), .ZN(n10887) );
  NAND2_X1 U13535 ( .A1(n10887), .A2(n10886), .ZN(n10888) );
  NAND2_X1 U13536 ( .A1(n10890), .A2(n14872), .ZN(n10893) );
  NAND2_X1 U13537 ( .A1(n10891), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10892) );
  NAND2_X1 U13538 ( .A1(n10893), .A2(n10892), .ZN(n10985) );
  XNOR2_X1 U13539 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n10894) );
  XNOR2_X1 U13540 ( .A(n10985), .B(n10894), .ZN(n10895) );
  OAI21_X1 U13541 ( .B1(n10896), .B2(n10895), .A(n10994), .ZN(n10897) );
  INV_X1 U13542 ( .A(n10897), .ZN(SUB_1596_U57) );
  INV_X1 U13543 ( .A(n11462), .ZN(n10900) );
  INV_X1 U13544 ( .A(n10898), .ZN(n10902) );
  OAI222_X1 U13545 ( .A1(n10900), .A2(P2_U3088), .B1(n14644), .B2(n10902), 
        .C1(n10899), .C2(n14646), .ZN(P2_U3317) );
  INV_X1 U13546 ( .A(n14924), .ZN(n10903) );
  OAI222_X1 U13547 ( .A1(n10903), .A2(P1_U3086), .B1(n15426), .B2(n10902), 
        .C1(n10901), .C2(n15435), .ZN(P1_U3345) );
  INV_X1 U13548 ( .A(n12453), .ZN(n12462) );
  INV_X1 U13549 ( .A(n10904), .ZN(n10907) );
  OAI222_X1 U13550 ( .A1(n12462), .A2(P2_U3088), .B1(n14644), .B2(n10907), 
        .C1(n10905), .C2(n14646), .ZN(P2_U3316) );
  INV_X1 U13551 ( .A(n11269), .ZN(n11003) );
  OAI222_X1 U13552 ( .A1(n11003), .A2(P1_U3086), .B1(n15433), .B2(n10907), 
        .C1(n10906), .C2(n15435), .ZN(P1_U3344) );
  AND2_X1 U13553 ( .A1(n10908), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U13554 ( .A1(n10908), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U13555 ( .A1(n10908), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U13556 ( .A1(n10908), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U13557 ( .A1(n10908), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U13558 ( .A1(n10908), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U13559 ( .A1(n10908), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U13560 ( .A1(n10908), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U13561 ( .A1(n10908), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U13562 ( .A1(n10908), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U13563 ( .A1(n10908), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U13564 ( .A1(n10908), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U13565 ( .A1(n10908), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U13566 ( .A1(n10908), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  OAI222_X1 U13567 ( .A1(n13430), .A2(P3_U3151), .B1(n13808), .B2(n10910), 
        .C1(n10909), .C2(n13805), .ZN(P3_U3282) );
  OR2_X1 U13568 ( .A1(n10963), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10956) );
  NAND2_X1 U13569 ( .A1(n10963), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10911) );
  NAND2_X1 U13570 ( .A1(n10956), .A2(n10911), .ZN(n10929) );
  INV_X1 U13571 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10912) );
  AND2_X1 U13572 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10913) );
  INV_X1 U13573 ( .A(n14828), .ZN(n14825) );
  NAND2_X1 U13574 ( .A1(n14825), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10914) );
  NAND2_X1 U13575 ( .A1(n14831), .A2(n10914), .ZN(n14842) );
  INV_X1 U13576 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10915) );
  INV_X1 U13577 ( .A(n14843), .ZN(n14849) );
  NAND2_X1 U13578 ( .A1(n14849), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14865) );
  MUX2_X1 U13579 ( .A(n10917), .B(P1_REG1_REG_3__SCAN_IN), .S(n14863), .Z(
        n10916) );
  OR2_X1 U13580 ( .A1(n14863), .A2(n10917), .ZN(n15502) );
  MUX2_X1 U13581 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10918), .S(n15507), .Z(
        n10919) );
  NAND2_X1 U13582 ( .A1(n15507), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10920) );
  MUX2_X1 U13583 ( .A(n9661), .B(P1_REG1_REG_5__SCAN_IN), .S(n14879), .Z(
        n14876) );
  NAND2_X1 U13584 ( .A1(n14879), .A2(n9661), .ZN(n10921) );
  MUX2_X1 U13585 ( .A(n14895), .B(P1_REG1_REG_6__SCAN_IN), .S(n14894), .Z(
        n10922) );
  NAND2_X1 U13586 ( .A1(n14894), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n14907) );
  MUX2_X1 U13587 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10923), .S(n14911), .Z(
        n10924) );
  AND2_X1 U13588 ( .A1(n14911), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10926) );
  INV_X1 U13589 ( .A(n10926), .ZN(n10925) );
  NAND2_X1 U13590 ( .A1(n14910), .A2(n10925), .ZN(n10928) );
  NOR2_X1 U13591 ( .A1(n10929), .A2(n10926), .ZN(n10927) );
  AOI21_X1 U13592 ( .B1(n10929), .B2(n10928), .A(n10958), .ZN(n10955) );
  NAND2_X1 U13593 ( .A1(n10931), .A2(n10930), .ZN(n15494) );
  NOR2_X2 U13594 ( .A1(n15494), .A2(n15489), .ZN(n15506) );
  INV_X1 U13595 ( .A(n15506), .ZN(n14942) );
  NOR2_X2 U13596 ( .A1(n15494), .A2(n14839), .ZN(n15500) );
  INV_X1 U13597 ( .A(n15492), .ZN(n15497) );
  INV_X1 U13598 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n11653) );
  NAND2_X1 U13599 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n12218) );
  OAI21_X1 U13600 ( .B1(n15497), .B2(n11653), .A(n12218), .ZN(n10932) );
  AOI21_X1 U13601 ( .B1(n10963), .B2(n15500), .A(n10932), .ZN(n10954) );
  INV_X1 U13602 ( .A(n15494), .ZN(n10934) );
  NOR2_X1 U13603 ( .A1(n14836), .A2(n15436), .ZN(n10933) );
  NAND2_X1 U13604 ( .A1(n10934), .A2(n10933), .ZN(n14989) );
  MUX2_X1 U13605 ( .A(n11501), .B(P1_REG2_REG_1__SCAN_IN), .S(n14828), .Z(
        n14827) );
  AND2_X1 U13606 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14838) );
  NAND2_X1 U13607 ( .A1(n14827), .A2(n14838), .ZN(n14826) );
  NAND2_X1 U13608 ( .A1(n14825), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10935) );
  NAND2_X1 U13609 ( .A1(n14826), .A2(n10935), .ZN(n14850) );
  MUX2_X1 U13610 ( .A(n10936), .B(P1_REG2_REG_2__SCAN_IN), .S(n14843), .Z(
        n14851) );
  NAND2_X1 U13611 ( .A1(n14850), .A2(n14851), .ZN(n14861) );
  NAND2_X1 U13612 ( .A1(n14849), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14860) );
  NAND2_X1 U13613 ( .A1(n14861), .A2(n14860), .ZN(n10938) );
  MUX2_X1 U13614 ( .A(n10939), .B(P1_REG2_REG_3__SCAN_IN), .S(n14863), .Z(
        n10937) );
  NAND2_X1 U13615 ( .A1(n10938), .A2(n10937), .ZN(n15510) );
  OR2_X1 U13616 ( .A1(n14863), .A2(n10939), .ZN(n15509) );
  NAND2_X1 U13617 ( .A1(n15510), .A2(n15509), .ZN(n10941) );
  MUX2_X1 U13618 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11563), .S(n15507), .Z(
        n10940) );
  NAND2_X1 U13619 ( .A1(n10941), .A2(n10940), .ZN(n15512) );
  NAND2_X1 U13620 ( .A1(n15507), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n14881) );
  NAND2_X1 U13621 ( .A1(n15512), .A2(n14881), .ZN(n10943) );
  INV_X1 U13622 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11808) );
  MUX2_X1 U13623 ( .A(n11808), .B(P1_REG2_REG_5__SCAN_IN), .S(n14879), .Z(
        n10942) );
  NAND2_X1 U13624 ( .A1(n10943), .A2(n10942), .ZN(n14892) );
  NAND2_X1 U13625 ( .A1(n14874), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n14891) );
  NAND2_X1 U13626 ( .A1(n14892), .A2(n14891), .ZN(n10945) );
  INV_X1 U13627 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n14889) );
  MUX2_X1 U13628 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n14889), .S(n14894), .Z(
        n10944) );
  NAND2_X1 U13629 ( .A1(n10945), .A2(n10944), .ZN(n14902) );
  NAND2_X1 U13630 ( .A1(n14894), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n14901) );
  NAND2_X1 U13631 ( .A1(n14902), .A2(n14901), .ZN(n10947) );
  INV_X1 U13632 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n12034) );
  MUX2_X1 U13633 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n12034), .S(n14911), .Z(
        n10946) );
  NAND2_X1 U13634 ( .A1(n10947), .A2(n10946), .ZN(n14904) );
  NAND2_X1 U13635 ( .A1(n14911), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10951) );
  NAND2_X1 U13636 ( .A1(n14904), .A2(n10951), .ZN(n10949) );
  INV_X1 U13637 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n12302) );
  MUX2_X1 U13638 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n12302), .S(n10963), .Z(
        n10948) );
  NAND2_X1 U13639 ( .A1(n10949), .A2(n10948), .ZN(n10968) );
  MUX2_X1 U13640 ( .A(n12302), .B(P1_REG2_REG_8__SCAN_IN), .S(n10963), .Z(
        n10950) );
  NAND3_X1 U13641 ( .A1(n14904), .A2(n10951), .A3(n10950), .ZN(n10952) );
  NAND3_X1 U13642 ( .A1(n15513), .A2(n10968), .A3(n10952), .ZN(n10953) );
  OAI211_X1 U13643 ( .C1(n10955), .C2(n14942), .A(n10954), .B(n10953), .ZN(
        P1_U3251) );
  INV_X1 U13644 ( .A(n10956), .ZN(n10957) );
  XNOR2_X1 U13645 ( .A(n11005), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n10959) );
  AOI21_X1 U13646 ( .B1(n10960), .B2(n10959), .A(n14919), .ZN(n10972) );
  INV_X1 U13647 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14468) );
  NAND2_X1 U13648 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n10961) );
  OAI21_X1 U13649 ( .B1(n15497), .B2(n14468), .A(n10961), .ZN(n10962) );
  AOI21_X1 U13650 ( .B1(n11005), .B2(n15500), .A(n10962), .ZN(n10971) );
  NAND2_X1 U13651 ( .A1(n10963), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10967) );
  NAND2_X1 U13652 ( .A1(n10968), .A2(n10967), .ZN(n10965) );
  INV_X1 U13653 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n12311) );
  MUX2_X1 U13654 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n12311), .S(n11005), .Z(
        n10964) );
  NAND2_X1 U13655 ( .A1(n10965), .A2(n10964), .ZN(n14927) );
  MUX2_X1 U13656 ( .A(n12311), .B(P1_REG2_REG_9__SCAN_IN), .S(n11005), .Z(
        n10966) );
  NAND3_X1 U13657 ( .A1(n10968), .A2(n10967), .A3(n10966), .ZN(n10969) );
  NAND3_X1 U13658 ( .A1(n15513), .A2(n14927), .A3(n10969), .ZN(n10970) );
  OAI211_X1 U13659 ( .C1(n10972), .C2(n14942), .A(n10971), .B(n10970), .ZN(
        P1_U3252) );
  OAI222_X1 U13660 ( .A1(P3_U3151), .A2(n13449), .B1(n13808), .B2(n10974), 
        .C1(n10973), .C2(n13805), .ZN(P3_U3280) );
  OAI222_X1 U13661 ( .A1(n10977), .A2(P3_U3151), .B1(n13808), .B2(n10976), 
        .C1(n10975), .C2(n13805), .ZN(P3_U3281) );
  INV_X1 U13662 ( .A(n14940), .ZN(n12127) );
  INV_X1 U13663 ( .A(n10978), .ZN(n10981) );
  OAI222_X1 U13664 ( .A1(n12127), .A2(P1_U3086), .B1(n15433), .B2(n10981), 
        .C1(n10979), .C2(n15435), .ZN(P1_U3340) );
  INV_X1 U13665 ( .A(n12640), .ZN(n12469) );
  OAI222_X1 U13666 ( .A1(n12469), .A2(P2_U3088), .B1(n14637), .B2(n10981), 
        .C1(n10980), .C2(n14646), .ZN(P2_U3312) );
  INV_X1 U13667 ( .A(n10982), .ZN(n10998) );
  INV_X1 U13668 ( .A(n15580), .ZN(n12455) );
  OAI222_X1 U13669 ( .A1(n14637), .A2(n10998), .B1(n14646), .B2(n10983), .C1(
        n12455), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U13670 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14886) );
  AND2_X1 U13671 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14886), .ZN(n10984) );
  INV_X1 U13672 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n10986) );
  NAND2_X1 U13673 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n10986), .ZN(n10987) );
  INV_X1 U13674 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n10989) );
  XNOR2_X1 U13675 ( .A(n11308), .B(n10989), .ZN(n11307) );
  INV_X1 U13676 ( .A(n11307), .ZN(n10990) );
  XNOR2_X1 U13677 ( .A(n10990), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n10996) );
  INV_X1 U13678 ( .A(n10991), .ZN(n10992) );
  NAND2_X1 U13679 ( .A1(n10992), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10993) );
  INV_X1 U13680 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n11226) );
  OAI21_X1 U13681 ( .B1(n10996), .B2(n10995), .A(n11305), .ZN(n10997) );
  INV_X1 U13682 ( .A(n10997), .ZN(SUB_1596_U56) );
  INV_X1 U13683 ( .A(n11609), .ZN(n11267) );
  OAI222_X1 U13684 ( .A1(P1_U3086), .A2(n11267), .B1(n15435), .B2(n10999), 
        .C1(n15433), .C2(n10998), .ZN(P1_U3343) );
  NAND2_X1 U13685 ( .A1(n11003), .A2(n14437), .ZN(n11262) );
  OAI21_X1 U13686 ( .B1(n11003), .B2(n14437), .A(n11262), .ZN(n11002) );
  NOR2_X1 U13687 ( .A1(n11005), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n14918) );
  XNOR2_X1 U13688 ( .A(n14924), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n14917) );
  AND2_X1 U13689 ( .A1(n14924), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11000) );
  OR2_X1 U13690 ( .A1(n14916), .A2(n11000), .ZN(n11001) );
  AOI21_X1 U13691 ( .B1(n11002), .B2(n11001), .A(n11264), .ZN(n11015) );
  AND2_X1 U13692 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n12592) );
  INV_X1 U13693 ( .A(n15500), .ZN(n14975) );
  NOR2_X1 U13694 ( .A1(n14975), .A2(n11003), .ZN(n11004) );
  AOI211_X1 U13695 ( .C1(n15492), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n12592), 
        .B(n11004), .ZN(n11014) );
  NAND2_X1 U13696 ( .A1(n11005), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n14926) );
  NAND2_X1 U13697 ( .A1(n14927), .A2(n14926), .ZN(n11007) );
  INV_X1 U13698 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n12330) );
  MUX2_X1 U13699 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n12330), .S(n14924), .Z(
        n11006) );
  NAND2_X1 U13700 ( .A1(n11007), .A2(n11006), .ZN(n14929) );
  NAND2_X1 U13701 ( .A1(n14924), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11011) );
  NAND2_X1 U13702 ( .A1(n14929), .A2(n11011), .ZN(n11009) );
  INV_X1 U13703 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n12424) );
  MUX2_X1 U13704 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n12424), .S(n11269), .Z(
        n11008) );
  NAND2_X1 U13705 ( .A1(n11009), .A2(n11008), .ZN(n11271) );
  MUX2_X1 U13706 ( .A(n12424), .B(P1_REG2_REG_11__SCAN_IN), .S(n11269), .Z(
        n11010) );
  NAND3_X1 U13707 ( .A1(n14929), .A2(n11011), .A3(n11010), .ZN(n11012) );
  NAND3_X1 U13708 ( .A1(n11271), .A2(n15513), .A3(n11012), .ZN(n11013) );
  OAI211_X1 U13709 ( .C1(n11015), .C2(n14942), .A(n11014), .B(n11013), .ZN(
        P1_U3254) );
  INV_X1 U13710 ( .A(n11016), .ZN(n11018) );
  INV_X1 U13711 ( .A(n11017), .ZN(n13470) );
  OAI222_X1 U13712 ( .A1(n13805), .A2(n11019), .B1(n13808), .B2(n11018), .C1(
        P3_U3151), .C2(n13470), .ZN(P3_U3279) );
  INV_X1 U13713 ( .A(n12466), .ZN(n15607) );
  INV_X1 U13714 ( .A(n11020), .ZN(n11023) );
  OAI222_X1 U13715 ( .A1(n15607), .A2(P2_U3088), .B1(n14644), .B2(n11023), 
        .C1(n11021), .C2(n14646), .ZN(P2_U3313) );
  INV_X1 U13716 ( .A(n12124), .ZN(n12122) );
  OAI222_X1 U13717 ( .A1(n12122), .A2(P1_U3086), .B1(n15433), .B2(n11023), 
        .C1(n11022), .C2(n15435), .ZN(P1_U3341) );
  INV_X1 U13718 ( .A(n11024), .ZN(n11102) );
  OAI222_X1 U13719 ( .A1(n14637), .A2(n11102), .B1(n14646), .B2(n11025), .C1(
        n12457), .C2(P2_U3088), .ZN(P2_U3314) );
  OAI21_X1 U13720 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n11027), .A(n11026), .ZN(
        n11028) );
  NAND2_X1 U13721 ( .A1(n13495), .A2(n11028), .ZN(n11034) );
  OAI21_X1 U13722 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n11030), .A(n11029), .ZN(
        n11031) );
  NAND2_X1 U13723 ( .A1(n13504), .A2(n11031), .ZN(n11033) );
  AND2_X1 U13724 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11784) );
  AOI21_X1 U13725 ( .B1(n15671), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11784), .ZN(
        n11032) );
  AND3_X1 U13726 ( .A1(n11034), .A2(n11033), .A3(n11032), .ZN(n11040) );
  AND3_X1 U13727 ( .A1(n11214), .A2(n11036), .A3(n11035), .ZN(n11037) );
  OAI21_X1 U13728 ( .B1(n6994), .B2(n11037), .A(n13509), .ZN(n11039) );
  OAI211_X1 U13729 ( .C1(n13486), .C2(n11041), .A(n11040), .B(n11039), .ZN(
        P3_U3187) );
  OAI21_X1 U13730 ( .B1(n11044), .B2(n11043), .A(n11042), .ZN(n11045) );
  INV_X1 U13731 ( .A(n11045), .ZN(n11047) );
  AND2_X1 U13732 ( .A1(n8885), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11048) );
  INV_X1 U13733 ( .A(n15587), .ZN(n15608) );
  INV_X1 U13734 ( .A(n13983), .ZN(n13982) );
  MUX2_X1 U13735 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n8964), .S(n13983), .Z(
        n13990) );
  INV_X1 U13736 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n13991) );
  MUX2_X1 U13737 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n8971), .S(n11071), .Z(
        n11050) );
  NOR2_X1 U13738 ( .A1(n8885), .A2(P2_U3088), .ZN(n14639) );
  AND2_X1 U13739 ( .A1(n11064), .A2(n14639), .ZN(n11058) );
  INV_X1 U13740 ( .A(n15610), .ZN(n15597) );
  AOI211_X1 U13741 ( .C1(n11051), .C2(n11050), .A(n11072), .B(n15597), .ZN(
        n11063) );
  MUX2_X1 U13742 ( .A(n13984), .B(P2_REG2_REG_1__SCAN_IN), .S(n13983), .Z(
        n11053) );
  AND2_X1 U13743 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n11052) );
  NAND2_X1 U13744 ( .A1(n11053), .A2(n11052), .ZN(n13988) );
  NAND2_X1 U13745 ( .A1(n13982), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n11054) );
  NAND2_X1 U13746 ( .A1(n13988), .A2(n11054), .ZN(n11056) );
  INV_X1 U13747 ( .A(n11056), .ZN(n11061) );
  INV_X1 U13748 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11976) );
  MUX2_X1 U13749 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n11976), .S(n11071), .Z(
        n11060) );
  MUX2_X1 U13750 ( .A(n11976), .B(P2_REG2_REG_2__SCAN_IN), .S(n11071), .Z(
        n11055) );
  NAND2_X1 U13751 ( .A1(n11056), .A2(n11055), .ZN(n11082) );
  INV_X1 U13752 ( .A(n11082), .ZN(n11059) );
  INV_X1 U13753 ( .A(n14647), .ZN(n11057) );
  NAND2_X1 U13754 ( .A1(n11058), .A2(n11057), .ZN(n15591) );
  AOI211_X1 U13755 ( .C1(n11061), .C2(n11060), .A(n11059), .B(n15591), .ZN(
        n11062) );
  NOR2_X1 U13756 ( .A1(n11063), .A2(n11062), .ZN(n11067) );
  NOR2_X2 U13757 ( .A1(n11064), .A2(P2_U3088), .ZN(n15585) );
  NOR2_X1 U13758 ( .A1(n11975), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11065) );
  AOI21_X1 U13759 ( .B1(n15585), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n11065), .ZN(
        n11066) );
  OAI211_X1 U13760 ( .C1(n11071), .C2(n15608), .A(n11067), .B(n11066), .ZN(
        P2_U3216) );
  INV_X1 U13761 ( .A(n11068), .ZN(n11123) );
  INV_X1 U13762 ( .A(n12645), .ZN(n14043) );
  OAI222_X1 U13763 ( .A1(n14637), .A2(n11123), .B1(n14646), .B2(n11069), .C1(
        n14043), .C2(P2_U3088), .ZN(P2_U3311) );
  XNOR2_X1 U13764 ( .A(n11422), .B(n11070), .ZN(n11078) );
  INV_X1 U13765 ( .A(n11071), .ZN(n11080) );
  INV_X1 U13766 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n11714) );
  MUX2_X1 U13767 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n11714), .S(n15560), .Z(
        n15566) );
  NOR2_X1 U13768 ( .A1(n15560), .A2(n11714), .ZN(n14006) );
  INV_X1 U13769 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n11073) );
  MUX2_X1 U13770 ( .A(n11073), .B(P2_REG1_REG_4__SCAN_IN), .S(n14005), .Z(
        n11074) );
  NAND2_X1 U13771 ( .A1(n14000), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n11133) );
  INV_X1 U13772 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n11919) );
  MUX2_X1 U13773 ( .A(n11919), .B(P2_REG1_REG_5__SCAN_IN), .S(n11087), .Z(
        n11132) );
  NOR2_X1 U13774 ( .A1(n11142), .A2(n11919), .ZN(n14014) );
  MUX2_X1 U13775 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n11075), .S(n14023), .Z(
        n11076) );
  NAND2_X1 U13776 ( .A1(n14023), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n11224) );
  INV_X1 U13777 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n12254) );
  MUX2_X1 U13778 ( .A(n12254), .B(P2_REG1_REG_7__SCAN_IN), .S(n11228), .Z(
        n11223) );
  INV_X1 U13779 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n12441) );
  XNOR2_X1 U13780 ( .A(n11243), .B(n12441), .ZN(n11237) );
  OAI22_X1 U13781 ( .A1(n11238), .A2(n11237), .B1(n11243), .B2(n12441), .ZN(
        n11077) );
  AOI21_X1 U13782 ( .B1(n11078), .B2(n11077), .A(n11418), .ZN(n11100) );
  NAND2_X1 U13783 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n12140) );
  OAI21_X1 U13784 ( .B1(n15608), .B2(n11422), .A(n12140), .ZN(n11079) );
  AOI21_X1 U13785 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(n15585), .A(n11079), .ZN(
        n11099) );
  NAND2_X1 U13786 ( .A1(n11080), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n11081) );
  NAND2_X1 U13787 ( .A1(n11082), .A2(n11081), .ZN(n15563) );
  MUX2_X1 U13788 ( .A(n12262), .B(P2_REG2_REG_3__SCAN_IN), .S(n15560), .Z(
        n15564) );
  NAND2_X1 U13789 ( .A1(n15563), .A2(n15564), .ZN(n15562) );
  OR2_X1 U13790 ( .A1(n15560), .A2(n12262), .ZN(n14001) );
  NAND2_X1 U13791 ( .A1(n15562), .A2(n14001), .ZN(n11085) );
  MUX2_X1 U13792 ( .A(n11083), .B(P2_REG2_REG_4__SCAN_IN), .S(n14005), .Z(
        n11084) );
  NAND2_X1 U13793 ( .A1(n11085), .A2(n11084), .ZN(n14004) );
  NAND2_X1 U13794 ( .A1(n14000), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n11086) );
  NAND2_X1 U13795 ( .A1(n14004), .A2(n11086), .ZN(n11136) );
  MUX2_X1 U13796 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11957), .S(n11087), .Z(
        n11137) );
  NAND2_X1 U13797 ( .A1(n11136), .A2(n11137), .ZN(n14026) );
  NAND2_X1 U13798 ( .A1(n11087), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n14025) );
  NAND2_X1 U13799 ( .A1(n14026), .A2(n14025), .ZN(n11089) );
  INV_X1 U13800 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n12061) );
  MUX2_X1 U13801 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n12061), .S(n14023), .Z(
        n11088) );
  NAND2_X1 U13802 ( .A1(n11089), .A2(n11088), .ZN(n14028) );
  NAND2_X1 U13803 ( .A1(n14023), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n11230) );
  NAND2_X1 U13804 ( .A1(n14028), .A2(n11230), .ZN(n11091) );
  MUX2_X1 U13805 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n15621), .S(n11228), .Z(
        n11090) );
  NAND2_X1 U13806 ( .A1(n11091), .A2(n11090), .ZN(n11232) );
  NAND2_X1 U13807 ( .A1(n11228), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n11092) );
  NAND2_X1 U13808 ( .A1(n11232), .A2(n11092), .ZN(n11240) );
  MUX2_X1 U13809 ( .A(n12382), .B(P2_REG2_REG_8__SCAN_IN), .S(n11243), .Z(
        n11241) );
  NAND2_X1 U13810 ( .A1(n11240), .A2(n11241), .ZN(n11239) );
  NAND2_X1 U13811 ( .A1(n11093), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n11094) );
  INV_X1 U13812 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11421) );
  MUX2_X1 U13813 ( .A(n11421), .B(P2_REG2_REG_9__SCAN_IN), .S(n11422), .Z(
        n11095) );
  NAND2_X1 U13814 ( .A1(n11096), .A2(n11095), .ZN(n11424) );
  OAI21_X1 U13815 ( .B1(n11096), .B2(n11095), .A(n11424), .ZN(n11097) );
  NAND2_X1 U13816 ( .A1(n11097), .A2(n15613), .ZN(n11098) );
  OAI211_X1 U13817 ( .C1(n11100), .C2(n15597), .A(n11099), .B(n11098), .ZN(
        P2_U3223) );
  OAI222_X1 U13818 ( .A1(n13485), .A2(P3_U3151), .B1(n13808), .B2(n11101), 
        .C1(n14461), .C2(n13805), .ZN(P3_U3278) );
  INV_X1 U13819 ( .A(n11663), .ZN(n11619) );
  OAI222_X1 U13820 ( .A1(P1_U3086), .A2(n11619), .B1(n15435), .B2(n11103), 
        .C1(n15433), .C2(n11102), .ZN(P1_U3342) );
  OAI21_X1 U13821 ( .B1(n11106), .B2(n11105), .A(n11104), .ZN(n11120) );
  INV_X1 U13822 ( .A(n11107), .ZN(n11109) );
  NAND3_X1 U13823 ( .A1(n11109), .A2(n11108), .A3(n11396), .ZN(n11110) );
  NAND2_X1 U13824 ( .A1(n11332), .A2(n11110), .ZN(n11111) );
  AOI22_X1 U13825 ( .A1(n13509), .A2(n11111), .B1(P3_REG3_REG_2__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11118) );
  OAI21_X1 U13826 ( .B1(n11114), .B2(n11113), .A(n11112), .ZN(n11115) );
  NAND2_X1 U13827 ( .A1(n13504), .A2(n11115), .ZN(n11117) );
  NAND2_X1 U13828 ( .A1(n15671), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n11116) );
  NAND3_X1 U13829 ( .A1(n11118), .A2(n11117), .A3(n11116), .ZN(n11119) );
  AOI21_X1 U13830 ( .B1(n13495), .B2(n11120), .A(n11119), .ZN(n11121) );
  OAI21_X1 U13831 ( .B1(n11122), .B2(n13486), .A(n11121), .ZN(P3_U3184) );
  OAI222_X1 U13832 ( .A1(P1_U3086), .A2(n14951), .B1(n15435), .B2(n11124), 
        .C1(n15433), .C2(n11123), .ZN(P1_U3339) );
  INV_X1 U13833 ( .A(n15260), .ZN(n15160) );
  AOI21_X1 U13834 ( .B1(n15160), .B2(n15354), .A(n11125), .ZN(n11126) );
  AOI21_X1 U13835 ( .B1(n15258), .B2(n10096), .A(n11126), .ZN(n11892) );
  NAND3_X1 U13836 ( .A1(n11128), .A2(n11825), .A3(n11127), .ZN(n11895) );
  NAND2_X1 U13837 ( .A1(n11892), .A2(n11895), .ZN(n11130) );
  NAND2_X1 U13838 ( .A1(n11130), .A2(n15554), .ZN(n11129) );
  OAI21_X1 U13839 ( .B1(n15554), .B2(n10087), .A(n11129), .ZN(P1_U3528) );
  NAND2_X1 U13840 ( .A1(n11130), .A2(n15550), .ZN(n11131) );
  OAI21_X1 U13841 ( .B1(n15550), .B2(n9588), .A(n11131), .ZN(P1_U3459) );
  INV_X1 U13842 ( .A(n14019), .ZN(n11135) );
  NAND3_X1 U13843 ( .A1(n14009), .A2(n11133), .A3(n11132), .ZN(n11134) );
  NAND3_X1 U13844 ( .A1(n11135), .A2(n15610), .A3(n11134), .ZN(n11141) );
  NAND2_X1 U13845 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n11570) );
  OAI211_X1 U13846 ( .C1(n11137), .C2(n11136), .A(n15613), .B(n14026), .ZN(
        n11138) );
  NAND2_X1 U13847 ( .A1(n11570), .A2(n11138), .ZN(n11139) );
  AOI21_X1 U13848 ( .B1(n15585), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n11139), .ZN(
        n11140) );
  OAI211_X1 U13849 ( .C1(n15608), .C2(n11142), .A(n11141), .B(n11140), .ZN(
        P2_U3219) );
  INV_X1 U13850 ( .A(n14795), .ZN(n14763) );
  NAND2_X1 U13851 ( .A1(n14771), .A2(n11143), .ZN(n12973) );
  INV_X1 U13852 ( .A(n11144), .ZN(n11145) );
  AOI21_X1 U13853 ( .B1(n11147), .B2(n11146), .A(n11145), .ZN(n14837) );
  OR2_X1 U13854 ( .A1(n14778), .A2(n15241), .ZN(n14790) );
  OAI22_X1 U13855 ( .A1(n14837), .A2(n14797), .B1(n9991), .B2(n14790), .ZN(
        n11148) );
  AOI21_X1 U13856 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n12973), .A(n11148), .ZN(
        n11149) );
  OAI21_X1 U13857 ( .B1(n11151), .B2(n14763), .A(n11149), .ZN(P1_U3232) );
  XNOR2_X1 U13858 ( .A(n11153), .B(n11150), .ZN(n11505) );
  INV_X1 U13859 ( .A(n11505), .ZN(n11163) );
  OR2_X1 U13860 ( .A1(n11498), .A2(n11151), .ZN(n11152) );
  NAND2_X1 U13861 ( .A1(n11253), .A2(n11152), .ZN(n11155) );
  NOR2_X1 U13862 ( .A1(n11155), .A2(n15270), .ZN(n11500) );
  INV_X1 U13863 ( .A(n15257), .ZN(n15239) );
  OAI21_X1 U13864 ( .B1(n11153), .B2(n15160), .A(n15239), .ZN(n11161) );
  XNOR2_X1 U13865 ( .A(n11155), .B(n10096), .ZN(n11157) );
  NAND3_X1 U13866 ( .A1(n11157), .A2(n11156), .A3(n15260), .ZN(n11158) );
  OAI21_X1 U13867 ( .B1(n11159), .B2(n15241), .A(n11158), .ZN(n11160) );
  AOI21_X1 U13868 ( .B1(n11161), .B2(n11154), .A(n11160), .ZN(n11502) );
  INV_X1 U13869 ( .A(n11502), .ZN(n11162) );
  AOI211_X1 U13870 ( .C1(n15370), .C2(n11163), .A(n11500), .B(n11162), .ZN(
        n11168) );
  OAI22_X1 U13871 ( .A1(n10072), .A2(n11498), .B1(n15550), .B2(n9609), .ZN(
        n11164) );
  INV_X1 U13872 ( .A(n11164), .ZN(n11165) );
  OAI21_X1 U13873 ( .B1(n11168), .B2(n15549), .A(n11165), .ZN(P1_U3462) );
  AOI22_X1 U13874 ( .A1(n12686), .A2(n11166), .B1(n15552), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n11167) );
  OAI21_X1 U13875 ( .B1(n11168), .B2(n15552), .A(n11167), .ZN(P1_U3529) );
  INV_X1 U13876 ( .A(n11182), .ZN(n11175) );
  AND3_X1 U13877 ( .A1(n11171), .A2(n11170), .A3(n11169), .ZN(n11174) );
  OR2_X1 U13878 ( .A1(n11185), .A2(n11172), .ZN(n11173) );
  OAI211_X1 U13879 ( .C1(n11189), .C2(n11175), .A(n11174), .B(n11173), .ZN(
        n11176) );
  NAND2_X1 U13880 ( .A1(n11176), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11179) );
  INV_X1 U13881 ( .A(n13189), .ZN(n11177) );
  OR2_X1 U13882 ( .A1(n11177), .A2(n11185), .ZN(n11178) );
  NOR2_X1 U13883 ( .A1(n13362), .A2(P3_U3151), .ZN(n11383) );
  NAND2_X1 U13884 ( .A1(n11185), .A2(n13189), .ZN(n11282) );
  INV_X1 U13885 ( .A(n11282), .ZN(n11180) );
  NAND4_X1 U13886 ( .A1(n11189), .A2(n11183), .A3(n11182), .A4(n15715), .ZN(
        n11187) );
  NAND2_X1 U13887 ( .A1(n11185), .A2(n11184), .ZN(n11186) );
  NAND2_X1 U13888 ( .A1(n6432), .A2(n11390), .ZN(n13055) );
  INV_X1 U13889 ( .A(n13055), .ZN(n11188) );
  NOR2_X1 U13890 ( .A1(n13716), .A2(n11188), .ZN(n13008) );
  OR2_X1 U13891 ( .A1(n11189), .A2(n15674), .ZN(n11192) );
  INV_X1 U13892 ( .A(n11190), .ZN(n11191) );
  NAND2_X1 U13893 ( .A1(n11192), .A2(n11191), .ZN(n13367) );
  OAI22_X1 U13894 ( .A1(n13351), .A2(n13008), .B1(n13367), .B2(n11390), .ZN(
        n11193) );
  AOI21_X1 U13895 ( .B1(n13357), .B2(n11181), .A(n11193), .ZN(n11194) );
  OAI21_X1 U13896 ( .B1(n11383), .B2(n11366), .A(n11194), .ZN(P3_U3172) );
  INV_X1 U13897 ( .A(n11195), .ZN(n11248) );
  OAI222_X1 U13898 ( .A1(n14637), .A2(n11248), .B1(n14646), .B2(n11196), .C1(
        n12648), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U13899 ( .A(n11197), .ZN(n11199) );
  NAND3_X1 U13900 ( .A1(n11328), .A2(n11199), .A3(n11198), .ZN(n11200) );
  NAND2_X1 U13901 ( .A1(n11201), .A2(n11200), .ZN(n11217) );
  INV_X1 U13902 ( .A(n11202), .ZN(n11204) );
  NAND3_X1 U13903 ( .A1(n11335), .A2(n11204), .A3(n11203), .ZN(n11205) );
  NAND2_X1 U13904 ( .A1(n11206), .A2(n11205), .ZN(n11207) );
  NAND2_X1 U13905 ( .A1(n13504), .A2(n11207), .ZN(n11210) );
  NAND2_X1 U13906 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n11589) );
  INV_X1 U13907 ( .A(n11589), .ZN(n11208) );
  AOI21_X1 U13908 ( .B1(n15671), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n11208), .ZN(
        n11209) );
  NAND2_X1 U13909 ( .A1(n11210), .A2(n11209), .ZN(n11216) );
  OR3_X1 U13910 ( .A1(n11329), .A2(n11212), .A3(n11211), .ZN(n11213) );
  AOI21_X1 U13911 ( .B1(n11214), .B2(n11213), .A(n13407), .ZN(n11215) );
  AOI211_X1 U13912 ( .C1(n13495), .C2(n11217), .A(n11216), .B(n11215), .ZN(
        n11218) );
  OAI21_X1 U13913 ( .B1(n11219), .B2(n13486), .A(n11218), .ZN(P3_U3186) );
  OAI222_X1 U13914 ( .A1(P3_U3151), .A2(n11222), .B1(n13808), .B2(n11221), 
        .C1(n11220), .C2(n13805), .ZN(P3_U3277) );
  NAND3_X1 U13915 ( .A1(n14017), .A2(n11224), .A3(n11223), .ZN(n11225) );
  NAND2_X1 U13916 ( .A1(n11225), .A2(n15610), .ZN(n11235) );
  INV_X1 U13917 ( .A(n15585), .ZN(n15618) );
  NAND2_X1 U13918 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n11752) );
  OAI21_X1 U13919 ( .B1(n15618), .B2(n11226), .A(n11752), .ZN(n11227) );
  AOI21_X1 U13920 ( .B1(n11228), .B2(n15587), .A(n11227), .ZN(n11234) );
  MUX2_X1 U13921 ( .A(n15621), .B(P2_REG2_REG_7__SCAN_IN), .S(n11228), .Z(
        n11229) );
  NAND3_X1 U13922 ( .A1(n14028), .A2(n11230), .A3(n11229), .ZN(n11231) );
  NAND3_X1 U13923 ( .A1(n15613), .A2(n11232), .A3(n11231), .ZN(n11233) );
  OAI211_X1 U13924 ( .C1(n11236), .C2(n11235), .A(n11234), .B(n11233), .ZN(
        P2_U3221) );
  XNOR2_X1 U13925 ( .A(n11238), .B(n11237), .ZN(n11247) );
  NAND2_X1 U13926 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n12008) );
  OAI211_X1 U13927 ( .C1(n11241), .C2(n11240), .A(n15613), .B(n11239), .ZN(
        n11242) );
  NAND2_X1 U13928 ( .A1(n12008), .A2(n11242), .ZN(n11245) );
  NOR2_X1 U13929 ( .A1(n15608), .A2(n11243), .ZN(n11244) );
  AOI211_X1 U13930 ( .C1(n15585), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n11245), .B(
        n11244), .ZN(n11246) );
  OAI21_X1 U13931 ( .B1(n11247), .B2(n15597), .A(n11246), .ZN(P2_U3222) );
  INV_X1 U13932 ( .A(n14965), .ZN(n14968) );
  OAI222_X1 U13933 ( .A1(P1_U3086), .A2(n14968), .B1(n15435), .B2(n11249), 
        .C1(n15433), .C2(n11248), .ZN(P1_U3338) );
  INV_X1 U13934 ( .A(n11317), .ZN(n11252) );
  AOI211_X1 U13935 ( .C1(n11259), .C2(n11253), .A(n15270), .B(n11252), .ZN(
        n11674) );
  XNOR2_X1 U13936 ( .A(n11255), .B(n11254), .ZN(n11256) );
  OAI22_X1 U13937 ( .A1(n9991), .A2(n15239), .B1(n9995), .B2(n15241), .ZN(
        n12972) );
  AOI21_X1 U13938 ( .B1(n11256), .B2(n15260), .A(n12972), .ZN(n11682) );
  INV_X1 U13939 ( .A(n11682), .ZN(n11257) );
  AOI211_X1 U13940 ( .C1(n15370), .C2(n11680), .A(n11674), .B(n11257), .ZN(
        n11261) );
  AOI22_X1 U13941 ( .A1(n12478), .A2(n11259), .B1(n15549), .B2(
        P1_REG0_REG_2__SCAN_IN), .ZN(n11258) );
  OAI21_X1 U13942 ( .B1(n11261), .B2(n15549), .A(n11258), .ZN(P1_U3465) );
  AOI22_X1 U13943 ( .A1(n12686), .A2(n11259), .B1(n15552), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n11260) );
  OAI21_X1 U13944 ( .B1(n11261), .B2(n15552), .A(n11260), .ZN(P1_U3530) );
  INV_X1 U13945 ( .A(n11262), .ZN(n11263) );
  XNOR2_X1 U13946 ( .A(n11609), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n11265) );
  AOI21_X1 U13947 ( .B1(n11266), .B2(n11265), .A(n11606), .ZN(n11280) );
  AND2_X1 U13948 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n12631) );
  NOR2_X1 U13949 ( .A1(n14975), .A2(n11267), .ZN(n11268) );
  AOI211_X1 U13950 ( .C1(n15492), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n12631), 
        .B(n11268), .ZN(n11279) );
  NAND2_X1 U13951 ( .A1(n11269), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11270) );
  NAND2_X1 U13952 ( .A1(n11271), .A2(n11270), .ZN(n11274) );
  INV_X1 U13953 ( .A(n11274), .ZN(n11276) );
  INV_X1 U13954 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11272) );
  MUX2_X1 U13955 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n11272), .S(n11609), .Z(
        n11275) );
  MUX2_X1 U13956 ( .A(n11272), .B(P1_REG2_REG_12__SCAN_IN), .S(n11609), .Z(
        n11273) );
  OAI21_X1 U13957 ( .B1(n11276), .B2(n11275), .A(n11611), .ZN(n11277) );
  NAND2_X1 U13958 ( .A1(n11277), .A2(n15513), .ZN(n11278) );
  OAI211_X1 U13959 ( .C1(n11280), .C2(n14942), .A(n11279), .B(n11278), .ZN(
        P1_U3255) );
  INV_X1 U13960 ( .A(n13359), .ZN(n13328) );
  INV_X1 U13961 ( .A(n13385), .ZN(n11549) );
  OAI22_X1 U13962 ( .A1(n13331), .A2(n11549), .B1(n11448), .B2(n13367), .ZN(
        n11283) );
  AOI21_X1 U13963 ( .B1(n13328), .B2(n11181), .A(n11283), .ZN(n11294) );
  NAND2_X1 U13964 ( .A1(n13059), .A2(n11284), .ZN(n11285) );
  NAND2_X1 U13965 ( .A1(n11285), .A2(n11804), .ZN(n11286) );
  NAND2_X4 U13966 ( .A1(n11287), .A2(n11286), .ZN(n12935) );
  XNOR2_X1 U13967 ( .A(n12935), .B(n11448), .ZN(n11546) );
  XNOR2_X1 U13968 ( .A(n11546), .B(n6974), .ZN(n11291) );
  NAND2_X1 U13969 ( .A1(n11181), .A2(n6959), .ZN(n11289) );
  OAI21_X1 U13970 ( .B1(n11291), .B2(n11290), .A(n11553), .ZN(n11292) );
  NAND2_X1 U13971 ( .A1(n11292), .A2(n13353), .ZN(n11293) );
  OAI211_X1 U13972 ( .C1(n11383), .C2(n11295), .A(n11294), .B(n11293), .ZN(
        P3_U3177) );
  OAI21_X1 U13973 ( .B1(n7794), .B2(n11297), .A(n11296), .ZN(n11301) );
  INV_X1 U13974 ( .A(n14790), .ZN(n14748) );
  AND2_X1 U13975 ( .A1(n14766), .A2(n15257), .ZN(n14727) );
  AOI22_X1 U13976 ( .A1(n14748), .A2(n14820), .B1(n14727), .B2(n11154), .ZN(
        n11299) );
  NAND2_X1 U13977 ( .A1(n12973), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n11298) );
  OAI211_X1 U13978 ( .C1(n14763), .C2(n11498), .A(n11299), .B(n11298), .ZN(
        n11300) );
  AOI21_X1 U13979 ( .B1(n14754), .B2(n11301), .A(n11300), .ZN(n11302) );
  INV_X1 U13980 ( .A(n11302), .ZN(P1_U3222) );
  NAND2_X1 U13981 ( .A1(n11303), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n11304) );
  INV_X1 U13982 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n11306) );
  NAND2_X1 U13983 ( .A1(n11307), .A2(n11306), .ZN(n11310) );
  NAND2_X1 U13984 ( .A1(n11308), .A2(P3_ADDR_REG_7__SCAN_IN), .ZN(n11309) );
  NAND2_X1 U13985 ( .A1(n11310), .A2(n11309), .ZN(n11652) );
  XNOR2_X1 U13986 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(P3_ADDR_REG_8__SCAN_IN), 
        .ZN(n11651) );
  INV_X1 U13987 ( .A(n11651), .ZN(n11311) );
  XNOR2_X1 U13988 ( .A(n11652), .B(n11311), .ZN(n11646) );
  OAI21_X1 U13989 ( .B1(n11312), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n11650), .ZN(
        n11313) );
  INV_X1 U13990 ( .A(n11313), .ZN(SUB_1596_U55) );
  OR2_X1 U13991 ( .A1(n11315), .A2(n11314), .ZN(n11316) );
  NAND2_X1 U13992 ( .A1(n11317), .A2(n15523), .ZN(n11318) );
  INV_X1 U13993 ( .A(n15270), .ZN(n15168) );
  NAND2_X1 U13994 ( .A1(n11318), .A2(n15168), .ZN(n11319) );
  NOR2_X1 U13995 ( .A1(n11508), .A2(n11319), .ZN(n15521) );
  XNOR2_X1 U13996 ( .A(n11320), .B(n11321), .ZN(n11323) );
  AOI22_X1 U13997 ( .A1(n15257), .A2(n14820), .B1(n14818), .B2(n15258), .ZN(
        n11541) );
  INV_X1 U13998 ( .A(n11541), .ZN(n11322) );
  AOI21_X1 U13999 ( .B1(n11323), .B2(n15260), .A(n11322), .ZN(n15532) );
  INV_X1 U14000 ( .A(n15532), .ZN(n11324) );
  AOI211_X1 U14001 ( .C1(n15370), .C2(n15520), .A(n15521), .B(n11324), .ZN(
        n11327) );
  AOI22_X1 U14002 ( .A1(n12686), .A2(n15523), .B1(n15552), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n11325) );
  OAI21_X1 U14003 ( .B1(n11327), .B2(n15552), .A(n11325), .ZN(P1_U3531) );
  AOI22_X1 U14004 ( .A1(n12478), .A2(n15523), .B1(n15549), .B2(
        P1_REG0_REG_3__SCAN_IN), .ZN(n11326) );
  OAI21_X1 U14005 ( .B1(n11327), .B2(n15549), .A(n11326), .ZN(P1_U3468) );
  OAI21_X1 U14006 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(n6633), .A(n11328), .ZN(
        n11342) );
  INV_X1 U14007 ( .A(n11329), .ZN(n11334) );
  NAND3_X1 U14008 ( .A1(n11332), .A2(n11331), .A3(n11330), .ZN(n11333) );
  AOI21_X1 U14009 ( .B1(n11334), .B2(n11333), .A(n13407), .ZN(n11341) );
  INV_X1 U14010 ( .A(n11335), .ZN(n11336) );
  AOI21_X1 U14011 ( .B1(n11730), .B2(n11337), .A(n11336), .ZN(n11339) );
  AOI22_X1 U14012 ( .A1(n15671), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n11338) );
  OAI21_X1 U14013 ( .B1(n13490), .B2(n11339), .A(n11338), .ZN(n11340) );
  AOI211_X1 U14014 ( .C1(n13495), .C2(n11342), .A(n11341), .B(n11340), .ZN(
        n11343) );
  OAI21_X1 U14015 ( .B1(n11344), .B2(n13486), .A(n11343), .ZN(P3_U3185) );
  INV_X1 U14016 ( .A(n11345), .ZN(n11348) );
  INV_X1 U14017 ( .A(n11532), .ZN(n11347) );
  AOI21_X1 U14018 ( .B1(n15732), .B2(n11348), .A(n11347), .ZN(n11362) );
  OAI21_X1 U14019 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n11349), .A(n11350), .ZN(
        n11354) );
  AND2_X1 U14020 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n12359) );
  AOI21_X1 U14021 ( .B1(n15671), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n12359), .ZN(
        n11351) );
  OAI21_X1 U14022 ( .B1(n13486), .B2(n11352), .A(n11351), .ZN(n11353) );
  AOI21_X1 U14023 ( .B1(n11354), .B2(n13504), .A(n11353), .ZN(n11361) );
  AND3_X1 U14024 ( .A1(n11357), .A2(n11356), .A3(n11355), .ZN(n11358) );
  OAI21_X1 U14025 ( .B1(n11359), .B2(n11358), .A(n13509), .ZN(n11360) );
  OAI211_X1 U14026 ( .C1(n11362), .C2(n13461), .A(n11361), .B(n11360), .ZN(
        P3_U3189) );
  NOR3_X1 U14027 ( .A1(n13495), .A2(n13504), .A3(n13509), .ZN(n11373) );
  OAI21_X1 U14028 ( .B1(n13188), .B2(n13407), .A(n13490), .ZN(n11363) );
  NAND2_X1 U14029 ( .A1(n11363), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11364) );
  MUX2_X1 U14030 ( .A(n13486), .B(n11364), .S(n7802), .Z(n11372) );
  OAI21_X1 U14031 ( .B1(n11365), .B2(n13407), .A(n13461), .ZN(n11370) );
  INV_X1 U14032 ( .A(n15671), .ZN(n13499) );
  INV_X1 U14033 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n11367) );
  OAI22_X1 U14034 ( .A1(n13499), .A2(n11367), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11366), .ZN(n11368) );
  AOI21_X1 U14035 ( .B1(n11370), .B2(n11369), .A(n11368), .ZN(n11371) );
  OAI211_X1 U14036 ( .C1(n11373), .C2(n11394), .A(n11372), .B(n11371), .ZN(
        P3_U3182) );
  OAI22_X1 U14037 ( .A1(n13331), .A2(n6974), .B1(n13732), .B2(n13367), .ZN(
        n11374) );
  AOI21_X1 U14038 ( .B1(n13328), .B2(n6432), .A(n11374), .ZN(n11382) );
  INV_X1 U14039 ( .A(n13716), .ZN(n11376) );
  NAND3_X1 U14040 ( .A1(n12935), .A2(n11375), .A3(n11376), .ZN(n11377) );
  OAI211_X1 U14041 ( .C1(n11379), .C2(n13720), .A(n11378), .B(n11377), .ZN(
        n11380) );
  NAND2_X1 U14042 ( .A1(n11380), .A2(n13353), .ZN(n11381) );
  OAI211_X1 U14043 ( .C1(n11383), .C2(n11400), .A(n11382), .B(n11381), .ZN(
        P3_U3162) );
  NAND2_X1 U14044 ( .A1(n11384), .A2(n15715), .ZN(n11385) );
  OR2_X1 U14045 ( .A1(n13008), .A2(n11385), .ZN(n11387) );
  NAND2_X1 U14046 ( .A1(n13722), .A2(n11181), .ZN(n11386) );
  AND2_X1 U14047 ( .A1(n11387), .A2(n11386), .ZN(n11411) );
  MUX2_X1 U14048 ( .A(n11411), .B(n8117), .S(n15721), .Z(n11388) );
  OAI21_X1 U14049 ( .B1(n11390), .B2(n13790), .A(n11388), .ZN(P3_U3390) );
  MUX2_X1 U14050 ( .A(n7922), .B(n11411), .S(n15734), .Z(n11389) );
  OAI21_X1 U14051 ( .B1(n11390), .B2(n13709), .A(n11389), .ZN(P3_U3459) );
  NAND2_X1 U14052 ( .A1(n11391), .A2(n15689), .ZN(n11392) );
  NAND2_X1 U14053 ( .A1(n11393), .A2(n11392), .ZN(n11407) );
  NAND2_X1 U14054 ( .A1(n11396), .A2(n11395), .ZN(n11397) );
  NAND2_X1 U14055 ( .A1(n13509), .A2(n11397), .ZN(n11399) );
  NAND2_X1 U14056 ( .A1(n15671), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n11398) );
  OAI211_X1 U14057 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n11400), .A(n11399), .B(
        n11398), .ZN(n11406) );
  NAND2_X1 U14058 ( .A1(n11402), .A2(n11401), .ZN(n11403) );
  AOI21_X1 U14059 ( .B1(n11404), .B2(n11403), .A(n13461), .ZN(n11405) );
  AOI211_X1 U14060 ( .C1(n13504), .C2(n11407), .A(n11406), .B(n11405), .ZN(
        n11408) );
  OAI21_X1 U14061 ( .B1(n11409), .B2(n13486), .A(n11408), .ZN(P3_U3183) );
  MUX2_X1 U14062 ( .A(n11411), .B(n11410), .S(n15691), .Z(n11415) );
  AOI22_X1 U14063 ( .A1(n13659), .A2(n11413), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(n11412), .ZN(n11414) );
  NAND2_X1 U14064 ( .A1(n11415), .A2(n11414), .ZN(P3_U3233) );
  XNOR2_X1 U14065 ( .A(n11462), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n11420) );
  INV_X1 U14066 ( .A(n11422), .ZN(n11416) );
  NOR2_X1 U14067 ( .A1(n11416), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n11417) );
  OR2_X1 U14068 ( .A1(n11418), .A2(n11417), .ZN(n11419) );
  AOI211_X1 U14069 ( .C1(n11420), .C2(n11419), .A(n15597), .B(n11459), .ZN(
        n11432) );
  NAND2_X1 U14070 ( .A1(n11422), .A2(n11421), .ZN(n11423) );
  NAND2_X1 U14071 ( .A1(n11424), .A2(n11423), .ZN(n11428) );
  INV_X1 U14072 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11425) );
  MUX2_X1 U14073 ( .A(n11425), .B(P2_REG2_REG_10__SCAN_IN), .S(n11462), .Z(
        n11427) );
  INV_X1 U14074 ( .A(n11464), .ZN(n11426) );
  AOI211_X1 U14075 ( .C1(n11428), .C2(n11427), .A(n15591), .B(n11426), .ZN(
        n11431) );
  INV_X1 U14076 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n11945) );
  NAND2_X1 U14077 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n12234)
         );
  NAND2_X1 U14078 ( .A1(n15587), .A2(n11462), .ZN(n11429) );
  OAI211_X1 U14079 ( .C1(n15618), .C2(n11945), .A(n12234), .B(n11429), .ZN(
        n11430) );
  OR3_X1 U14080 ( .A1(n11432), .A2(n11431), .A3(n11430), .ZN(P2_U3224) );
  INV_X1 U14081 ( .A(n11433), .ZN(n11481) );
  INV_X1 U14082 ( .A(n14062), .ZN(n14055) );
  OAI222_X1 U14083 ( .A1(n14637), .A2(n11481), .B1(n14646), .B2(n11434), .C1(
        n14055), .C2(P2_U3088), .ZN(P2_U3309) );
  OAI222_X1 U14084 ( .A1(n13805), .A2(n11436), .B1(P3_U3151), .B2(n13031), 
        .C1(n13808), .C2(n11435), .ZN(P3_U3276) );
  OR2_X1 U14085 ( .A1(n13007), .A2(n11437), .ZN(n11438) );
  NAND2_X1 U14086 ( .A1(n11439), .A2(n11438), .ZN(n15672) );
  NAND2_X1 U14087 ( .A1(n15672), .A2(n13718), .ZN(n11447) );
  AOI22_X1 U14088 ( .A1(n13722), .A2(n13385), .B1(n13724), .B2(n11181), .ZN(
        n11446) );
  NAND3_X1 U14089 ( .A1(n13719), .A2(n13007), .A3(n11442), .ZN(n11443) );
  NAND2_X1 U14090 ( .A1(n11725), .A2(n11443), .ZN(n11444) );
  NAND2_X1 U14091 ( .A1(n11444), .A2(n13728), .ZN(n11445) );
  NAND3_X1 U14092 ( .A1(n11447), .A2(n11446), .A3(n11445), .ZN(n15678) );
  NAND2_X1 U14093 ( .A1(n15672), .A2(n15720), .ZN(n11449) );
  NAND2_X1 U14094 ( .A1(n15703), .A2(n6973), .ZN(n15673) );
  NAND2_X1 U14095 ( .A1(n11449), .A2(n15673), .ZN(n11450) );
  NOR2_X1 U14096 ( .A1(n15678), .A2(n11450), .ZN(n15694) );
  MUX2_X1 U14097 ( .A(n11451), .B(n15694), .S(n15734), .Z(n11452) );
  INV_X1 U14098 ( .A(n11452), .ZN(P3_U3461) );
  INV_X1 U14099 ( .A(n11453), .ZN(n11457) );
  OAI222_X1 U14100 ( .A1(n11455), .A2(P2_U3088), .B1(n14637), .B2(n11457), 
        .C1(n11454), .C2(n14646), .ZN(P2_U3308) );
  OAI222_X1 U14101 ( .A1(n11458), .A2(P1_U3086), .B1(n15433), .B2(n11457), 
        .C1(n11456), .C2(n15435), .ZN(P1_U3336) );
  XNOR2_X1 U14102 ( .A(n12453), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n12464) );
  XNOR2_X1 U14103 ( .A(n12465), .B(n12464), .ZN(n11470) );
  NOR2_X1 U14104 ( .A1(n11460), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12490) );
  NOR2_X1 U14105 ( .A1(n15608), .A2(n12462), .ZN(n11461) );
  AOI211_X1 U14106 ( .C1(n15585), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n12490), 
        .B(n11461), .ZN(n11469) );
  NAND2_X1 U14107 ( .A1(n11462), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11463) );
  MUX2_X1 U14108 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n9074), .S(n12453), .Z(
        n11465) );
  NAND2_X1 U14109 ( .A1(n11466), .A2(n11465), .ZN(n15574) );
  OAI21_X1 U14110 ( .B1(n11466), .B2(n11465), .A(n15574), .ZN(n11467) );
  NAND2_X1 U14111 ( .A1(n11467), .A2(n15613), .ZN(n11468) );
  OAI211_X1 U14112 ( .C1(n11470), .C2(n15597), .A(n11469), .B(n11468), .ZN(
        P2_U3225) );
  INV_X1 U14113 ( .A(n13860), .ZN(n11472) );
  NOR2_X1 U14114 ( .A1(n11472), .A2(n11471), .ZN(n11476) );
  INV_X1 U14115 ( .A(n13822), .ZN(n11474) );
  NAND2_X1 U14116 ( .A1(n11474), .A2(n11473), .ZN(n11475) );
  NOR2_X1 U14117 ( .A1(n11476), .A2(n11475), .ZN(n13823) );
  AOI21_X1 U14118 ( .B1(n11476), .B2(n11475), .A(n13823), .ZN(n11480) );
  OR2_X1 U14119 ( .A1(n11477), .A2(n15642), .ZN(n13858) );
  AOI22_X1 U14120 ( .A1(n13954), .A2(n11979), .B1(n13858), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n11479) );
  INV_X1 U14121 ( .A(n13941), .ZN(n13857) );
  AOI22_X1 U14122 ( .A1(n13857), .A2(n9353), .B1(n13937), .B2(n13978), .ZN(
        n11478) );
  OAI211_X1 U14123 ( .C1(n11480), .C2(n13956), .A(n11479), .B(n11478), .ZN(
        P2_U3209) );
  INV_X1 U14124 ( .A(n14983), .ZN(n14974) );
  OAI222_X1 U14125 ( .A1(P1_U3086), .A2(n14974), .B1(n15435), .B2(n11482), 
        .C1(n15433), .C2(n11481), .ZN(P1_U3337) );
  AOI21_X1 U14126 ( .B1(n11484), .B2(n14320), .A(n11483), .ZN(n11488) );
  AOI22_X1 U14127 ( .A1(n13937), .A2(n9353), .B1(n11485), .B2(n13954), .ZN(
        n11487) );
  NAND2_X1 U14128 ( .A1(n13858), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n11486) );
  OAI211_X1 U14129 ( .C1(n11488), .C2(n13956), .A(n11487), .B(n11486), .ZN(
        P2_U3204) );
  AND2_X1 U14130 ( .A1(n11490), .A2(n11489), .ZN(n11493) );
  INV_X1 U14131 ( .A(n11491), .ZN(n11492) );
  NAND2_X1 U14132 ( .A1(n11493), .A2(n11492), .ZN(n13202) );
  INV_X1 U14133 ( .A(n11494), .ZN(n11495) );
  NAND2_X1 U14134 ( .A1(n11496), .A2(n11495), .ZN(n15217) );
  OAI22_X1 U14135 ( .A1(n15234), .A2(n11498), .B1(n15217), .B2(n14822), .ZN(
        n11499) );
  AOI21_X1 U14136 ( .B1(n15522), .B2(n11500), .A(n11499), .ZN(n11504) );
  MUX2_X1 U14137 ( .A(n11502), .B(n11501), .S(n15533), .Z(n11503) );
  OAI211_X1 U14138 ( .C1(n15248), .C2(n11505), .A(n11504), .B(n11503), .ZN(
        P1_U3292) );
  OAI21_X1 U14139 ( .B1(n11507), .B2(n11512), .A(n11506), .ZN(n11560) );
  INV_X1 U14140 ( .A(n11508), .ZN(n11510) );
  AOI211_X1 U14141 ( .C1(n11830), .C2(n11510), .A(n15270), .B(n11509), .ZN(
        n11566) );
  XNOR2_X1 U14142 ( .A(n11511), .B(n11512), .ZN(n11516) );
  NAND2_X1 U14143 ( .A1(n14817), .A2(n15258), .ZN(n11514) );
  NAND2_X1 U14144 ( .A1(n14819), .A2(n15257), .ZN(n11513) );
  NAND2_X1 U14145 ( .A1(n11514), .A2(n11513), .ZN(n11831) );
  INV_X1 U14146 ( .A(n11831), .ZN(n11515) );
  OAI21_X1 U14147 ( .B1(n11516), .B2(n15160), .A(n11515), .ZN(n11561) );
  AOI211_X1 U14148 ( .C1(n15370), .C2(n11560), .A(n11566), .B(n11561), .ZN(
        n11519) );
  AOI22_X1 U14149 ( .A1(n12478), .A2(n11830), .B1(n15549), .B2(
        P1_REG0_REG_4__SCAN_IN), .ZN(n11517) );
  OAI21_X1 U14150 ( .B1(n11519), .B2(n15549), .A(n11517), .ZN(P1_U3471) );
  AOI22_X1 U14151 ( .A1(n12686), .A2(n11830), .B1(n15552), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n11518) );
  OAI21_X1 U14152 ( .B1(n11519), .B2(n15552), .A(n11518), .ZN(P1_U3532) );
  AOI21_X1 U14153 ( .B1(n11522), .B2(n11521), .A(n11520), .ZN(n11536) );
  INV_X1 U14154 ( .A(n13486), .ZN(n13501) );
  INV_X1 U14155 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n11523) );
  NAND2_X1 U14156 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n12345) );
  OAI21_X1 U14157 ( .B1(n13499), .B2(n11523), .A(n12345), .ZN(n11528) );
  NAND3_X1 U14158 ( .A1(n11350), .A2(n11525), .A3(n11524), .ZN(n11526) );
  AOI21_X1 U14159 ( .B1(n6619), .B2(n11526), .A(n13490), .ZN(n11527) );
  AOI211_X1 U14160 ( .C1(n13501), .C2(n11529), .A(n11528), .B(n11527), .ZN(
        n11535) );
  AND3_X1 U14161 ( .A1(n11532), .A2(n11531), .A3(n11530), .ZN(n11533) );
  OAI21_X1 U14162 ( .B1(n7493), .B2(n11533), .A(n13495), .ZN(n11534) );
  OAI211_X1 U14163 ( .C1(n11536), .C2(n13407), .A(n11535), .B(n11534), .ZN(
        P3_U3190) );
  AOI21_X1 U14164 ( .B1(n11538), .B2(n11537), .A(n14797), .ZN(n11540) );
  NAND2_X1 U14165 ( .A1(n11540), .A2(n11539), .ZN(n11544) );
  INV_X1 U14166 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n15525) );
  NAND2_X1 U14167 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n14855) );
  OAI21_X1 U14168 ( .B1(n14778), .B2(n11541), .A(n14855), .ZN(n11542) );
  AOI21_X1 U14169 ( .B1(n14776), .B2(n15525), .A(n11542), .ZN(n11543) );
  OAI211_X1 U14170 ( .C1(n11545), .C2(n14763), .A(n11544), .B(n11543), .ZN(
        P1_U3218) );
  INV_X1 U14171 ( .A(n11546), .ZN(n11547) );
  NAND2_X1 U14172 ( .A1(n11547), .A2(n6974), .ZN(n11550) );
  XNOR2_X1 U14173 ( .A(n12935), .B(n11548), .ZN(n11580) );
  XNOR2_X1 U14174 ( .A(n11580), .B(n13385), .ZN(n11551) );
  AOI21_X1 U14175 ( .B1(n11553), .B2(n11550), .A(n11551), .ZN(n11559) );
  AND2_X1 U14176 ( .A1(n11551), .A2(n11550), .ZN(n11552) );
  NAND2_X1 U14177 ( .A1(n11583), .A2(n13353), .ZN(n11558) );
  MUX2_X1 U14178 ( .A(P3_U3151), .B(n13362), .S(n11732), .Z(n11556) );
  OAI22_X1 U14179 ( .A1(n13331), .A2(n11782), .B1(n13367), .B2(n11731), .ZN(
        n11555) );
  AOI211_X1 U14180 ( .C1(n13328), .C2(n13721), .A(n11556), .B(n11555), .ZN(
        n11557) );
  OAI21_X1 U14181 ( .B1(n11559), .B2(n11558), .A(n11557), .ZN(P3_U3158) );
  INV_X1 U14182 ( .A(n11560), .ZN(n11569) );
  INV_X1 U14183 ( .A(n11561), .ZN(n11562) );
  INV_X2 U14184 ( .A(n15533), .ZN(n15220) );
  MUX2_X1 U14185 ( .A(n11563), .B(n11562), .S(n15220), .Z(n11568) );
  OAI22_X1 U14186 ( .A1(n15234), .A2(n11564), .B1(n15217), .B2(n11834), .ZN(
        n11565) );
  AOI21_X1 U14187 ( .B1(n11566), .B2(n15522), .A(n11565), .ZN(n11567) );
  OAI211_X1 U14188 ( .C1(n11569), .C2(n15248), .A(n11568), .B(n11567), .ZN(
        P1_U3289) );
  INV_X1 U14189 ( .A(n11570), .ZN(n11573) );
  OAI22_X1 U14190 ( .A1(n13952), .A2(n11958), .B1(n11571), .B2(n13908), .ZN(
        n11572) );
  AOI211_X1 U14191 ( .C1(n13857), .C2(n13977), .A(n11573), .B(n11572), .ZN(
        n11579) );
  OAI21_X1 U14192 ( .B1(n11576), .B2(n11575), .A(n11574), .ZN(n11577) );
  NAND2_X1 U14193 ( .A1(n11577), .A2(n13915), .ZN(n11578) );
  OAI211_X1 U14194 ( .C1(n7628), .C2(n13925), .A(n11579), .B(n11578), .ZN(
        P2_U3199) );
  AOI21_X1 U14195 ( .B1(n11588), .B2(n11587), .A(n6623), .ZN(n11594) );
  INV_X1 U14196 ( .A(n11696), .ZN(n11592) );
  AOI22_X1 U14197 ( .A1(n13328), .A2(n13385), .B1(n13357), .B2(n13384), .ZN(
        n11590) );
  OAI211_X1 U14198 ( .C1(n13367), .C2(n15699), .A(n11590), .B(n11589), .ZN(
        n11591) );
  AOI21_X1 U14199 ( .B1(n11592), .B2(n13362), .A(n11591), .ZN(n11593) );
  OAI21_X1 U14200 ( .B1(n11594), .B2(n13351), .A(n11593), .ZN(P3_U3170) );
  NOR2_X1 U14201 ( .A1(n9354), .A2(n11595), .ZN(n11621) );
  INV_X1 U14202 ( .A(n11596), .ZN(n11598) );
  OAI21_X1 U14203 ( .B1(n12060), .B2(n14339), .A(n11622), .ZN(n11597) );
  AOI21_X1 U14204 ( .B1(n11621), .B2(n11598), .A(n11620), .ZN(n11603) );
  INV_X1 U14205 ( .A(n12069), .ZN(n11601) );
  INV_X1 U14206 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n13986) );
  OAI22_X1 U14207 ( .A1(n15622), .A2(n13986), .B1(n11599), .B2(n15619), .ZN(
        n11600) );
  AOI21_X1 U14208 ( .B1(n11601), .B2(n11622), .A(n11600), .ZN(n11602) );
  OAI21_X1 U14209 ( .B1(n14341), .B2(n11603), .A(n11602), .ZN(P2_U3265) );
  NOR2_X1 U14210 ( .A1(n11609), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11605) );
  XNOR2_X1 U14211 ( .A(n11663), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n11604) );
  INV_X1 U14212 ( .A(n11658), .ZN(n11608) );
  OAI21_X1 U14213 ( .B1(n11606), .B2(n11605), .A(n11604), .ZN(n11607) );
  NAND3_X1 U14214 ( .A1(n11608), .A2(n15506), .A3(n11607), .ZN(n11618) );
  NAND2_X1 U14215 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14743)
         );
  MUX2_X1 U14216 ( .A(n12717), .B(P1_REG2_REG_13__SCAN_IN), .S(n11663), .Z(
        n11612) );
  OR2_X1 U14217 ( .A1(n11609), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11610) );
  NAND2_X1 U14218 ( .A1(n11611), .A2(n11610), .ZN(n11613) );
  AOI21_X1 U14219 ( .B1(n11612), .B2(n11613), .A(n14989), .ZN(n11614) );
  NAND2_X1 U14220 ( .A1(n11614), .A2(n11669), .ZN(n11615) );
  NAND2_X1 U14221 ( .A1(n14743), .A2(n11615), .ZN(n11616) );
  AOI21_X1 U14222 ( .B1(n15492), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11616), 
        .ZN(n11617) );
  OAI211_X1 U14223 ( .C1(n14975), .C2(n11619), .A(n11618), .B(n11617), .ZN(
        P1_U3256) );
  INV_X1 U14224 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n11624) );
  AOI211_X1 U14225 ( .C1(n15653), .C2(n11622), .A(n11621), .B(n11620), .ZN(
        n11625) );
  OR2_X1 U14226 ( .A1(n11625), .A2(n15664), .ZN(n11623) );
  OAI21_X1 U14227 ( .B1(n15666), .B2(n11624), .A(n11623), .ZN(P2_U3430) );
  OR2_X1 U14228 ( .A1(n11625), .A2(n15668), .ZN(n11626) );
  OAI21_X1 U14229 ( .B1(n15670), .B2(n11049), .A(n11626), .ZN(P2_U3499) );
  XNOR2_X1 U14230 ( .A(n11628), .B(n11627), .ZN(n11636) );
  INV_X1 U14231 ( .A(n12065), .ZN(n11633) );
  NAND2_X1 U14232 ( .A1(n13974), .A2(n14286), .ZN(n11630) );
  NAND2_X1 U14233 ( .A1(n13976), .A2(n14285), .ZN(n11629) );
  NAND2_X1 U14234 ( .A1(n11630), .A2(n11629), .ZN(n12058) );
  INV_X1 U14235 ( .A(n12058), .ZN(n11631) );
  NAND2_X1 U14236 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n14020) );
  OAI21_X1 U14237 ( .B1(n13891), .B2(n11631), .A(n14020), .ZN(n11632) );
  AOI21_X1 U14238 ( .B1(n11633), .B2(n13938), .A(n11632), .ZN(n11635) );
  NAND2_X1 U14239 ( .A1(n13954), .A2(n12064), .ZN(n11634) );
  OAI211_X1 U14240 ( .C1(n11636), .C2(n13956), .A(n11635), .B(n11634), .ZN(
        P2_U3211) );
  INV_X1 U14241 ( .A(n11637), .ZN(n11638) );
  AOI21_X1 U14242 ( .B1(n11640), .B2(n11639), .A(n11638), .ZN(n11645) );
  INV_X1 U14243 ( .A(n11940), .ZN(n11641) );
  AOI22_X1 U14244 ( .A1(n13937), .A2(n13976), .B1(n13938), .B2(n11641), .ZN(
        n11642) );
  NAND2_X1 U14245 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n13997) );
  OAI211_X1 U14246 ( .C1(n11982), .C2(n13941), .A(n11642), .B(n13997), .ZN(
        n11643) );
  AOI21_X1 U14247 ( .B1(n15657), .B2(n13954), .A(n11643), .ZN(n11644) );
  OAI21_X1 U14248 ( .B1(n11645), .B2(n13956), .A(n11644), .ZN(P2_U3202) );
  INV_X1 U14249 ( .A(n11646), .ZN(n11647) );
  NAND2_X1 U14250 ( .A1(n11648), .A2(n11647), .ZN(n11649) );
  NAND2_X1 U14251 ( .A1(n11652), .A2(n11651), .ZN(n11655) );
  NAND2_X1 U14252 ( .A1(n11653), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n11654) );
  NAND2_X1 U14253 ( .A1(n11655), .A2(n11654), .ZN(n11796) );
  NAND2_X1 U14254 ( .A1(n14468), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n11797) );
  OAI21_X1 U14255 ( .B1(n14468), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11797), .ZN(
        n11656) );
  XNOR2_X1 U14256 ( .A(n11796), .B(n11656), .ZN(n11791) );
  INV_X1 U14257 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n11789) );
  XNOR2_X1 U14258 ( .A(n11790), .B(n11789), .ZN(SUB_1596_U54) );
  XNOR2_X1 U14259 ( .A(n12124), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n11660) );
  AND2_X1 U14260 ( .A1(n11663), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11657) );
  OR2_X1 U14261 ( .A1(n11658), .A2(n11657), .ZN(n11659) );
  AOI21_X1 U14262 ( .B1(n11660), .B2(n11659), .A(n12121), .ZN(n11673) );
  INV_X1 U14263 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n11661) );
  NAND2_X1 U14264 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n14652)
         );
  OAI21_X1 U14265 ( .B1(n15497), .B2(n11661), .A(n14652), .ZN(n11662) );
  AOI21_X1 U14266 ( .B1(n12124), .B2(n15500), .A(n11662), .ZN(n11672) );
  NAND2_X1 U14267 ( .A1(n11663), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11668) );
  NAND2_X1 U14268 ( .A1(n11669), .A2(n11668), .ZN(n11666) );
  INV_X1 U14269 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11664) );
  MUX2_X1 U14270 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11664), .S(n12124), .Z(
        n11665) );
  NAND2_X1 U14271 ( .A1(n11666), .A2(n11665), .ZN(n12126) );
  MUX2_X1 U14272 ( .A(n11664), .B(P1_REG2_REG_14__SCAN_IN), .S(n12124), .Z(
        n11667) );
  NAND3_X1 U14273 ( .A1(n11669), .A2(n11668), .A3(n11667), .ZN(n11670) );
  NAND3_X1 U14274 ( .A1(n12126), .A2(n15513), .A3(n11670), .ZN(n11671) );
  OAI211_X1 U14275 ( .C1(n11673), .C2(n14942), .A(n11672), .B(n11671), .ZN(
        P1_U3257) );
  INV_X1 U14276 ( .A(n15248), .ZN(n15519) );
  NAND2_X1 U14277 ( .A1(n15522), .A2(n11674), .ZN(n11678) );
  NOR2_X1 U14278 ( .A1(n15217), .A2(n11675), .ZN(n11676) );
  AOI21_X1 U14279 ( .B1(n15533), .B2(P1_REG2_REG_2__SCAN_IN), .A(n11676), .ZN(
        n11677) );
  OAI211_X1 U14280 ( .C1(n7048), .C2(n15234), .A(n11678), .B(n11677), .ZN(
        n11679) );
  AOI21_X1 U14281 ( .B1(n15519), .B2(n11680), .A(n11679), .ZN(n11681) );
  OAI21_X1 U14282 ( .B1(n15533), .B2(n11682), .A(n11681), .ZN(P1_U3291) );
  INV_X1 U14283 ( .A(n11683), .ZN(n11685) );
  OAI211_X1 U14284 ( .C1(n11686), .C2(n15660), .A(n11685), .B(n11684), .ZN(
        n11692) );
  INV_X1 U14285 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n11687) );
  OAI22_X1 U14286 ( .A1(n14627), .A2(n11690), .B1(n15666), .B2(n11687), .ZN(
        n11688) );
  AOI21_X1 U14287 ( .B1(n11692), .B2(n15666), .A(n11688), .ZN(n11689) );
  INV_X1 U14288 ( .A(n11689), .ZN(P2_U3433) );
  OAI22_X1 U14289 ( .A1(n14582), .A2(n11690), .B1(n15670), .B2(n8964), .ZN(
        n11691) );
  AOI21_X1 U14290 ( .B1(n11692), .B2(n15670), .A(n11691), .ZN(n11693) );
  INV_X1 U14291 ( .A(n11693), .ZN(P2_U3500) );
  XNOR2_X1 U14292 ( .A(n11694), .B(n13074), .ZN(n15702) );
  INV_X1 U14293 ( .A(n11695), .ZN(n15675) );
  OR2_X1 U14294 ( .A1(n15691), .A2(n15675), .ZN(n12230) );
  INV_X1 U14295 ( .A(n12230), .ZN(n15687) );
  OAI22_X1 U14296 ( .A1(n13588), .A2(n15699), .B1(n11696), .B2(n13645), .ZN(
        n11703) );
  XNOR2_X1 U14297 ( .A(n11698), .B(n11697), .ZN(n11701) );
  NAND2_X1 U14298 ( .A1(n15702), .A2(n13718), .ZN(n11700) );
  AOI22_X1 U14299 ( .A1(n13722), .A2(n13384), .B1(n13724), .B2(n13385), .ZN(
        n11699) );
  OAI211_X1 U14300 ( .C1(n13638), .C2(n11701), .A(n11700), .B(n11699), .ZN(
        n15700) );
  MUX2_X1 U14301 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n15700), .S(n9345), .Z(
        n11702) );
  AOI211_X1 U14302 ( .C1(n15702), .C2(n15687), .A(n11703), .B(n11702), .ZN(
        n11704) );
  INV_X1 U14303 ( .A(n11704), .ZN(P3_U3229) );
  NAND2_X1 U14304 ( .A1(n10753), .A2(n11705), .ZN(n11968) );
  NAND2_X1 U14305 ( .A1(n11968), .A2(n10331), .ZN(n11969) );
  NAND3_X1 U14306 ( .A1(n11969), .A2(n11710), .A3(n11706), .ZN(n11708) );
  NAND2_X1 U14307 ( .A1(n11708), .A2(n11707), .ZN(n12267) );
  INV_X1 U14308 ( .A(n12267), .ZN(n11713) );
  OAI21_X1 U14309 ( .B1(n11711), .B2(n11710), .A(n11709), .ZN(n11712) );
  AOI222_X1 U14310 ( .A1(n14339), .A2(n11712), .B1(n13977), .B2(n14286), .C1(
        n9514), .C2(n14285), .ZN(n12261) );
  OAI211_X1 U14311 ( .C1(n11972), .C2(n12264), .A(n14310), .B(n11937), .ZN(
        n12263) );
  OAI211_X1 U14312 ( .C1(n14575), .C2(n11713), .A(n12261), .B(n12263), .ZN(
        n11719) );
  OAI22_X1 U14313 ( .A1(n14582), .A2(n12264), .B1(n15670), .B2(n11714), .ZN(
        n11715) );
  AOI21_X1 U14314 ( .B1(n11719), .B2(n15670), .A(n11715), .ZN(n11716) );
  INV_X1 U14315 ( .A(n11716), .ZN(P2_U3502) );
  INV_X1 U14316 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11717) );
  OAI22_X1 U14317 ( .A1(n14627), .A2(n12264), .B1(n15666), .B2(n11717), .ZN(
        n11718) );
  AOI21_X1 U14318 ( .B1(n11719), .B2(n15666), .A(n11718), .ZN(n11720) );
  INV_X1 U14319 ( .A(n11720), .ZN(P2_U3439) );
  XNOR2_X1 U14320 ( .A(n11721), .B(n11722), .ZN(n15698) );
  INV_X1 U14321 ( .A(n15698), .ZN(n11736) );
  OAI22_X1 U14322 ( .A1(n6974), .A2(n13641), .B1(n13643), .B2(n11782), .ZN(
        n11729) );
  INV_X1 U14323 ( .A(n11723), .ZN(n11727) );
  AOI21_X1 U14324 ( .B1(n11725), .B2(n11724), .A(n13009), .ZN(n11726) );
  NOR3_X1 U14325 ( .A1(n11727), .A2(n11726), .A3(n13638), .ZN(n11728) );
  AOI211_X1 U14326 ( .C1(n15698), .C2(n13718), .A(n11729), .B(n11728), .ZN(
        n15695) );
  MUX2_X1 U14327 ( .A(n11730), .B(n15695), .S(n9345), .Z(n11735) );
  INV_X1 U14328 ( .A(n11989), .ZN(n11733) );
  NOR2_X1 U14329 ( .A1(n15715), .A2(n11731), .ZN(n15697) );
  AOI22_X1 U14330 ( .A1(n11733), .A2(n15697), .B1(n15685), .B2(n11732), .ZN(
        n11734) );
  OAI211_X1 U14331 ( .C1(n11736), .C2(n12230), .A(n11735), .B(n11734), .ZN(
        P3_U3230) );
  OR2_X1 U14332 ( .A1(n11737), .A2(n13079), .ZN(n11738) );
  NAND2_X1 U14333 ( .A1(n11739), .A2(n11738), .ZN(n15705) );
  INV_X1 U14334 ( .A(n15705), .ZN(n11747) );
  INV_X1 U14335 ( .A(n13383), .ZN(n12357) );
  OAI22_X1 U14336 ( .A1(n12357), .A2(n13643), .B1(n13641), .B2(n11782), .ZN(
        n11743) );
  OR2_X1 U14337 ( .A1(n11740), .A2(n13079), .ZN(n11994) );
  NAND2_X1 U14338 ( .A1(n11740), .A2(n13079), .ZN(n11741) );
  AOI21_X1 U14339 ( .B1(n11994), .B2(n11741), .A(n13638), .ZN(n11742) );
  AOI211_X1 U14340 ( .C1(n13718), .C2(n15705), .A(n11743), .B(n11742), .ZN(
        n15707) );
  MUX2_X1 U14341 ( .A(n14433), .B(n15707), .S(n9345), .Z(n11746) );
  INV_X1 U14342 ( .A(n11779), .ZN(n15704) );
  INV_X1 U14343 ( .A(n11744), .ZN(n11785) );
  AOI22_X1 U14344 ( .A1(n13659), .A2(n15704), .B1(n15685), .B2(n11785), .ZN(
        n11745) );
  OAI211_X1 U14345 ( .C1(n11747), .C2(n12230), .A(n11746), .B(n11745), .ZN(
        P3_U3228) );
  XNOR2_X1 U14346 ( .A(n11749), .B(n11748), .ZN(n11758) );
  INV_X1 U14347 ( .A(n15620), .ZN(n11755) );
  NAND2_X1 U14348 ( .A1(n13973), .A2(n14286), .ZN(n11751) );
  NAND2_X1 U14349 ( .A1(n13975), .A2(n14285), .ZN(n11750) );
  NAND2_X1 U14350 ( .A1(n11751), .A2(n11750), .ZN(n12249) );
  INV_X1 U14351 ( .A(n12249), .ZN(n11753) );
  OAI21_X1 U14352 ( .B1(n13891), .B2(n11753), .A(n11752), .ZN(n11754) );
  AOI21_X1 U14353 ( .B1(n11755), .B2(n13938), .A(n11754), .ZN(n11757) );
  NAND2_X1 U14354 ( .A1(n13954), .A2(n15624), .ZN(n11756) );
  OAI211_X1 U14355 ( .C1(n11758), .C2(n13956), .A(n11757), .B(n11756), .ZN(
        P2_U3185) );
  INV_X1 U14356 ( .A(n11759), .ZN(n11769) );
  OAI22_X1 U14357 ( .A1(n11865), .A2(n15239), .B1(n11903), .B2(n15241), .ZN(
        n11768) );
  INV_X1 U14358 ( .A(n11760), .ZN(n11763) );
  NAND3_X1 U14359 ( .A1(n11506), .A2(n15370), .A3(n11761), .ZN(n11762) );
  OAI21_X1 U14360 ( .B1(n11763), .B2(n15160), .A(n11762), .ZN(n11766) );
  NOR2_X1 U14361 ( .A1(n11760), .A2(n15160), .ZN(n11765) );
  MUX2_X1 U14362 ( .A(n11766), .B(n11765), .S(n11764), .Z(n11767) );
  AOI211_X1 U14363 ( .C1(n15370), .C2(n11769), .A(n11768), .B(n11767), .ZN(
        n11807) );
  OAI211_X1 U14364 ( .C1(n11509), .C2(n11770), .A(n15168), .B(n11871), .ZN(
        n11812) );
  AND2_X1 U14365 ( .A1(n11807), .A2(n11812), .ZN(n11773) );
  AOI22_X1 U14366 ( .A1(n12686), .A2(n11868), .B1(n15552), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n11771) );
  OAI21_X1 U14367 ( .B1(n11773), .B2(n15552), .A(n11771), .ZN(P1_U3533) );
  AOI22_X1 U14368 ( .A1(n12478), .A2(n11868), .B1(n15549), .B2(
        P1_REG0_REG_5__SCAN_IN), .ZN(n11772) );
  OAI21_X1 U14369 ( .B1(n11773), .B2(n15549), .A(n11772), .ZN(P1_U3474) );
  INV_X1 U14370 ( .A(n11774), .ZN(n11813) );
  OAI222_X1 U14371 ( .A1(n15435), .A2(n11776), .B1(n15433), .B2(n11813), .C1(
        n11775), .C2(P1_U3086), .ZN(P1_U3335) );
  INV_X1 U14372 ( .A(n11777), .ZN(n11778) );
  XNOR2_X1 U14373 ( .A(n12932), .B(n11779), .ZN(n12159) );
  XNOR2_X1 U14374 ( .A(n12159), .B(n13384), .ZN(n11780) );
  AOI21_X1 U14375 ( .B1(n11781), .B2(n11780), .A(n12161), .ZN(n11788) );
  INV_X1 U14376 ( .A(n13367), .ZN(n13349) );
  OAI22_X1 U14377 ( .A1(n13331), .A2(n12357), .B1(n11782), .B2(n13359), .ZN(
        n11783) );
  AOI211_X1 U14378 ( .C1(n13349), .C2(n15704), .A(n11784), .B(n11783), .ZN(
        n11787) );
  NAND2_X1 U14379 ( .A1(n13362), .A2(n11785), .ZN(n11786) );
  OAI211_X1 U14380 ( .C1(n11788), .C2(n13351), .A(n11787), .B(n11786), .ZN(
        P3_U3167) );
  INV_X1 U14381 ( .A(n11791), .ZN(n11792) );
  OR2_X1 U14382 ( .A1(n14468), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n11795) );
  NAND2_X1 U14383 ( .A1(n11796), .A2(n11795), .ZN(n11798) );
  NAND2_X1 U14384 ( .A1(n11798), .A2(n11797), .ZN(n11948) );
  INV_X1 U14385 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14922) );
  NAND2_X1 U14386 ( .A1(n14922), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n11949) );
  INV_X1 U14387 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n11799) );
  NAND2_X1 U14388 ( .A1(n11799), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n11800) );
  AND2_X1 U14389 ( .A1(n11949), .A2(n11800), .ZN(n11947) );
  INV_X1 U14390 ( .A(n11947), .ZN(n11801) );
  XNOR2_X1 U14391 ( .A(n11948), .B(n11801), .ZN(n11944) );
  XNOR2_X1 U14392 ( .A(n11944), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(n11802) );
  XNOR2_X1 U14393 ( .A(n11946), .B(n11802), .ZN(SUB_1596_U70) );
  INV_X1 U14394 ( .A(n11803), .ZN(n11805) );
  OAI222_X1 U14395 ( .A1(n13805), .A2(n11806), .B1(n13808), .B2(n11805), .C1(
        n11804), .C2(P3_U3151), .ZN(P3_U3275) );
  MUX2_X1 U14396 ( .A(n11808), .B(n11807), .S(n15220), .Z(n11811) );
  INV_X1 U14397 ( .A(n15217), .ZN(n15526) );
  INV_X1 U14398 ( .A(n11864), .ZN(n11809) );
  AOI22_X1 U14399 ( .A1(n15524), .A2(n11868), .B1(n15526), .B2(n11809), .ZN(
        n11810) );
  OAI211_X1 U14400 ( .C1(n15174), .C2(n11812), .A(n11811), .B(n11810), .ZN(
        P1_U3288) );
  OAI222_X1 U14401 ( .A1(P2_U3088), .A2(n11815), .B1(n14646), .B2(n11814), 
        .C1(n14637), .C2(n11813), .ZN(P2_U3307) );
  OAI211_X1 U14402 ( .C1(n11818), .C2(n11817), .A(n11816), .B(n14754), .ZN(
        n11822) );
  AND2_X1 U14403 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n14888) );
  INV_X1 U14404 ( .A(n14727), .ZN(n14789) );
  OAI22_X1 U14405 ( .A1(n11819), .A2(n14789), .B1(n14792), .B2(n11886), .ZN(
        n11820) );
  AOI211_X1 U14406 ( .C1(n14748), .C2(n14815), .A(n14888), .B(n11820), .ZN(
        n11821) );
  OAI211_X1 U14407 ( .C1(n7768), .C2(n14763), .A(n11822), .B(n11821), .ZN(
        P1_U3239) );
  INV_X1 U14408 ( .A(n11823), .ZN(n12980) );
  OAI222_X1 U14409 ( .A1(n11825), .A2(P1_U3086), .B1(n15433), .B2(n12980), 
        .C1(n11824), .C2(n15435), .ZN(P1_U3334) );
  XNOR2_X1 U14410 ( .A(n11827), .B(n11828), .ZN(n11857) );
  XNOR2_X1 U14411 ( .A(n11857), .B(n11829), .ZN(n11836) );
  NAND2_X1 U14412 ( .A1(n14795), .A2(n11830), .ZN(n11833) );
  AND2_X1 U14413 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n15499) );
  AOI21_X1 U14414 ( .B1(n14766), .B2(n11831), .A(n15499), .ZN(n11832) );
  OAI211_X1 U14415 ( .C1(n14792), .C2(n11834), .A(n11833), .B(n11832), .ZN(
        n11835) );
  AOI21_X1 U14416 ( .B1(n11836), .B2(n14754), .A(n11835), .ZN(n11837) );
  INV_X1 U14417 ( .A(n11837), .ZN(P1_U3230) );
  INV_X1 U14418 ( .A(n13395), .ZN(n11838) );
  AOI21_X1 U14419 ( .B1(n12297), .B2(n6628), .A(n11838), .ZN(n11854) );
  OAI21_X1 U14420 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n11840), .A(n11839), .ZN(
        n11852) );
  INV_X1 U14421 ( .A(n11845), .ZN(n11841) );
  NAND2_X1 U14422 ( .A1(n11842), .A2(n11841), .ZN(n11847) );
  OAI21_X1 U14423 ( .B1(n11845), .B2(n11844), .A(n11843), .ZN(n11846) );
  AOI21_X1 U14424 ( .B1(n11847), .B2(n11846), .A(n13407), .ZN(n11851) );
  NAND2_X1 U14425 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n12535) );
  NAND2_X1 U14426 ( .A1(n15671), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n11848) );
  OAI211_X1 U14427 ( .C1(n13486), .C2(n11849), .A(n12535), .B(n11848), .ZN(
        n11850) );
  AOI211_X1 U14428 ( .C1(n11852), .C2(n13504), .A(n11851), .B(n11850), .ZN(
        n11853) );
  OAI21_X1 U14429 ( .B1(n11854), .B2(n13461), .A(n11853), .ZN(P3_U3191) );
  AOI22_X1 U14430 ( .A1(n11857), .A2(n11856), .B1(n11827), .B2(n11855), .ZN(
        n11862) );
  OAI21_X1 U14431 ( .B1(n11860), .B2(n11859), .A(n11858), .ZN(n11861) );
  XNOR2_X1 U14432 ( .A(n11862), .B(n11861), .ZN(n11870) );
  OAI22_X1 U14433 ( .A1(n14790), .A2(n11903), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11863), .ZN(n11867) );
  OAI22_X1 U14434 ( .A1(n11865), .A2(n14789), .B1(n14792), .B2(n11864), .ZN(
        n11866) );
  AOI211_X1 U14435 ( .C1(n14795), .C2(n11868), .A(n11867), .B(n11866), .ZN(
        n11869) );
  OAI21_X1 U14436 ( .B1(n11870), .B2(n14797), .A(n11869), .ZN(P1_U3227) );
  INV_X1 U14437 ( .A(n11871), .ZN(n11872) );
  OAI211_X1 U14438 ( .C1(n11872), .C2(n7768), .A(n15168), .B(n12020), .ZN(
        n15540) );
  NOR2_X1 U14439 ( .A1(n11873), .A2(n15160), .ZN(n11878) );
  NAND3_X1 U14440 ( .A1(n11759), .A2(n15370), .A3(n11879), .ZN(n11875) );
  NAND2_X1 U14441 ( .A1(n11873), .A2(n15260), .ZN(n11874) );
  NAND2_X1 U14442 ( .A1(n11875), .A2(n11874), .ZN(n11877) );
  MUX2_X1 U14443 ( .A(n11878), .B(n11877), .S(n11876), .Z(n11884) );
  NAND2_X1 U14444 ( .A1(n11759), .A2(n11879), .ZN(n11881) );
  NAND2_X1 U14445 ( .A1(n11881), .A2(n11880), .ZN(n12025) );
  AOI22_X1 U14446 ( .A1(n15257), .A2(n14817), .B1(n14815), .B2(n15258), .ZN(
        n11882) );
  OAI21_X1 U14447 ( .B1(n12025), .B2(n15354), .A(n11882), .ZN(n11883) );
  OR2_X1 U14448 ( .A1(n11884), .A2(n11883), .ZN(n15541) );
  INV_X1 U14449 ( .A(n15541), .ZN(n11885) );
  MUX2_X1 U14450 ( .A(n11885), .B(n14889), .S(n15533), .Z(n11889) );
  INV_X1 U14451 ( .A(n11886), .ZN(n11887) );
  AOI22_X1 U14452 ( .A1(n15524), .A2(n15543), .B1(n11887), .B2(n15526), .ZN(
        n11888) );
  OAI211_X1 U14453 ( .C1(n15174), .C2(n15540), .A(n11889), .B(n11888), .ZN(
        P1_U3287) );
  AOI21_X1 U14454 ( .B1(n11890), .B2(n15220), .A(n15522), .ZN(n11896) );
  INV_X1 U14455 ( .A(n15220), .ZN(n15274) );
  OAI22_X1 U14456 ( .A1(n11892), .A2(n15274), .B1(n11891), .B2(n15217), .ZN(
        n11893) );
  AOI21_X1 U14457 ( .B1(n15533), .B2(P1_REG2_REG_0__SCAN_IN), .A(n11893), .ZN(
        n11894) );
  OAI21_X1 U14458 ( .B1(n11896), .B2(n11895), .A(n11894), .ZN(P1_U3293) );
  INV_X1 U14459 ( .A(SI_21_), .ZN(n11899) );
  INV_X1 U14460 ( .A(n11897), .ZN(n11898) );
  OAI222_X1 U14461 ( .A1(n13805), .A2(n11899), .B1(n13808), .B2(n11898), .C1(
        n13059), .C2(P3_U3151), .ZN(P3_U3274) );
  OAI211_X1 U14462 ( .C1(n11902), .C2(n11901), .A(n11900), .B(n14754), .ZN(
        n11906) );
  AND2_X1 U14463 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n14905) );
  OAI22_X1 U14464 ( .A1(n11903), .A2(n14789), .B1(n14792), .B2(n12036), .ZN(
        n11904) );
  AOI211_X1 U14465 ( .C1(n14748), .C2(n14814), .A(n14905), .B(n11904), .ZN(
        n11905) );
  OAI211_X1 U14466 ( .C1(n7767), .C2(n14763), .A(n11906), .B(n11905), .ZN(
        P1_U3213) );
  OAI21_X1 U14467 ( .B1(n11909), .B2(n11908), .A(n11907), .ZN(n11910) );
  INV_X1 U14468 ( .A(n11910), .ZN(n11963) );
  OAI21_X1 U14469 ( .B1(n11912), .B2(n11911), .A(n12054), .ZN(n11913) );
  AOI222_X1 U14470 ( .A1(n14339), .A2(n11913), .B1(n13975), .B2(n14286), .C1(
        n13977), .C2(n14285), .ZN(n11956) );
  AOI211_X1 U14471 ( .C1(n11914), .C2(n11938), .A(n14320), .B(n12062), .ZN(
        n11960) );
  INV_X1 U14472 ( .A(n11960), .ZN(n11915) );
  OAI211_X1 U14473 ( .C1(n14575), .C2(n11963), .A(n11956), .B(n11915), .ZN(
        n11921) );
  INV_X1 U14474 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11916) );
  OAI22_X1 U14475 ( .A1(n14627), .A2(n7628), .B1(n15666), .B2(n11916), .ZN(
        n11917) );
  AOI21_X1 U14476 ( .B1(n11921), .B2(n15666), .A(n11917), .ZN(n11918) );
  INV_X1 U14477 ( .A(n11918), .ZN(P2_U3445) );
  OAI22_X1 U14478 ( .A1(n14582), .A2(n7628), .B1(n15670), .B2(n11919), .ZN(
        n11920) );
  AOI21_X1 U14479 ( .B1(n11921), .B2(n15670), .A(n11920), .ZN(n11922) );
  INV_X1 U14480 ( .A(n11922), .ZN(P2_U3504) );
  INV_X1 U14481 ( .A(n11923), .ZN(n11925) );
  OAI222_X1 U14482 ( .A1(n14646), .A2(n11926), .B1(n14637), .B2(n11925), .C1(
        P2_U3088), .C2(n11924), .ZN(P2_U3305) );
  OR2_X1 U14483 ( .A1(n11927), .A2(n6872), .ZN(n11929) );
  AND2_X1 U14484 ( .A1(n11928), .A2(n11929), .ZN(n15661) );
  OAI21_X1 U14485 ( .B1(n11932), .B2(n11931), .A(n11930), .ZN(n11933) );
  NAND2_X1 U14486 ( .A1(n11933), .A2(n14339), .ZN(n11935) );
  AOI22_X1 U14487 ( .A1(n14285), .A2(n13978), .B1(n13976), .B2(n14286), .ZN(
        n11934) );
  OAI211_X1 U14488 ( .C1(n15661), .C2(n11986), .A(n11935), .B(n11934), .ZN(
        n15663) );
  MUX2_X1 U14489 ( .A(n15663), .B(P2_REG2_REG_4__SCAN_IN), .S(n14341), .Z(
        n11936) );
  INV_X1 U14490 ( .A(n11936), .ZN(n11943) );
  AOI21_X1 U14491 ( .B1(n11937), .B2(n15657), .A(n14320), .ZN(n11939) );
  AND2_X1 U14492 ( .A1(n11939), .A2(n11938), .ZN(n15655) );
  AOI21_X1 U14493 ( .B1(n14344), .B2(n15655), .A(n11941), .ZN(n11942) );
  OAI211_X1 U14494 ( .C1(n15661), .C2(n12069), .A(n11943), .B(n11942), .ZN(
        P2_U3261) );
  NAND2_X1 U14495 ( .A1(n11948), .A2(n11947), .ZN(n11950) );
  NAND2_X1 U14496 ( .A1(n11950), .A2(n11949), .ZN(n12322) );
  INV_X1 U14497 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n11951) );
  NAND2_X1 U14498 ( .A1(n11951), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n12323) );
  INV_X1 U14499 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n11952) );
  NAND2_X1 U14500 ( .A1(n11952), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n11953) );
  AND2_X1 U14501 ( .A1(n12323), .A2(n11953), .ZN(n12321) );
  INV_X1 U14502 ( .A(n12321), .ZN(n11954) );
  XNOR2_X1 U14503 ( .A(n12322), .B(n11954), .ZN(n12316) );
  XNOR2_X1 U14504 ( .A(n12316), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(n11955) );
  XNOR2_X1 U14505 ( .A(n12318), .B(n11955), .ZN(SUB_1596_U69) );
  MUX2_X1 U14506 ( .A(n11957), .B(n11956), .S(n15622), .Z(n11962) );
  OAI22_X1 U14507 ( .A1(n14326), .A2(n7628), .B1(n15619), .B2(n11958), .ZN(
        n11959) );
  AOI21_X1 U14508 ( .B1(n11960), .B2(n14344), .A(n11959), .ZN(n11961) );
  OAI211_X1 U14509 ( .C1(n11963), .C2(n14346), .A(n11962), .B(n11961), .ZN(
        P2_U3260) );
  AOI22_X1 U14510 ( .A1(n11964), .A2(P3_STATE_REG_SCAN_IN), .B1(n8804), .B2(
        n13799), .ZN(n11965) );
  OAI21_X1 U14511 ( .B1(n11966), .B2(n13808), .A(n11965), .ZN(n11967) );
  INV_X1 U14512 ( .A(n11967), .ZN(P3_U3273) );
  OR2_X1 U14513 ( .A1(n11968), .A2(n10331), .ZN(n11970) );
  AND2_X1 U14514 ( .A1(n11970), .A2(n11969), .ZN(n15646) );
  INV_X1 U14515 ( .A(n14326), .ZN(n15625) );
  INV_X1 U14516 ( .A(n11971), .ZN(n11974) );
  INV_X1 U14517 ( .A(n11972), .ZN(n11973) );
  OAI211_X1 U14518 ( .C1(n15649), .C2(n11974), .A(n11973), .B(n14310), .ZN(
        n15647) );
  NOR2_X1 U14519 ( .A1(n15627), .A2(n15647), .ZN(n11978) );
  OAI22_X1 U14520 ( .A1(n15622), .A2(n11976), .B1(n11975), .B2(n15619), .ZN(
        n11977) );
  AOI211_X1 U14521 ( .C1(n15625), .C2(n11979), .A(n11978), .B(n11977), .ZN(
        n11988) );
  OAI21_X1 U14522 ( .B1(n10332), .B2(n11980), .A(n11981), .ZN(n11984) );
  AOI21_X1 U14523 ( .B1(n11984), .B2(n14339), .A(n11983), .ZN(n11985) );
  OAI21_X1 U14524 ( .B1(n15646), .B2(n11986), .A(n11985), .ZN(n15650) );
  NAND2_X1 U14525 ( .A1(n15650), .A2(n15622), .ZN(n11987) );
  OAI211_X1 U14526 ( .C1(n15646), .C2(n12069), .A(n11988), .B(n11987), .ZN(
        P2_U3263) );
  NAND2_X1 U14527 ( .A1(n12168), .A2(n15703), .ZN(n15710) );
  OAI22_X1 U14528 ( .A1(n15710), .A2(n11989), .B1(n13645), .B2(n12171), .ZN(
        n12000) );
  AOI21_X1 U14529 ( .B1(n11994), .B2(n11991), .A(n11990), .ZN(n11998) );
  INV_X1 U14530 ( .A(n11992), .ZN(n11993) );
  NAND2_X1 U14531 ( .A1(n11994), .A2(n11993), .ZN(n12084) );
  NAND2_X1 U14532 ( .A1(n12084), .A2(n13728), .ZN(n11997) );
  NAND2_X1 U14533 ( .A1(n15709), .A2(n13718), .ZN(n11996) );
  AOI22_X1 U14534 ( .A1(n13724), .A2(n13384), .B1(n13722), .B2(n13382), .ZN(
        n11995) );
  OAI211_X1 U14535 ( .C1(n11998), .C2(n11997), .A(n11996), .B(n11995), .ZN(
        n15713) );
  MUX2_X1 U14536 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n15713), .S(n9345), .Z(
        n11999) );
  AOI211_X1 U14537 ( .C1(n15709), .C2(n15687), .A(n12000), .B(n11999), .ZN(
        n12001) );
  INV_X1 U14538 ( .A(n12001), .ZN(P3_U3227) );
  OAI21_X1 U14539 ( .B1(n12004), .B2(n12003), .A(n12002), .ZN(n12005) );
  NAND2_X1 U14540 ( .A1(n12005), .A2(n13915), .ZN(n12012) );
  INV_X1 U14541 ( .A(n12384), .ZN(n12010) );
  NAND2_X1 U14542 ( .A1(n13971), .A2(n14286), .ZN(n12007) );
  NAND2_X1 U14543 ( .A1(n13974), .A2(n14285), .ZN(n12006) );
  AND2_X1 U14544 ( .A1(n12007), .A2(n12006), .ZN(n12379) );
  OAI21_X1 U14545 ( .B1(n13891), .B2(n12379), .A(n12008), .ZN(n12009) );
  AOI21_X1 U14546 ( .B1(n12010), .B2(n13938), .A(n12009), .ZN(n12011) );
  OAI211_X1 U14547 ( .C1(n12442), .C2(n13925), .A(n12012), .B(n12011), .ZN(
        P2_U3193) );
  AND2_X1 U14548 ( .A1(n12087), .A2(n13094), .ZN(n12172) );
  INV_X1 U14549 ( .A(n13015), .ZN(n13097) );
  XNOR2_X1 U14550 ( .A(n12172), .B(n13097), .ZN(n12120) );
  INV_X1 U14551 ( .A(n12120), .ZN(n12018) );
  INV_X1 U14552 ( .A(n13718), .ZN(n12179) );
  INV_X1 U14553 ( .A(n12013), .ZN(n12014) );
  OR2_X1 U14554 ( .A1(n12013), .A2(n13097), .ZN(n12074) );
  OAI21_X1 U14555 ( .B1(n12014), .B2(n13015), .A(n12074), .ZN(n12016) );
  INV_X1 U14556 ( .A(n13382), .ZN(n12346) );
  OAI22_X1 U14557 ( .A1(n12702), .A2(n13643), .B1(n13641), .B2(n12346), .ZN(
        n12015) );
  AOI21_X1 U14558 ( .B1(n12016), .B2(n13728), .A(n12015), .ZN(n12017) );
  OAI21_X1 U14559 ( .B1(n12120), .B2(n12179), .A(n12017), .ZN(n12114) );
  AOI21_X1 U14560 ( .B1(n15720), .B2(n12018), .A(n12114), .ZN(n12183) );
  AOI22_X1 U14561 ( .A1(n13774), .A2(n12351), .B1(n15721), .B2(
        P3_REG0_REG_8__SCAN_IN), .ZN(n12019) );
  OAI21_X1 U14562 ( .B1(n12183), .B2(n15721), .A(n12019), .ZN(P3_U3414) );
  INV_X1 U14563 ( .A(n12020), .ZN(n12022) );
  INV_X1 U14564 ( .A(n12021), .ZN(n12148) );
  OAI211_X1 U14565 ( .C1(n7767), .C2(n12022), .A(n12148), .B(n15168), .ZN(
        n15544) );
  NOR2_X1 U14566 ( .A1(n12023), .A2(n15160), .ZN(n12030) );
  NAND3_X1 U14567 ( .A1(n12025), .A2(n15370), .A3(n12024), .ZN(n12027) );
  NAND2_X1 U14568 ( .A1(n12023), .A2(n15260), .ZN(n12026) );
  NAND2_X1 U14569 ( .A1(n12027), .A2(n12026), .ZN(n12029) );
  MUX2_X1 U14570 ( .A(n12030), .B(n12029), .S(n12028), .Z(n12033) );
  AOI22_X1 U14571 ( .A1(n15257), .A2(n14816), .B1(n14814), .B2(n15258), .ZN(
        n12031) );
  INV_X1 U14572 ( .A(n15545), .ZN(n12035) );
  MUX2_X1 U14573 ( .A(n12035), .B(n12034), .S(n15533), .Z(n12039) );
  INV_X1 U14574 ( .A(n12036), .ZN(n12037) );
  AOI22_X1 U14575 ( .A1(n15524), .A2(n15548), .B1(n12037), .B2(n15526), .ZN(
        n12038) );
  OAI211_X1 U14576 ( .C1(n15174), .C2(n15544), .A(n12039), .B(n12038), .ZN(
        P1_U3286) );
  NAND2_X1 U14577 ( .A1(n12045), .A2(n12040), .ZN(n12042) );
  OAI211_X1 U14578 ( .C1(n12043), .C2(n14646), .A(n12042), .B(n12041), .ZN(
        P2_U3304) );
  NAND2_X1 U14579 ( .A1(n12045), .A2(n12044), .ZN(n12047) );
  OAI211_X1 U14580 ( .C1(n12048), .C2(n15435), .A(n12047), .B(n12046), .ZN(
        P1_U3332) );
  OR2_X1 U14581 ( .A1(n12049), .A2(n12053), .ZN(n12050) );
  NAND2_X1 U14582 ( .A1(n12051), .A2(n12050), .ZN(n12059) );
  INV_X1 U14583 ( .A(n12059), .ZN(n12100) );
  NAND3_X1 U14584 ( .A1(n12054), .A2(n12053), .A3(n12052), .ZN(n12055) );
  INV_X1 U14585 ( .A(n14339), .ZN(n14288) );
  AOI21_X1 U14586 ( .B1(n12056), .B2(n12055), .A(n14288), .ZN(n12057) );
  AOI211_X1 U14587 ( .C1(n12060), .C2(n12059), .A(n12058), .B(n12057), .ZN(
        n12099) );
  MUX2_X1 U14588 ( .A(n12061), .B(n12099), .S(n15622), .Z(n12068) );
  INV_X1 U14589 ( .A(n12062), .ZN(n12063) );
  AOI211_X1 U14590 ( .C1(n12064), .C2(n12063), .A(n14320), .B(n12252), .ZN(
        n12097) );
  OAI22_X1 U14591 ( .A1(n14326), .A2(n12104), .B1(n15619), .B2(n12065), .ZN(
        n12066) );
  AOI21_X1 U14592 ( .B1(n12097), .B2(n14344), .A(n12066), .ZN(n12067) );
  OAI211_X1 U14593 ( .C1(n12100), .C2(n12069), .A(n12068), .B(n12067), .ZN(
        P2_U3259) );
  NAND2_X1 U14594 ( .A1(n12070), .A2(n12076), .ZN(n12071) );
  AND2_X1 U14595 ( .A1(n12202), .A2(n12071), .ZN(n12451) );
  INV_X1 U14596 ( .A(n12451), .ZN(n12287) );
  INV_X1 U14597 ( .A(n13110), .ZN(n12072) );
  AOI22_X1 U14598 ( .A1(n13774), .A2(n12072), .B1(P3_REG0_REG_10__SCAN_IN), 
        .B2(n15721), .ZN(n12082) );
  NAND2_X1 U14599 ( .A1(n12074), .A2(n12073), .ZN(n12174) );
  INV_X1 U14600 ( .A(n13013), .ZN(n13102) );
  OR2_X1 U14601 ( .A1(n12174), .A2(n13102), .ZN(n12175) );
  NAND2_X1 U14602 ( .A1(n12175), .A2(n12075), .ZN(n12077) );
  XNOR2_X1 U14603 ( .A(n12077), .B(n8479), .ZN(n12078) );
  NAND2_X1 U14604 ( .A1(n12078), .A2(n13728), .ZN(n12080) );
  AOI22_X1 U14605 ( .A1(n13722), .A2(n13378), .B1(n13724), .B2(n13380), .ZN(
        n12079) );
  NAND2_X1 U14606 ( .A1(n12080), .A2(n12079), .ZN(n12448) );
  INV_X2 U14607 ( .A(n15721), .ZN(n15722) );
  NAND2_X1 U14608 ( .A1(n12448), .A2(n15722), .ZN(n12081) );
  OAI211_X1 U14609 ( .C1(n12287), .C2(n13793), .A(n12082), .B(n12081), .ZN(
        P3_U3420) );
  INV_X1 U14610 ( .A(n12363), .ZN(n12092) );
  NAND2_X1 U14611 ( .A1(n12084), .A2(n12083), .ZN(n12086) );
  XNOR2_X1 U14612 ( .A(n12086), .B(n12085), .ZN(n12091) );
  OAI21_X1 U14613 ( .B1(n12088), .B2(n13092), .A(n12087), .ZN(n15719) );
  OAI22_X1 U14614 ( .A1(n12537), .A2(n13643), .B1(n13641), .B2(n12357), .ZN(
        n12089) );
  AOI21_X1 U14615 ( .B1(n15719), .B2(n13718), .A(n12089), .ZN(n12090) );
  OAI21_X1 U14616 ( .B1(n13638), .B2(n12091), .A(n12090), .ZN(n15717) );
  AOI21_X1 U14617 ( .B1(n15685), .B2(n12092), .A(n15717), .ZN(n12093) );
  MUX2_X1 U14618 ( .A(n12094), .B(n12093), .S(n9345), .Z(n12096) );
  AOI22_X1 U14619 ( .A1(n15719), .A2(n15687), .B1(n12360), .B2(n13659), .ZN(
        n12095) );
  NAND2_X1 U14620 ( .A1(n12096), .A2(n12095), .ZN(P3_U3226) );
  INV_X1 U14621 ( .A(n12097), .ZN(n12098) );
  OAI211_X1 U14622 ( .C1(n12100), .C2(n15660), .A(n12099), .B(n12098), .ZN(
        n12106) );
  OAI22_X1 U14623 ( .A1(n14582), .A2(n12104), .B1(n15670), .B2(n11075), .ZN(
        n12101) );
  AOI21_X1 U14624 ( .B1(n12106), .B2(n15670), .A(n12101), .ZN(n12102) );
  INV_X1 U14625 ( .A(n12102), .ZN(P2_U3505) );
  INV_X1 U14626 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n12103) );
  OAI22_X1 U14627 ( .A1(n14627), .A2(n12104), .B1(n15666), .B2(n12103), .ZN(
        n12105) );
  AOI21_X1 U14628 ( .B1(n12106), .B2(n15666), .A(n12105), .ZN(n12107) );
  INV_X1 U14629 ( .A(n12107), .ZN(P2_U3448) );
  INV_X1 U14630 ( .A(n12108), .ZN(n12112) );
  OAI222_X1 U14631 ( .A1(n15435), .A2(n12110), .B1(n15433), .B2(n12112), .C1(
        P1_U3086), .C2(n12109), .ZN(P1_U3331) );
  OAI222_X1 U14632 ( .A1(n12113), .A2(P2_U3088), .B1(n14637), .B2(n12112), 
        .C1(n12111), .C2(n14646), .ZN(P2_U3303) );
  INV_X1 U14633 ( .A(n12114), .ZN(n12115) );
  MUX2_X1 U14634 ( .A(n12116), .B(n12115), .S(n9345), .Z(n12119) );
  INV_X1 U14635 ( .A(n12349), .ZN(n12117) );
  AOI22_X1 U14636 ( .A1(n13659), .A2(n12351), .B1(n15685), .B2(n12117), .ZN(
        n12118) );
  OAI211_X1 U14637 ( .C1(n12120), .C2(n12230), .A(n12119), .B(n12118), .ZN(
        P3_U3225) );
  INV_X1 U14638 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15358) );
  XNOR2_X1 U14639 ( .A(n14939), .B(n15358), .ZN(n12133) );
  INV_X1 U14640 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15445) );
  NAND2_X1 U14641 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14787)
         );
  OAI21_X1 U14642 ( .B1(n15497), .B2(n15445), .A(n14787), .ZN(n12123) );
  AOI21_X1 U14643 ( .B1(n14940), .B2(n15500), .A(n12123), .ZN(n12132) );
  NAND2_X1 U14644 ( .A1(n12124), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n12125) );
  NAND2_X1 U14645 ( .A1(n12126), .A2(n12125), .ZN(n14933) );
  XNOR2_X1 U14646 ( .A(n14933), .B(n12127), .ZN(n12129) );
  INV_X1 U14647 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n12128) );
  NAND2_X1 U14648 ( .A1(n12129), .A2(n12128), .ZN(n14936) );
  OAI21_X1 U14649 ( .B1(n12129), .B2(n12128), .A(n14936), .ZN(n12130) );
  NAND2_X1 U14650 ( .A1(n12130), .A2(n15513), .ZN(n12131) );
  OAI211_X1 U14651 ( .C1(n12133), .C2(n14942), .A(n12132), .B(n12131), .ZN(
        P1_U3258) );
  INV_X1 U14652 ( .A(n12409), .ZN(n12596) );
  OAI21_X1 U14653 ( .B1(n12136), .B2(n12135), .A(n12134), .ZN(n12137) );
  NAND2_X1 U14654 ( .A1(n12137), .A2(n13915), .ZN(n12144) );
  INV_X1 U14655 ( .A(n12595), .ZN(n12142) );
  NAND2_X1 U14656 ( .A1(n14329), .A2(n14286), .ZN(n12139) );
  NAND2_X1 U14657 ( .A1(n13973), .A2(n14285), .ZN(n12138) );
  AND2_X1 U14658 ( .A1(n12139), .A2(n12138), .ZN(n12405) );
  OAI21_X1 U14659 ( .B1(n13891), .B2(n12405), .A(n12140), .ZN(n12141) );
  AOI21_X1 U14660 ( .B1(n12142), .B2(n13938), .A(n12141), .ZN(n12143) );
  OAI211_X1 U14661 ( .C1(n12596), .C2(n13925), .A(n12144), .B(n12143), .ZN(
        P2_U3203) );
  OAI21_X1 U14662 ( .B1(n12146), .B2(n12152), .A(n12145), .ZN(n12299) );
  AOI211_X1 U14663 ( .C1(n12220), .C2(n12148), .A(n15270), .B(n7051), .ZN(
        n12306) );
  INV_X1 U14664 ( .A(n12149), .ZN(n12150) );
  AOI211_X1 U14665 ( .C1(n12152), .C2(n12151), .A(n15160), .B(n12150), .ZN(
        n12155) );
  OAI22_X1 U14666 ( .A1(n12154), .A2(n15239), .B1(n12153), .B2(n15241), .ZN(
        n12216) );
  OR2_X1 U14667 ( .A1(n12155), .A2(n12216), .ZN(n12300) );
  AOI211_X1 U14668 ( .C1(n15370), .C2(n12299), .A(n12306), .B(n12300), .ZN(
        n12158) );
  AOI22_X1 U14669 ( .A1(n12686), .A2(n12220), .B1(P1_REG1_REG_8__SCAN_IN), 
        .B2(n15552), .ZN(n12156) );
  OAI21_X1 U14670 ( .B1(n12158), .B2(n15552), .A(n12156), .ZN(P1_U3536) );
  AOI22_X1 U14671 ( .A1(n12478), .A2(n12220), .B1(P1_REG0_REG_8__SCAN_IN), 
        .B2(n15549), .ZN(n12157) );
  OAI21_X1 U14672 ( .B1(n12158), .B2(n15549), .A(n12157), .ZN(P1_U3483) );
  INV_X1 U14673 ( .A(n13362), .ZN(n12704) );
  INV_X1 U14674 ( .A(n12159), .ZN(n12160) );
  XNOR2_X1 U14675 ( .A(n12932), .B(n12168), .ZN(n12341) );
  XNOR2_X1 U14676 ( .A(n12341), .B(n13383), .ZN(n12163) );
  INV_X1 U14677 ( .A(n12342), .ZN(n12162) );
  OAI211_X1 U14678 ( .C1(n12164), .C2(n12163), .A(n12162), .B(n13353), .ZN(
        n12170) );
  OAI22_X1 U14679 ( .A1(n13331), .A2(n12346), .B1(n12165), .B2(n13359), .ZN(
        n12166) );
  AOI211_X1 U14680 ( .C1(n13349), .C2(n12168), .A(n12167), .B(n12166), .ZN(
        n12169) );
  OAI211_X1 U14681 ( .C1(n12171), .C2(n12704), .A(n12170), .B(n12169), .ZN(
        P3_U3179) );
  OAI21_X1 U14682 ( .B1(n12172), .B2(n13015), .A(n13100), .ZN(n12173) );
  XNOR2_X1 U14683 ( .A(n12173), .B(n13013), .ZN(n12231) );
  INV_X1 U14684 ( .A(n12231), .ZN(n12180) );
  AOI22_X1 U14685 ( .A1(n13724), .A2(n13381), .B1(n13722), .B2(n13379), .ZN(
        n12178) );
  INV_X1 U14686 ( .A(n12174), .ZN(n12176) );
  OAI211_X1 U14687 ( .C1(n12176), .C2(n13013), .A(n13728), .B(n12175), .ZN(
        n12177) );
  OAI211_X1 U14688 ( .C1(n12231), .C2(n12179), .A(n12178), .B(n12177), .ZN(
        n12223) );
  AOI21_X1 U14689 ( .B1(n15720), .B2(n12180), .A(n12223), .ZN(n12296) );
  INV_X1 U14690 ( .A(n12534), .ZN(n12227) );
  AOI22_X1 U14691 ( .A1(n13774), .A2(n12227), .B1(P3_REG0_REG_9__SCAN_IN), 
        .B2(n15721), .ZN(n12181) );
  OAI21_X1 U14692 ( .B1(n12296), .B2(n15721), .A(n12181), .ZN(P3_U3417) );
  INV_X1 U14693 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n14471) );
  NAND2_X1 U14694 ( .A1(n13541), .A2(P3_U3897), .ZN(n12182) );
  OAI21_X1 U14695 ( .B1(P3_U3897), .B2(n14471), .A(n12182), .ZN(P3_U3516) );
  INV_X1 U14696 ( .A(n12351), .ZN(n12186) );
  MUX2_X1 U14697 ( .A(n12184), .B(n12183), .S(n15734), .Z(n12185) );
  OAI21_X1 U14698 ( .B1(n12186), .B2(n13709), .A(n12185), .ZN(P3_U3467) );
  OAI21_X1 U14699 ( .B1(n12189), .B2(n12188), .A(n12187), .ZN(n12195) );
  OAI22_X1 U14700 ( .A1(n12522), .A2(n15239), .B1(n12590), .B2(n15241), .ZN(
        n12194) );
  NAND2_X1 U14701 ( .A1(n12190), .A2(n12189), .ZN(n12191) );
  AOI21_X1 U14702 ( .B1(n12192), .B2(n12191), .A(n15160), .ZN(n12193) );
  AOI211_X1 U14703 ( .C1(n15370), .C2(n12195), .A(n12194), .B(n12193), .ZN(
        n12310) );
  AOI21_X1 U14704 ( .B1(n12196), .B2(n12516), .A(n15270), .ZN(n12197) );
  NAND2_X1 U14705 ( .A1(n12197), .A2(n12334), .ZN(n12315) );
  AND2_X1 U14706 ( .A1(n12310), .A2(n12315), .ZN(n12200) );
  AOI22_X1 U14707 ( .A1(n12478), .A2(n12516), .B1(P1_REG0_REG_9__SCAN_IN), 
        .B2(n15549), .ZN(n12198) );
  OAI21_X1 U14708 ( .B1(n12200), .B2(n15549), .A(n12198), .ZN(P1_U3486) );
  AOI22_X1 U14709 ( .A1(n12686), .A2(n12516), .B1(P1_REG1_REG_9__SCAN_IN), 
        .B2(n15552), .ZN(n12199) );
  OAI21_X1 U14710 ( .B1(n12200), .B2(n15552), .A(n12199), .ZN(P1_U3537) );
  NAND2_X1 U14711 ( .A1(n12202), .A2(n12201), .ZN(n12274) );
  INV_X1 U14712 ( .A(n13051), .ZN(n12203) );
  NOR2_X1 U14713 ( .A1(n13049), .A2(n12203), .ZN(n13114) );
  INV_X1 U14714 ( .A(n13114), .ZN(n12275) );
  NOR2_X1 U14715 ( .A1(n12274), .A2(n12275), .ZN(n12273) );
  NOR2_X1 U14716 ( .A1(n12273), .A2(n13049), .ZN(n12204) );
  XNOR2_X1 U14717 ( .A(n12204), .B(n13018), .ZN(n12367) );
  AOI22_X1 U14718 ( .A1(n13774), .A2(n13278), .B1(P3_REG0_REG_12__SCAN_IN), 
        .B2(n15721), .ZN(n12211) );
  NAND2_X1 U14719 ( .A1(n12205), .A2(n13018), .ZN(n12206) );
  NAND3_X1 U14720 ( .A1(n12207), .A2(n13728), .A3(n12206), .ZN(n12209) );
  AOI22_X1 U14721 ( .A1(n13724), .A2(n13378), .B1(n13722), .B2(n13376), .ZN(
        n12208) );
  NAND2_X1 U14722 ( .A1(n12209), .A2(n12208), .ZN(n12364) );
  NAND2_X1 U14723 ( .A1(n12364), .A2(n15722), .ZN(n12210) );
  OAI211_X1 U14724 ( .C1(n12367), .C2(n13793), .A(n12211), .B(n12210), .ZN(
        P3_U3426) );
  INV_X1 U14725 ( .A(n12212), .ZN(n12213) );
  AOI21_X1 U14726 ( .B1(n12215), .B2(n12214), .A(n12213), .ZN(n12222) );
  NAND2_X1 U14727 ( .A1(n14766), .A2(n12216), .ZN(n12217) );
  OAI211_X1 U14728 ( .C1(n14792), .C2(n12303), .A(n12218), .B(n12217), .ZN(
        n12219) );
  AOI21_X1 U14729 ( .B1(n14795), .B2(n12220), .A(n12219), .ZN(n12221) );
  OAI21_X1 U14730 ( .B1(n12222), .B2(n14797), .A(n12221), .ZN(P1_U3221) );
  INV_X1 U14731 ( .A(n12223), .ZN(n12224) );
  MUX2_X1 U14732 ( .A(n12225), .B(n12224), .S(n9345), .Z(n12229) );
  INV_X1 U14733 ( .A(n12226), .ZN(n12540) );
  AOI22_X1 U14734 ( .A1(n13659), .A2(n12227), .B1(n15685), .B2(n12540), .ZN(
        n12228) );
  OAI211_X1 U14735 ( .C1(n12231), .C2(n12230), .A(n12229), .B(n12228), .ZN(
        P3_U3224) );
  XNOR2_X1 U14736 ( .A(n12483), .B(n12482), .ZN(n12240) );
  INV_X1 U14737 ( .A(n12736), .ZN(n12237) );
  NAND2_X1 U14738 ( .A1(n13971), .A2(n14285), .ZN(n12233) );
  NAND2_X1 U14739 ( .A1(n13970), .A2(n14286), .ZN(n12232) );
  NAND2_X1 U14740 ( .A1(n12233), .A2(n12232), .ZN(n12729) );
  INV_X1 U14741 ( .A(n12729), .ZN(n12235) );
  OAI21_X1 U14742 ( .B1(n13891), .B2(n12235), .A(n12234), .ZN(n12236) );
  AOI21_X1 U14743 ( .B1(n12237), .B2(n13938), .A(n12236), .ZN(n12239) );
  NAND2_X1 U14744 ( .A1(n12735), .A2(n13954), .ZN(n12238) );
  OAI211_X1 U14745 ( .C1(n12240), .C2(n13956), .A(n12239), .B(n12238), .ZN(
        P2_U3189) );
  INV_X1 U14746 ( .A(n12241), .ZN(n12245) );
  OAI222_X1 U14747 ( .A1(n12243), .A2(P1_U3086), .B1(n15433), .B2(n12245), 
        .C1(n12242), .C2(n15435), .ZN(P1_U3330) );
  OAI222_X1 U14748 ( .A1(n12246), .A2(P2_U3088), .B1(n14637), .B2(n12245), 
        .C1(n12244), .C2(n14646), .ZN(P2_U3302) );
  OAI21_X1 U14749 ( .B1(n12247), .B2(n12248), .A(n12369), .ZN(n15631) );
  INV_X1 U14750 ( .A(n15631), .ZN(n12253) );
  INV_X1 U14751 ( .A(n12373), .ZN(n12376) );
  XNOR2_X1 U14752 ( .A(n12376), .B(n12248), .ZN(n12250) );
  AOI21_X1 U14753 ( .B1(n12250), .B2(n14339), .A(n12249), .ZN(n15633) );
  OAI211_X1 U14754 ( .C1(n12252), .C2(n12375), .A(n14310), .B(n12251), .ZN(
        n15628) );
  OAI211_X1 U14755 ( .C1(n14575), .C2(n12253), .A(n15633), .B(n15628), .ZN(
        n12259) );
  OAI22_X1 U14756 ( .A1(n14582), .A2(n12375), .B1(n15670), .B2(n12254), .ZN(
        n12255) );
  AOI21_X1 U14757 ( .B1(n12259), .B2(n15670), .A(n12255), .ZN(n12256) );
  INV_X1 U14758 ( .A(n12256), .ZN(P2_U3506) );
  INV_X1 U14759 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n12257) );
  OAI22_X1 U14760 ( .A1(n14627), .A2(n12375), .B1(n15666), .B2(n12257), .ZN(
        n12258) );
  AOI21_X1 U14761 ( .B1(n12259), .B2(n15666), .A(n12258), .ZN(n12260) );
  INV_X1 U14762 ( .A(n12260), .ZN(P2_U3451) );
  MUX2_X1 U14763 ( .A(n12262), .B(n12261), .S(n15622), .Z(n12269) );
  NOR2_X1 U14764 ( .A1(n15627), .A2(n12263), .ZN(n12266) );
  OAI22_X1 U14765 ( .A1(n14326), .A2(n12264), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n15619), .ZN(n12265) );
  AOI211_X1 U14766 ( .C1(n15630), .C2(n12267), .A(n12266), .B(n12265), .ZN(
        n12268) );
  NAND2_X1 U14767 ( .A1(n12269), .A2(n12268), .ZN(P2_U3262) );
  NAND2_X1 U14768 ( .A1(n12270), .A2(n13801), .ZN(n12271) );
  OAI211_X1 U14769 ( .C1(n12272), .C2(n13805), .A(n12271), .B(n13193), .ZN(
        P3_U3272) );
  AOI21_X1 U14770 ( .B1(n12275), .B2(n12274), .A(n12273), .ZN(n12290) );
  AOI22_X1 U14771 ( .A1(n13659), .A2(n12280), .B1(n15685), .B2(n12860), .ZN(
        n12279) );
  XNOR2_X1 U14772 ( .A(n12276), .B(n13114), .ZN(n12277) );
  AOI222_X1 U14773 ( .A1(n13379), .A2(n13724), .B1(n13728), .B2(n12277), .C1(
        n13377), .C2(n13722), .ZN(n12295) );
  MUX2_X1 U14774 ( .A(n12662), .B(n12295), .S(n9345), .Z(n12278) );
  OAI211_X1 U14775 ( .C1(n12290), .C2(n13663), .A(n12279), .B(n12278), .ZN(
        P3_U3222) );
  MUX2_X1 U14776 ( .A(n12656), .B(n12295), .S(n15734), .Z(n12282) );
  INV_X1 U14777 ( .A(n13709), .ZN(n13698) );
  NAND2_X1 U14778 ( .A1(n13698), .A2(n12280), .ZN(n12281) );
  OAI211_X1 U14779 ( .C1(n12290), .C2(n13715), .A(n12282), .B(n12281), .ZN(
        P3_U3470) );
  AOI22_X1 U14780 ( .A1(n13278), .A2(n13659), .B1(n15685), .B2(n13277), .ZN(
        n12286) );
  INV_X1 U14781 ( .A(n12364), .ZN(n12283) );
  MUX2_X1 U14782 ( .A(n12284), .B(n12283), .S(n9345), .Z(n12285) );
  OAI211_X1 U14783 ( .C1(n12367), .C2(n13663), .A(n12286), .B(n12285), .ZN(
        P3_U3221) );
  MUX2_X1 U14784 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n12448), .S(n15734), .Z(
        n12289) );
  OAI22_X1 U14785 ( .A1(n12287), .A2(n13715), .B1(n13110), .B2(n13709), .ZN(
        n12288) );
  OR2_X1 U14786 ( .A1(n12289), .A2(n12288), .ZN(P3_U3469) );
  INV_X1 U14787 ( .A(n12290), .ZN(n12293) );
  INV_X1 U14788 ( .A(n13793), .ZN(n13785) );
  OAI22_X1 U14789 ( .A1(n12855), .A2(n13790), .B1(n15722), .B2(n12291), .ZN(
        n12292) );
  AOI21_X1 U14790 ( .B1(n12293), .B2(n13785), .A(n12292), .ZN(n12294) );
  OAI21_X1 U14791 ( .B1(n15721), .B2(n12295), .A(n12294), .ZN(P3_U3423) );
  MUX2_X1 U14792 ( .A(n12297), .B(n12296), .S(n15734), .Z(n12298) );
  OAI21_X1 U14793 ( .B1(n13709), .B2(n12534), .A(n12298), .ZN(P3_U3468) );
  INV_X1 U14794 ( .A(n12299), .ZN(n12309) );
  INV_X1 U14795 ( .A(n12300), .ZN(n12301) );
  MUX2_X1 U14796 ( .A(n12302), .B(n12301), .S(n15220), .Z(n12308) );
  OAI22_X1 U14797 ( .A1(n15234), .A2(n12304), .B1(n15217), .B2(n12303), .ZN(
        n12305) );
  AOI21_X1 U14798 ( .B1(n12306), .B2(n15522), .A(n12305), .ZN(n12307) );
  OAI211_X1 U14799 ( .C1(n12309), .C2(n15248), .A(n12308), .B(n12307), .ZN(
        P1_U3285) );
  MUX2_X1 U14800 ( .A(n12311), .B(n12310), .S(n15220), .Z(n12314) );
  INV_X1 U14801 ( .A(n12521), .ZN(n12312) );
  AOI22_X1 U14802 ( .A1(n15524), .A2(n12516), .B1(n15526), .B2(n12312), .ZN(
        n12313) );
  OAI211_X1 U14803 ( .C1(n15174), .C2(n12315), .A(n12314), .B(n12313), .ZN(
        P1_U3284) );
  INV_X1 U14804 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n12317) );
  NAND2_X1 U14805 ( .A1(n12318), .A2(n12317), .ZN(n12319) );
  NAND2_X1 U14806 ( .A1(n12320), .A2(n12319), .ZN(n12498) );
  NAND2_X1 U14807 ( .A1(n12322), .A2(n12321), .ZN(n12324) );
  NAND2_X1 U14808 ( .A1(n12324), .A2(n12323), .ZN(n12501) );
  INV_X1 U14809 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n12325) );
  NAND2_X1 U14810 ( .A1(n12325), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n12502) );
  INV_X1 U14811 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n12326) );
  NAND2_X1 U14812 ( .A1(n12326), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n12327) );
  AND2_X1 U14813 ( .A1(n12502), .A2(n12327), .ZN(n12500) );
  XNOR2_X1 U14814 ( .A(n12501), .B(n12500), .ZN(n12496) );
  INV_X1 U14815 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15584) );
  XNOR2_X1 U14816 ( .A(n12495), .B(n15584), .ZN(SUB_1596_U68) );
  AOI21_X1 U14817 ( .B1(n12328), .B2(n12332), .A(n15160), .ZN(n12329) );
  OR2_X1 U14818 ( .A1(n12328), .A2(n12332), .ZN(n12428) );
  AOI22_X1 U14819 ( .A1(n12329), .A2(n12428), .B1(n15257), .B2(n14813), .ZN(
        n12475) );
  MUX2_X1 U14820 ( .A(n12330), .B(n12475), .S(n15220), .Z(n12340) );
  OAI21_X1 U14821 ( .B1(n12333), .B2(n12332), .A(n12331), .ZN(n12477) );
  AOI21_X1 U14822 ( .B1(n12334), .B2(n14674), .A(n15270), .ZN(n12335) );
  AND2_X1 U14823 ( .A1(n14811), .A2(n15258), .ZN(n14671) );
  AOI21_X1 U14824 ( .B1(n12335), .B2(n12422), .A(n14671), .ZN(n12474) );
  INV_X1 U14825 ( .A(n12336), .ZN(n14675) );
  AOI22_X1 U14826 ( .A1(n15524), .A2(n14674), .B1(n15526), .B2(n14675), .ZN(
        n12337) );
  OAI21_X1 U14827 ( .B1(n12474), .B2(n15174), .A(n12337), .ZN(n12338) );
  AOI21_X1 U14828 ( .B1(n12477), .B2(n15519), .A(n12338), .ZN(n12339) );
  NAND2_X1 U14829 ( .A1(n12340), .A2(n12339), .ZN(P1_U3283) );
  INV_X1 U14830 ( .A(n12341), .ZN(n12343) );
  XNOR2_X1 U14831 ( .A(n12935), .B(n15716), .ZN(n12344) );
  XNOR2_X1 U14832 ( .A(n12344), .B(n13382), .ZN(n12355) );
  XNOR2_X1 U14833 ( .A(n12935), .B(n12351), .ZN(n12527) );
  XNOR2_X1 U14834 ( .A(n12527), .B(n13381), .ZN(n12529) );
  XNOR2_X1 U14835 ( .A(n12530), .B(n12529), .ZN(n12353) );
  OAI21_X1 U14836 ( .B1(n13359), .B2(n12346), .A(n12345), .ZN(n12347) );
  AOI21_X1 U14837 ( .B1(n13357), .B2(n13380), .A(n12347), .ZN(n12348) );
  OAI21_X1 U14838 ( .B1(n12349), .B2(n12704), .A(n12348), .ZN(n12350) );
  AOI21_X1 U14839 ( .B1(n13349), .B2(n12351), .A(n12350), .ZN(n12352) );
  OAI21_X1 U14840 ( .B1(n12353), .B2(n13351), .A(n12352), .ZN(P3_U3161) );
  XOR2_X1 U14841 ( .A(n12355), .B(n12354), .Z(n12356) );
  NAND2_X1 U14842 ( .A1(n12356), .A2(n13353), .ZN(n12362) );
  OAI22_X1 U14843 ( .A1(n13331), .A2(n12537), .B1(n12357), .B2(n13359), .ZN(
        n12358) );
  AOI211_X1 U14844 ( .C1(n13349), .C2(n12360), .A(n12359), .B(n12358), .ZN(
        n12361) );
  OAI211_X1 U14845 ( .C1(n12363), .C2(n12704), .A(n12362), .B(n12361), .ZN(
        P3_U3153) );
  MUX2_X1 U14846 ( .A(n12364), .B(P3_REG1_REG_12__SCAN_IN), .S(n15731), .Z(
        n12365) );
  AOI21_X1 U14847 ( .B1(n13698), .B2(n13278), .A(n12365), .ZN(n12366) );
  OAI21_X1 U14848 ( .B1(n12367), .B2(n13715), .A(n12366), .ZN(P3_U3471) );
  NAND2_X1 U14849 ( .A1(n12369), .A2(n12368), .ZN(n12370) );
  NOR2_X1 U14850 ( .A1(n12370), .A2(n12371), .ZN(n12399) );
  AOI21_X1 U14851 ( .B1(n12371), .B2(n12370), .A(n12399), .ZN(n12440) );
  INV_X1 U14852 ( .A(n12440), .ZN(n12388) );
  OAI21_X1 U14853 ( .B1(n12373), .B2(n15624), .A(n12372), .ZN(n12374) );
  OAI21_X1 U14854 ( .B1(n12376), .B2(n12375), .A(n12374), .ZN(n12378) );
  XNOR2_X1 U14855 ( .A(n12378), .B(n12377), .ZN(n12380) );
  OAI21_X1 U14856 ( .B1(n12380), .B2(n14288), .A(n12379), .ZN(n12438) );
  INV_X1 U14857 ( .A(n12438), .ZN(n12381) );
  MUX2_X1 U14858 ( .A(n12382), .B(n12381), .S(n15622), .Z(n12387) );
  AOI21_X1 U14859 ( .B1(n12251), .B2(n12445), .A(n14320), .ZN(n12383) );
  AND2_X1 U14860 ( .A1(n12383), .A2(n12401), .ZN(n12439) );
  OAI22_X1 U14861 ( .A1(n14326), .A2(n12442), .B1(n15619), .B2(n12384), .ZN(
        n12385) );
  AOI21_X1 U14862 ( .B1(n12439), .B2(n14344), .A(n12385), .ZN(n12386) );
  OAI211_X1 U14863 ( .C1(n14346), .C2(n12388), .A(n12387), .B(n12386), .ZN(
        P2_U3257) );
  XOR2_X1 U14864 ( .A(n13126), .B(n12389), .Z(n12414) );
  INV_X1 U14865 ( .A(n12793), .ZN(n12390) );
  OAI22_X1 U14866 ( .A1(n12790), .A2(n13588), .B1(n12390), .B2(n13645), .ZN(
        n12391) );
  AOI21_X1 U14867 ( .B1(n12414), .B2(n13563), .A(n12391), .ZN(n12397) );
  OAI211_X1 U14868 ( .C1(n12393), .C2(n13126), .A(n12392), .B(n13728), .ZN(
        n12395) );
  AOI22_X1 U14869 ( .A1(n13724), .A2(n13377), .B1(n13722), .B2(n13375), .ZN(
        n12394) );
  AND2_X1 U14870 ( .A1(n12395), .A2(n12394), .ZN(n12416) );
  MUX2_X1 U14871 ( .A(n12416), .B(n13431), .S(n15691), .Z(n12396) );
  NAND2_X1 U14872 ( .A1(n12397), .A2(n12396), .ZN(P3_U3220) );
  NOR2_X1 U14873 ( .A1(n12399), .A2(n12398), .ZN(n12400) );
  XNOR2_X1 U14874 ( .A(n12400), .B(n12402), .ZN(n12602) );
  INV_X1 U14875 ( .A(n12602), .ZN(n12407) );
  AOI211_X1 U14876 ( .C1(n12409), .C2(n12401), .A(n14320), .B(n12732), .ZN(
        n12600) );
  OAI21_X1 U14877 ( .B1(n12403), .B2(n12402), .A(n14339), .ZN(n12404) );
  OR2_X1 U14878 ( .A1(n14330), .A2(n12404), .ZN(n12406) );
  NAND2_X1 U14879 ( .A1(n12406), .A2(n12405), .ZN(n12597) );
  AOI211_X1 U14880 ( .C1(n12407), .C2(n14579), .A(n12600), .B(n12597), .ZN(
        n12411) );
  AOI22_X1 U14881 ( .A1(n8939), .A2(n12409), .B1(P2_REG1_REG_9__SCAN_IN), .B2(
        n15668), .ZN(n12408) );
  OAI21_X1 U14882 ( .B1(n12411), .B2(n15668), .A(n12408), .ZN(P2_U3508) );
  AOI22_X1 U14883 ( .A1(n10703), .A2(n12409), .B1(P2_REG0_REG_9__SCAN_IN), 
        .B2(n15664), .ZN(n12410) );
  OAI21_X1 U14884 ( .B1(n12411), .B2(n15664), .A(n12410), .ZN(P2_U3457) );
  INV_X1 U14885 ( .A(n13715), .ZN(n13706) );
  NAND2_X1 U14886 ( .A1(n12414), .A2(n13706), .ZN(n12413) );
  MUX2_X1 U14887 ( .A(n12416), .B(n13424), .S(n15731), .Z(n12412) );
  OAI211_X1 U14888 ( .C1(n13709), .C2(n12790), .A(n12413), .B(n12412), .ZN(
        P3_U3472) );
  NAND2_X1 U14889 ( .A1(n12414), .A2(n13785), .ZN(n12418) );
  INV_X1 U14890 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12415) );
  MUX2_X1 U14891 ( .A(n12416), .B(n12415), .S(n15721), .Z(n12417) );
  OAI211_X1 U14892 ( .C1(n13790), .C2(n12790), .A(n12418), .B(n12417), .ZN(
        P3_U3429) );
  OAI21_X1 U14893 ( .B1(n12421), .B2(n12420), .A(n12419), .ZN(n12689) );
  INV_X1 U14894 ( .A(n12689), .ZN(n12436) );
  AOI211_X1 U14895 ( .C1(n12423), .C2(n12422), .A(n15270), .B(n12565), .ZN(
        n12688) );
  INV_X1 U14896 ( .A(n12423), .ZN(n12694) );
  NOR2_X1 U14897 ( .A1(n12694), .A2(n15234), .ZN(n12426) );
  OAI22_X1 U14898 ( .A1(n15220), .A2(n12424), .B1(n12589), .B2(n15217), .ZN(
        n12425) );
  AOI211_X1 U14899 ( .C1(n12688), .C2(n15522), .A(n12426), .B(n12425), .ZN(
        n12435) );
  NAND2_X1 U14900 ( .A1(n12428), .A2(n12427), .ZN(n12431) );
  OAI211_X1 U14901 ( .C1(n12431), .C2(n12430), .A(n12429), .B(n15260), .ZN(
        n12433) );
  AOI22_X1 U14902 ( .A1(n15257), .A2(n14812), .B1(n14810), .B2(n15258), .ZN(
        n12432) );
  NAND2_X1 U14903 ( .A1(n12433), .A2(n12432), .ZN(n12687) );
  NAND2_X1 U14904 ( .A1(n12687), .A2(n15220), .ZN(n12434) );
  OAI211_X1 U14905 ( .C1(n12436), .C2(n15248), .A(n12435), .B(n12434), .ZN(
        P1_U3282) );
  INV_X1 U14906 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n14459) );
  NAND2_X1 U14907 ( .A1(n13542), .A2(P3_U3897), .ZN(n12437) );
  OAI21_X1 U14908 ( .B1(P3_U3897), .B2(n14459), .A(n12437), .ZN(P3_U3518) );
  AOI211_X1 U14909 ( .C1(n12440), .C2(n14579), .A(n12439), .B(n12438), .ZN(
        n12447) );
  OAI22_X1 U14910 ( .A1(n14582), .A2(n12442), .B1(n15670), .B2(n12441), .ZN(
        n12443) );
  INV_X1 U14911 ( .A(n12443), .ZN(n12444) );
  OAI21_X1 U14912 ( .B1(n12447), .B2(n15668), .A(n12444), .ZN(P2_U3507) );
  AOI22_X1 U14913 ( .A1(n10703), .A2(n12445), .B1(P2_REG0_REG_8__SCAN_IN), 
        .B2(n15664), .ZN(n12446) );
  OAI21_X1 U14914 ( .B1(n12447), .B2(n15664), .A(n12446), .ZN(P2_U3454) );
  OAI22_X1 U14915 ( .A1(n13588), .A2(n13110), .B1(n12703), .B2(n13645), .ZN(
        n12450) );
  MUX2_X1 U14916 ( .A(n12448), .B(P3_REG2_REG_10__SCAN_IN), .S(n15691), .Z(
        n12449) );
  AOI211_X1 U14917 ( .C1(n12451), .C2(n13563), .A(n12450), .B(n12449), .ZN(
        n12452) );
  INV_X1 U14918 ( .A(n12452), .ZN(P3_U3223) );
  OR2_X1 U14919 ( .A1(n12453), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n15572) );
  NAND2_X1 U14920 ( .A1(n15574), .A2(n15572), .ZN(n12454) );
  MUX2_X1 U14921 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n12605), .S(n15580), .Z(
        n15571) );
  NAND2_X1 U14922 ( .A1(n12454), .A2(n15571), .ZN(n15576) );
  NAND2_X1 U14923 ( .A1(n12455), .A2(n12605), .ZN(n12456) );
  NAND2_X1 U14924 ( .A1(n15576), .A2(n12456), .ZN(n15593) );
  MUX2_X1 U14925 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n12680), .S(n12457), .Z(
        n15592) );
  NAND2_X1 U14926 ( .A1(n15586), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n12458) );
  NAND2_X1 U14927 ( .A1(n15612), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n12461) );
  NAND2_X1 U14928 ( .A1(n12459), .A2(n12466), .ZN(n12460) );
  NAND2_X1 U14929 ( .A1(n12461), .A2(n12460), .ZN(n12641) );
  XNOR2_X1 U14930 ( .A(n12641), .B(n12469), .ZN(n12639) );
  XNOR2_X1 U14931 ( .A(n12639), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n12473) );
  INV_X1 U14932 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n12463) );
  XNOR2_X1 U14933 ( .A(n15580), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n15577) );
  XNOR2_X1 U14934 ( .A(n15586), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n15599) );
  AOI21_X1 U14935 ( .B1(n15586), .B2(P2_REG1_REG_13__SCAN_IN), .A(n15596), 
        .ZN(n15604) );
  XNOR2_X1 U14936 ( .A(n12466), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n15605) );
  INV_X1 U14937 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n12467) );
  XNOR2_X1 U14938 ( .A(n12636), .B(n14558), .ZN(n12471) );
  NAND2_X1 U14939 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n13951)
         );
  NAND2_X1 U14940 ( .A1(n15585), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n12468) );
  OAI211_X1 U14941 ( .C1(n15608), .C2(n12469), .A(n13951), .B(n12468), .ZN(
        n12470) );
  AOI21_X1 U14942 ( .B1(n12471), .B2(n15610), .A(n12470), .ZN(n12472) );
  OAI21_X1 U14943 ( .B1(n12473), .B2(n15591), .A(n12472), .ZN(P2_U3229) );
  NAND2_X1 U14944 ( .A1(n12475), .A2(n12474), .ZN(n12476) );
  AOI21_X1 U14945 ( .B1(n15370), .B2(n12477), .A(n12476), .ZN(n12481) );
  AOI22_X1 U14946 ( .A1(n14674), .A2(n12478), .B1(P1_REG0_REG_10__SCAN_IN), 
        .B2(n15549), .ZN(n12479) );
  OAI21_X1 U14947 ( .B1(n12481), .B2(n15549), .A(n12479), .ZN(P1_U3489) );
  AOI22_X1 U14948 ( .A1(n14674), .A2(n12686), .B1(P1_REG1_REG_10__SCAN_IN), 
        .B2(n15552), .ZN(n12480) );
  OAI21_X1 U14949 ( .B1(n12481), .B2(n15552), .A(n12480), .ZN(P1_U3538) );
  OR2_X1 U14950 ( .A1(n12483), .A2(n12482), .ZN(n12485) );
  NAND2_X1 U14951 ( .A1(n12485), .A2(n12484), .ZN(n12487) );
  AOI21_X1 U14952 ( .B1(n12487), .B2(n12486), .A(n7798), .ZN(n12494) );
  NAND2_X1 U14953 ( .A1(n14329), .A2(n14285), .ZN(n12489) );
  NAND2_X1 U14954 ( .A1(n13969), .A2(n14286), .ZN(n12488) );
  NAND2_X1 U14955 ( .A1(n12489), .A2(n12488), .ZN(n14338) );
  AOI21_X1 U14956 ( .B1(n13949), .B2(n14338), .A(n12490), .ZN(n12491) );
  OAI21_X1 U14957 ( .B1(n13952), .B2(n14322), .A(n12491), .ZN(n12492) );
  AOI21_X1 U14958 ( .B1(n14571), .B2(n13954), .A(n12492), .ZN(n12493) );
  OAI21_X1 U14959 ( .B1(n12494), .B2(n13956), .A(n12493), .ZN(P2_U3208) );
  INV_X1 U14960 ( .A(n12496), .ZN(n12497) );
  NAND2_X1 U14961 ( .A1(n12498), .A2(n12497), .ZN(n12499) );
  NAND2_X1 U14962 ( .A1(n12501), .A2(n12500), .ZN(n12503) );
  NAND2_X1 U14963 ( .A1(n12503), .A2(n12502), .ZN(n12832) );
  XNOR2_X1 U14964 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(P3_ADDR_REG_13__SCAN_IN), 
        .ZN(n12504) );
  XNOR2_X1 U14965 ( .A(n12832), .B(n12504), .ZN(n12825) );
  INV_X1 U14966 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n12826) );
  XNOR2_X1 U14967 ( .A(n12825), .B(n12826), .ZN(n12505) );
  XNOR2_X1 U14968 ( .A(n12824), .B(n12505), .ZN(SUB_1596_U67) );
  OAI21_X1 U14969 ( .B1(n12508), .B2(n12507), .A(n12506), .ZN(n12509) );
  NAND2_X1 U14970 ( .A1(n12509), .A2(n13915), .ZN(n12515) );
  NAND2_X1 U14971 ( .A1(n13970), .A2(n14285), .ZN(n12511) );
  NAND2_X1 U14972 ( .A1(n13968), .A2(n14286), .ZN(n12510) );
  NAND2_X1 U14973 ( .A1(n12511), .A2(n12510), .ZN(n12575) );
  NAND2_X1 U14974 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n15582)
         );
  INV_X1 U14975 ( .A(n15582), .ZN(n12513) );
  NOR2_X1 U14976 ( .A1(n13952), .A2(n12604), .ZN(n12512) );
  AOI211_X1 U14977 ( .C1(n13949), .C2(n12575), .A(n12513), .B(n12512), .ZN(
        n12514) );
  OAI211_X1 U14978 ( .C1(n7612), .C2(n13925), .A(n12515), .B(n12514), .ZN(
        P2_U3196) );
  XNOR2_X1 U14979 ( .A(n12517), .B(n12518), .ZN(n12520) );
  NAND2_X1 U14980 ( .A1(n12520), .A2(n12519), .ZN(n14664) );
  OAI211_X1 U14981 ( .C1(n12520), .C2(n12519), .A(n14664), .B(n14754), .ZN(
        n12526) );
  NOR2_X1 U14982 ( .A1(n14790), .A2(n12590), .ZN(n12524) );
  OAI22_X1 U14983 ( .A1(n12522), .A2(n14789), .B1(n14792), .B2(n12521), .ZN(
        n12523) );
  AOI211_X1 U14984 ( .C1(P1_REG3_REG_9__SCAN_IN), .C2(P1_U3086), .A(n12524), 
        .B(n12523), .ZN(n12525) );
  OAI211_X1 U14985 ( .C1(n7050), .C2(n14763), .A(n12526), .B(n12525), .ZN(
        P1_U3231) );
  XNOR2_X1 U14986 ( .A(n12935), .B(n12534), .ZN(n12695) );
  XNOR2_X1 U14987 ( .A(n12695), .B(n12702), .ZN(n12532) );
  INV_X1 U14988 ( .A(n12527), .ZN(n12528) );
  OAI21_X1 U14989 ( .B1(n12532), .B2(n12531), .A(n12700), .ZN(n12533) );
  NAND2_X1 U14990 ( .A1(n12533), .A2(n13353), .ZN(n12542) );
  NOR2_X1 U14991 ( .A1(n13367), .A2(n12534), .ZN(n12539) );
  NAND2_X1 U14992 ( .A1(n13357), .A2(n13379), .ZN(n12536) );
  OAI211_X1 U14993 ( .C1(n12537), .C2(n13359), .A(n12536), .B(n12535), .ZN(
        n12538) );
  AOI211_X1 U14994 ( .C1(n12540), .C2(n13362), .A(n12539), .B(n12538), .ZN(
        n12541) );
  NAND2_X1 U14995 ( .A1(n12542), .A2(n12541), .ZN(P3_U3171) );
  INV_X1 U14996 ( .A(n12543), .ZN(n12546) );
  OAI222_X1 U14997 ( .A1(P2_U3088), .A2(n12545), .B1(n14646), .B2(n12544), 
        .C1(n14644), .C2(n12546), .ZN(P2_U3301) );
  OAI222_X1 U14998 ( .A1(P1_U3086), .A2(n12548), .B1(n15435), .B2(n12547), 
        .C1(n15433), .C2(n12546), .ZN(P1_U3329) );
  XNOR2_X1 U14999 ( .A(n12550), .B(n12549), .ZN(n12554) );
  NAND2_X1 U15000 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n15589)
         );
  OAI21_X1 U15001 ( .B1(n13941), .B2(n12674), .A(n15589), .ZN(n12552) );
  OAI22_X1 U15002 ( .A1(n13952), .A2(n12679), .B1(n12675), .B2(n13908), .ZN(
        n12551) );
  AOI211_X1 U15003 ( .C1(n12678), .C2(n13954), .A(n12552), .B(n12551), .ZN(
        n12553) );
  OAI21_X1 U15004 ( .B1(n12554), .B2(n13956), .A(n12553), .ZN(P2_U3206) );
  OAI21_X1 U15005 ( .B1(n12557), .B2(n12556), .A(n12555), .ZN(n12558) );
  NAND2_X1 U15006 ( .A1(n12558), .A2(n15370), .ZN(n12564) );
  AOI22_X1 U15007 ( .A1(n15257), .A2(n14811), .B1(n14809), .B2(n15258), .ZN(
        n12563) );
  OAI211_X1 U15008 ( .C1(n12561), .C2(n12560), .A(n12559), .B(n15260), .ZN(
        n12562) );
  NAND3_X1 U15009 ( .A1(n12564), .A2(n12563), .A3(n12562), .ZN(n12749) );
  INV_X1 U15010 ( .A(n12749), .ZN(n12571) );
  INV_X1 U15011 ( .A(n12565), .ZN(n12566) );
  AOI211_X1 U15012 ( .C1(n12567), .C2(n12566), .A(n15270), .B(n6601), .ZN(
        n12748) );
  NOR2_X1 U15013 ( .A1(n12755), .A2(n15234), .ZN(n12569) );
  OAI22_X1 U15014 ( .A1(n15220), .A2(n11272), .B1(n12628), .B2(n15217), .ZN(
        n12568) );
  AOI211_X1 U15015 ( .C1(n12748), .C2(n15522), .A(n12569), .B(n12568), .ZN(
        n12570) );
  OAI21_X1 U15016 ( .B1(n12571), .B2(n15274), .A(n12570), .ZN(P1_U3281) );
  XNOR2_X1 U15017 ( .A(n12572), .B(n12573), .ZN(n12603) );
  XNOR2_X1 U15018 ( .A(n12574), .B(n12573), .ZN(n12576) );
  AOI21_X1 U15019 ( .B1(n12576), .B2(n14339), .A(n12575), .ZN(n12612) );
  OAI211_X1 U15020 ( .C1(n6600), .C2(n7612), .A(n14310), .B(n12677), .ZN(
        n12606) );
  OAI211_X1 U15021 ( .C1(n7612), .C2(n15648), .A(n12612), .B(n12606), .ZN(
        n12577) );
  AOI21_X1 U15022 ( .B1(n12603), .B2(n14579), .A(n12577), .ZN(n12580) );
  NAND2_X1 U15023 ( .A1(n15664), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n12578) );
  OAI21_X1 U15024 ( .B1(n12580), .B2(n15664), .A(n12578), .ZN(P2_U3466) );
  NAND2_X1 U15025 ( .A1(n15668), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n12579) );
  OAI21_X1 U15026 ( .B1(n12580), .B2(n15668), .A(n12579), .ZN(P2_U3511) );
  OR2_X1 U15027 ( .A1(n12517), .A2(n12581), .ZN(n12584) );
  AND2_X1 U15028 ( .A1(n12584), .A2(n12582), .ZN(n12586) );
  NAND2_X1 U15029 ( .A1(n12584), .A2(n12583), .ZN(n12585) );
  OAI21_X1 U15030 ( .B1(n12587), .B2(n12586), .A(n12585), .ZN(n12588) );
  NAND2_X1 U15031 ( .A1(n12588), .A2(n14754), .ZN(n12594) );
  OAI22_X1 U15032 ( .A1(n12590), .A2(n14789), .B1(n14792), .B2(n12589), .ZN(
        n12591) );
  AOI211_X1 U15033 ( .C1(n14748), .C2(n14810), .A(n12592), .B(n12591), .ZN(
        n12593) );
  OAI211_X1 U15034 ( .C1(n12694), .C2(n14763), .A(n12594), .B(n12593), .ZN(
        P1_U3236) );
  OAI22_X1 U15035 ( .A1(n12596), .A2(n14326), .B1(n12595), .B2(n15619), .ZN(
        n12599) );
  MUX2_X1 U15036 ( .A(n12597), .B(P2_REG2_REG_9__SCAN_IN), .S(n14341), .Z(
        n12598) );
  AOI211_X1 U15037 ( .C1(n12600), .C2(n14344), .A(n12599), .B(n12598), .ZN(
        n12601) );
  OAI21_X1 U15038 ( .B1(n14346), .B2(n12602), .A(n12601), .ZN(P2_U3256) );
  NAND2_X1 U15039 ( .A1(n12603), .A2(n15630), .ZN(n12611) );
  OAI22_X1 U15040 ( .A1(n15622), .A2(n12605), .B1(n12604), .B2(n15619), .ZN(
        n12608) );
  NOR2_X1 U15041 ( .A1(n12606), .A2(n15627), .ZN(n12607) );
  AOI211_X1 U15042 ( .C1(n15625), .C2(n12609), .A(n12608), .B(n12607), .ZN(
        n12610) );
  OAI211_X1 U15043 ( .C1(n14341), .C2(n12612), .A(n12611), .B(n12610), .ZN(
        P2_U3253) );
  INV_X1 U15044 ( .A(n12615), .ZN(n13124) );
  XNOR2_X1 U15045 ( .A(n12613), .B(n13124), .ZN(n12741) );
  OAI211_X1 U15046 ( .C1(n12616), .C2(n12615), .A(n12614), .B(n13728), .ZN(
        n12618) );
  NAND2_X1 U15047 ( .A1(n13724), .A2(n13376), .ZN(n12617) );
  OAI211_X1 U15048 ( .C1(n13293), .C2(n13643), .A(n12618), .B(n12617), .ZN(
        n12743) );
  INV_X1 U15049 ( .A(n12743), .ZN(n12619) );
  MUX2_X1 U15050 ( .A(n12620), .B(n12619), .S(n15722), .Z(n12623) );
  INV_X1 U15051 ( .A(n13236), .ZN(n12621) );
  NAND2_X1 U15052 ( .A1(n12621), .A2(n13774), .ZN(n12622) );
  OAI211_X1 U15053 ( .C1(n12741), .C2(n13793), .A(n12623), .B(n12622), .ZN(
        P3_U3432) );
  AOI21_X1 U15054 ( .B1(n12625), .B2(n12624), .A(n14797), .ZN(n12627) );
  NAND2_X1 U15055 ( .A1(n12627), .A2(n12626), .ZN(n12633) );
  OAI22_X1 U15056 ( .A1(n12629), .A2(n14789), .B1(n14792), .B2(n12628), .ZN(
        n12630) );
  AOI211_X1 U15057 ( .C1(n14748), .C2(n14809), .A(n12631), .B(n12630), .ZN(
        n12632) );
  OAI211_X1 U15058 ( .C1(n12755), .C2(n14763), .A(n12633), .B(n12632), .ZN(
        P1_U3224) );
  OAI22_X1 U15059 ( .A1(n12741), .A2(n13715), .B1(n13236), .B2(n13709), .ZN(
        n12635) );
  MUX2_X1 U15060 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n12743), .S(n15734), .Z(
        n12634) );
  OR2_X1 U15061 ( .A1(n12635), .A2(n12634), .ZN(P3_U3473) );
  XNOR2_X1 U15062 ( .A(n12645), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14035) );
  XNOR2_X1 U15063 ( .A(n12648), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14051) );
  XNOR2_X1 U15064 ( .A(n14052), .B(n14051), .ZN(n12654) );
  INV_X1 U15065 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15463) );
  NAND2_X1 U15066 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13890)
         );
  OAI21_X1 U15067 ( .B1(n15618), .B2(n15463), .A(n13890), .ZN(n12638) );
  AOI21_X1 U15068 ( .B1(n14050), .B2(n15587), .A(n12638), .ZN(n12653) );
  NAND2_X1 U15069 ( .A1(n12639), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n12643) );
  NAND2_X1 U15070 ( .A1(n12641), .A2(n12640), .ZN(n12642) );
  NAND2_X1 U15071 ( .A1(n12643), .A2(n12642), .ZN(n14033) );
  INV_X1 U15072 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12644) );
  MUX2_X1 U15073 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n12644), .S(n12645), .Z(
        n14034) );
  NAND2_X1 U15074 ( .A1(n14033), .A2(n14034), .ZN(n14032) );
  NAND2_X1 U15075 ( .A1(n12645), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n12650) );
  NAND2_X1 U15076 ( .A1(n14032), .A2(n12650), .ZN(n12647) );
  MUX2_X1 U15077 ( .A(n14277), .B(P2_REG2_REG_17__SCAN_IN), .S(n12648), .Z(
        n12646) );
  NAND2_X1 U15078 ( .A1(n12647), .A2(n12646), .ZN(n14045) );
  MUX2_X1 U15079 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n14277), .S(n12648), .Z(
        n12649) );
  NAND3_X1 U15080 ( .A1(n14032), .A2(n12650), .A3(n12649), .ZN(n12651) );
  NAND3_X1 U15081 ( .A1(n14045), .A2(n15613), .A3(n12651), .ZN(n12652) );
  OAI211_X1 U15082 ( .C1(n12654), .C2(n15597), .A(n12653), .B(n12652), .ZN(
        P2_U3231) );
  AOI21_X1 U15083 ( .B1(n12656), .B2(n12655), .A(n6464), .ZN(n12668) );
  XNOR2_X1 U15084 ( .A(n12658), .B(n12657), .ZN(n12666) );
  NAND2_X1 U15085 ( .A1(n13501), .A2(n12659), .ZN(n12660) );
  NAND2_X1 U15086 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12856)
         );
  OAI211_X1 U15087 ( .C1(n11952), .C2(n13499), .A(n12660), .B(n12856), .ZN(
        n12665) );
  AOI21_X1 U15088 ( .B1(n12662), .B2(n12661), .A(n6466), .ZN(n12663) );
  NOR2_X1 U15089 ( .A1(n12663), .A2(n13490), .ZN(n12664) );
  AOI211_X1 U15090 ( .C1(n13509), .C2(n12666), .A(n12665), .B(n12664), .ZN(
        n12667) );
  OAI21_X1 U15091 ( .B1(n12668), .B2(n13461), .A(n12667), .ZN(P3_U3193) );
  XNOR2_X1 U15092 ( .A(n12670), .B(n12669), .ZN(n14567) );
  INV_X1 U15093 ( .A(n14567), .ZN(n12685) );
  AOI21_X1 U15094 ( .B1(n12672), .B2(n12671), .A(n6450), .ZN(n12673) );
  OAI222_X1 U15095 ( .A1(n14192), .A2(n12675), .B1(n14190), .B2(n12674), .C1(
        n14288), .C2(n12673), .ZN(n14565) );
  NAND2_X1 U15096 ( .A1(n14565), .A2(n15622), .ZN(n12684) );
  INV_X1 U15097 ( .A(n12817), .ZN(n12676) );
  AOI211_X1 U15098 ( .C1(n12678), .C2(n12677), .A(n14320), .B(n12676), .ZN(
        n14566) );
  INV_X1 U15099 ( .A(n12678), .ZN(n14622) );
  NOR2_X1 U15100 ( .A1(n14622), .A2(n14326), .ZN(n12682) );
  OAI22_X1 U15101 ( .A1(n15622), .A2(n12680), .B1(n12679), .B2(n15619), .ZN(
        n12681) );
  AOI211_X1 U15102 ( .C1(n14566), .C2(n14344), .A(n12682), .B(n12681), .ZN(
        n12683) );
  OAI211_X1 U15103 ( .C1(n12685), .C2(n14346), .A(n12684), .B(n12683), .ZN(
        P2_U3252) );
  AOI211_X1 U15104 ( .C1(n15370), .C2(n12689), .A(n12688), .B(n12687), .ZN(
        n12691) );
  MUX2_X1 U15105 ( .A(n14437), .B(n12691), .S(n15554), .Z(n12690) );
  OAI21_X1 U15106 ( .B1(n12694), .B2(n10080), .A(n12690), .ZN(P1_U3539) );
  MUX2_X1 U15107 ( .A(n12692), .B(n12691), .S(n15550), .Z(n12693) );
  OAI21_X1 U15108 ( .B1(n12694), .B2(n10072), .A(n12693), .ZN(P1_U3492) );
  XNOR2_X1 U15109 ( .A(n13110), .B(n12932), .ZN(n12777) );
  XNOR2_X1 U15110 ( .A(n12777), .B(n13109), .ZN(n12698) );
  INV_X1 U15111 ( .A(n12695), .ZN(n12696) );
  NAND2_X1 U15112 ( .A1(n12696), .A2(n12702), .ZN(n12699) );
  AND2_X1 U15113 ( .A1(n12698), .A2(n12699), .ZN(n12697) );
  INV_X1 U15114 ( .A(n12784), .ZN(n12851) );
  AOI21_X1 U15115 ( .B1(n12700), .B2(n12699), .A(n12698), .ZN(n12701) );
  OR3_X1 U15116 ( .A1(n12851), .A2(n13351), .A3(n12701), .ZN(n12708) );
  NAND2_X1 U15117 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n13386)
         );
  OAI21_X1 U15118 ( .B1(n13359), .B2(n12702), .A(n13386), .ZN(n12706) );
  NOR2_X1 U15119 ( .A1(n12704), .A2(n12703), .ZN(n12705) );
  AOI211_X1 U15120 ( .C1(n13357), .C2(n13378), .A(n12706), .B(n12705), .ZN(
        n12707) );
  OAI211_X1 U15121 ( .C1(n13367), .C2(n13110), .A(n12708), .B(n12707), .ZN(
        P3_U3157) );
  OAI21_X1 U15122 ( .B1(n12711), .B2(n12710), .A(n12709), .ZN(n15369) );
  INV_X1 U15123 ( .A(n15369), .ZN(n12723) );
  OAI211_X1 U15124 ( .C1(n12714), .C2(n12713), .A(n12712), .B(n15260), .ZN(
        n12715) );
  OAI21_X1 U15125 ( .B1(n14745), .B2(n15239), .A(n12715), .ZN(n15367) );
  NAND2_X1 U15126 ( .A1(n15256), .A2(n15258), .ZN(n15365) );
  INV_X1 U15127 ( .A(n15365), .ZN(n12716) );
  OAI21_X1 U15128 ( .B1(n15367), .B2(n12716), .A(n15220), .ZN(n12722) );
  OAI22_X1 U15129 ( .A1(n15220), .A2(n12717), .B1(n14744), .B2(n15217), .ZN(
        n12719) );
  INV_X1 U15130 ( .A(n12720), .ZN(n15421) );
  OAI211_X1 U15131 ( .C1(n15421), .C2(n6601), .A(n12769), .B(n15168), .ZN(
        n15366) );
  NOR2_X1 U15132 ( .A1(n15366), .A2(n15174), .ZN(n12718) );
  AOI211_X1 U15133 ( .C1(n15524), .C2(n12720), .A(n12719), .B(n12718), .ZN(
        n12721) );
  OAI211_X1 U15134 ( .C1(n12723), .C2(n15248), .A(n12722), .B(n12721), .ZN(
        P1_U3280) );
  OAI21_X1 U15135 ( .B1(n12726), .B2(n10344), .A(n12725), .ZN(n14578) );
  INV_X1 U15136 ( .A(n14578), .ZN(n12740) );
  NOR2_X1 U15137 ( .A1(n14330), .A2(n12727), .ZN(n12728) );
  NOR2_X1 U15138 ( .A1(n12728), .A2(n10344), .ZN(n14328) );
  AOI211_X1 U15139 ( .C1(n10344), .C2(n12728), .A(n14288), .B(n14328), .ZN(
        n12730) );
  OR2_X1 U15140 ( .A1(n12730), .A2(n12729), .ZN(n14576) );
  INV_X1 U15141 ( .A(n14576), .ZN(n12731) );
  MUX2_X1 U15142 ( .A(n11425), .B(n12731), .S(n15622), .Z(n12739) );
  INV_X1 U15143 ( .A(n12732), .ZN(n12734) );
  AOI211_X1 U15144 ( .C1(n12735), .C2(n12734), .A(n14320), .B(n12733), .ZN(
        n14577) );
  OAI22_X1 U15145 ( .A1(n14628), .A2(n14326), .B1(n15619), .B2(n12736), .ZN(
        n12737) );
  AOI21_X1 U15146 ( .B1(n14577), .B2(n14344), .A(n12737), .ZN(n12738) );
  OAI211_X1 U15147 ( .C1(n14346), .C2(n12740), .A(n12739), .B(n12738), .ZN(
        P2_U3255) );
  INV_X1 U15148 ( .A(n12741), .ZN(n12746) );
  INV_X1 U15149 ( .A(n13233), .ZN(n12742) );
  OAI22_X1 U15150 ( .A1(n13236), .A2(n13588), .B1(n12742), .B2(n13645), .ZN(
        n12745) );
  MUX2_X1 U15151 ( .A(P3_REG2_REG_14__SCAN_IN), .B(n12743), .S(n9345), .Z(
        n12744) );
  AOI211_X1 U15152 ( .C1(n13563), .C2(n12746), .A(n12745), .B(n12744), .ZN(
        n12747) );
  INV_X1 U15153 ( .A(n12747), .ZN(P3_U3219) );
  NOR2_X1 U15154 ( .A1(n12749), .A2(n12748), .ZN(n12752) );
  MUX2_X1 U15155 ( .A(n12750), .B(n12752), .S(n15554), .Z(n12751) );
  OAI21_X1 U15156 ( .B1(n12755), .B2(n10080), .A(n12751), .ZN(P1_U3540) );
  MUX2_X1 U15157 ( .A(n12753), .B(n12752), .S(n15550), .Z(n12754) );
  OAI21_X1 U15158 ( .B1(n12755), .B2(n10072), .A(n12754), .ZN(P1_U3495) );
  XOR2_X1 U15159 ( .A(n13021), .B(n12756), .Z(n12757) );
  OAI222_X1 U15160 ( .A1(n13643), .A2(n13640), .B1(n13641), .B2(n13293), .C1(
        n12757), .C2(n13638), .ZN(n13711) );
  INV_X1 U15161 ( .A(n13711), .ZN(n12762) );
  OAI21_X1 U15162 ( .B1(n12758), .B2(n13021), .A(n13630), .ZN(n13710) );
  INV_X1 U15163 ( .A(n13712), .ZN(n13298) );
  AOI22_X1 U15164 ( .A1(n15691), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15685), 
        .B2(n13295), .ZN(n12759) );
  OAI21_X1 U15165 ( .B1(n13298), .B2(n13588), .A(n12759), .ZN(n12760) );
  AOI21_X1 U15166 ( .B1(n13710), .B2(n13563), .A(n12760), .ZN(n12761) );
  OAI21_X1 U15167 ( .B1(n12762), .B2(n15691), .A(n12761), .ZN(P3_U3217) );
  AOI21_X1 U15168 ( .B1(n12764), .B2(n12763), .A(n15250), .ZN(n15362) );
  INV_X1 U15169 ( .A(n15362), .ZN(n12776) );
  NAND3_X1 U15170 ( .A1(n12712), .A2(n7521), .A3(n12765), .ZN(n12766) );
  NAND3_X1 U15171 ( .A1(n12767), .A2(n15260), .A3(n12766), .ZN(n12768) );
  AOI22_X1 U15172 ( .A1(n14808), .A2(n15258), .B1(n15257), .B2(n14809), .ZN(
        n14653) );
  NAND2_X1 U15173 ( .A1(n12768), .A2(n14653), .ZN(n15360) );
  AOI211_X1 U15174 ( .C1(n7761), .C2(n12769), .A(n15270), .B(n15268), .ZN(
        n15361) );
  NAND2_X1 U15175 ( .A1(n15361), .A2(n15522), .ZN(n12773) );
  INV_X1 U15176 ( .A(n12771), .ZN(n14655) );
  AOI22_X1 U15177 ( .A1(n15533), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n14655), 
        .B2(n15526), .ZN(n12772) );
  OAI211_X1 U15178 ( .C1(n7762), .C2(n15234), .A(n12773), .B(n12772), .ZN(
        n12774) );
  AOI21_X1 U15179 ( .B1(n15360), .B2(n15220), .A(n12774), .ZN(n12775) );
  OAI21_X1 U15180 ( .B1(n12776), .B2(n15248), .A(n12775), .ZN(P1_U3279) );
  XNOR2_X1 U15181 ( .A(n13278), .B(n7063), .ZN(n13271) );
  NAND2_X1 U15182 ( .A1(n12777), .A2(n13379), .ZN(n12853) );
  NAND2_X1 U15183 ( .A1(n12853), .A2(n13275), .ZN(n12778) );
  XNOR2_X1 U15184 ( .A(n12855), .B(n7063), .ZN(n12852) );
  NAND2_X1 U15185 ( .A1(n12852), .A2(n12853), .ZN(n12850) );
  AOI22_X1 U15186 ( .A1(n13271), .A2(n13377), .B1(n12778), .B2(n12850), .ZN(
        n12783) );
  AOI21_X1 U15187 ( .B1(n12852), .B2(n13275), .A(n13270), .ZN(n12781) );
  NAND2_X1 U15188 ( .A1(n13270), .A2(n13275), .ZN(n12780) );
  INV_X1 U15189 ( .A(n12852), .ZN(n12779) );
  OAI22_X1 U15190 ( .A1(n13271), .A2(n12781), .B1(n12780), .B2(n12779), .ZN(
        n12782) );
  XNOR2_X1 U15191 ( .A(n12790), .B(n12932), .ZN(n12786) );
  INV_X1 U15192 ( .A(n12786), .ZN(n12785) );
  NAND2_X1 U15193 ( .A1(n12785), .A2(n13231), .ZN(n12896) );
  INV_X1 U15194 ( .A(n12896), .ZN(n12787) );
  AND2_X1 U15195 ( .A1(n12786), .A2(n13376), .ZN(n12895) );
  NOR2_X1 U15196 ( .A1(n12787), .A2(n12895), .ZN(n12788) );
  XNOR2_X1 U15197 ( .A(n12897), .B(n12788), .ZN(n12795) );
  NAND2_X1 U15198 ( .A1(n13357), .A2(n13375), .ZN(n12789) );
  NAND2_X1 U15199 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n13429)
         );
  OAI211_X1 U15200 ( .C1(n13270), .C2(n13359), .A(n12789), .B(n13429), .ZN(
        n12792) );
  NOR2_X1 U15201 ( .A1(n12790), .A2(n13367), .ZN(n12791) );
  AOI211_X1 U15202 ( .C1(n12793), .C2(n13362), .A(n12792), .B(n12791), .ZN(
        n12794) );
  OAI21_X1 U15203 ( .B1(n12795), .B2(n13351), .A(n12794), .ZN(P3_U3174) );
  XNOR2_X1 U15204 ( .A(n12796), .B(n13130), .ZN(n12797) );
  AOI222_X1 U15205 ( .A1(n13375), .A2(n13724), .B1(n13728), .B2(n12797), .C1(
        n13654), .C2(n13722), .ZN(n12845) );
  MUX2_X1 U15206 ( .A(n7338), .B(n12845), .S(n9345), .Z(n12802) );
  XNOR2_X1 U15207 ( .A(n12798), .B(n13130), .ZN(n12847) );
  INV_X1 U15208 ( .A(n13363), .ZN(n12799) );
  OAI22_X1 U15209 ( .A1(n13366), .A2(n13588), .B1(n12799), .B2(n13645), .ZN(
        n12800) );
  AOI21_X1 U15210 ( .B1(n12847), .B2(n13563), .A(n12800), .ZN(n12801) );
  NAND2_X1 U15211 ( .A1(n12802), .A2(n12801), .ZN(P3_U3218) );
  OAI21_X1 U15212 ( .B1(n12805), .B2(n12804), .A(n12803), .ZN(n12806) );
  NAND2_X1 U15213 ( .A1(n12806), .A2(n13915), .ZN(n12811) );
  INV_X1 U15214 ( .A(n12807), .ZN(n12818) );
  AOI22_X1 U15215 ( .A1(n13937), .A2(n14284), .B1(n13938), .B2(n12818), .ZN(
        n12808) );
  NAND2_X1 U15216 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n15606)
         );
  OAI211_X1 U15217 ( .C1(n12816), .C2(n13941), .A(n12808), .B(n15606), .ZN(
        n12809) );
  AOI21_X1 U15218 ( .B1(n14562), .B2(n13954), .A(n12809), .ZN(n12810) );
  NAND2_X1 U15219 ( .A1(n12811), .A2(n12810), .ZN(P2_U3187) );
  XNOR2_X1 U15220 ( .A(n12812), .B(n12813), .ZN(n14564) );
  XNOR2_X1 U15221 ( .A(n12814), .B(n12813), .ZN(n12815) );
  OAI222_X1 U15222 ( .A1(n14192), .A2(n13882), .B1(n14190), .B2(n12816), .C1(
        n14288), .C2(n12815), .ZN(n14560) );
  INV_X1 U15223 ( .A(n14562), .ZN(n12821) );
  AOI211_X1 U15224 ( .C1(n14562), .C2(n12817), .A(n14320), .B(n14311), .ZN(
        n14561) );
  NAND2_X1 U15225 ( .A1(n14561), .A2(n14344), .ZN(n12820) );
  AOI22_X1 U15226 ( .A1(n14341), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12818), 
        .B2(n14323), .ZN(n12819) );
  OAI211_X1 U15227 ( .C1(n12821), .C2(n14326), .A(n12820), .B(n12819), .ZN(
        n12822) );
  AOI21_X1 U15228 ( .B1(n14560), .B2(n15622), .A(n12822), .ZN(n12823) );
  OAI21_X1 U15229 ( .B1(n14564), .B2(n14346), .A(n12823), .ZN(P2_U3251) );
  INV_X1 U15230 ( .A(n12825), .ZN(n12827) );
  NAND2_X1 U15231 ( .A1(n12827), .A2(n12826), .ZN(n12828) );
  INV_X1 U15232 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n12829) );
  NAND2_X1 U15233 ( .A1(n12829), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n12831) );
  NOR2_X1 U15234 ( .A1(n12829), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n12830) );
  AOI21_X1 U15235 ( .B1(n12832), .B2(n12831), .A(n12830), .ZN(n12868) );
  INV_X1 U15236 ( .A(n12868), .ZN(n12836) );
  INV_X1 U15237 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n12833) );
  NAND2_X1 U15238 ( .A1(n12833), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n12865) );
  NAND2_X1 U15239 ( .A1(n11661), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n12834) );
  AND2_X1 U15240 ( .A1(n12865), .A2(n12834), .ZN(n12867) );
  INV_X1 U15241 ( .A(n12867), .ZN(n12835) );
  XNOR2_X1 U15242 ( .A(n12836), .B(n12835), .ZN(n12837) );
  NOR2_X1 U15243 ( .A1(n12839), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n12864) );
  INV_X1 U15244 ( .A(n12864), .ZN(n12841) );
  OAI21_X1 U15245 ( .B1(n12839), .B2(n12863), .A(P2_ADDR_REG_14__SCAN_IN), 
        .ZN(n12840) );
  OAI21_X1 U15246 ( .B1(n12841), .B2(n12863), .A(n12840), .ZN(SUB_1596_U66) );
  INV_X1 U15247 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12842) );
  MUX2_X1 U15248 ( .A(n12842), .B(n12845), .S(n15734), .Z(n12844) );
  NAND2_X1 U15249 ( .A1(n12847), .A2(n13706), .ZN(n12843) );
  OAI211_X1 U15250 ( .C1(n13709), .C2(n13366), .A(n12844), .B(n12843), .ZN(
        P3_U3474) );
  INV_X1 U15251 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12846) );
  MUX2_X1 U15252 ( .A(n12846), .B(n12845), .S(n15722), .Z(n12849) );
  NAND2_X1 U15253 ( .A1(n12847), .A2(n13785), .ZN(n12848) );
  OAI211_X1 U15254 ( .C1(n13790), .C2(n13366), .A(n12849), .B(n12848), .ZN(
        P3_U3435) );
  NOR2_X1 U15255 ( .A1(n12851), .A2(n12850), .ZN(n13269) );
  AOI21_X1 U15256 ( .B1(n12784), .B2(n12853), .A(n12852), .ZN(n13267) );
  NOR2_X1 U15257 ( .A1(n13269), .A2(n13267), .ZN(n12854) );
  XNOR2_X1 U15258 ( .A(n12854), .B(n13378), .ZN(n12862) );
  NOR2_X1 U15259 ( .A1(n12855), .A2(n13367), .ZN(n12859) );
  NAND2_X1 U15260 ( .A1(n13357), .A2(n13377), .ZN(n12857) );
  OAI211_X1 U15261 ( .C1(n13109), .C2(n13359), .A(n12857), .B(n12856), .ZN(
        n12858) );
  AOI211_X1 U15262 ( .C1(n12860), .C2(n13362), .A(n12859), .B(n12858), .ZN(
        n12861) );
  OAI21_X1 U15263 ( .B1(n12862), .B2(n13351), .A(n12861), .ZN(P3_U3176) );
  INV_X1 U15264 ( .A(n12865), .ZN(n12866) );
  AOI21_X1 U15265 ( .B1(n12868), .B2(n12867), .A(n12866), .ZN(n15447) );
  XNOR2_X1 U15266 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n12869) );
  XNOR2_X1 U15267 ( .A(n15447), .B(n12869), .ZN(n15441) );
  XNOR2_X1 U15268 ( .A(n15441), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(n12870) );
  XNOR2_X1 U15269 ( .A(n15442), .B(n12870), .ZN(SUB_1596_U65) );
  INV_X1 U15270 ( .A(n12871), .ZN(n12873) );
  NAND2_X1 U15271 ( .A1(n15431), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12872) );
  XNOR2_X1 U15272 ( .A(n13213), .B(P1_DATAO_REG_30__SCAN_IN), .ZN(n12946) );
  XNOR2_X1 U15273 ( .A(n12948), .B(n12946), .ZN(n13195) );
  INV_X1 U15274 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12879) );
  NAND2_X1 U15275 ( .A1(n12875), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12878) );
  INV_X1 U15276 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12876) );
  OR2_X1 U15277 ( .A1(n8153), .A2(n12876), .ZN(n12877) );
  OAI211_X1 U15278 ( .C1(n12880), .C2(n12879), .A(n12878), .B(n12877), .ZN(
        n12881) );
  INV_X1 U15279 ( .A(n12881), .ZN(n12882) );
  NAND2_X1 U15280 ( .A1(n13368), .A2(n12884), .ZN(n12888) );
  NOR2_X1 U15281 ( .A1(n12888), .A2(n15721), .ZN(n13735) );
  AOI21_X1 U15282 ( .B1(n15721), .B2(P3_REG0_REG_30__SCAN_IN), .A(n13735), 
        .ZN(n12885) );
  OAI21_X1 U15283 ( .B1(n12996), .B2(n13790), .A(n12885), .ZN(P3_U3457) );
  NOR2_X1 U15284 ( .A1(n12888), .A2(n15731), .ZN(n13665) );
  AOI21_X1 U15285 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n15731), .A(n13665), 
        .ZN(n12886) );
  OAI21_X1 U15286 ( .B1(n12996), .B2(n13709), .A(n12886), .ZN(P3_U3489) );
  OAI21_X1 U15287 ( .B1(n12888), .B2(n15691), .A(n12887), .ZN(n13517) );
  AOI21_X1 U15288 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(n15691), .A(n13517), 
        .ZN(n12889) );
  OAI21_X1 U15289 ( .B1(n12996), .B2(n13588), .A(n12889), .ZN(P3_U3203) );
  INV_X1 U15290 ( .A(n12890), .ZN(n14642) );
  OAI222_X1 U15291 ( .A1(P1_U3086), .A2(n14836), .B1(n15435), .B2(n12891), 
        .C1(n15433), .C2(n14642), .ZN(P1_U3327) );
  INV_X1 U15292 ( .A(n12892), .ZN(n12894) );
  OAI222_X1 U15293 ( .A1(n13805), .A2(n14491), .B1(n13808), .B2(n12894), .C1(
        n12893), .C2(P3_U3151), .ZN(P3_U3266) );
  XNOR2_X1 U15294 ( .A(n13236), .B(n12932), .ZN(n12898) );
  XNOR2_X1 U15295 ( .A(n12898), .B(n13375), .ZN(n13225) );
  NAND2_X1 U15296 ( .A1(n12898), .A2(n13375), .ZN(n12899) );
  XNOR2_X1 U15297 ( .A(n13366), .B(n12932), .ZN(n12900) );
  XNOR2_X1 U15298 ( .A(n12900), .B(n13293), .ZN(n13355) );
  XNOR2_X1 U15299 ( .A(n13712), .B(n12932), .ZN(n12901) );
  XNOR2_X1 U15300 ( .A(n12901), .B(n13654), .ZN(n13290) );
  NAND2_X1 U15301 ( .A1(n13291), .A2(n13290), .ZN(n13289) );
  INV_X1 U15302 ( .A(n12901), .ZN(n12902) );
  NAND2_X1 U15303 ( .A1(n12902), .A2(n13654), .ZN(n12903) );
  NAND2_X1 U15304 ( .A1(n13289), .A2(n12903), .ZN(n13301) );
  XNOR2_X1 U15305 ( .A(n13789), .B(n12932), .ZN(n12904) );
  XNOR2_X1 U15306 ( .A(n12904), .B(n13640), .ZN(n13300) );
  NAND2_X1 U15307 ( .A1(n12904), .A2(n13373), .ZN(n12905) );
  XNOR2_X1 U15308 ( .A(n13702), .B(n12932), .ZN(n12906) );
  XNOR2_X1 U15309 ( .A(n12906), .B(n13655), .ZN(n13336) );
  INV_X1 U15310 ( .A(n12906), .ZN(n12907) );
  NAND2_X1 U15311 ( .A1(n12907), .A2(n13655), .ZN(n12908) );
  XNOR2_X1 U15312 ( .A(n13775), .B(n12932), .ZN(n12909) );
  XNOR2_X1 U15313 ( .A(n12909), .B(n13615), .ZN(n13247) );
  INV_X1 U15314 ( .A(n12909), .ZN(n12910) );
  XNOR2_X1 U15315 ( .A(n13768), .B(n12932), .ZN(n12911) );
  XNOR2_X1 U15316 ( .A(n12911), .B(n13623), .ZN(n13317) );
  INV_X1 U15317 ( .A(n12911), .ZN(n12912) );
  NAND2_X1 U15318 ( .A1(n12912), .A2(n13623), .ZN(n12913) );
  XNOR2_X1 U15319 ( .A(n13762), .B(n12932), .ZN(n12914) );
  XNOR2_X1 U15320 ( .A(n12914), .B(n13320), .ZN(n13260) );
  NAND2_X1 U15321 ( .A1(n12914), .A2(n13320), .ZN(n13237) );
  XNOR2_X1 U15322 ( .A(n8488), .B(n7063), .ZN(n13310) );
  XNOR2_X1 U15323 ( .A(n13243), .B(n7063), .ZN(n13308) );
  AND2_X1 U15324 ( .A1(n13308), .A2(n13595), .ZN(n12915) );
  AOI21_X1 U15325 ( .B1(n13310), .B2(n13582), .A(n12915), .ZN(n12916) );
  XNOR2_X1 U15326 ( .A(n13756), .B(n7063), .ZN(n13325) );
  NAND2_X1 U15327 ( .A1(n13325), .A2(n13604), .ZN(n13239) );
  INV_X1 U15328 ( .A(n12916), .ZN(n12923) );
  INV_X1 U15329 ( .A(n13325), .ZN(n12917) );
  NAND2_X1 U15330 ( .A1(n12917), .A2(n13263), .ZN(n13238) );
  INV_X1 U15331 ( .A(n13310), .ZN(n12921) );
  OAI21_X1 U15332 ( .B1(n13308), .B2(n13595), .A(n13582), .ZN(n12920) );
  NOR2_X1 U15333 ( .A1(n13582), .A2(n13595), .ZN(n12919) );
  INV_X1 U15334 ( .A(n13308), .ZN(n12918) );
  AOI22_X1 U15335 ( .A1(n12921), .A2(n12920), .B1(n12919), .B2(n12918), .ZN(
        n12922) );
  XNOR2_X1 U15336 ( .A(n13675), .B(n12932), .ZN(n12926) );
  XNOR2_X1 U15337 ( .A(n12926), .B(n13541), .ZN(n13283) );
  NAND2_X1 U15338 ( .A1(n13282), .A2(n13283), .ZN(n12928) );
  NAND2_X1 U15339 ( .A1(n12926), .A2(n13570), .ZN(n12927) );
  NAND2_X1 U15340 ( .A1(n12928), .A2(n12927), .ZN(n13344) );
  XNOR2_X1 U15341 ( .A(n13671), .B(n12932), .ZN(n12929) );
  XNOR2_X1 U15342 ( .A(n12929), .B(n13371), .ZN(n13345) );
  NAND2_X1 U15343 ( .A1(n13344), .A2(n13345), .ZN(n12931) );
  NAND2_X1 U15344 ( .A1(n12929), .A2(n13552), .ZN(n12930) );
  NAND2_X1 U15345 ( .A1(n12931), .A2(n12930), .ZN(n13219) );
  XNOR2_X1 U15346 ( .A(n12933), .B(n12932), .ZN(n12934) );
  XNOR2_X1 U15347 ( .A(n12934), .B(n13542), .ZN(n13218) );
  XOR2_X1 U15348 ( .A(n12935), .B(n13520), .Z(n12936) );
  XNOR2_X1 U15349 ( .A(n12937), .B(n12936), .ZN(n12943) );
  AOI22_X1 U15350 ( .A1(n13525), .A2(n13362), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12938) );
  OAI21_X1 U15351 ( .B1(n12939), .B2(n13359), .A(n12938), .ZN(n12941) );
  NOR2_X1 U15352 ( .A1(n13741), .A2(n13367), .ZN(n12940) );
  AOI211_X1 U15353 ( .C1(n13357), .C2(n13522), .A(n12941), .B(n12940), .ZN(
        n12942) );
  OAI21_X1 U15354 ( .B1(n12943), .B2(n13351), .A(n12942), .ZN(P3_U3160) );
  NAND3_X1 U15355 ( .A1(n12945), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n12953) );
  INV_X1 U15356 ( .A(n12946), .ZN(n12947) );
  NAND2_X1 U15357 ( .A1(n13213), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12986) );
  NAND2_X1 U15358 ( .A1(n12992), .A2(n12986), .ZN(n12949) );
  XNOR2_X1 U15359 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12987) );
  INV_X1 U15360 ( .A(n12987), .ZN(n12982) );
  XNOR2_X1 U15361 ( .A(n12949), .B(n12982), .ZN(n12950) );
  NAND2_X1 U15362 ( .A1(n12950), .A2(n13801), .ZN(n12952) );
  NAND2_X1 U15363 ( .A1(n13799), .A2(SI_31_), .ZN(n12951) );
  OAI211_X1 U15364 ( .C1(n12944), .C2(n12953), .A(n12952), .B(n12951), .ZN(
        P3_U3264) );
  INV_X1 U15365 ( .A(n12954), .ZN(n12955) );
  OAI222_X1 U15366 ( .A1(n13805), .A2(n14412), .B1(n13808), .B2(n12955), .C1(
        n13188), .C2(P3_U3151), .ZN(P3_U3268) );
  INV_X1 U15367 ( .A(n12956), .ZN(n12958) );
  OAI222_X1 U15368 ( .A1(P3_U3151), .A2(n12959), .B1(n13808), .B2(n12958), 
        .C1(n12957), .C2(n13805), .ZN(P3_U3269) );
  XNOR2_X1 U15369 ( .A(n12961), .B(n12960), .ZN(n12967) );
  AOI22_X1 U15370 ( .A1(n15037), .A2(n14727), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12963) );
  NAND2_X1 U15371 ( .A1(n15043), .A2(n14776), .ZN(n12962) );
  OAI211_X1 U15372 ( .C1(n12964), .C2(n14790), .A(n12963), .B(n12962), .ZN(
        n12965) );
  AOI21_X1 U15373 ( .B1(n15042), .B2(n14795), .A(n12965), .ZN(n12966) );
  OAI21_X1 U15374 ( .B1(n12967), .B2(n14797), .A(n12966), .ZN(P1_U3214) );
  OAI21_X1 U15375 ( .B1(n12970), .B2(n12969), .A(n12968), .ZN(n12971) );
  NAND2_X1 U15376 ( .A1(n12971), .A2(n14754), .ZN(n12975) );
  AOI22_X1 U15377 ( .A1(n12973), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n14766), 
        .B2(n12972), .ZN(n12974) );
  OAI211_X1 U15378 ( .C1(n7048), .C2(n14763), .A(n12975), .B(n12974), .ZN(
        P1_U3237) );
  INV_X1 U15379 ( .A(SI_24_), .ZN(n12978) );
  INV_X1 U15380 ( .A(n12976), .ZN(n12977) );
  OAI222_X1 U15381 ( .A1(n13805), .A2(n12978), .B1(n13808), .B2(n12977), .C1(
        P3_U3151), .C2(n8510), .ZN(P3_U3271) );
  OAI222_X1 U15382 ( .A1(n9533), .A2(P2_U3088), .B1(n14637), .B2(n12980), .C1(
        n12979), .C2(n14646), .ZN(P2_U3306) );
  INV_X1 U15383 ( .A(n13522), .ZN(n12993) );
  NAND2_X1 U15384 ( .A1(n12988), .A2(n12982), .ZN(n12991) );
  NOR2_X1 U15385 ( .A1(n12987), .A2(n12986), .ZN(n12984) );
  AOI22_X1 U15386 ( .A1(n12985), .A2(n12984), .B1(n12983), .B2(SI_31_), .ZN(
        n12990) );
  NAND4_X1 U15387 ( .A1(n12992), .A2(n12988), .A3(n12987), .A4(n12986), .ZN(
        n12989) );
  OAI22_X1 U15388 ( .A1(n12996), .A2(n13369), .B1(n12997), .B2(n13516), .ZN(
        n13181) );
  NAND2_X1 U15389 ( .A1(n12994), .A2(n12993), .ZN(n13174) );
  OAI21_X1 U15390 ( .B1(n12996), .B2(n13368), .A(n13174), .ZN(n12995) );
  NAND2_X1 U15391 ( .A1(n13177), .A2(n13516), .ZN(n12999) );
  INV_X1 U15392 ( .A(n13147), .ZN(n13001) );
  INV_X1 U15393 ( .A(n13602), .ZN(n13024) );
  INV_X1 U15394 ( .A(n13004), .ZN(n13005) );
  OR2_X1 U15395 ( .A1(n13006), .A2(n13005), .ZN(n13621) );
  AND4_X1 U15396 ( .A1(n13008), .A2(n13074), .A3(n13007), .A4(n13079), .ZN(
        n13012) );
  NOR2_X1 U15397 ( .A1(n11375), .A2(n13009), .ZN(n13010) );
  NAND4_X1 U15398 ( .A1(n13012), .A2(n13092), .A3(n13011), .A4(n13010), .ZN(
        n13014) );
  OR2_X1 U15399 ( .A1(n13014), .A2(n13013), .ZN(n13016) );
  NOR2_X1 U15400 ( .A1(n13016), .A2(n13015), .ZN(n13017) );
  NAND4_X1 U15401 ( .A1(n13018), .A2(n8479), .A3(n13114), .A4(n13017), .ZN(
        n13019) );
  NOR2_X1 U15402 ( .A1(n13126), .A2(n13019), .ZN(n13020) );
  AND4_X1 U15403 ( .A1(n13653), .A2(n13124), .A3(n13130), .A4(n13020), .ZN(
        n13022) );
  NAND4_X1 U15404 ( .A1(n13621), .A2(n13637), .A3(n13022), .A4(n13021), .ZN(
        n13023) );
  OR4_X1 U15405 ( .A1(n13593), .A2(n13024), .A3(n13611), .A4(n13023), .ZN(
        n13025) );
  NOR2_X1 U15406 ( .A1(n13025), .A2(n13580), .ZN(n13026) );
  NAND4_X1 U15407 ( .A1(n13557), .A2(n13165), .A3(n8489), .A4(n13026), .ZN(
        n13027) );
  NOR4_X1 U15408 ( .A1(n13180), .A2(n13520), .A3(n13539), .A4(n13027), .ZN(
        n13030) );
  INV_X1 U15409 ( .A(n13181), .ZN(n13029) );
  NAND4_X1 U15410 ( .A1(n13030), .A2(n13029), .A3(n13028), .A4(n7036), .ZN(
        n13032) );
  INV_X1 U15411 ( .A(n13243), .ZN(n13754) );
  MUX2_X1 U15412 ( .A(n13033), .B(n6497), .S(n13172), .Z(n13143) );
  MUX2_X1 U15413 ( .A(n13035), .B(n13034), .S(n13168), .Z(n13142) );
  INV_X1 U15414 ( .A(n13038), .ZN(n13036) );
  MUX2_X1 U15415 ( .A(n13046), .B(n13036), .S(n13168), .Z(n13141) );
  INV_X1 U15416 ( .A(n13037), .ZN(n13631) );
  NAND2_X1 U15417 ( .A1(n13637), .A2(n13631), .ZN(n13039) );
  NAND3_X1 U15418 ( .A1(n13039), .A2(n13042), .A3(n13038), .ZN(n13048) );
  INV_X1 U15419 ( .A(n13040), .ZN(n13041) );
  NAND2_X1 U15420 ( .A1(n13042), .A2(n13041), .ZN(n13044) );
  NAND2_X1 U15421 ( .A1(n13044), .A2(n13043), .ZN(n13045) );
  OR2_X1 U15422 ( .A1(n13046), .A2(n13045), .ZN(n13047) );
  MUX2_X1 U15423 ( .A(n13048), .B(n13047), .S(n13168), .Z(n13140) );
  INV_X1 U15424 ( .A(n13049), .ZN(n13050) );
  AND2_X1 U15425 ( .A1(n13118), .A2(n13050), .ZN(n13053) );
  AND2_X1 U15426 ( .A1(n13117), .A2(n13051), .ZN(n13052) );
  MUX2_X1 U15427 ( .A(n13053), .B(n13052), .S(n13168), .Z(n13116) );
  NAND2_X1 U15428 ( .A1(n13055), .A2(n13191), .ZN(n13058) );
  NAND2_X1 U15429 ( .A1(n13055), .A2(n13054), .ZN(n13056) );
  NAND3_X1 U15430 ( .A1(n13064), .A2(n13056), .A3(n13172), .ZN(n13057) );
  OAI21_X1 U15431 ( .B1(n11375), .B2(n13058), .A(n13057), .ZN(n13062) );
  NAND2_X1 U15432 ( .A1(n13716), .A2(n13059), .ZN(n13061) );
  AOI21_X1 U15433 ( .B1(n13062), .B2(n13061), .A(n13060), .ZN(n13071) );
  MUX2_X1 U15434 ( .A(n13064), .B(n13063), .S(n13172), .Z(n13070) );
  NAND2_X1 U15435 ( .A1(n13073), .A2(n13065), .ZN(n13068) );
  NAND2_X1 U15436 ( .A1(n13072), .A2(n13066), .ZN(n13067) );
  MUX2_X1 U15437 ( .A(n13068), .B(n13067), .S(n13168), .Z(n13069) );
  MUX2_X1 U15438 ( .A(n13073), .B(n13072), .S(n13172), .Z(n13075) );
  NAND2_X1 U15439 ( .A1(n13075), .A2(n13074), .ZN(n13080) );
  MUX2_X1 U15440 ( .A(n13077), .B(n13076), .S(n13168), .Z(n13078) );
  OAI211_X1 U15441 ( .C1(n13081), .C2(n13080), .A(n13079), .B(n13078), .ZN(
        n13088) );
  NAND2_X1 U15442 ( .A1(n13090), .A2(n13082), .ZN(n13085) );
  NAND2_X1 U15443 ( .A1(n13089), .A2(n13083), .ZN(n13084) );
  MUX2_X1 U15444 ( .A(n13085), .B(n13084), .S(n13172), .Z(n13086) );
  INV_X1 U15445 ( .A(n13086), .ZN(n13087) );
  NAND2_X1 U15446 ( .A1(n13088), .A2(n13087), .ZN(n13093) );
  MUX2_X1 U15447 ( .A(n13090), .B(n13089), .S(n13168), .Z(n13091) );
  NAND3_X1 U15448 ( .A1(n13093), .A2(n13092), .A3(n13091), .ZN(n13098) );
  NAND2_X1 U15449 ( .A1(n15716), .A2(n13382), .ZN(n13095) );
  MUX2_X1 U15450 ( .A(n13095), .B(n13094), .S(n13168), .Z(n13096) );
  NAND3_X1 U15451 ( .A1(n13098), .A2(n13097), .A3(n13096), .ZN(n13103) );
  MUX2_X1 U15452 ( .A(n13100), .B(n13099), .S(n13168), .Z(n13101) );
  NAND3_X1 U15453 ( .A1(n13103), .A2(n13102), .A3(n13101), .ZN(n13107) );
  MUX2_X1 U15454 ( .A(n13105), .B(n13104), .S(n13168), .Z(n13106) );
  NAND2_X1 U15455 ( .A1(n13107), .A2(n13106), .ZN(n13108) );
  NAND2_X1 U15456 ( .A1(n13108), .A2(n8479), .ZN(n13115) );
  NAND2_X1 U15457 ( .A1(n13168), .A2(n13109), .ZN(n13112) );
  NAND2_X1 U15458 ( .A1(n13172), .A2(n13379), .ZN(n13111) );
  MUX2_X1 U15459 ( .A(n13112), .B(n13111), .S(n13110), .Z(n13113) );
  MUX2_X1 U15460 ( .A(n13118), .B(n13117), .S(n13172), .Z(n13119) );
  NAND2_X1 U15461 ( .A1(n13120), .A2(n13119), .ZN(n13125) );
  MUX2_X1 U15462 ( .A(n13122), .B(n13121), .S(n13172), .Z(n13123) );
  MUX2_X1 U15463 ( .A(n13128), .B(n13127), .S(n13168), .Z(n13129) );
  OAI21_X1 U15464 ( .B1(n13712), .B2(n13303), .A(n13131), .ZN(n13132) );
  NAND2_X1 U15465 ( .A1(n13132), .A2(n13172), .ZN(n13133) );
  INV_X1 U15466 ( .A(n13134), .ZN(n13629) );
  AOI21_X1 U15467 ( .B1(n13629), .B2(n13135), .A(n13172), .ZN(n13137) );
  NAND2_X1 U15468 ( .A1(n13654), .A2(n13168), .ZN(n13136) );
  OAI22_X1 U15469 ( .A1(n13138), .A2(n13137), .B1(n13712), .B2(n13136), .ZN(
        n13139) );
  INV_X1 U15470 ( .A(n13145), .ZN(n13146) );
  MUX2_X1 U15471 ( .A(n13147), .B(n13146), .S(n13168), .Z(n13148) );
  INV_X1 U15472 ( .A(n13150), .ZN(n13155) );
  OR2_X1 U15473 ( .A1(n13155), .A2(n13151), .ZN(n13153) );
  NAND2_X1 U15474 ( .A1(n13153), .A2(n13152), .ZN(n13154) );
  NAND2_X1 U15475 ( .A1(n13154), .A2(n13172), .ZN(n13157) );
  NAND2_X1 U15476 ( .A1(n13155), .A2(n13168), .ZN(n13156) );
  NAND2_X1 U15477 ( .A1(n13157), .A2(n13156), .ZN(n13158) );
  MUX2_X1 U15478 ( .A(n13160), .B(n13159), .S(n13172), .Z(n13161) );
  OAI211_X1 U15479 ( .C1(n13162), .C2(n7213), .A(n13537), .B(n13161), .ZN(
        n13166) );
  NAND3_X1 U15480 ( .A1(n13169), .A2(n13168), .A3(n13167), .ZN(n13170) );
  NOR3_X1 U15481 ( .A1(n13173), .A2(n13520), .A3(n13172), .ZN(n13176) );
  INV_X1 U15482 ( .A(n13174), .ZN(n13175) );
  NOR2_X1 U15483 ( .A1(n13176), .A2(n13175), .ZN(n13178) );
  OAI21_X1 U15484 ( .B1(n13182), .B2(n13181), .A(n12998), .ZN(n13185) );
  NOR2_X1 U15485 ( .A1(n13185), .A2(n13183), .ZN(n13184) );
  NAND3_X1 U15486 ( .A1(n13189), .A2(n13800), .A3(n13188), .ZN(n13190) );
  OAI211_X1 U15487 ( .C1(n13191), .C2(n13193), .A(n13190), .B(P3_B_REG_SCAN_IN), .ZN(n13192) );
  INV_X1 U15488 ( .A(SI_30_), .ZN(n13197) );
  INV_X1 U15489 ( .A(n13195), .ZN(n13196) );
  NAND2_X1 U15490 ( .A1(n13199), .A2(n15220), .ZN(n13211) );
  INV_X1 U15491 ( .A(n13200), .ZN(n13209) );
  INV_X1 U15492 ( .A(n13201), .ZN(n13206) );
  OAI22_X1 U15493 ( .A1(n15220), .A2(n13204), .B1(n13203), .B2(n13202), .ZN(
        n13205) );
  AOI21_X1 U15494 ( .B1(n13206), .B2(n15526), .A(n13205), .ZN(n13207) );
  OAI21_X1 U15495 ( .B1(n10070), .B2(n15234), .A(n13207), .ZN(n13208) );
  AOI21_X1 U15496 ( .B1(n13209), .B2(n15522), .A(n13208), .ZN(n13210) );
  OAI211_X1 U15497 ( .C1(n13198), .C2(n15248), .A(n13211), .B(n13210), .ZN(
        P1_U3356) );
  INV_X1 U15498 ( .A(n13212), .ZN(n13215) );
  OAI222_X1 U15499 ( .A1(n13214), .A2(P1_U3086), .B1(n15426), .B2(n13215), 
        .C1(n13213), .C2(n15435), .ZN(P1_U3325) );
  OAI222_X1 U15500 ( .A1(n14646), .A2(n13217), .B1(n13216), .B2(P2_U3088), 
        .C1(n14644), .C2(n13215), .ZN(P2_U3297) );
  XNOR2_X1 U15501 ( .A(n13219), .B(n13218), .ZN(n13220) );
  NAND2_X1 U15502 ( .A1(n13220), .A2(n13353), .ZN(n13224) );
  AOI22_X1 U15503 ( .A1(n13531), .A2(n13362), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13221) );
  OAI21_X1 U15504 ( .B1(n13552), .B2(n13359), .A(n13221), .ZN(n13222) );
  AOI21_X1 U15505 ( .B1(n13370), .B2(n13357), .A(n13222), .ZN(n13223) );
  OAI211_X1 U15506 ( .C1(n13744), .C2(n13367), .A(n13224), .B(n13223), .ZN(
        P3_U3154) );
  AOI21_X1 U15507 ( .B1(n13226), .B2(n13225), .A(n13351), .ZN(n13228) );
  NAND2_X1 U15508 ( .A1(n13228), .A2(n13227), .ZN(n13235) );
  NAND2_X1 U15509 ( .A1(n13357), .A2(n13374), .ZN(n13230) );
  OAI211_X1 U15510 ( .C1(n13231), .C2(n13359), .A(n13230), .B(n13229), .ZN(
        n13232) );
  AOI21_X1 U15511 ( .B1(n13233), .B2(n13362), .A(n13232), .ZN(n13234) );
  OAI211_X1 U15512 ( .C1(n13367), .C2(n13236), .A(n13235), .B(n13234), .ZN(
        P3_U3155) );
  XNOR2_X1 U15513 ( .A(n13309), .B(n13569), .ZN(n13245) );
  AOI22_X1 U15514 ( .A1(n13604), .A2(n13328), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13241) );
  NAND2_X1 U15515 ( .A1(n13586), .A2(n13362), .ZN(n13240) );
  OAI211_X1 U15516 ( .C1(n13551), .C2(n13331), .A(n13241), .B(n13240), .ZN(
        n13242) );
  AOI21_X1 U15517 ( .B1(n13243), .B2(n13349), .A(n13242), .ZN(n13244) );
  OAI21_X1 U15518 ( .B1(n13245), .B2(n13351), .A(n13244), .ZN(P3_U3156) );
  INV_X1 U15519 ( .A(n13775), .ZN(n13256) );
  OAI211_X1 U15520 ( .C1(n13248), .C2(n13247), .A(n13246), .B(n13353), .ZN(
        n13255) );
  NOR2_X1 U15521 ( .A1(n13359), .A2(n13249), .ZN(n13253) );
  OAI21_X1 U15522 ( .B1(n13251), .B2(n13331), .A(n13250), .ZN(n13252) );
  AOI211_X1 U15523 ( .C1(n13626), .C2(n13362), .A(n13253), .B(n13252), .ZN(
        n13254) );
  OAI211_X1 U15524 ( .C1(n13256), .C2(n13367), .A(n13255), .B(n13254), .ZN(
        P3_U3159) );
  INV_X1 U15525 ( .A(n13257), .ZN(n13258) );
  AOI21_X1 U15526 ( .B1(n13260), .B2(n13259), .A(n13258), .ZN(n13266) );
  AOI22_X1 U15527 ( .A1(n13623), .A2(n13328), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13262) );
  NAND2_X1 U15528 ( .A1(n13607), .A2(n13362), .ZN(n13261) );
  OAI211_X1 U15529 ( .C1(n13263), .C2(n13331), .A(n13262), .B(n13261), .ZN(
        n13264) );
  AOI21_X1 U15530 ( .B1(n13762), .B2(n13349), .A(n13264), .ZN(n13265) );
  OAI21_X1 U15531 ( .B1(n13266), .B2(n13351), .A(n13265), .ZN(P3_U3163) );
  INV_X1 U15532 ( .A(n13267), .ZN(n13268) );
  OAI21_X1 U15533 ( .B1(n13269), .B2(n13275), .A(n13268), .ZN(n13273) );
  XNOR2_X1 U15534 ( .A(n13271), .B(n13270), .ZN(n13272) );
  XNOR2_X1 U15535 ( .A(n13273), .B(n13272), .ZN(n13281) );
  NAND2_X1 U15536 ( .A1(n13357), .A2(n13376), .ZN(n13274) );
  NAND2_X1 U15537 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n13405)
         );
  OAI211_X1 U15538 ( .C1(n13275), .C2(n13359), .A(n13274), .B(n13405), .ZN(
        n13276) );
  AOI21_X1 U15539 ( .B1(n13277), .B2(n13362), .A(n13276), .ZN(n13280) );
  NAND2_X1 U15540 ( .A1(n13278), .A2(n13349), .ZN(n13279) );
  OAI211_X1 U15541 ( .C1(n13281), .C2(n13351), .A(n13280), .B(n13279), .ZN(
        P3_U3164) );
  XOR2_X1 U15542 ( .A(n13283), .B(n13282), .Z(n13288) );
  NAND2_X1 U15543 ( .A1(n13371), .A2(n13357), .ZN(n13285) );
  AOI22_X1 U15544 ( .A1(n13559), .A2(n13362), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13284) );
  OAI211_X1 U15545 ( .C1(n13551), .C2(n13359), .A(n13285), .B(n13284), .ZN(
        n13286) );
  AOI21_X1 U15546 ( .B1(n13675), .B2(n13349), .A(n13286), .ZN(n13287) );
  OAI21_X1 U15547 ( .B1(n13288), .B2(n13351), .A(n13287), .ZN(P3_U3165) );
  OAI211_X1 U15548 ( .C1(n13291), .C2(n13290), .A(n13289), .B(n13353), .ZN(
        n13297) );
  AND2_X1 U15549 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13467) );
  AOI21_X1 U15550 ( .B1(n13357), .B2(n13373), .A(n13467), .ZN(n13292) );
  OAI21_X1 U15551 ( .B1(n13293), .B2(n13359), .A(n13292), .ZN(n13294) );
  AOI21_X1 U15552 ( .B1(n13295), .B2(n13362), .A(n13294), .ZN(n13296) );
  OAI211_X1 U15553 ( .C1(n13298), .C2(n13367), .A(n13297), .B(n13296), .ZN(
        P3_U3166) );
  OAI211_X1 U15554 ( .C1(n13301), .C2(n13300), .A(n13299), .B(n13353), .ZN(
        n13306) );
  AND2_X1 U15555 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13482) );
  AOI21_X1 U15556 ( .B1(n13357), .B2(n13655), .A(n13482), .ZN(n13302) );
  OAI21_X1 U15557 ( .B1(n13303), .B2(n13359), .A(n13302), .ZN(n13304) );
  AOI21_X1 U15558 ( .B1(n13658), .B2(n13362), .A(n13304), .ZN(n13305) );
  OAI211_X1 U15559 ( .C1(n13367), .C2(n13789), .A(n13306), .B(n13305), .ZN(
        P3_U3168) );
  XNOR2_X1 U15560 ( .A(n13310), .B(n13582), .ZN(n13311) );
  NAND2_X1 U15561 ( .A1(n13541), .A2(n13357), .ZN(n13313) );
  AOI22_X1 U15562 ( .A1(n13574), .A2(n13362), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13312) );
  OAI211_X1 U15563 ( .C1(n13569), .C2(n13359), .A(n13313), .B(n13312), .ZN(
        n13314) );
  AOI21_X1 U15564 ( .B1(n8488), .B2(n13349), .A(n13314), .ZN(n13315) );
  INV_X1 U15565 ( .A(n13768), .ZN(n13324) );
  OAI211_X1 U15566 ( .C1(n13318), .C2(n13317), .A(n13316), .B(n13353), .ZN(
        n13323) );
  AOI22_X1 U15567 ( .A1(n13328), .A2(n13615), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13319) );
  OAI21_X1 U15568 ( .B1(n13320), .B2(n13331), .A(n13319), .ZN(n13321) );
  AOI21_X1 U15569 ( .B1(n13617), .B2(n13362), .A(n13321), .ZN(n13322) );
  OAI211_X1 U15570 ( .C1(n13324), .C2(n13367), .A(n13323), .B(n13322), .ZN(
        P3_U3173) );
  XNOR2_X1 U15571 ( .A(n13325), .B(n13604), .ZN(n13326) );
  XNOR2_X1 U15572 ( .A(n13327), .B(n13326), .ZN(n13334) );
  AOI22_X1 U15573 ( .A1(n13613), .A2(n13328), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13330) );
  NAND2_X1 U15574 ( .A1(n13598), .A2(n13362), .ZN(n13329) );
  OAI211_X1 U15575 ( .C1(n13569), .C2(n13331), .A(n13330), .B(n13329), .ZN(
        n13332) );
  AOI21_X1 U15576 ( .B1(n13756), .B2(n13349), .A(n13332), .ZN(n13333) );
  OAI21_X1 U15577 ( .B1(n13334), .B2(n13351), .A(n13333), .ZN(P3_U3175) );
  INV_X1 U15578 ( .A(n13702), .ZN(n13343) );
  OAI211_X1 U15579 ( .C1(n13337), .C2(n13336), .A(n13335), .B(n13353), .ZN(
        n13342) );
  NAND2_X1 U15580 ( .A1(n13615), .A2(n13357), .ZN(n13339) );
  NAND2_X1 U15581 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13498)
         );
  OAI211_X1 U15582 ( .C1(n13640), .C2(n13359), .A(n13339), .B(n13498), .ZN(
        n13340) );
  AOI21_X1 U15583 ( .B1(n13644), .B2(n13362), .A(n13340), .ZN(n13341) );
  OAI211_X1 U15584 ( .C1(n13343), .C2(n13367), .A(n13342), .B(n13341), .ZN(
        P3_U3178) );
  XOR2_X1 U15585 ( .A(n13345), .B(n13344), .Z(n13352) );
  NAND2_X1 U15586 ( .A1(n13542), .A2(n13357), .ZN(n13347) );
  AOI22_X1 U15587 ( .A1(n13546), .A2(n13362), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13346) );
  OAI211_X1 U15588 ( .C1(n13570), .C2(n13359), .A(n13347), .B(n13346), .ZN(
        n13348) );
  AOI21_X1 U15589 ( .B1(n13671), .B2(n13349), .A(n13348), .ZN(n13350) );
  OAI21_X1 U15590 ( .B1(n13352), .B2(n13351), .A(n13350), .ZN(P3_U3180) );
  OAI211_X1 U15591 ( .C1(n13356), .C2(n13355), .A(n13354), .B(n13353), .ZN(
        n13365) );
  AND2_X1 U15592 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13446) );
  AOI21_X1 U15593 ( .B1(n13357), .B2(n13654), .A(n13446), .ZN(n13358) );
  OAI21_X1 U15594 ( .B1(n13360), .B2(n13359), .A(n13358), .ZN(n13361) );
  AOI21_X1 U15595 ( .B1(n13363), .B2(n13362), .A(n13361), .ZN(n13364) );
  OAI211_X1 U15596 ( .C1(n13367), .C2(n13366), .A(n13365), .B(n13364), .ZN(
        P3_U3181) );
  MUX2_X1 U15597 ( .A(n13368), .B(P3_DATAO_REG_31__SCAN_IN), .S(n13372), .Z(
        P3_U3522) );
  MUX2_X1 U15598 ( .A(n13369), .B(P3_DATAO_REG_30__SCAN_IN), .S(n13372), .Z(
        P3_U3521) );
  MUX2_X1 U15599 ( .A(n13522), .B(P3_DATAO_REG_29__SCAN_IN), .S(n13372), .Z(
        P3_U3520) );
  MUX2_X1 U15600 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n13370), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15601 ( .A(n13371), .B(P3_DATAO_REG_26__SCAN_IN), .S(n13372), .Z(
        P3_U3517) );
  MUX2_X1 U15602 ( .A(n13582), .B(P3_DATAO_REG_24__SCAN_IN), .S(n13372), .Z(
        P3_U3515) );
  MUX2_X1 U15603 ( .A(n13595), .B(P3_DATAO_REG_23__SCAN_IN), .S(n13372), .Z(
        P3_U3514) );
  MUX2_X1 U15604 ( .A(n13604), .B(P3_DATAO_REG_22__SCAN_IN), .S(n13372), .Z(
        P3_U3513) );
  MUX2_X1 U15605 ( .A(n13613), .B(P3_DATAO_REG_21__SCAN_IN), .S(n13372), .Z(
        P3_U3512) );
  MUX2_X1 U15606 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13623), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15607 ( .A(n13615), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13372), .Z(
        P3_U3510) );
  MUX2_X1 U15608 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13655), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15609 ( .A(n13373), .B(P3_DATAO_REG_17__SCAN_IN), .S(n13372), .Z(
        P3_U3508) );
  MUX2_X1 U15610 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13654), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15611 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n13374), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15612 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n13375), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15613 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n13376), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15614 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13377), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15615 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13378), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15616 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n13379), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15617 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n13380), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15618 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13381), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15619 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n13382), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15620 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13383), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15621 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13384), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15622 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n13385), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15623 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13721), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15624 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n11181), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15625 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n6432), .S(P3_U3897), .Z(
        P3_U3491) );
  OAI21_X1 U15626 ( .B1(n13499), .B2(n11799), .A(n13386), .ZN(n13392) );
  AOI21_X1 U15627 ( .B1(n13389), .B2(n13388), .A(n13387), .ZN(n13390) );
  NOR2_X1 U15628 ( .A1(n13390), .A2(n13407), .ZN(n13391) );
  AOI211_X1 U15629 ( .C1(n13501), .C2(n13393), .A(n13392), .B(n13391), .ZN(
        n13404) );
  AND3_X1 U15630 ( .A1(n13395), .A2(n13394), .A3(n7487), .ZN(n13396) );
  OAI21_X1 U15631 ( .B1(n13397), .B2(n13396), .A(n13495), .ZN(n13403) );
  AND3_X1 U15632 ( .A1(n11839), .A2(n13399), .A3(n13398), .ZN(n13400) );
  OAI21_X1 U15633 ( .B1(n13401), .B2(n13400), .A(n13504), .ZN(n13402) );
  NAND3_X1 U15634 ( .A1(n13404), .A2(n13403), .A3(n13402), .ZN(P3_U3192) );
  OAI21_X1 U15635 ( .B1(n13499), .B2(n12326), .A(n13405), .ZN(n13411) );
  AOI211_X1 U15636 ( .C1(n13409), .C2(n13408), .A(n13407), .B(n13406), .ZN(
        n13410) );
  AOI211_X1 U15637 ( .C1(n13501), .C2(n13412), .A(n13411), .B(n13410), .ZN(
        n13420) );
  NOR3_X1 U15638 ( .A1(n13414), .A2(n6466), .A3(n13413), .ZN(n13415) );
  OAI21_X1 U15639 ( .B1(n6609), .B2(n13415), .A(n13504), .ZN(n13419) );
  NOR3_X1 U15640 ( .A1(n7511), .A2(n6464), .A3(n13416), .ZN(n13417) );
  OAI21_X1 U15641 ( .B1(n6608), .B2(n13417), .A(n13495), .ZN(n13418) );
  NAND3_X1 U15642 ( .A1(n13420), .A2(n13419), .A3(n13418), .ZN(P3_U3194) );
  INV_X1 U15643 ( .A(n13421), .ZN(n13422) );
  AOI21_X1 U15644 ( .B1(n13424), .B2(n13423), .A(n13422), .ZN(n13439) );
  OAI21_X1 U15645 ( .B1(n13427), .B2(n13426), .A(n13425), .ZN(n13437) );
  NAND2_X1 U15646 ( .A1(n15671), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n13428) );
  OAI211_X1 U15647 ( .C1(n13486), .C2(n13430), .A(n13429), .B(n13428), .ZN(
        n13436) );
  NAND2_X1 U15648 ( .A1(n13432), .A2(n13431), .ZN(n13433) );
  AOI21_X1 U15649 ( .B1(n13434), .B2(n13433), .A(n13490), .ZN(n13435) );
  AOI211_X1 U15650 ( .C1(n13509), .C2(n13437), .A(n13436), .B(n13435), .ZN(
        n13438) );
  OAI21_X1 U15651 ( .B1(n13439), .B2(n13461), .A(n13438), .ZN(P3_U3195) );
  AOI21_X1 U15652 ( .B1(n7338), .B2(n6500), .A(n13440), .ZN(n13453) );
  INV_X1 U15653 ( .A(n13460), .ZN(n13441) );
  OAI21_X1 U15654 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n13442), .A(n13441), 
        .ZN(n13451) );
  OAI211_X1 U15655 ( .C1(n13445), .C2(n13444), .A(n13443), .B(n13509), .ZN(
        n13448) );
  AOI21_X1 U15656 ( .B1(n15671), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n13446), 
        .ZN(n13447) );
  OAI211_X1 U15657 ( .C1(n13486), .C2(n13449), .A(n13448), .B(n13447), .ZN(
        n13450) );
  AOI21_X1 U15658 ( .B1(n13451), .B2(n13495), .A(n13450), .ZN(n13452) );
  OAI21_X1 U15659 ( .B1(n13453), .B2(n13490), .A(n13452), .ZN(P3_U3197) );
  OR3_X1 U15660 ( .A1(n13440), .A2(n13455), .A3(n13454), .ZN(n13456) );
  AOI21_X1 U15661 ( .B1(n13457), .B2(n13456), .A(n13490), .ZN(n13473) );
  OR3_X1 U15662 ( .A1(n13460), .A2(n7093), .A3(n13458), .ZN(n13462) );
  AOI21_X1 U15663 ( .B1(n13463), .B2(n13462), .A(n13461), .ZN(n13472) );
  OAI211_X1 U15664 ( .C1(n13466), .C2(n13465), .A(n13464), .B(n13509), .ZN(
        n13469) );
  AOI21_X1 U15665 ( .B1(n15671), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n13467), 
        .ZN(n13468) );
  OAI211_X1 U15666 ( .C1(n13486), .C2(n13470), .A(n13469), .B(n13468), .ZN(
        n13471) );
  OR3_X1 U15667 ( .A1(n13473), .A2(n13472), .A3(n13471), .ZN(P3_U3198) );
  INV_X1 U15668 ( .A(n13474), .ZN(n13475) );
  AOI21_X1 U15669 ( .B1(n13657), .B2(n13476), .A(n13475), .ZN(n13491) );
  OAI21_X1 U15670 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n7485), .A(n13478), .ZN(
        n13488) );
  OAI211_X1 U15671 ( .C1(n13481), .C2(n13480), .A(n13479), .B(n13509), .ZN(
        n13484) );
  AOI21_X1 U15672 ( .B1(n15671), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n13482), 
        .ZN(n13483) );
  OAI211_X1 U15673 ( .C1(n13486), .C2(n13485), .A(n13484), .B(n13483), .ZN(
        n13487) );
  AOI21_X1 U15674 ( .B1(n13488), .B2(n13495), .A(n13487), .ZN(n13489) );
  OAI21_X1 U15675 ( .B1(n13491), .B2(n13490), .A(n13489), .ZN(P3_U3199) );
  INV_X1 U15676 ( .A(n13492), .ZN(n13497) );
  OAI21_X1 U15677 ( .B1(n13497), .B2(n13496), .A(n13495), .ZN(n13515) );
  INV_X1 U15678 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15475) );
  OAI21_X1 U15679 ( .B1(n13499), .B2(n15475), .A(n13498), .ZN(n13500) );
  AOI21_X1 U15680 ( .B1(n13501), .B2(n6599), .A(n13500), .ZN(n13514) );
  AND3_X1 U15681 ( .A1(n13503), .A2(n13474), .A3(n13502), .ZN(n13505) );
  OAI21_X1 U15682 ( .B1(n13506), .B2(n13505), .A(n13504), .ZN(n13513) );
  AND2_X1 U15683 ( .A1(n13508), .A2(n13507), .ZN(n13510) );
  OAI21_X1 U15684 ( .B1(n13511), .B2(n13510), .A(n13509), .ZN(n13512) );
  NAND4_X1 U15685 ( .A1(n13515), .A2(n13514), .A3(n13513), .A4(n13512), .ZN(
        P3_U3200) );
  INV_X1 U15686 ( .A(n13516), .ZN(n13737) );
  AOI21_X1 U15687 ( .B1(n15691), .B2(P3_REG2_REG_31__SCAN_IN), .A(n13517), 
        .ZN(n13518) );
  OAI21_X1 U15688 ( .B1(n13737), .B2(n13588), .A(n13518), .ZN(P3_U3202) );
  INV_X1 U15689 ( .A(n13668), .ZN(n13529) );
  OAI211_X1 U15690 ( .C1(n13521), .C2(n13520), .A(n13519), .B(n13728), .ZN(
        n13524) );
  AOI22_X1 U15691 ( .A1(n13522), .A2(n13722), .B1(n13724), .B2(n13542), .ZN(
        n13523) );
  AOI22_X1 U15692 ( .A1(n13525), .A2(n15685), .B1(n15691), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13526) );
  OAI21_X1 U15693 ( .B1(n13741), .B2(n13588), .A(n13526), .ZN(n13527) );
  AOI21_X1 U15694 ( .B1(n13667), .B2(n9345), .A(n13527), .ZN(n13528) );
  OAI21_X1 U15695 ( .B1(n13663), .B2(n13529), .A(n13528), .ZN(P3_U3205) );
  INV_X1 U15696 ( .A(n13530), .ZN(n13536) );
  AOI22_X1 U15697 ( .A1(n13531), .A2(n15685), .B1(n15691), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13532) );
  OAI21_X1 U15698 ( .B1(n13744), .B2(n13588), .A(n13532), .ZN(n13533) );
  AOI21_X1 U15699 ( .B1(n13534), .B2(n15687), .A(n13533), .ZN(n13535) );
  OAI21_X1 U15700 ( .B1(n13536), .B2(n15691), .A(n13535), .ZN(P3_U3206) );
  XNOR2_X1 U15701 ( .A(n13540), .B(n13539), .ZN(n13544) );
  AOI22_X1 U15702 ( .A1(n13542), .A2(n13722), .B1(n13724), .B2(n13541), .ZN(
        n13543) );
  OAI21_X1 U15703 ( .B1(n13544), .B2(n13638), .A(n13543), .ZN(n13545) );
  AOI22_X1 U15704 ( .A1(n13546), .A2(n15685), .B1(n15691), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13547) );
  OAI21_X1 U15705 ( .B1(n7159), .B2(n13588), .A(n13547), .ZN(n13548) );
  AOI21_X1 U15706 ( .B1(n13672), .B2(n15687), .A(n13548), .ZN(n13549) );
  OAI21_X1 U15707 ( .B1(n13674), .B2(n15691), .A(n13549), .ZN(P3_U3207) );
  AOI21_X1 U15708 ( .B1(n13550), .B2(n13557), .A(n13638), .ZN(n13555) );
  OAI22_X1 U15709 ( .A1(n13552), .A2(n13643), .B1(n13551), .B2(n13641), .ZN(
        n13553) );
  AOI21_X1 U15710 ( .B1(n13555), .B2(n13554), .A(n13553), .ZN(n13678) );
  OAI21_X1 U15711 ( .B1(n13558), .B2(n13557), .A(n13556), .ZN(n13677) );
  INV_X1 U15712 ( .A(n13675), .ZN(n13561) );
  AOI22_X1 U15713 ( .A1(n13559), .A2(n15685), .B1(n15691), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13560) );
  OAI21_X1 U15714 ( .B1(n13561), .B2(n13588), .A(n13560), .ZN(n13562) );
  AOI21_X1 U15715 ( .B1(n13677), .B2(n13563), .A(n13562), .ZN(n13564) );
  OAI21_X1 U15716 ( .B1(n13678), .B2(n15691), .A(n13564), .ZN(P3_U3208) );
  XNOR2_X1 U15717 ( .A(n13566), .B(n13565), .ZN(n13573) );
  OAI21_X1 U15718 ( .B1(n13568), .B2(n8489), .A(n13567), .ZN(n13681) );
  OAI22_X1 U15719 ( .A1(n13570), .A2(n13643), .B1(n13569), .B2(n13641), .ZN(
        n13571) );
  AOI21_X1 U15720 ( .B1(n13681), .B2(n13718), .A(n13571), .ZN(n13572) );
  OAI21_X1 U15721 ( .B1(n13638), .B2(n13573), .A(n13572), .ZN(n13680) );
  INV_X1 U15722 ( .A(n13680), .ZN(n13578) );
  INV_X1 U15723 ( .A(n8488), .ZN(n13750) );
  AOI22_X1 U15724 ( .A1(n13574), .A2(n15685), .B1(n15691), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13575) );
  OAI21_X1 U15725 ( .B1(n13750), .B2(n13588), .A(n13575), .ZN(n13576) );
  AOI21_X1 U15726 ( .B1(n13681), .B2(n15687), .A(n13576), .ZN(n13577) );
  OAI21_X1 U15727 ( .B1(n13578), .B2(n15691), .A(n13577), .ZN(P3_U3209) );
  XNOR2_X1 U15728 ( .A(n13579), .B(n13580), .ZN(n13585) );
  XNOR2_X1 U15729 ( .A(n13581), .B(n13580), .ZN(n13685) );
  NAND2_X1 U15730 ( .A1(n13685), .A2(n13718), .ZN(n13584) );
  AOI22_X1 U15731 ( .A1(n13582), .A2(n13722), .B1(n13724), .B2(n13604), .ZN(
        n13583) );
  OAI211_X1 U15732 ( .C1(n13585), .C2(n13638), .A(n13584), .B(n13583), .ZN(
        n13684) );
  INV_X1 U15733 ( .A(n13684), .ZN(n13591) );
  AOI22_X1 U15734 ( .A1(n13586), .A2(n15685), .B1(n15691), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n13587) );
  OAI21_X1 U15735 ( .B1(n13754), .B2(n13588), .A(n13587), .ZN(n13589) );
  AOI21_X1 U15736 ( .B1(n13685), .B2(n15687), .A(n13589), .ZN(n13590) );
  OAI21_X1 U15737 ( .B1(n13591), .B2(n15691), .A(n13590), .ZN(P3_U3210) );
  XNOR2_X1 U15738 ( .A(n13592), .B(n13593), .ZN(n13759) );
  INV_X1 U15739 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13597) );
  XNOR2_X1 U15740 ( .A(n13594), .B(n13593), .ZN(n13596) );
  AOI222_X1 U15741 ( .A1(n13596), .A2(n13728), .B1(n13595), .B2(n13722), .C1(
        n13613), .C2(n13724), .ZN(n13755) );
  MUX2_X1 U15742 ( .A(n13597), .B(n13755), .S(n9345), .Z(n13600) );
  AOI22_X1 U15743 ( .A1(n13756), .A2(n13659), .B1(n15685), .B2(n13598), .ZN(
        n13599) );
  OAI211_X1 U15744 ( .C1(n13759), .C2(n13663), .A(n13600), .B(n13599), .ZN(
        P3_U3211) );
  XNOR2_X1 U15745 ( .A(n13601), .B(n13602), .ZN(n13765) );
  XNOR2_X1 U15746 ( .A(n13603), .B(n13602), .ZN(n13605) );
  AOI222_X1 U15747 ( .A1(n13605), .A2(n13728), .B1(n13604), .B2(n13722), .C1(
        n13623), .C2(n13724), .ZN(n13760) );
  MUX2_X1 U15748 ( .A(n13606), .B(n13760), .S(n9345), .Z(n13609) );
  AOI22_X1 U15749 ( .A1(n13762), .A2(n13659), .B1(n15685), .B2(n13607), .ZN(
        n13608) );
  OAI211_X1 U15750 ( .C1(n13765), .C2(n13663), .A(n13609), .B(n13608), .ZN(
        P3_U3212) );
  XNOR2_X1 U15751 ( .A(n13610), .B(n13611), .ZN(n13771) );
  XOR2_X1 U15752 ( .A(n13612), .B(n13611), .Z(n13614) );
  AOI222_X1 U15753 ( .A1(n13615), .A2(n13724), .B1(n13728), .B2(n13614), .C1(
        n13613), .C2(n13722), .ZN(n13766) );
  MUX2_X1 U15754 ( .A(n13616), .B(n13766), .S(n9345), .Z(n13619) );
  AOI22_X1 U15755 ( .A1(n13768), .A2(n13659), .B1(n15685), .B2(n13617), .ZN(
        n13618) );
  OAI211_X1 U15756 ( .C1(n13771), .C2(n13663), .A(n13619), .B(n13618), .ZN(
        P3_U3213) );
  XNOR2_X1 U15757 ( .A(n13620), .B(n13621), .ZN(n13778) );
  XOR2_X1 U15758 ( .A(n13622), .B(n13621), .Z(n13624) );
  AOI222_X1 U15759 ( .A1(n13655), .A2(n13724), .B1(n13728), .B2(n13624), .C1(
        n13623), .C2(n13722), .ZN(n13772) );
  MUX2_X1 U15760 ( .A(n13625), .B(n13772), .S(n9345), .Z(n13628) );
  AOI22_X1 U15761 ( .A1(n13775), .A2(n13659), .B1(n15685), .B2(n13626), .ZN(
        n13627) );
  OAI211_X1 U15762 ( .C1(n13778), .C2(n13663), .A(n13628), .B(n13627), .ZN(
        P3_U3214) );
  NAND2_X1 U15763 ( .A1(n13630), .A2(n13629), .ZN(n13651) );
  AOI21_X1 U15764 ( .B1(n13651), .B2(n13653), .A(n13631), .ZN(n13633) );
  OAI21_X1 U15765 ( .B1(n13633), .B2(n13637), .A(n13632), .ZN(n13782) );
  INV_X1 U15766 ( .A(n6988), .ZN(n13635) );
  AOI21_X1 U15767 ( .B1(n13637), .B2(n13636), .A(n13635), .ZN(n13639) );
  OAI222_X1 U15768 ( .A1(n13643), .A2(n13642), .B1(n13641), .B2(n13640), .C1(
        n13639), .C2(n13638), .ZN(n13701) );
  NAND2_X1 U15769 ( .A1(n13701), .A2(n9345), .ZN(n13650) );
  INV_X1 U15770 ( .A(n13644), .ZN(n13646) );
  OAI22_X1 U15771 ( .A1(n9345), .A2(n13647), .B1(n13646), .B2(n13645), .ZN(
        n13648) );
  AOI21_X1 U15772 ( .B1(n13702), .B2(n13659), .A(n13648), .ZN(n13649) );
  OAI211_X1 U15773 ( .C1(n13782), .C2(n13663), .A(n13650), .B(n13649), .ZN(
        P3_U3215) );
  XNOR2_X1 U15774 ( .A(n13651), .B(n13653), .ZN(n13786) );
  INV_X1 U15775 ( .A(n13786), .ZN(n13664) );
  XOR2_X1 U15776 ( .A(n13653), .B(n13652), .Z(n13656) );
  AOI222_X1 U15777 ( .A1(n13656), .A2(n13728), .B1(n13655), .B2(n13722), .C1(
        n13654), .C2(n13724), .ZN(n13783) );
  MUX2_X1 U15778 ( .A(n13657), .B(n13783), .S(n9345), .Z(n13662) );
  INV_X1 U15779 ( .A(n13789), .ZN(n13660) );
  AOI22_X1 U15780 ( .A1(n13660), .A2(n13659), .B1(n15685), .B2(n13658), .ZN(
        n13661) );
  OAI211_X1 U15781 ( .C1(n13664), .C2(n13663), .A(n13662), .B(n13661), .ZN(
        P3_U3216) );
  AOI21_X1 U15782 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n15731), .A(n13665), 
        .ZN(n13666) );
  OAI21_X1 U15783 ( .B1(n13737), .B2(n13709), .A(n13666), .ZN(P3_U3490) );
  INV_X1 U15784 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13669) );
  MUX2_X1 U15785 ( .A(n13669), .B(n13738), .S(n15734), .Z(n13670) );
  AOI22_X1 U15786 ( .A1(n13672), .A2(n15720), .B1(n15703), .B2(n13671), .ZN(
        n13673) );
  NAND2_X1 U15787 ( .A1(n13674), .A2(n13673), .ZN(n13745) );
  MUX2_X1 U15788 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n13745), .S(n15734), .Z(
        P3_U3485) );
  AOI22_X1 U15789 ( .A1(n13677), .A2(n13676), .B1(n15703), .B2(n13675), .ZN(
        n13679) );
  NAND2_X1 U15790 ( .A1(n13679), .A2(n13678), .ZN(n13746) );
  MUX2_X1 U15791 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13746), .S(n15734), .Z(
        P3_U3484) );
  INV_X1 U15792 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13682) );
  AOI21_X1 U15793 ( .B1(n15720), .B2(n13681), .A(n13680), .ZN(n13747) );
  MUX2_X1 U15794 ( .A(n13682), .B(n13747), .S(n15734), .Z(n13683) );
  OAI21_X1 U15795 ( .B1(n13750), .B2(n13709), .A(n13683), .ZN(P3_U3483) );
  INV_X1 U15796 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13686) );
  AOI21_X1 U15797 ( .B1(n15720), .B2(n13685), .A(n13684), .ZN(n13751) );
  MUX2_X1 U15798 ( .A(n13686), .B(n13751), .S(n15734), .Z(n13687) );
  OAI21_X1 U15799 ( .B1(n13754), .B2(n13709), .A(n13687), .ZN(P3_U3482) );
  INV_X1 U15800 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13688) );
  MUX2_X1 U15801 ( .A(n13688), .B(n13755), .S(n15734), .Z(n13690) );
  NAND2_X1 U15802 ( .A1(n13756), .A2(n13698), .ZN(n13689) );
  OAI211_X1 U15803 ( .C1(n13715), .C2(n13759), .A(n13690), .B(n13689), .ZN(
        P3_U3481) );
  INV_X1 U15804 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13691) );
  MUX2_X1 U15805 ( .A(n13691), .B(n13760), .S(n15734), .Z(n13693) );
  NAND2_X1 U15806 ( .A1(n13762), .A2(n13698), .ZN(n13692) );
  OAI211_X1 U15807 ( .C1(n13715), .C2(n13765), .A(n13693), .B(n13692), .ZN(
        P3_U3480) );
  INV_X1 U15808 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13694) );
  MUX2_X1 U15809 ( .A(n13694), .B(n13766), .S(n15734), .Z(n13696) );
  NAND2_X1 U15810 ( .A1(n13768), .A2(n13698), .ZN(n13695) );
  OAI211_X1 U15811 ( .C1(n13715), .C2(n13771), .A(n13696), .B(n13695), .ZN(
        P3_U3479) );
  INV_X1 U15812 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13697) );
  MUX2_X1 U15813 ( .A(n13697), .B(n13772), .S(n15734), .Z(n13700) );
  NAND2_X1 U15814 ( .A1(n13775), .A2(n13698), .ZN(n13699) );
  OAI211_X1 U15815 ( .C1(n13715), .C2(n13778), .A(n13700), .B(n13699), .ZN(
        P3_U3478) );
  AOI21_X1 U15816 ( .B1(n15703), .B2(n13702), .A(n13701), .ZN(n13779) );
  MUX2_X1 U15817 ( .A(n13703), .B(n13779), .S(n15734), .Z(n13704) );
  OAI21_X1 U15818 ( .B1(n13715), .B2(n13782), .A(n13704), .ZN(P3_U3477) );
  MUX2_X1 U15819 ( .A(n13705), .B(n13783), .S(n15734), .Z(n13708) );
  NAND2_X1 U15820 ( .A1(n13786), .A2(n13706), .ZN(n13707) );
  OAI211_X1 U15821 ( .C1(n13709), .C2(n13789), .A(n13708), .B(n13707), .ZN(
        P3_U3476) );
  INV_X1 U15822 ( .A(n13710), .ZN(n13794) );
  AOI21_X1 U15823 ( .B1(n15703), .B2(n13712), .A(n13711), .ZN(n13791) );
  MUX2_X1 U15824 ( .A(n13713), .B(n13791), .S(n15734), .Z(n13714) );
  OAI21_X1 U15825 ( .B1(n13794), .B2(n13715), .A(n13714), .ZN(P3_U3475) );
  INV_X1 U15826 ( .A(n11375), .ZN(n13717) );
  XNOR2_X1 U15827 ( .A(n13716), .B(n13717), .ZN(n15686) );
  NAND2_X1 U15828 ( .A1(n15686), .A2(n13718), .ZN(n13731) );
  OAI21_X1 U15829 ( .B1(n13720), .B2(n11375), .A(n13719), .ZN(n13729) );
  NAND2_X1 U15830 ( .A1(n13722), .A2(n13721), .ZN(n13726) );
  NAND2_X1 U15831 ( .A1(n13724), .A2(n6432), .ZN(n13725) );
  NAND2_X1 U15832 ( .A1(n13726), .A2(n13725), .ZN(n13727) );
  AOI21_X1 U15833 ( .B1(n13729), .B2(n13728), .A(n13727), .ZN(n13730) );
  AND2_X1 U15834 ( .A1(n13731), .A2(n13730), .ZN(n15681) );
  NOR2_X1 U15835 ( .A1(n15715), .A2(n13732), .ZN(n15684) );
  AOI21_X1 U15836 ( .B1(n15686), .B2(n15720), .A(n15684), .ZN(n13733) );
  AND2_X1 U15837 ( .A1(n15681), .A2(n13733), .ZN(n15692) );
  INV_X1 U15838 ( .A(n15692), .ZN(n13734) );
  MUX2_X1 U15839 ( .A(P3_REG1_REG_1__SCAN_IN), .B(n13734), .S(n15734), .Z(
        P3_U3460) );
  AOI21_X1 U15840 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n15721), .A(n13735), 
        .ZN(n13736) );
  OAI21_X1 U15841 ( .B1(n13737), .B2(n13790), .A(n13736), .ZN(P3_U3458) );
  INV_X1 U15842 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13739) );
  MUX2_X1 U15843 ( .A(n13739), .B(n13738), .S(n15722), .Z(n13740) );
  INV_X1 U15844 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13743) );
  MUX2_X1 U15845 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n13745), .S(n15722), .Z(
        P3_U3453) );
  MUX2_X1 U15846 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n13746), .S(n15722), .Z(
        P3_U3452) );
  INV_X1 U15847 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13748) );
  MUX2_X1 U15848 ( .A(n13748), .B(n13747), .S(n15722), .Z(n13749) );
  OAI21_X1 U15849 ( .B1(n13750), .B2(n13790), .A(n13749), .ZN(P3_U3451) );
  INV_X1 U15850 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13752) );
  MUX2_X1 U15851 ( .A(n13752), .B(n13751), .S(n15722), .Z(n13753) );
  OAI21_X1 U15852 ( .B1(n13754), .B2(n13790), .A(n13753), .ZN(P3_U3450) );
  MUX2_X1 U15853 ( .A(n14453), .B(n13755), .S(n15722), .Z(n13758) );
  NAND2_X1 U15854 ( .A1(n13756), .A2(n13774), .ZN(n13757) );
  OAI211_X1 U15855 ( .C1(n13759), .C2(n13793), .A(n13758), .B(n13757), .ZN(
        P3_U3449) );
  INV_X1 U15856 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13761) );
  MUX2_X1 U15857 ( .A(n13761), .B(n13760), .S(n15722), .Z(n13764) );
  NAND2_X1 U15858 ( .A1(n13762), .A2(n13774), .ZN(n13763) );
  OAI211_X1 U15859 ( .C1(n13765), .C2(n13793), .A(n13764), .B(n13763), .ZN(
        P3_U3448) );
  INV_X1 U15860 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13767) );
  MUX2_X1 U15861 ( .A(n13767), .B(n13766), .S(n15722), .Z(n13770) );
  NAND2_X1 U15862 ( .A1(n13768), .A2(n13774), .ZN(n13769) );
  OAI211_X1 U15863 ( .C1(n13771), .C2(n13793), .A(n13770), .B(n13769), .ZN(
        P3_U3447) );
  INV_X1 U15864 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13773) );
  MUX2_X1 U15865 ( .A(n13773), .B(n13772), .S(n15722), .Z(n13777) );
  NAND2_X1 U15866 ( .A1(n13775), .A2(n13774), .ZN(n13776) );
  OAI211_X1 U15867 ( .C1(n13778), .C2(n13793), .A(n13777), .B(n13776), .ZN(
        P3_U3446) );
  INV_X1 U15868 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13780) );
  MUX2_X1 U15869 ( .A(n13780), .B(n13779), .S(n15722), .Z(n13781) );
  OAI21_X1 U15870 ( .B1(n13782), .B2(n13793), .A(n13781), .ZN(P3_U3444) );
  INV_X1 U15871 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13784) );
  MUX2_X1 U15872 ( .A(n13784), .B(n13783), .S(n15722), .Z(n13788) );
  NAND2_X1 U15873 ( .A1(n13786), .A2(n13785), .ZN(n13787) );
  OAI211_X1 U15874 ( .C1(n13790), .C2(n13789), .A(n13788), .B(n13787), .ZN(
        P3_U3441) );
  MUX2_X1 U15875 ( .A(n14482), .B(n13791), .S(n15722), .Z(n13792) );
  OAI21_X1 U15876 ( .B1(n13794), .B2(n13793), .A(n13792), .ZN(P3_U3438) );
  MUX2_X1 U15877 ( .A(P3_D_REG_1__SCAN_IN), .B(n13795), .S(n13797), .Z(
        P3_U3377) );
  INV_X1 U15878 ( .A(n13796), .ZN(n13798) );
  MUX2_X1 U15879 ( .A(P3_D_REG_0__SCAN_IN), .B(n13798), .S(n13797), .Z(
        P3_U3376) );
  AOI222_X1 U15880 ( .A1(n13802), .A2(n13801), .B1(n13800), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_28_), .C2(n13799), .ZN(n13803) );
  INV_X1 U15881 ( .A(n13803), .ZN(P3_U3267) );
  INV_X1 U15882 ( .A(n13804), .ZN(n13807) );
  OAI222_X1 U15883 ( .A1(P3_U3151), .A2(n13809), .B1(n13808), .B2(n13807), 
        .C1(n13806), .C2(n13805), .ZN(P3_U3270) );
  MUX2_X1 U15884 ( .A(n13810), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  AND2_X1 U15885 ( .A1(n13811), .A2(n13917), .ZN(n13914) );
  NOR2_X1 U15886 ( .A1(n13914), .A2(n13812), .ZN(n13816) );
  XNOR2_X1 U15887 ( .A(n13814), .B(n13813), .ZN(n13815) );
  XNOR2_X1 U15888 ( .A(n13816), .B(n13815), .ZN(n13821) );
  OAI22_X1 U15889 ( .A1(n14191), .A2(n13941), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13817), .ZN(n13819) );
  OAI22_X1 U15890 ( .A1(n14127), .A2(n13908), .B1(n14162), .B2(n13952), .ZN(
        n13818) );
  AOI211_X1 U15891 ( .C1(n14378), .C2(n13954), .A(n13819), .B(n13818), .ZN(
        n13820) );
  OAI21_X1 U15892 ( .B1(n13821), .B2(n13956), .A(n13820), .ZN(P2_U3188) );
  NOR2_X1 U15893 ( .A1(n13823), .A2(n13822), .ZN(n13824) );
  XOR2_X1 U15894 ( .A(n13825), .B(n13824), .Z(n13826) );
  NAND2_X1 U15895 ( .A1(n13826), .A2(n13915), .ZN(n13831) );
  AOI22_X1 U15896 ( .A1(n13857), .A2(n9514), .B1(n13937), .B2(n13977), .ZN(
        n13830) );
  AOI22_X1 U15897 ( .A1(n13954), .A2(n13827), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13829) );
  INV_X1 U15898 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n15559) );
  NAND2_X1 U15899 ( .A1(n13938), .A2(n15559), .ZN(n13828) );
  NAND4_X1 U15900 ( .A1(n13831), .A2(n13830), .A3(n13829), .A4(n13828), .ZN(
        P2_U3190) );
  NOR2_X1 U15901 ( .A1(n6801), .A2(n13833), .ZN(n13834) );
  XNOR2_X1 U15902 ( .A(n13835), .B(n13834), .ZN(n13840) );
  OAI22_X1 U15903 ( .A1(n14189), .A2(n14192), .B1(n13836), .B2(n14190), .ZN(
        n14225) );
  NAND2_X1 U15904 ( .A1(n14225), .A2(n13949), .ZN(n13837) );
  NAND2_X1 U15905 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14071)
         );
  OAI211_X1 U15906 ( .C1(n13952), .C2(n14233), .A(n13837), .B(n14071), .ZN(
        n13838) );
  AOI21_X1 U15907 ( .B1(n14232), .B2(n13954), .A(n13838), .ZN(n13839) );
  OAI21_X1 U15908 ( .B1(n13840), .B2(n13956), .A(n13839), .ZN(P2_U3191) );
  NAND2_X1 U15909 ( .A1(n14093), .A2(n14320), .ZN(n13841) );
  XNOR2_X1 U15910 ( .A(n13841), .B(n8969), .ZN(n13842) );
  XNOR2_X1 U15911 ( .A(n14087), .B(n13842), .ZN(n13849) );
  INV_X1 U15912 ( .A(n13849), .ZN(n13843) );
  NAND2_X1 U15913 ( .A1(n13843), .A2(n13915), .ZN(n13855) );
  INV_X1 U15914 ( .A(n13844), .ZN(n13848) );
  NAND2_X1 U15915 ( .A1(n13854), .A2(n7783), .ZN(n13853) );
  INV_X1 U15916 ( .A(n13845), .ZN(n14086) );
  AOI22_X1 U15917 ( .A1(n14086), .A2(n13938), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13846) );
  OAI21_X1 U15918 ( .B1(n13847), .B2(n13891), .A(n13846), .ZN(n13851) );
  NOR3_X1 U15919 ( .A1(n13849), .A2(n13848), .A3(n13956), .ZN(n13850) );
  AOI211_X1 U15920 ( .C1(n14087), .C2(n13954), .A(n13851), .B(n13850), .ZN(
        n13852) );
  OAI211_X1 U15921 ( .C1(n13855), .C2(n13854), .A(n13853), .B(n13852), .ZN(
        P2_U3192) );
  AOI22_X1 U15922 ( .A1(n13857), .A2(n9355), .B1(n13937), .B2(n9514), .ZN(
        n13866) );
  AOI22_X1 U15923 ( .A1(n13954), .A2(n13859), .B1(n13858), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n13865) );
  OAI21_X1 U15924 ( .B1(n13862), .B2(n13861), .A(n13860), .ZN(n13863) );
  NAND2_X1 U15925 ( .A1(n13863), .A2(n13915), .ZN(n13864) );
  NAND3_X1 U15926 ( .A1(n13866), .A2(n13865), .A3(n13864), .ZN(P2_U3194) );
  OAI211_X1 U15927 ( .C1(n13869), .C2(n13868), .A(n13867), .B(n13915), .ZN(
        n13875) );
  OAI22_X1 U15928 ( .A1(n14127), .A2(n13941), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13870), .ZN(n13873) );
  NOR2_X1 U15929 ( .A1(n13871), .A2(n13908), .ZN(n13872) );
  AOI211_X1 U15930 ( .C1(n13938), .C2(n14134), .A(n13873), .B(n13872), .ZN(
        n13874) );
  OAI211_X1 U15931 ( .C1(n7631), .C2(n13925), .A(n13875), .B(n13874), .ZN(
        P2_U3197) );
  NAND2_X1 U15932 ( .A1(n13877), .A2(n13876), .ZN(n13881) );
  XNOR2_X1 U15933 ( .A(n13878), .B(n13879), .ZN(n13946) );
  OAI22_X1 U15934 ( .A1(n13946), .A2(n13945), .B1(n13879), .B2(n13878), .ZN(
        n13880) );
  XOR2_X1 U15935 ( .A(n13881), .B(n13880), .Z(n13886) );
  NAND2_X1 U15936 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n14039)
         );
  OAI21_X1 U15937 ( .B1(n13941), .B2(n13882), .A(n14039), .ZN(n13884) );
  OAI22_X1 U15938 ( .A1(n13952), .A2(n14283), .B1(n13928), .B2(n13908), .ZN(
        n13883) );
  AOI211_X1 U15939 ( .C1(n14546), .C2(n13954), .A(n13884), .B(n13883), .ZN(
        n13885) );
  OAI21_X1 U15940 ( .B1(n13886), .B2(n13956), .A(n13885), .ZN(P2_U3198) );
  AOI21_X1 U15941 ( .B1(n13887), .B2(n13888), .A(n6536), .ZN(n13895) );
  NOR2_X1 U15942 ( .A1(n13952), .A2(n14276), .ZN(n13893) );
  AND2_X1 U15943 ( .A1(n13966), .A2(n14285), .ZN(n13889) );
  AOI21_X1 U15944 ( .B1(n13965), .B2(n14286), .A(n13889), .ZN(n14272) );
  OAI21_X1 U15945 ( .B1(n14272), .B2(n13891), .A(n13890), .ZN(n13892) );
  AOI211_X1 U15946 ( .C1(n14275), .C2(n13954), .A(n13893), .B(n13892), .ZN(
        n13894) );
  OAI21_X1 U15947 ( .B1(n13895), .B2(n13956), .A(n13894), .ZN(P2_U3200) );
  INV_X1 U15948 ( .A(n14149), .ZN(n14594) );
  OAI211_X1 U15949 ( .C1(n13898), .C2(n13897), .A(n13896), .B(n13915), .ZN(
        n13904) );
  AND2_X1 U15950 ( .A1(n13963), .A2(n14285), .ZN(n13899) );
  AOI21_X1 U15951 ( .B1(n13962), .B2(n14286), .A(n13899), .ZN(n14141) );
  INV_X1 U15952 ( .A(n14141), .ZN(n13902) );
  OAI22_X1 U15953 ( .A1(n14150), .A2(n13952), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13900), .ZN(n13901) );
  AOI21_X1 U15954 ( .B1(n13902), .B2(n13949), .A(n13901), .ZN(n13903) );
  OAI211_X1 U15955 ( .C1(n14594), .C2(n13925), .A(n13904), .B(n13903), .ZN(
        P2_U3201) );
  XOR2_X1 U15956 ( .A(n13906), .B(n13905), .Z(n13913) );
  OAI22_X1 U15957 ( .A1(n13918), .A2(n13908), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13907), .ZN(n13911) );
  INV_X1 U15958 ( .A(n14210), .ZN(n13909) );
  OAI22_X1 U15959 ( .A1(n13952), .A2(n13909), .B1(n13941), .B2(n13929), .ZN(
        n13910) );
  AOI211_X1 U15960 ( .C1(n14393), .C2(n13954), .A(n13911), .B(n13910), .ZN(
        n13912) );
  OAI21_X1 U15961 ( .B1(n13913), .B2(n13956), .A(n13912), .ZN(P2_U3205) );
  INV_X1 U15962 ( .A(n13914), .ZN(n13916) );
  OAI211_X1 U15963 ( .C1(n13811), .C2(n13917), .A(n13916), .B(n13915), .ZN(
        n13924) );
  OAI22_X1 U15964 ( .A1(n13919), .A2(n14192), .B1(n13918), .B2(n14190), .ZN(
        n14173) );
  INV_X1 U15965 ( .A(n14181), .ZN(n13921) );
  OAI22_X1 U15966 ( .A1(n13952), .A2(n13921), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13920), .ZN(n13922) );
  AOI21_X1 U15967 ( .B1(n14173), .B2(n13949), .A(n13922), .ZN(n13923) );
  OAI211_X1 U15968 ( .C1(n14599), .C2(n13925), .A(n13924), .B(n13923), .ZN(
        P2_U3207) );
  XNOR2_X1 U15969 ( .A(n13926), .B(n13927), .ZN(n13933) );
  OAI22_X1 U15970 ( .A1(n13929), .A2(n14192), .B1(n13928), .B2(n14190), .ZN(
        n14249) );
  AOI22_X1 U15971 ( .A1(n14249), .A2(n13949), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13930) );
  OAI21_X1 U15972 ( .B1(n14254), .B2(n13952), .A(n13930), .ZN(n13931) );
  AOI21_X1 U15973 ( .B1(n14537), .B2(n13954), .A(n13931), .ZN(n13932) );
  OAI21_X1 U15974 ( .B1(n13933), .B2(n13956), .A(n13932), .ZN(P2_U3210) );
  AOI21_X1 U15975 ( .B1(n13936), .B2(n13935), .A(n13934), .ZN(n13944) );
  NAND2_X1 U15976 ( .A1(n13961), .A2(n13937), .ZN(n13940) );
  AOI22_X1 U15977 ( .A1(n14114), .A2(n13938), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13939) );
  OAI211_X1 U15978 ( .C1(n14109), .C2(n13941), .A(n13940), .B(n13939), .ZN(
        n13942) );
  AOI21_X1 U15979 ( .B1(n14113), .B2(n13954), .A(n13942), .ZN(n13943) );
  OAI21_X1 U15980 ( .B1(n13944), .B2(n13956), .A(n13943), .ZN(P2_U3212) );
  XNOR2_X1 U15981 ( .A(n13946), .B(n13945), .ZN(n13957) );
  NAND2_X1 U15982 ( .A1(n13966), .A2(n14286), .ZN(n13948) );
  NAND2_X1 U15983 ( .A1(n13967), .A2(n14285), .ZN(n13947) );
  NAND2_X1 U15984 ( .A1(n13948), .A2(n13947), .ZN(n14308) );
  NAND2_X1 U15985 ( .A1(n13949), .A2(n14308), .ZN(n13950) );
  OAI211_X1 U15986 ( .C1(n13952), .C2(n14309), .A(n13951), .B(n13950), .ZN(
        n13953) );
  AOI21_X1 U15987 ( .B1(n14313), .B2(n13954), .A(n13953), .ZN(n13955) );
  OAI21_X1 U15988 ( .B1(n13957), .B2(n13956), .A(n13955), .ZN(P2_U3213) );
  INV_X2 U15989 ( .A(P2_U3947), .ZN(n13972) );
  MUX2_X1 U15990 ( .A(n13958), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13972), .Z(
        P2_U3562) );
  MUX2_X1 U15991 ( .A(n13959), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13972), .Z(
        P2_U3561) );
  MUX2_X1 U15992 ( .A(n13960), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13972), .Z(
        P2_U3560) );
  MUX2_X1 U15993 ( .A(n14093), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13972), .Z(
        P2_U3559) );
  MUX2_X1 U15994 ( .A(n13961), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13972), .Z(
        P2_U3558) );
  MUX2_X1 U15995 ( .A(n14125), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13972), .Z(
        P2_U3557) );
  MUX2_X1 U15996 ( .A(n13962), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13972), .Z(
        P2_U3556) );
  MUX2_X1 U15997 ( .A(n14160), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13972), .Z(
        P2_U3555) );
  MUX2_X1 U15998 ( .A(n13963), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13972), .Z(
        P2_U3554) );
  MUX2_X1 U15999 ( .A(n14159), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13972), .Z(
        P2_U3553) );
  MUX2_X1 U16000 ( .A(n14206), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13972), .Z(
        P2_U3552) );
  MUX2_X1 U16001 ( .A(n13964), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13972), .Z(
        P2_U3551) );
  MUX2_X1 U16002 ( .A(n14207), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13972), .Z(
        P2_U3550) );
  MUX2_X1 U16003 ( .A(n13965), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13972), .Z(
        P2_U3549) );
  MUX2_X1 U16004 ( .A(n14287), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13972), .Z(
        P2_U3548) );
  MUX2_X1 U16005 ( .A(n13966), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13972), .Z(
        P2_U3547) );
  MUX2_X1 U16006 ( .A(n14284), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13972), .Z(
        P2_U3546) );
  MUX2_X1 U16007 ( .A(n13967), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13972), .Z(
        P2_U3545) );
  MUX2_X1 U16008 ( .A(n13968), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13972), .Z(
        P2_U3544) );
  MUX2_X1 U16009 ( .A(n13969), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13972), .Z(
        P2_U3543) );
  MUX2_X1 U16010 ( .A(n13970), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13972), .Z(
        P2_U3542) );
  MUX2_X1 U16011 ( .A(n14329), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13972), .Z(
        P2_U3541) );
  MUX2_X1 U16012 ( .A(n13971), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13972), .Z(
        P2_U3540) );
  MUX2_X1 U16013 ( .A(n13973), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13972), .Z(
        P2_U3539) );
  MUX2_X1 U16014 ( .A(n13974), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13972), .Z(
        P2_U3538) );
  MUX2_X1 U16015 ( .A(n13975), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13972), .Z(
        P2_U3537) );
  MUX2_X1 U16016 ( .A(n13976), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13972), .Z(
        P2_U3536) );
  MUX2_X1 U16017 ( .A(n13977), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13972), .Z(
        P2_U3535) );
  MUX2_X1 U16018 ( .A(n13978), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13972), .Z(
        P2_U3534) );
  MUX2_X1 U16019 ( .A(n9514), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13972), .Z(
        P2_U3533) );
  MUX2_X1 U16020 ( .A(n9353), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13972), .Z(
        P2_U3532) );
  MUX2_X1 U16021 ( .A(n9355), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13972), .Z(
        P2_U3531) );
  NAND2_X1 U16022 ( .A1(n15585), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n13979) );
  OAI21_X1 U16023 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n13980), .A(n13979), .ZN(
        n13981) );
  AOI21_X1 U16024 ( .B1(n13982), .B2(n15587), .A(n13981), .ZN(n13996) );
  INV_X1 U16025 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n13984) );
  MUX2_X1 U16026 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n13984), .S(n13983), .Z(
        n13985) );
  OAI21_X1 U16027 ( .B1(n13986), .B2(n13991), .A(n13985), .ZN(n13987) );
  NAND3_X1 U16028 ( .A1(n15613), .A2(n13988), .A3(n13987), .ZN(n13995) );
  INV_X1 U16029 ( .A(n13989), .ZN(n13993) );
  OAI21_X1 U16030 ( .B1(n11049), .B2(n13991), .A(n13990), .ZN(n13992) );
  NAND3_X1 U16031 ( .A1(n15610), .A2(n13993), .A3(n13992), .ZN(n13994) );
  NAND3_X1 U16032 ( .A1(n13996), .A2(n13995), .A3(n13994), .ZN(P2_U3215) );
  OAI21_X1 U16033 ( .B1(n15618), .B2(n13998), .A(n13997), .ZN(n13999) );
  AOI21_X1 U16034 ( .B1(n14000), .B2(n15587), .A(n13999), .ZN(n14013) );
  MUX2_X1 U16035 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11083), .S(n14005), .Z(
        n14002) );
  NAND3_X1 U16036 ( .A1(n14002), .A2(n15562), .A3(n14001), .ZN(n14003) );
  NAND3_X1 U16037 ( .A1(n15613), .A2(n14004), .A3(n14003), .ZN(n14012) );
  MUX2_X1 U16038 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n11073), .S(n14005), .Z(
        n14008) );
  INV_X1 U16039 ( .A(n14006), .ZN(n14007) );
  NAND2_X1 U16040 ( .A1(n14008), .A2(n14007), .ZN(n14010) );
  OAI211_X1 U16041 ( .C1(n6476), .C2(n14010), .A(n15610), .B(n14009), .ZN(
        n14011) );
  NAND3_X1 U16042 ( .A1(n14013), .A2(n14012), .A3(n14011), .ZN(P2_U3218) );
  INV_X1 U16043 ( .A(n14014), .ZN(n14016) );
  MUX2_X1 U16044 ( .A(n11075), .B(P2_REG1_REG_6__SCAN_IN), .S(n14023), .Z(
        n14015) );
  NAND2_X1 U16045 ( .A1(n14016), .A2(n14015), .ZN(n14018) );
  OAI211_X1 U16046 ( .C1(n14019), .C2(n14018), .A(n14017), .B(n15610), .ZN(
        n14031) );
  INV_X1 U16047 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n14021) );
  OAI21_X1 U16048 ( .B1(n15618), .B2(n14021), .A(n14020), .ZN(n14022) );
  AOI21_X1 U16049 ( .B1(n14023), .B2(n15587), .A(n14022), .ZN(n14030) );
  MUX2_X1 U16050 ( .A(n12061), .B(P2_REG2_REG_6__SCAN_IN), .S(n14023), .Z(
        n14024) );
  NAND3_X1 U16051 ( .A1(n14026), .A2(n14025), .A3(n14024), .ZN(n14027) );
  NAND3_X1 U16052 ( .A1(n15613), .A2(n14028), .A3(n14027), .ZN(n14029) );
  NAND3_X1 U16053 ( .A1(n14031), .A2(n14030), .A3(n14029), .ZN(P2_U3220) );
  OAI211_X1 U16054 ( .C1(n14034), .C2(n14033), .A(n14032), .B(n15613), .ZN(
        n14042) );
  XOR2_X1 U16055 ( .A(n14036), .B(n14035), .Z(n14037) );
  NAND2_X1 U16056 ( .A1(n15610), .A2(n14037), .ZN(n14038) );
  NAND2_X1 U16057 ( .A1(n14039), .A2(n14038), .ZN(n14040) );
  AOI21_X1 U16058 ( .B1(n15585), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n14040), 
        .ZN(n14041) );
  OAI211_X1 U16059 ( .C1(n15608), .C2(n14043), .A(n14042), .B(n14041), .ZN(
        P2_U3230) );
  NAND2_X1 U16060 ( .A1(n14050), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n14044) );
  NAND2_X1 U16061 ( .A1(n14045), .A2(n14044), .ZN(n14046) );
  NAND2_X1 U16062 ( .A1(n14046), .A2(n14062), .ZN(n14047) );
  INV_X1 U16063 ( .A(n14066), .ZN(n14048) );
  AOI21_X1 U16064 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n14049), .A(n14048), 
        .ZN(n14059) );
  XNOR2_X1 U16065 ( .A(n14060), .B(n14062), .ZN(n14063) );
  XOR2_X1 U16066 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14063), .Z(n14057) );
  NAND2_X1 U16067 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3088), .ZN(n14054)
         );
  NAND2_X1 U16068 ( .A1(n15585), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n14053) );
  OAI211_X1 U16069 ( .C1(n15608), .C2(n14055), .A(n14054), .B(n14053), .ZN(
        n14056) );
  AOI21_X1 U16070 ( .B1(n14057), .B2(n15610), .A(n14056), .ZN(n14058) );
  OAI21_X1 U16071 ( .B1(n14059), .B2(n15591), .A(n14058), .ZN(P2_U3232) );
  INV_X1 U16072 ( .A(n14060), .ZN(n14061) );
  AOI22_X1 U16073 ( .A1(n14063), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n14062), 
        .B2(n14061), .ZN(n14064) );
  INV_X1 U16074 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14534) );
  XNOR2_X1 U16075 ( .A(n14064), .B(n14534), .ZN(n14069) );
  NAND2_X1 U16076 ( .A1(n14066), .A2(n14065), .ZN(n14067) );
  XNOR2_X1 U16077 ( .A(n14067), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n14068) );
  NAND2_X1 U16078 ( .A1(n14073), .A2(n14344), .ZN(n14076) );
  INV_X1 U16079 ( .A(n14347), .ZN(n14074) );
  NOR2_X1 U16080 ( .A1(n14341), .A2(n14074), .ZN(n14082) );
  AOI21_X1 U16081 ( .B1(n14341), .B2(P2_REG2_REG_31__SCAN_IN), .A(n14082), 
        .ZN(n14075) );
  OAI211_X1 U16082 ( .C1(n14077), .C2(n14326), .A(n14076), .B(n14075), .ZN(
        P2_U3234) );
  INV_X1 U16083 ( .A(n14078), .ZN(n14080) );
  NAND2_X1 U16084 ( .A1(n14348), .A2(n14344), .ZN(n14084) );
  AOI21_X1 U16085 ( .B1(n14341), .B2(P2_REG2_REG_30__SCAN_IN), .A(n14082), 
        .ZN(n14083) );
  OAI211_X1 U16086 ( .C1(n14585), .C2(n14326), .A(n14084), .B(n14083), .ZN(
        P2_U3235) );
  AOI21_X1 U16087 ( .B1(n14086), .B2(n14323), .A(n14085), .ZN(n14092) );
  AOI22_X1 U16088 ( .A1(n14087), .A2(n15625), .B1(n14341), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n14088) );
  OAI21_X1 U16089 ( .B1(n14089), .B2(n15627), .A(n14088), .ZN(n14090) );
  OAI21_X1 U16090 ( .B1(n14092), .B2(n14312), .A(n14091), .ZN(P2_U3237) );
  AOI222_X1 U16091 ( .A1(n14339), .A2(n14094), .B1(n14093), .B2(n14286), .C1(
        n14125), .C2(n14285), .ZN(n14361) );
  OAI211_X1 U16092 ( .C1(n14095), .C2(n14099), .A(n14310), .B(n14096), .ZN(
        n14358) );
  INV_X1 U16093 ( .A(n14358), .ZN(n14101) );
  AOI22_X1 U16094 ( .A1(n14097), .A2(n14323), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14312), .ZN(n14098) );
  OAI21_X1 U16095 ( .B1(n14099), .B2(n14326), .A(n14098), .ZN(n14100) );
  AOI21_X1 U16096 ( .B1(n14101), .B2(n14344), .A(n14100), .ZN(n14105) );
  NAND2_X1 U16097 ( .A1(n10372), .A2(n14102), .ZN(n14357) );
  NAND3_X1 U16098 ( .A1(n14357), .A2(n15630), .A3(n14103), .ZN(n14104) );
  OAI211_X1 U16099 ( .C1(n14361), .C2(n14312), .A(n14105), .B(n14104), .ZN(
        P2_U3238) );
  XNOR2_X1 U16100 ( .A(n14107), .B(n14106), .ZN(n14108) );
  OAI222_X1 U16101 ( .A1(n14192), .A2(n14110), .B1(n14190), .B2(n14109), .C1(
        n14288), .C2(n14108), .ZN(n14362) );
  INV_X1 U16102 ( .A(n14362), .ZN(n14119) );
  XNOR2_X1 U16103 ( .A(n14112), .B(n14111), .ZN(n14364) );
  AOI211_X1 U16104 ( .C1(n14113), .C2(n14132), .A(n14320), .B(n14095), .ZN(
        n14363) );
  NAND2_X1 U16105 ( .A1(n14363), .A2(n14344), .ZN(n14116) );
  AOI22_X1 U16106 ( .A1(n14114), .A2(n14323), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14312), .ZN(n14115) );
  OAI211_X1 U16107 ( .C1(n7629), .C2(n14326), .A(n14116), .B(n14115), .ZN(
        n14117) );
  AOI21_X1 U16108 ( .B1(n14364), .B2(n15630), .A(n14117), .ZN(n14118) );
  OAI21_X1 U16109 ( .B1(n14119), .B2(n14312), .A(n14118), .ZN(P2_U3239) );
  NAND2_X1 U16110 ( .A1(n14120), .A2(n14121), .ZN(n14140) );
  NAND2_X1 U16111 ( .A1(n14140), .A2(n14143), .ZN(n14123) );
  NAND2_X1 U16112 ( .A1(n14123), .A2(n14122), .ZN(n14124) );
  XNOR2_X1 U16113 ( .A(n14124), .B(n14130), .ZN(n14129) );
  NAND2_X1 U16114 ( .A1(n14125), .A2(n14286), .ZN(n14126) );
  OAI21_X1 U16115 ( .B1(n14127), .B2(n14190), .A(n14126), .ZN(n14128) );
  AOI21_X1 U16116 ( .B1(n14129), .B2(n14339), .A(n14128), .ZN(n14371) );
  XNOR2_X1 U16117 ( .A(n14131), .B(n14130), .ZN(n14369) );
  AOI21_X1 U16118 ( .B1(n14147), .B2(n14135), .A(n14320), .ZN(n14133) );
  NAND2_X1 U16119 ( .A1(n14133), .A2(n14132), .ZN(n14367) );
  AOI22_X1 U16120 ( .A1(n14134), .A2(n14323), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14312), .ZN(n14137) );
  NAND2_X1 U16121 ( .A1(n14135), .A2(n15625), .ZN(n14136) );
  OAI211_X1 U16122 ( .C1(n14367), .C2(n15627), .A(n14137), .B(n14136), .ZN(
        n14138) );
  AOI21_X1 U16123 ( .B1(n14369), .B2(n15630), .A(n14138), .ZN(n14139) );
  OAI21_X1 U16124 ( .B1(n14371), .B2(n14312), .A(n14139), .ZN(P2_U3240) );
  XOR2_X1 U16125 ( .A(n14140), .B(n14143), .Z(n14142) );
  OAI21_X1 U16126 ( .B1(n14142), .B2(n14288), .A(n14141), .ZN(n14372) );
  INV_X1 U16127 ( .A(n14372), .ZN(n14156) );
  NAND2_X1 U16128 ( .A1(n14144), .A2(n14143), .ZN(n14145) );
  AND2_X1 U16129 ( .A1(n14146), .A2(n14145), .ZN(n14374) );
  INV_X1 U16130 ( .A(n14147), .ZN(n14148) );
  AOI211_X1 U16131 ( .C1(n14149), .C2(n14164), .A(n14320), .B(n14148), .ZN(
        n14373) );
  NAND2_X1 U16132 ( .A1(n14373), .A2(n14344), .ZN(n14153) );
  INV_X1 U16133 ( .A(n14150), .ZN(n14151) );
  AOI22_X1 U16134 ( .A1(n14151), .A2(n14323), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n14312), .ZN(n14152) );
  OAI211_X1 U16135 ( .C1(n14594), .C2(n14326), .A(n14153), .B(n14152), .ZN(
        n14154) );
  AOI21_X1 U16136 ( .B1(n14374), .B2(n15630), .A(n14154), .ZN(n14155) );
  OAI21_X1 U16137 ( .B1(n14156), .B2(n14312), .A(n14155), .ZN(P2_U3241) );
  XNOR2_X1 U16138 ( .A(n14158), .B(n14157), .ZN(n14381) );
  OAI21_X1 U16139 ( .B1(n6510), .B2(n7571), .A(n14120), .ZN(n14161) );
  AOI222_X1 U16140 ( .A1(n14339), .A2(n14161), .B1(n14160), .B2(n14286), .C1(
        n14159), .C2(n14285), .ZN(n14380) );
  OAI21_X1 U16141 ( .B1(n14162), .B2(n15619), .A(n14380), .ZN(n14163) );
  NAND2_X1 U16142 ( .A1(n14163), .A2(n15622), .ZN(n14171) );
  INV_X1 U16143 ( .A(n14178), .ZN(n14166) );
  INV_X1 U16144 ( .A(n14164), .ZN(n14165) );
  AOI211_X1 U16145 ( .C1(n14378), .C2(n14166), .A(n14320), .B(n14165), .ZN(
        n14377) );
  INV_X1 U16146 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n14167) );
  OAI22_X1 U16147 ( .A1(n14168), .A2(n14326), .B1(n14167), .B2(n15622), .ZN(
        n14169) );
  AOI21_X1 U16148 ( .B1(n14377), .B2(n14344), .A(n14169), .ZN(n14170) );
  OAI211_X1 U16149 ( .C1(n14381), .C2(n14346), .A(n14171), .B(n14170), .ZN(
        P2_U3242) );
  XNOR2_X1 U16150 ( .A(n14172), .B(n14177), .ZN(n14175) );
  INV_X1 U16151 ( .A(n14173), .ZN(n14174) );
  OAI21_X1 U16152 ( .B1(n14175), .B2(n14288), .A(n14174), .ZN(n14382) );
  INV_X1 U16153 ( .A(n14382), .ZN(n14186) );
  XOR2_X1 U16154 ( .A(n14176), .B(n14177), .Z(n14384) );
  INV_X1 U16155 ( .A(n14195), .ZN(n14179) );
  AOI211_X1 U16156 ( .C1(n14180), .C2(n14179), .A(n14320), .B(n14178), .ZN(
        n14383) );
  NAND2_X1 U16157 ( .A1(n14383), .A2(n14344), .ZN(n14183) );
  AOI22_X1 U16158 ( .A1(n14181), .A2(n14323), .B1(n14341), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n14182) );
  OAI211_X1 U16159 ( .C1(n14599), .C2(n14326), .A(n14183), .B(n14182), .ZN(
        n14184) );
  AOI21_X1 U16160 ( .B1(n14384), .B2(n15630), .A(n14184), .ZN(n14185) );
  OAI21_X1 U16161 ( .B1(n14186), .B2(n14312), .A(n14185), .ZN(P2_U3243) );
  XNOR2_X1 U16162 ( .A(n14187), .B(n14193), .ZN(n14188) );
  OAI222_X1 U16163 ( .A1(n14192), .A2(n14191), .B1(n14190), .B2(n14189), .C1(
        n14288), .C2(n14188), .ZN(n14387) );
  INV_X1 U16164 ( .A(n14387), .ZN(n14203) );
  XOR2_X1 U16165 ( .A(n14194), .B(n14193), .Z(n14389) );
  AOI211_X1 U16166 ( .C1(n14196), .C2(n14208), .A(n14320), .B(n14195), .ZN(
        n14388) );
  NAND2_X1 U16167 ( .A1(n14388), .A2(n14344), .ZN(n14200) );
  INV_X1 U16168 ( .A(n14197), .ZN(n14198) );
  AOI22_X1 U16169 ( .A1(P2_REG2_REG_21__SCAN_IN), .A2(n14312), .B1(n14198), 
        .B2(n14323), .ZN(n14199) );
  OAI211_X1 U16170 ( .C1(n14603), .C2(n14326), .A(n14200), .B(n14199), .ZN(
        n14201) );
  AOI21_X1 U16171 ( .B1(n14389), .B2(n15630), .A(n14201), .ZN(n14202) );
  OAI21_X1 U16172 ( .B1(n14203), .B2(n14312), .A(n14202), .ZN(P2_U3244) );
  XNOR2_X1 U16173 ( .A(n14204), .B(n14217), .ZN(n14205) );
  AOI222_X1 U16174 ( .A1(n14207), .A2(n14285), .B1(n14206), .B2(n14286), .C1(
        n14339), .C2(n14205), .ZN(n14395) );
  INV_X1 U16175 ( .A(n14208), .ZN(n14209) );
  AOI211_X1 U16176 ( .C1(n14393), .C2(n14230), .A(n14320), .B(n14209), .ZN(
        n14392) );
  INV_X1 U16177 ( .A(n14393), .ZN(n14212) );
  AOI22_X1 U16178 ( .A1(n14312), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14210), 
        .B2(n14323), .ZN(n14211) );
  OAI21_X1 U16179 ( .B1(n14212), .B2(n14326), .A(n14211), .ZN(n14219) );
  NAND2_X1 U16180 ( .A1(n14213), .A2(n14214), .ZN(n14228) );
  NOR2_X1 U16181 ( .A1(n14228), .A2(n14229), .ZN(n14227) );
  NOR2_X1 U16182 ( .A1(n14227), .A2(n14215), .ZN(n14216) );
  XOR2_X1 U16183 ( .A(n14217), .B(n14216), .Z(n14396) );
  NOR2_X1 U16184 ( .A1(n14396), .A2(n14346), .ZN(n14218) );
  AOI211_X1 U16185 ( .C1(n14392), .C2(n14344), .A(n14219), .B(n14218), .ZN(
        n14220) );
  OAI21_X1 U16186 ( .B1(n14341), .B2(n14395), .A(n14220), .ZN(P2_U3245) );
  INV_X1 U16187 ( .A(n14221), .ZN(n14222) );
  AOI211_X1 U16188 ( .C1(n14224), .C2(n14223), .A(n14288), .B(n14222), .ZN(
        n14226) );
  OR2_X1 U16189 ( .A1(n14226), .A2(n14225), .ZN(n14531) );
  INV_X1 U16190 ( .A(n14531), .ZN(n14239) );
  AOI21_X1 U16191 ( .B1(n14229), .B2(n14228), .A(n14227), .ZN(n14533) );
  INV_X1 U16192 ( .A(n14252), .ZN(n14231) );
  AOI211_X1 U16193 ( .C1(n14232), .C2(n14231), .A(n14320), .B(n7616), .ZN(
        n14532) );
  NAND2_X1 U16194 ( .A1(n14532), .A2(n14344), .ZN(n14236) );
  INV_X1 U16195 ( .A(n14233), .ZN(n14234) );
  AOI22_X1 U16196 ( .A1(n14341), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14234), 
        .B2(n14323), .ZN(n14235) );
  OAI211_X1 U16197 ( .C1(n14608), .C2(n14326), .A(n14236), .B(n14235), .ZN(
        n14237) );
  AOI21_X1 U16198 ( .B1(n14533), .B2(n15630), .A(n14237), .ZN(n14238) );
  OAI21_X1 U16199 ( .B1(n14239), .B2(n14312), .A(n14238), .ZN(P2_U3246) );
  NAND2_X1 U16200 ( .A1(n14241), .A2(n14240), .ZN(n14306) );
  NAND2_X1 U16201 ( .A1(n14306), .A2(n14305), .ZN(n14243) );
  NAND2_X1 U16202 ( .A1(n14243), .A2(n14242), .ZN(n14290) );
  OR2_X1 U16203 ( .A1(n14290), .A2(n14244), .ZN(n14268) );
  AND2_X1 U16204 ( .A1(n14268), .A2(n14245), .ZN(n14248) );
  OAI21_X1 U16205 ( .B1(n14248), .B2(n14247), .A(n14246), .ZN(n14250) );
  AOI21_X1 U16206 ( .B1(n14250), .B2(n14339), .A(n14249), .ZN(n14539) );
  INV_X1 U16207 ( .A(n14251), .ZN(n14253) );
  AOI211_X1 U16208 ( .C1(n14537), .C2(n14253), .A(n14320), .B(n14252), .ZN(
        n14536) );
  INV_X1 U16209 ( .A(n14254), .ZN(n14255) );
  AOI22_X1 U16210 ( .A1(n14341), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14255), 
        .B2(n14323), .ZN(n14256) );
  OAI21_X1 U16211 ( .B1(n14257), .B2(n14326), .A(n14256), .ZN(n14265) );
  INV_X1 U16212 ( .A(n14258), .ZN(n14295) );
  NOR2_X1 U16213 ( .A1(n14295), .A2(n14259), .ZN(n14274) );
  AOI211_X1 U16214 ( .C1(n14274), .C2(n10381), .A(n14261), .B(n14260), .ZN(
        n14263) );
  INV_X1 U16215 ( .A(n14213), .ZN(n14262) );
  NOR2_X1 U16216 ( .A1(n14263), .A2(n14262), .ZN(n14540) );
  NOR2_X1 U16217 ( .A1(n14540), .A2(n14346), .ZN(n14264) );
  AOI211_X1 U16218 ( .C1(n14536), .C2(n14344), .A(n14265), .B(n14264), .ZN(
        n14266) );
  OAI21_X1 U16219 ( .B1(n14341), .B2(n14539), .A(n14266), .ZN(P2_U3247) );
  AND2_X1 U16220 ( .A1(n14268), .A2(n14267), .ZN(n14271) );
  OR2_X1 U16221 ( .A1(n14290), .A2(n14289), .ZN(n14291) );
  NAND3_X1 U16222 ( .A1(n14291), .A2(n10381), .A3(n14269), .ZN(n14270) );
  NAND3_X1 U16223 ( .A1(n14271), .A2(n14339), .A3(n14270), .ZN(n14273) );
  NAND2_X1 U16224 ( .A1(n14273), .A2(n14272), .ZN(n14541) );
  INV_X1 U16225 ( .A(n14541), .ZN(n14282) );
  XNOR2_X1 U16226 ( .A(n14274), .B(n10381), .ZN(n14543) );
  NAND2_X1 U16227 ( .A1(n14543), .A2(n15630), .ZN(n14281) );
  AOI211_X1 U16228 ( .C1(n14275), .C2(n14298), .A(n14320), .B(n14251), .ZN(
        n14542) );
  NOR2_X1 U16229 ( .A1(n7618), .A2(n14326), .ZN(n14279) );
  OAI22_X1 U16230 ( .A1(n15622), .A2(n14277), .B1(n14276), .B2(n15619), .ZN(
        n14278) );
  AOI211_X1 U16231 ( .C1(n14542), .C2(n14344), .A(n14279), .B(n14278), .ZN(
        n14280) );
  OAI211_X1 U16232 ( .C1(n14341), .C2(n14282), .A(n14281), .B(n14280), .ZN(
        P2_U3248) );
  INV_X1 U16233 ( .A(n14283), .ZN(n14294) );
  AOI22_X1 U16234 ( .A1(n14287), .A2(n14286), .B1(n14285), .B2(n14284), .ZN(
        n14547) );
  INV_X1 U16235 ( .A(n14547), .ZN(n14293) );
  AOI21_X1 U16236 ( .B1(n14290), .B2(n14289), .A(n14288), .ZN(n14292) );
  AND2_X1 U16237 ( .A1(n14292), .A2(n14291), .ZN(n14550) );
  AOI211_X1 U16238 ( .C1(n14323), .C2(n14294), .A(n14293), .B(n14550), .ZN(
        n14303) );
  AOI21_X1 U16239 ( .B1(n9523), .B2(n14296), .A(n14295), .ZN(n14551) );
  AOI21_X1 U16240 ( .B1(n14297), .B2(n14546), .A(n14320), .ZN(n14299) );
  NAND2_X1 U16241 ( .A1(n14299), .A2(n14298), .ZN(n14548) );
  AOI22_X1 U16242 ( .A1(n14546), .A2(n15625), .B1(n14341), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n14300) );
  OAI21_X1 U16243 ( .B1(n14548), .B2(n15627), .A(n14300), .ZN(n14301) );
  AOI21_X1 U16244 ( .B1(n14551), .B2(n15630), .A(n14301), .ZN(n14302) );
  OAI21_X1 U16245 ( .B1(n14341), .B2(n14303), .A(n14302), .ZN(P2_U3249) );
  XNOR2_X1 U16246 ( .A(n14304), .B(n14305), .ZN(n14557) );
  INV_X1 U16247 ( .A(n14557), .ZN(n14318) );
  XNOR2_X1 U16248 ( .A(n14306), .B(n14305), .ZN(n14307) );
  NAND2_X1 U16249 ( .A1(n14307), .A2(n14339), .ZN(n14555) );
  INV_X1 U16250 ( .A(n14308), .ZN(n14554) );
  OAI211_X1 U16251 ( .C1(n15619), .C2(n14309), .A(n14555), .B(n14554), .ZN(
        n14316) );
  OAI211_X1 U16252 ( .C1(n14311), .C2(n14617), .A(n14310), .B(n14297), .ZN(
        n14553) );
  AOI22_X1 U16253 ( .A1(n14313), .A2(n15625), .B1(P2_REG2_REG_15__SCAN_IN), 
        .B2(n14312), .ZN(n14314) );
  OAI21_X1 U16254 ( .B1(n14553), .B2(n15627), .A(n14314), .ZN(n14315) );
  AOI21_X1 U16255 ( .B1(n14316), .B2(n15622), .A(n14315), .ZN(n14317) );
  OAI21_X1 U16256 ( .B1(n14318), .B2(n14346), .A(n14317), .ZN(P2_U3250) );
  XNOR2_X1 U16257 ( .A(n14319), .B(n14336), .ZN(n14574) );
  INV_X1 U16258 ( .A(n12733), .ZN(n14321) );
  AOI211_X1 U16259 ( .C1(n14571), .C2(n14321), .A(n14320), .B(n6600), .ZN(
        n14570) );
  INV_X1 U16260 ( .A(n14322), .ZN(n14324) );
  AOI22_X1 U16261 ( .A1(n14312), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n14324), 
        .B2(n14323), .ZN(n14325) );
  OAI21_X1 U16262 ( .B1(n14327), .B2(n14326), .A(n14325), .ZN(n14343) );
  AOI21_X1 U16263 ( .B1(n14628), .B2(n14329), .A(n14328), .ZN(n14337) );
  INV_X1 U16264 ( .A(n14330), .ZN(n14333) );
  INV_X1 U16265 ( .A(n14331), .ZN(n14332) );
  NOR2_X1 U16266 ( .A1(n14333), .A2(n14332), .ZN(n14335) );
  OAI22_X1 U16267 ( .A1(n14337), .A2(n14336), .B1(n14335), .B2(n14334), .ZN(
        n14340) );
  AOI21_X1 U16268 ( .B1(n14340), .B2(n14339), .A(n14338), .ZN(n14573) );
  NOR2_X1 U16269 ( .A1(n14573), .A2(n14341), .ZN(n14342) );
  AOI211_X1 U16270 ( .C1(n14570), .C2(n14344), .A(n14343), .B(n14342), .ZN(
        n14345) );
  OAI21_X1 U16271 ( .B1(n14346), .B2(n14574), .A(n14345), .ZN(P2_U3254) );
  NOR2_X1 U16272 ( .A1(n14348), .A2(n14347), .ZN(n14583) );
  OAI21_X1 U16273 ( .B1(n14585), .B2(n14582), .A(n14350), .ZN(P2_U3529) );
  AOI21_X1 U16274 ( .B1(n15656), .B2(n7611), .A(n14351), .ZN(n14353) );
  NAND2_X1 U16275 ( .A1(n14356), .A2(n15656), .ZN(n14360) );
  NAND3_X1 U16276 ( .A1(n14357), .A2(n14579), .A3(n14103), .ZN(n14359) );
  NAND4_X1 U16277 ( .A1(n14361), .A2(n14360), .A3(n14359), .A4(n14358), .ZN(
        n14586) );
  MUX2_X1 U16278 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14586), .S(n15670), .Z(
        P2_U3526) );
  INV_X1 U16279 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n14365) );
  AOI211_X1 U16280 ( .C1(n14579), .C2(n14364), .A(n14363), .B(n14362), .ZN(
        n14587) );
  MUX2_X1 U16281 ( .A(n14365), .B(n14587), .S(n15670), .Z(n14366) );
  OAI21_X1 U16282 ( .B1(n7629), .B2(n14582), .A(n14366), .ZN(P2_U3525) );
  OAI21_X1 U16283 ( .B1(n7631), .B2(n15648), .A(n14367), .ZN(n14368) );
  AOI21_X1 U16284 ( .B1(n14369), .B2(n14579), .A(n14368), .ZN(n14370) );
  NAND2_X1 U16285 ( .A1(n14371), .A2(n14370), .ZN(n14590) );
  MUX2_X1 U16286 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14590), .S(n15670), .Z(
        P2_U3524) );
  AOI211_X1 U16287 ( .C1(n14374), .C2(n14579), .A(n14373), .B(n14372), .ZN(
        n14591) );
  MUX2_X1 U16288 ( .A(n14375), .B(n14591), .S(n15670), .Z(n14376) );
  OAI21_X1 U16289 ( .B1(n14594), .B2(n14582), .A(n14376), .ZN(P2_U3523) );
  AOI21_X1 U16290 ( .B1(n15656), .B2(n14378), .A(n14377), .ZN(n14379) );
  OAI211_X1 U16291 ( .C1(n14575), .C2(n14381), .A(n14380), .B(n14379), .ZN(
        n14595) );
  MUX2_X1 U16292 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14595), .S(n15670), .Z(
        P2_U3522) );
  AOI211_X1 U16293 ( .C1(n14579), .C2(n14384), .A(n14383), .B(n14382), .ZN(
        n14596) );
  MUX2_X1 U16294 ( .A(n14385), .B(n14596), .S(n15670), .Z(n14386) );
  OAI21_X1 U16295 ( .B1(n14599), .B2(n14582), .A(n14386), .ZN(P2_U3521) );
  AOI211_X1 U16296 ( .C1(n14579), .C2(n14389), .A(n14388), .B(n14387), .ZN(
        n14600) );
  MUX2_X1 U16297 ( .A(n14390), .B(n14600), .S(n15670), .Z(n14391) );
  OAI21_X1 U16298 ( .B1(n14603), .B2(n14582), .A(n14391), .ZN(P2_U3520) );
  AOI21_X1 U16299 ( .B1(n15656), .B2(n14393), .A(n14392), .ZN(n14394) );
  OAI211_X1 U16300 ( .C1(n14575), .C2(n14396), .A(n14395), .B(n14394), .ZN(
        n14604) );
  MUX2_X1 U16301 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14604), .S(n15670), .Z(
        n14530) );
  OR4_X1 U16302 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(P1_REG1_REG_23__SCAN_IN), 
        .A3(P1_REG2_REG_26__SCAN_IN), .A4(P3_D_REG_1__SCAN_IN), .ZN(n14408) );
  NAND3_X1 U16303 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .A3(
        n14433), .ZN(n14407) );
  NAND4_X1 U16304 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P3_DATAO_REG_27__SCAN_IN), 
        .A3(n14558), .A4(n14702), .ZN(n14406) );
  NAND4_X1 U16305 ( .A1(P2_REG2_REG_26__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), 
        .A3(P1_IR_REG_24__SCAN_IN), .A4(n8964), .ZN(n14398) );
  NAND3_X1 U16306 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n14453), .A3(n10067), 
        .ZN(n14397) );
  NOR2_X1 U16307 ( .A1(n14398), .A2(n14397), .ZN(n14400) );
  INV_X1 U16308 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14451) );
  NOR3_X1 U16309 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P1_DATAO_REG_29__SCAN_IN), 
        .A3(P1_REG1_REG_19__SCAN_IN), .ZN(n14399) );
  NAND4_X1 U16310 ( .A1(n14401), .A2(n14400), .A3(n14451), .A4(n14399), .ZN(
        n14403) );
  NOR3_X1 U16311 ( .A1(n14403), .A2(n14461), .A3(n14402), .ZN(n14404) );
  NAND3_X1 U16312 ( .A1(n14404), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .ZN(n14405) );
  OR4_X1 U16313 ( .A1(n14408), .A2(n14407), .A3(n14406), .A4(n14405), .ZN(
        n14424) );
  NOR4_X1 U16314 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_REG1_REG_2__SCAN_IN), 
        .A3(P3_REG0_REG_10__SCAN_IN), .A4(n14409), .ZN(n14410) );
  NAND4_X1 U16315 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14411), .A3(n14410), 
        .A4(n14872), .ZN(n14423) );
  OR4_X1 U16316 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_REG1_REG_11__SCAN_IN), .A4(P1_REG2_REG_6__SCAN_IN), .ZN(n14422) );
  NOR4_X1 U16317 ( .A1(n14645), .A2(n14413), .A3(n14412), .A4(
        P2_REG3_REG_0__SCAN_IN), .ZN(n14420) );
  INV_X1 U16318 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n14415) );
  NOR4_X1 U16319 ( .A1(n14485), .A2(n14415), .A3(n14414), .A4(
        P3_REG1_REG_3__SCAN_IN), .ZN(n14419) );
  NOR4_X1 U16320 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .A3(
        SI_29_), .A4(P2_DATAO_REG_31__SCAN_IN), .ZN(n14418) );
  NOR4_X1 U16321 ( .A1(n14416), .A2(n9588), .A3(P1_REG0_REG_10__SCAN_IN), .A4(
        P1_REG3_REG_26__SCAN_IN), .ZN(n14417) );
  NAND4_X1 U16322 ( .A1(n14420), .A2(n14419), .A3(n14418), .A4(n14417), .ZN(
        n14421) );
  NOR4_X1 U16323 ( .A1(n14424), .A2(n14423), .A3(n14422), .A4(n14421), .ZN(
        n14428) );
  NAND3_X1 U16324 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .A3(P3_DATAO_REG_4__SCAN_IN), .ZN(n14426) );
  NAND3_X1 U16325 ( .A1(P3_REG0_REG_16__SCAN_IN), .A2(P3_DATAO_REG_25__SCAN_IN), .A3(n14444), .ZN(n14425) );
  NOR4_X1 U16326 ( .A1(P2_REG0_REG_10__SCAN_IN), .A2(P3_REG0_REG_3__SCAN_IN), 
        .A3(n14426), .A4(n14425), .ZN(n14427) );
  AOI21_X1 U16327 ( .B1(n14428), .B2(n14427), .A(keyinput42), .ZN(n14429) );
  MUX2_X1 U16328 ( .A(n14429), .B(keyinput42), .S(P3_ADDR_REG_19__SCAN_IN), 
        .Z(n14528) );
  INV_X1 U16329 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15638) );
  INV_X1 U16330 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15534) );
  AOI22_X1 U16331 ( .A1(n15638), .A2(keyinput28), .B1(keyinput55), .B2(n15534), 
        .ZN(n14430) );
  OAI221_X1 U16332 ( .B1(n15638), .B2(keyinput28), .C1(n15534), .C2(keyinput55), .A(n14430), .ZN(n14441) );
  AOI22_X1 U16333 ( .A1(n14433), .A2(keyinput53), .B1(keyinput20), .B2(n14432), 
        .ZN(n14431) );
  OAI221_X1 U16334 ( .B1(n14433), .B2(keyinput53), .C1(n14432), .C2(keyinput20), .A(n14431), .ZN(n14440) );
  AOI22_X1 U16335 ( .A1(n14889), .A2(keyinput40), .B1(n14435), .B2(keyinput30), 
        .ZN(n14434) );
  OAI221_X1 U16336 ( .B1(n14889), .B2(keyinput40), .C1(n14435), .C2(keyinput30), .A(n14434), .ZN(n14439) );
  INV_X1 U16337 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n15636) );
  AOI22_X1 U16338 ( .A1(n14437), .A2(keyinput52), .B1(n15636), .B2(keyinput29), 
        .ZN(n14436) );
  OAI221_X1 U16339 ( .B1(n14437), .B2(keyinput52), .C1(n15636), .C2(keyinput29), .A(n14436), .ZN(n14438) );
  NOR4_X1 U16340 ( .A1(n14441), .A2(n14440), .A3(n14439), .A4(n14438), .ZN(
        n14527) );
  INV_X1 U16341 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15536) );
  INV_X1 U16342 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15635) );
  AOI22_X1 U16343 ( .A1(n15536), .A2(keyinput59), .B1(n15635), .B2(keyinput10), 
        .ZN(n14442) );
  OAI221_X1 U16344 ( .B1(n15536), .B2(keyinput59), .C1(n15635), .C2(keyinput10), .A(n14442), .ZN(n14448) );
  AOI22_X1 U16345 ( .A1(n14625), .A2(keyinput35), .B1(n14444), .B2(keyinput60), 
        .ZN(n14443) );
  OAI221_X1 U16346 ( .B1(n14625), .B2(keyinput35), .C1(n14444), .C2(keyinput60), .A(n14443), .ZN(n14447) );
  XNOR2_X1 U16347 ( .A(keyinput15), .B(n8139), .ZN(n14446) );
  XNOR2_X1 U16348 ( .A(keyinput27), .B(n14413), .ZN(n14445) );
  OR4_X1 U16349 ( .A1(n14448), .A2(n14447), .A3(n14446), .A4(n14445), .ZN(
        n14457) );
  AOI22_X1 U16350 ( .A1(n14702), .A2(keyinput7), .B1(n14558), .B2(keyinput9), 
        .ZN(n14449) );
  OAI221_X1 U16351 ( .B1(n14702), .B2(keyinput7), .C1(n14558), .C2(keyinput9), 
        .A(n14449), .ZN(n14456) );
  AOI22_X1 U16352 ( .A1(n14645), .A2(keyinput33), .B1(keyinput12), .B2(n14451), 
        .ZN(n14450) );
  OAI221_X1 U16353 ( .B1(n14645), .B2(keyinput33), .C1(n14451), .C2(keyinput12), .A(n14450), .ZN(n14455) );
  AOI22_X1 U16354 ( .A1(n10067), .A2(keyinput54), .B1(n14453), .B2(keyinput62), 
        .ZN(n14452) );
  OAI221_X1 U16355 ( .B1(n10067), .B2(keyinput54), .C1(n14453), .C2(keyinput62), .A(n14452), .ZN(n14454) );
  OR4_X1 U16356 ( .A1(n14457), .A2(n14456), .A3(n14455), .A4(n14454), .ZN(
        n14466) );
  AOI22_X1 U16357 ( .A1(n14459), .A2(keyinput22), .B1(n9727), .B2(keyinput37), 
        .ZN(n14458) );
  OAI221_X1 U16358 ( .B1(n14459), .B2(keyinput22), .C1(n9727), .C2(keyinput37), 
        .A(n14458), .ZN(n14465) );
  INV_X1 U16359 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n14462) );
  AOI22_X1 U16360 ( .A1(n14462), .A2(keyinput46), .B1(n14461), .B2(keyinput16), 
        .ZN(n14460) );
  OAI221_X1 U16361 ( .B1(n14462), .B2(keyinput46), .C1(n14461), .C2(keyinput16), .A(n14460), .ZN(n14464) );
  INV_X1 U16362 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15537) );
  XNOR2_X1 U16363 ( .A(n15537), .B(keyinput56), .ZN(n14463) );
  NOR4_X1 U16364 ( .A1(n14466), .A2(n14465), .A3(n14464), .A4(n14463), .ZN(
        n14526) );
  AOI22_X1 U16365 ( .A1(n14469), .A2(keyinput48), .B1(keyinput6), .B2(n14468), 
        .ZN(n14467) );
  OAI221_X1 U16366 ( .B1(n14469), .B2(keyinput48), .C1(n14468), .C2(keyinput6), 
        .A(n14467), .ZN(n14479) );
  AOI22_X1 U16367 ( .A1(n14471), .A2(keyinput45), .B1(n14872), .B2(keyinput26), 
        .ZN(n14470) );
  OAI221_X1 U16368 ( .B1(n14471), .B2(keyinput45), .C1(n14872), .C2(keyinput26), .A(n14470), .ZN(n14478) );
  AOI22_X1 U16369 ( .A1(n9623), .A2(keyinput61), .B1(n14473), .B2(keyinput39), 
        .ZN(n14472) );
  OAI221_X1 U16370 ( .B1(n9623), .B2(keyinput61), .C1(n14473), .C2(keyinput39), 
        .A(n14472), .ZN(n14477) );
  AOI22_X1 U16371 ( .A1(n14475), .A2(keyinput38), .B1(n14638), .B2(keyinput47), 
        .ZN(n14474) );
  OAI221_X1 U16372 ( .B1(n14475), .B2(keyinput38), .C1(n14638), .C2(keyinput47), .A(n14474), .ZN(n14476) );
  OR4_X1 U16373 ( .A1(n14479), .A2(n14478), .A3(n14477), .A4(n14476), .ZN(
        n14489) );
  AOI22_X1 U16374 ( .A1(n8573), .A2(keyinput63), .B1(keyinput50), .B2(n8971), 
        .ZN(n14480) );
  OAI221_X1 U16375 ( .B1(n8573), .B2(keyinput63), .C1(n8971), .C2(keyinput50), 
        .A(n14480), .ZN(n14488) );
  AOI22_X1 U16376 ( .A1(n14483), .A2(keyinput36), .B1(n14482), .B2(keyinput25), 
        .ZN(n14481) );
  OAI221_X1 U16377 ( .B1(n14483), .B2(keyinput36), .C1(n14482), .C2(keyinput25), .A(n14481), .ZN(n14487) );
  INV_X1 U16378 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15535) );
  AOI22_X1 U16379 ( .A1(n15535), .A2(keyinput31), .B1(n14485), .B2(keyinput43), 
        .ZN(n14484) );
  OAI221_X1 U16380 ( .B1(n15535), .B2(keyinput31), .C1(n14485), .C2(keyinput43), .A(n14484), .ZN(n14486) );
  NOR4_X1 U16381 ( .A1(n14489), .A2(n14488), .A3(n14487), .A4(n14486), .ZN(
        n14524) );
  AOI22_X1 U16382 ( .A1(n10800), .A2(keyinput11), .B1(n14491), .B2(keyinput2), 
        .ZN(n14490) );
  OAI221_X1 U16383 ( .B1(n10800), .B2(keyinput11), .C1(n14491), .C2(keyinput2), 
        .A(n14490), .ZN(n14497) );
  XNOR2_X1 U16384 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput51), .ZN(n14495) );
  XNOR2_X1 U16385 ( .A(P1_REG0_REG_21__SCAN_IN), .B(keyinput4), .ZN(n14494) );
  XNOR2_X1 U16386 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput19), .ZN(n14493) );
  XNOR2_X1 U16387 ( .A(P1_REG2_REG_17__SCAN_IN), .B(keyinput17), .ZN(n14492)
         );
  NAND4_X1 U16388 ( .A1(n14495), .A2(n14494), .A3(n14493), .A4(n14492), .ZN(
        n14496) );
  NOR2_X1 U16389 ( .A1(n14497), .A2(n14496), .ZN(n14523) );
  XNOR2_X1 U16390 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput14), .ZN(n14501)
         );
  XNOR2_X1 U16391 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput34), .ZN(n14500) );
  XNOR2_X1 U16392 ( .A(SI_7_), .B(keyinput49), .ZN(n14499) );
  XNOR2_X1 U16393 ( .A(P1_REG1_REG_23__SCAN_IN), .B(keyinput41), .ZN(n14498)
         );
  NAND4_X1 U16394 ( .A1(n14501), .A2(n14500), .A3(n14499), .A4(n14498), .ZN(
        n14507) );
  XNOR2_X1 U16395 ( .A(SI_10_), .B(keyinput44), .ZN(n14505) );
  XNOR2_X1 U16396 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput23), .ZN(n14504) );
  XNOR2_X1 U16397 ( .A(SI_27_), .B(keyinput32), .ZN(n14503) );
  XNOR2_X1 U16398 ( .A(P3_IR_REG_15__SCAN_IN), .B(keyinput21), .ZN(n14502) );
  NAND4_X1 U16399 ( .A1(n14505), .A2(n14504), .A3(n14503), .A4(n14502), .ZN(
        n14506) );
  NOR2_X1 U16400 ( .A1(n14507), .A2(n14506), .ZN(n14522) );
  AOI22_X1 U16401 ( .A1(n9248), .A2(keyinput18), .B1(keyinput24), .B2(n8964), 
        .ZN(n14508) );
  OAI221_X1 U16402 ( .B1(n9248), .B2(keyinput18), .C1(n8964), .C2(keyinput24), 
        .A(n14508), .ZN(n14520) );
  XNOR2_X1 U16403 ( .A(P3_REG1_REG_3__SCAN_IN), .B(keyinput8), .ZN(n14512) );
  XNOR2_X1 U16404 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput13), .ZN(n14511) );
  XNOR2_X1 U16405 ( .A(P3_D_REG_0__SCAN_IN), .B(keyinput3), .ZN(n14510) );
  XNOR2_X1 U16406 ( .A(P1_REG3_REG_26__SCAN_IN), .B(keyinput5), .ZN(n14509) );
  AND4_X1 U16407 ( .A1(n14512), .A2(n14511), .A3(n14510), .A4(n14509), .ZN(
        n14518) );
  XNOR2_X1 U16408 ( .A(keyinput58), .B(n15057), .ZN(n14514) );
  XNOR2_X1 U16409 ( .A(keyinput57), .B(n9588), .ZN(n14513) );
  NOR2_X1 U16410 ( .A1(n14514), .A2(n14513), .ZN(n14517) );
  XNOR2_X1 U16411 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput0), .ZN(n14516) );
  XNOR2_X1 U16412 ( .A(P3_IR_REG_6__SCAN_IN), .B(keyinput1), .ZN(n14515) );
  NAND4_X1 U16413 ( .A1(n14518), .A2(n14517), .A3(n14516), .A4(n14515), .ZN(
        n14519) );
  NOR2_X1 U16414 ( .A1(n14520), .A2(n14519), .ZN(n14521) );
  AND4_X1 U16415 ( .A1(n14524), .A2(n14523), .A3(n14522), .A4(n14521), .ZN(
        n14525) );
  NAND4_X1 U16416 ( .A1(n14528), .A2(n14527), .A3(n14526), .A4(n14525), .ZN(
        n14529) );
  XNOR2_X1 U16417 ( .A(n14530), .B(n14529), .ZN(P2_U3519) );
  AOI211_X1 U16418 ( .C1(n14533), .C2(n14579), .A(n14532), .B(n14531), .ZN(
        n14605) );
  MUX2_X1 U16419 ( .A(n14534), .B(n14605), .S(n15670), .Z(n14535) );
  OAI21_X1 U16420 ( .B1(n14608), .B2(n14582), .A(n14535), .ZN(P2_U3518) );
  AOI21_X1 U16421 ( .B1(n15656), .B2(n14537), .A(n14536), .ZN(n14538) );
  OAI211_X1 U16422 ( .C1(n14540), .C2(n14575), .A(n14539), .B(n14538), .ZN(
        n14609) );
  MUX2_X1 U16423 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14609), .S(n15670), .Z(
        P2_U3517) );
  INV_X1 U16424 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14544) );
  AOI211_X1 U16425 ( .C1(n14543), .C2(n14579), .A(n14542), .B(n14541), .ZN(
        n14610) );
  MUX2_X1 U16426 ( .A(n14544), .B(n14610), .S(n15670), .Z(n14545) );
  OAI21_X1 U16427 ( .B1(n7618), .B2(n14582), .A(n14545), .ZN(P2_U3516) );
  OAI211_X1 U16428 ( .C1(n6792), .C2(n15648), .A(n14548), .B(n14547), .ZN(
        n14549) );
  AOI211_X1 U16429 ( .C1(n14551), .C2(n14579), .A(n14550), .B(n14549), .ZN(
        n14552) );
  INV_X1 U16430 ( .A(n14552), .ZN(n14613) );
  MUX2_X1 U16431 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14613), .S(n15670), .Z(
        P2_U3515) );
  NAND3_X1 U16432 ( .A1(n14555), .A2(n14554), .A3(n14553), .ZN(n14556) );
  AOI21_X1 U16433 ( .B1(n14557), .B2(n14579), .A(n14556), .ZN(n14614) );
  MUX2_X1 U16434 ( .A(n14558), .B(n14614), .S(n15670), .Z(n14559) );
  OAI21_X1 U16435 ( .B1(n14617), .B2(n14582), .A(n14559), .ZN(P2_U3514) );
  AOI211_X1 U16436 ( .C1(n15656), .C2(n14562), .A(n14561), .B(n14560), .ZN(
        n14563) );
  OAI21_X1 U16437 ( .B1(n14575), .B2(n14564), .A(n14563), .ZN(n14618) );
  MUX2_X1 U16438 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14618), .S(n15670), .Z(
        P2_U3513) );
  INV_X1 U16439 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14568) );
  AOI211_X1 U16440 ( .C1(n14567), .C2(n14579), .A(n14566), .B(n14565), .ZN(
        n14619) );
  MUX2_X1 U16441 ( .A(n14568), .B(n14619), .S(n15670), .Z(n14569) );
  OAI21_X1 U16442 ( .B1(n14622), .B2(n14582), .A(n14569), .ZN(P2_U3512) );
  AOI21_X1 U16443 ( .B1(n15656), .B2(n14571), .A(n14570), .ZN(n14572) );
  OAI211_X1 U16444 ( .C1(n14575), .C2(n14574), .A(n14573), .B(n14572), .ZN(
        n14623) );
  MUX2_X1 U16445 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n14623), .S(n15670), .Z(
        P2_U3510) );
  INV_X1 U16446 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n14580) );
  AOI211_X1 U16447 ( .C1(n14579), .C2(n14578), .A(n14577), .B(n14576), .ZN(
        n14624) );
  MUX2_X1 U16448 ( .A(n14580), .B(n14624), .S(n15670), .Z(n14581) );
  OAI21_X1 U16449 ( .B1(n14628), .B2(n14582), .A(n14581), .ZN(P2_U3509) );
  OAI21_X1 U16450 ( .B1(n14585), .B2(n14627), .A(n14584), .ZN(P2_U3497) );
  MUX2_X1 U16451 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14586), .S(n15666), .Z(
        P2_U3494) );
  INV_X1 U16452 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n14588) );
  MUX2_X1 U16453 ( .A(n14588), .B(n14587), .S(n15666), .Z(n14589) );
  OAI21_X1 U16454 ( .B1(n7629), .B2(n14627), .A(n14589), .ZN(P2_U3493) );
  MUX2_X1 U16455 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14590), .S(n15666), .Z(
        P2_U3492) );
  INV_X1 U16456 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n14592) );
  MUX2_X1 U16457 ( .A(n14592), .B(n14591), .S(n15666), .Z(n14593) );
  OAI21_X1 U16458 ( .B1(n14594), .B2(n14627), .A(n14593), .ZN(P2_U3491) );
  MUX2_X1 U16459 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14595), .S(n15666), .Z(
        P2_U3490) );
  INV_X1 U16460 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14597) );
  MUX2_X1 U16461 ( .A(n14597), .B(n14596), .S(n15666), .Z(n14598) );
  OAI21_X1 U16462 ( .B1(n14599), .B2(n14627), .A(n14598), .ZN(P2_U3489) );
  INV_X1 U16463 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n14601) );
  MUX2_X1 U16464 ( .A(n14601), .B(n14600), .S(n15666), .Z(n14602) );
  OAI21_X1 U16465 ( .B1(n14603), .B2(n14627), .A(n14602), .ZN(P2_U3488) );
  MUX2_X1 U16466 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14604), .S(n15666), .Z(
        P2_U3487) );
  INV_X1 U16467 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14606) );
  MUX2_X1 U16468 ( .A(n14606), .B(n14605), .S(n15666), .Z(n14607) );
  OAI21_X1 U16469 ( .B1(n14608), .B2(n14627), .A(n14607), .ZN(P2_U3486) );
  MUX2_X1 U16470 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14609), .S(n15666), .Z(
        P2_U3484) );
  INV_X1 U16471 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14611) );
  MUX2_X1 U16472 ( .A(n14611), .B(n14610), .S(n15666), .Z(n14612) );
  OAI21_X1 U16473 ( .B1(n7618), .B2(n14627), .A(n14612), .ZN(P2_U3481) );
  MUX2_X1 U16474 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14613), .S(n15666), .Z(
        P2_U3478) );
  INV_X1 U16475 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14615) );
  MUX2_X1 U16476 ( .A(n14615), .B(n14614), .S(n15666), .Z(n14616) );
  OAI21_X1 U16477 ( .B1(n14617), .B2(n14627), .A(n14616), .ZN(P2_U3475) );
  MUX2_X1 U16478 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n14618), .S(n15666), .Z(
        P2_U3472) );
  INV_X1 U16479 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14620) );
  MUX2_X1 U16480 ( .A(n14620), .B(n14619), .S(n15666), .Z(n14621) );
  OAI21_X1 U16481 ( .B1(n14622), .B2(n14627), .A(n14621), .ZN(P2_U3469) );
  MUX2_X1 U16482 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n14623), .S(n15666), .Z(
        P2_U3463) );
  MUX2_X1 U16483 ( .A(n14625), .B(n14624), .S(n15666), .Z(n14626) );
  OAI21_X1 U16484 ( .B1(n14628), .B2(n14627), .A(n14626), .ZN(P2_U3460) );
  INV_X1 U16485 ( .A(n10639), .ZN(n15427) );
  INV_X1 U16486 ( .A(n14629), .ZN(n14631) );
  NOR4_X1 U16487 ( .A1(n14631), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14630), .A4(
        P2_U3088), .ZN(n14632) );
  AOI21_X1 U16488 ( .B1(n14640), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14632), 
        .ZN(n14633) );
  OAI21_X1 U16489 ( .B1(n15427), .B2(n14637), .A(n14633), .ZN(P2_U3296) );
  INV_X1 U16490 ( .A(n14634), .ZN(n15430) );
  OAI222_X1 U16491 ( .A1(n14646), .A2(n14638), .B1(n14637), .B2(n15430), .C1(
        P2_U3088), .C2(n14635), .ZN(P2_U3298) );
  AOI21_X1 U16492 ( .B1(n14640), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14639), 
        .ZN(n14641) );
  OAI21_X1 U16493 ( .B1(n14642), .B2(n14644), .A(n14641), .ZN(P2_U3299) );
  INV_X1 U16494 ( .A(n14643), .ZN(n15432) );
  OAI222_X1 U16495 ( .A1(P2_U3088), .A2(n14647), .B1(n14646), .B2(n14645), 
        .C1(n14644), .C2(n15432), .ZN(P2_U3300) );
  MUX2_X1 U16496 ( .A(n14648), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI21_X1 U16497 ( .B1(n14650), .B2(n6469), .A(n14649), .ZN(n14651) );
  NAND2_X1 U16498 ( .A1(n14651), .A2(n14754), .ZN(n14657) );
  OAI21_X1 U16499 ( .B1(n14778), .B2(n14653), .A(n14652), .ZN(n14654) );
  AOI21_X1 U16500 ( .B1(n14655), .B2(n14776), .A(n14654), .ZN(n14656) );
  OAI211_X1 U16501 ( .C1(n7762), .C2(n14763), .A(n14657), .B(n14656), .ZN(
        P1_U3215) );
  XOR2_X1 U16502 ( .A(n14659), .B(n14658), .Z(n14663) );
  AOI22_X1 U16503 ( .A1(n15258), .A2(n14802), .B1(n14803), .B2(n15257), .ZN(
        n15107) );
  AOI22_X1 U16504 ( .A1(n15114), .A2(n14776), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14660) );
  OAI21_X1 U16505 ( .B1(n15107), .B2(n14778), .A(n14660), .ZN(n14661) );
  AOI21_X1 U16506 ( .B1(n15113), .B2(n14795), .A(n14661), .ZN(n14662) );
  OAI21_X1 U16507 ( .B1(n14663), .B2(n14797), .A(n14662), .ZN(P1_U3216) );
  OAI21_X1 U16508 ( .B1(n14665), .B2(n12517), .A(n14664), .ZN(n14669) );
  XNOR2_X1 U16509 ( .A(n14667), .B(n14666), .ZN(n14668) );
  XNOR2_X1 U16510 ( .A(n14669), .B(n14668), .ZN(n14670) );
  NAND2_X1 U16511 ( .A1(n14670), .A2(n14754), .ZN(n14679) );
  NAND2_X1 U16512 ( .A1(n14766), .A2(n14671), .ZN(n14672) );
  NAND2_X1 U16513 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n14921)
         );
  NAND2_X1 U16514 ( .A1(n14672), .A2(n14921), .ZN(n14673) );
  AOI21_X1 U16515 ( .B1(n14727), .B2(n14813), .A(n14673), .ZN(n14678) );
  NAND2_X1 U16516 ( .A1(n14795), .A2(n14674), .ZN(n14677) );
  NAND2_X1 U16517 ( .A1(n14776), .A2(n14675), .ZN(n14676) );
  NAND4_X1 U16518 ( .A1(n14679), .A2(n14678), .A3(n14677), .A4(n14676), .ZN(
        P1_U3217) );
  OAI211_X1 U16519 ( .C1(n14682), .C2(n14681), .A(n14680), .B(n14754), .ZN(
        n14687) );
  INV_X1 U16520 ( .A(n15181), .ZN(n14685) );
  AND2_X1 U16521 ( .A1(n14806), .A2(n15257), .ZN(n14683) );
  AOI21_X1 U16522 ( .B1(n14804), .B2(n15258), .A(n14683), .ZN(n15329) );
  NAND2_X1 U16523 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14996)
         );
  OAI21_X1 U16524 ( .B1(n15329), .B2(n14778), .A(n14996), .ZN(n14684) );
  AOI21_X1 U16525 ( .B1(n14685), .B2(n14776), .A(n14684), .ZN(n14686) );
  OAI211_X1 U16526 ( .C1(n15186), .C2(n14763), .A(n14687), .B(n14686), .ZN(
        P1_U3219) );
  NAND2_X1 U16527 ( .A1(n15151), .A2(n15547), .ZN(n15323) );
  INV_X1 U16528 ( .A(n14771), .ZN(n14698) );
  OAI21_X1 U16529 ( .B1(n14689), .B2(n6543), .A(n14688), .ZN(n14690) );
  NAND2_X1 U16530 ( .A1(n14690), .A2(n14754), .ZN(n14697) );
  OR2_X1 U16531 ( .A1(n14691), .A2(n15241), .ZN(n14693) );
  NAND2_X1 U16532 ( .A1(n14804), .A2(n15257), .ZN(n14692) );
  NAND2_X1 U16533 ( .A1(n14693), .A2(n14692), .ZN(n15142) );
  OAI22_X1 U16534 ( .A1(n14792), .A2(n15149), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14694), .ZN(n14695) );
  AOI21_X1 U16535 ( .B1(n15142), .B2(n14766), .A(n14695), .ZN(n14696) );
  OAI211_X1 U16536 ( .C1(n15323), .C2(n14698), .A(n14697), .B(n14696), .ZN(
        P1_U3223) );
  XOR2_X1 U16537 ( .A(n14700), .B(n14699), .Z(n14706) );
  AND2_X1 U16538 ( .A1(n14802), .A2(n15257), .ZN(n14701) );
  AOI21_X1 U16539 ( .B1(n15037), .B2(n15258), .A(n14701), .ZN(n15300) );
  NOR2_X1 U16540 ( .A1(n15300), .A2(n14778), .ZN(n14704) );
  OAI22_X1 U16541 ( .A1(n15078), .A2(n14792), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14702), .ZN(n14703) );
  AOI211_X1 U16542 ( .C1(n15298), .C2(n14795), .A(n14704), .B(n14703), .ZN(
        n14705) );
  OAI21_X1 U16543 ( .B1(n14706), .B2(n14797), .A(n14705), .ZN(P1_U3225) );
  XOR2_X1 U16544 ( .A(n14708), .B(n14707), .Z(n14713) );
  INV_X1 U16545 ( .A(n14709), .ZN(n15243) );
  AOI22_X1 U16546 ( .A1(n14748), .A2(n14807), .B1(n14776), .B2(n15243), .ZN(
        n14710) );
  NAND2_X1 U16547 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14947)
         );
  OAI211_X1 U16548 ( .C1(n15240), .C2(n14789), .A(n14710), .B(n14947), .ZN(
        n14711) );
  AOI21_X1 U16549 ( .B1(n15351), .B2(n14795), .A(n14711), .ZN(n14712) );
  OAI21_X1 U16550 ( .B1(n14713), .B2(n14797), .A(n14712), .ZN(P1_U3226) );
  XOR2_X1 U16551 ( .A(n14714), .B(n14715), .Z(n14720) );
  NOR2_X1 U16552 ( .A1(n14792), .A2(n15216), .ZN(n14718) );
  AND2_X1 U16553 ( .A1(n15259), .A2(n15257), .ZN(n14716) );
  AOI21_X1 U16554 ( .B1(n14806), .B2(n15258), .A(n14716), .ZN(n15342) );
  NAND2_X1 U16555 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14958)
         );
  OAI21_X1 U16556 ( .B1(n15342), .B2(n14778), .A(n14958), .ZN(n14717) );
  AOI211_X1 U16557 ( .C1(n15345), .C2(n14795), .A(n14718), .B(n14717), .ZN(
        n14719) );
  OAI21_X1 U16558 ( .B1(n14720), .B2(n14797), .A(n14719), .ZN(P1_U3228) );
  XOR2_X1 U16559 ( .A(n14722), .B(n14721), .Z(n14730) );
  OAI22_X1 U16560 ( .A1(n15100), .A2(n14792), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14723), .ZN(n14726) );
  NOR2_X1 U16561 ( .A1(n14724), .A2(n14790), .ZN(n14725) );
  AOI211_X1 U16562 ( .C1(n14727), .C2(n15089), .A(n14726), .B(n14725), .ZN(
        n14729) );
  NAND2_X1 U16563 ( .A1(n15099), .A2(n14795), .ZN(n14728) );
  OAI211_X1 U16564 ( .C1(n14730), .C2(n14797), .A(n14729), .B(n14728), .ZN(
        P1_U3229) );
  INV_X1 U16565 ( .A(n14731), .ZN(n14732) );
  OAI211_X1 U16566 ( .C1(n14734), .C2(n14733), .A(n14732), .B(n14754), .ZN(
        n14739) );
  OAI22_X1 U16567 ( .A1(n14756), .A2(n15241), .B1(n14735), .B2(n15239), .ZN(
        n15164) );
  OAI22_X1 U16568 ( .A1(n14792), .A2(n15169), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14736), .ZN(n14737) );
  AOI21_X1 U16569 ( .B1(n15164), .B2(n14766), .A(n14737), .ZN(n14738) );
  OAI211_X1 U16570 ( .C1(n15328), .C2(n14763), .A(n14739), .B(n14738), .ZN(
        P1_U3233) );
  OAI211_X1 U16571 ( .C1(n14742), .C2(n14741), .A(n14740), .B(n14754), .ZN(
        n14750) );
  INV_X1 U16572 ( .A(n14743), .ZN(n14747) );
  OAI22_X1 U16573 ( .A1(n14745), .A2(n14789), .B1(n14792), .B2(n14744), .ZN(
        n14746) );
  AOI211_X1 U16574 ( .C1(n14748), .C2(n15256), .A(n14747), .B(n14746), .ZN(
        n14749) );
  OAI211_X1 U16575 ( .C1(n15421), .C2(n14763), .A(n14750), .B(n14749), .ZN(
        P1_U3234) );
  OAI21_X1 U16576 ( .B1(n14753), .B2(n14752), .A(n14751), .ZN(n14755) );
  NAND2_X1 U16577 ( .A1(n14755), .A2(n14754), .ZN(n14762) );
  OAI22_X1 U16578 ( .A1(n14757), .A2(n15241), .B1(n14756), .B2(n15239), .ZN(
        n15126) );
  INV_X1 U16579 ( .A(n15133), .ZN(n14759) );
  OAI22_X1 U16580 ( .A1(n14759), .A2(n14792), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14758), .ZN(n14760) );
  AOI21_X1 U16581 ( .B1(n15126), .B2(n14766), .A(n14760), .ZN(n14761) );
  OAI211_X1 U16582 ( .C1(n14763), .C2(n15404), .A(n14762), .B(n14761), .ZN(
        P1_U3235) );
  XOR2_X1 U16583 ( .A(n14765), .B(n14764), .Z(n14773) );
  AND2_X1 U16584 ( .A1(n15199), .A2(n15547), .ZN(n15336) );
  INV_X1 U16585 ( .A(n15200), .ZN(n14769) );
  NAND2_X1 U16586 ( .A1(n14805), .A2(n15258), .ZN(n15196) );
  NAND2_X1 U16587 ( .A1(n14807), .A2(n15257), .ZN(n15194) );
  NAND2_X1 U16588 ( .A1(n15196), .A2(n15194), .ZN(n14767) );
  NAND2_X1 U16589 ( .A1(n14767), .A2(n14766), .ZN(n14768) );
  NAND2_X1 U16590 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14973)
         );
  OAI211_X1 U16591 ( .C1(n14792), .C2(n14769), .A(n14768), .B(n14973), .ZN(
        n14770) );
  AOI21_X1 U16592 ( .B1(n15336), .B2(n14771), .A(n14770), .ZN(n14772) );
  OAI21_X1 U16593 ( .B1(n14773), .B2(n14797), .A(n14772), .ZN(P1_U3238) );
  AND2_X1 U16594 ( .A1(n15090), .A2(n15257), .ZN(n14775) );
  AOI21_X1 U16595 ( .B1(n14801), .B2(n15258), .A(n14775), .ZN(n15292) );
  AOI22_X1 U16596 ( .A1(n15052), .A2(n14776), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14777) );
  OAI21_X1 U16597 ( .B1(n15292), .B2(n14778), .A(n14777), .ZN(n14779) );
  AOI21_X1 U16598 ( .B1(n15053), .B2(n14795), .A(n14779), .ZN(n14780) );
  OAI21_X1 U16599 ( .B1(n14781), .B2(n14797), .A(n14780), .ZN(P1_U3240) );
  INV_X1 U16600 ( .A(n14782), .ZN(n14783) );
  NOR2_X1 U16601 ( .A1(n14784), .A2(n14783), .ZN(n14786) );
  XNOR2_X1 U16602 ( .A(n14786), .B(n14785), .ZN(n14798) );
  OAI21_X1 U16603 ( .B1(n14789), .B2(n14788), .A(n14787), .ZN(n14794) );
  OAI22_X1 U16604 ( .A1(n14792), .A2(n15249), .B1(n14791), .B2(n14790), .ZN(
        n14793) );
  AOI211_X1 U16605 ( .C1(n15271), .C2(n14795), .A(n14794), .B(n14793), .ZN(
        n14796) );
  OAI21_X1 U16606 ( .B1(n14798), .B2(n14797), .A(n14796), .ZN(P1_U3241) );
  MUX2_X1 U16607 ( .A(n15002), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14821), .Z(
        P1_U3591) );
  MUX2_X1 U16608 ( .A(n14799), .B(P1_DATAO_REG_30__SCAN_IN), .S(n14821), .Z(
        P1_U3590) );
  MUX2_X1 U16609 ( .A(n14800), .B(P1_DATAO_REG_29__SCAN_IN), .S(n14821), .Z(
        P1_U3589) );
  MUX2_X1 U16610 ( .A(n15038), .B(P1_DATAO_REG_28__SCAN_IN), .S(n14821), .Z(
        P1_U3588) );
  MUX2_X1 U16611 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14801), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16612 ( .A(n15037), .B(P1_DATAO_REG_26__SCAN_IN), .S(n14821), .Z(
        P1_U3586) );
  MUX2_X1 U16613 ( .A(n15090), .B(P1_DATAO_REG_25__SCAN_IN), .S(n14821), .Z(
        P1_U3585) );
  MUX2_X1 U16614 ( .A(n14802), .B(P1_DATAO_REG_24__SCAN_IN), .S(n14821), .Z(
        P1_U3584) );
  MUX2_X1 U16615 ( .A(n15089), .B(P1_DATAO_REG_23__SCAN_IN), .S(n14821), .Z(
        P1_U3583) );
  MUX2_X1 U16616 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14803), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16617 ( .A(n15122), .B(P1_DATAO_REG_21__SCAN_IN), .S(n14821), .Z(
        P1_U3581) );
  MUX2_X1 U16618 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14804), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16619 ( .A(n14805), .B(P1_DATAO_REG_19__SCAN_IN), .S(n14821), .Z(
        P1_U3579) );
  MUX2_X1 U16620 ( .A(n14806), .B(P1_DATAO_REG_18__SCAN_IN), .S(n14821), .Z(
        P1_U3578) );
  MUX2_X1 U16621 ( .A(n14807), .B(P1_DATAO_REG_17__SCAN_IN), .S(n14821), .Z(
        P1_U3577) );
  MUX2_X1 U16622 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n15259), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16623 ( .A(n14808), .B(P1_DATAO_REG_15__SCAN_IN), .S(n14821), .Z(
        P1_U3575) );
  MUX2_X1 U16624 ( .A(n15256), .B(P1_DATAO_REG_14__SCAN_IN), .S(n14821), .Z(
        P1_U3574) );
  MUX2_X1 U16625 ( .A(n14809), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14821), .Z(
        P1_U3573) );
  MUX2_X1 U16626 ( .A(n14810), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14821), .Z(
        P1_U3572) );
  MUX2_X1 U16627 ( .A(n14811), .B(P1_DATAO_REG_11__SCAN_IN), .S(n14821), .Z(
        P1_U3571) );
  MUX2_X1 U16628 ( .A(n14812), .B(P1_DATAO_REG_10__SCAN_IN), .S(n14821), .Z(
        P1_U3570) );
  MUX2_X1 U16629 ( .A(n14813), .B(P1_DATAO_REG_9__SCAN_IN), .S(n14821), .Z(
        P1_U3569) );
  MUX2_X1 U16630 ( .A(n14814), .B(P1_DATAO_REG_8__SCAN_IN), .S(n14821), .Z(
        P1_U3568) );
  MUX2_X1 U16631 ( .A(n14815), .B(P1_DATAO_REG_7__SCAN_IN), .S(n14821), .Z(
        P1_U3567) );
  MUX2_X1 U16632 ( .A(n14816), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14821), .Z(
        P1_U3566) );
  MUX2_X1 U16633 ( .A(n14817), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14821), .Z(
        P1_U3565) );
  MUX2_X1 U16634 ( .A(n14818), .B(P1_DATAO_REG_4__SCAN_IN), .S(n14821), .Z(
        P1_U3564) );
  MUX2_X1 U16635 ( .A(n14819), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14821), .Z(
        P1_U3563) );
  MUX2_X1 U16636 ( .A(n14820), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14821), .Z(
        P1_U3562) );
  MUX2_X1 U16637 ( .A(n10096), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14821), .Z(
        P1_U3561) );
  MUX2_X1 U16638 ( .A(n11154), .B(P1_DATAO_REG_0__SCAN_IN), .S(n14821), .Z(
        P1_U3560) );
  OAI22_X1 U16639 ( .A1(n15497), .A2(n14823), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14822), .ZN(n14824) );
  AOI21_X1 U16640 ( .B1(n14825), .B2(n15500), .A(n14824), .ZN(n14834) );
  OAI211_X1 U16641 ( .C1(n14838), .C2(n14827), .A(n15513), .B(n14826), .ZN(
        n14833) );
  MUX2_X1 U16642 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10912), .S(n14828), .Z(
        n14829) );
  OAI21_X1 U16643 ( .B1(n10087), .B2(n15490), .A(n14829), .ZN(n14830) );
  NAND3_X1 U16644 ( .A1(n15506), .A2(n14831), .A3(n14830), .ZN(n14832) );
  NAND3_X1 U16645 ( .A1(n14834), .A2(n14833), .A3(n14832), .ZN(P1_U3244) );
  NOR2_X1 U16646 ( .A1(n15436), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n14835) );
  NOR2_X1 U16647 ( .A1(n14836), .A2(n14835), .ZN(n15488) );
  MUX2_X1 U16648 ( .A(n14838), .B(n14837), .S(n15436), .Z(n14840) );
  NAND2_X1 U16649 ( .A1(n14840), .A2(n14839), .ZN(n14841) );
  OAI211_X1 U16650 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n15488), .A(n14841), .B(
        P1_U4016), .ZN(n15517) );
  INV_X1 U16651 ( .A(n14842), .ZN(n14845) );
  MUX2_X1 U16652 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10915), .S(n14843), .Z(
        n14844) );
  NAND2_X1 U16653 ( .A1(n14845), .A2(n14844), .ZN(n14846) );
  NAND3_X1 U16654 ( .A1(n15506), .A2(n14866), .A3(n14846), .ZN(n14848) );
  AOI22_X1 U16655 ( .A1(n15492), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n14847) );
  AND2_X1 U16656 ( .A1(n14848), .A2(n14847), .ZN(n14854) );
  NAND2_X1 U16657 ( .A1(n15500), .A2(n14849), .ZN(n14853) );
  OAI211_X1 U16658 ( .C1(n14851), .C2(n14850), .A(n15513), .B(n14861), .ZN(
        n14852) );
  NAND4_X1 U16659 ( .A1(n15517), .A2(n14854), .A3(n14853), .A4(n14852), .ZN(
        P1_U3245) );
  INV_X1 U16660 ( .A(n14863), .ZN(n14858) );
  OAI21_X1 U16661 ( .B1(n15497), .B2(n14856), .A(n14855), .ZN(n14857) );
  AOI21_X1 U16662 ( .B1(n14858), .B2(n15500), .A(n14857), .ZN(n14870) );
  MUX2_X1 U16663 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10939), .S(n14863), .Z(
        n14859) );
  NAND3_X1 U16664 ( .A1(n14861), .A2(n14860), .A3(n14859), .ZN(n14862) );
  NAND3_X1 U16665 ( .A1(n15513), .A2(n15510), .A3(n14862), .ZN(n14869) );
  MUX2_X1 U16666 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10917), .S(n14863), .Z(
        n14864) );
  NAND3_X1 U16667 ( .A1(n14866), .A2(n14865), .A3(n14864), .ZN(n14867) );
  NAND3_X1 U16668 ( .A1(n15506), .A2(n15503), .A3(n14867), .ZN(n14868) );
  NAND3_X1 U16669 ( .A1(n14870), .A2(n14869), .A3(n14868), .ZN(P1_U3246) );
  NAND2_X1 U16670 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n14871) );
  OAI21_X1 U16671 ( .B1(n15497), .B2(n14872), .A(n14871), .ZN(n14873) );
  AOI21_X1 U16672 ( .B1(n14874), .B2(n15500), .A(n14873), .ZN(n14885) );
  OAI21_X1 U16673 ( .B1(n14877), .B2(n14876), .A(n14875), .ZN(n14878) );
  NAND2_X1 U16674 ( .A1(n15506), .A2(n14878), .ZN(n14884) );
  MUX2_X1 U16675 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n11808), .S(n14879), .Z(
        n14880) );
  NAND3_X1 U16676 ( .A1(n15512), .A2(n14881), .A3(n14880), .ZN(n14882) );
  NAND3_X1 U16677 ( .A1(n15513), .A2(n14892), .A3(n14882), .ZN(n14883) );
  NAND3_X1 U16678 ( .A1(n14885), .A2(n14884), .A3(n14883), .ZN(P1_U3248) );
  NOR2_X1 U16679 ( .A1(n15497), .A2(n14886), .ZN(n14887) );
  AOI211_X1 U16680 ( .C1(n15500), .C2(n14894), .A(n14888), .B(n14887), .ZN(
        n14899) );
  MUX2_X1 U16681 ( .A(n14889), .B(P1_REG2_REG_6__SCAN_IN), .S(n14894), .Z(
        n14890) );
  NAND3_X1 U16682 ( .A1(n14892), .A2(n14891), .A3(n14890), .ZN(n14893) );
  NAND3_X1 U16683 ( .A1(n15513), .A2(n14902), .A3(n14893), .ZN(n14898) );
  MUX2_X1 U16684 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n14895), .S(n14894), .Z(
        n14896) );
  OAI211_X1 U16685 ( .C1(n6631), .C2(n14896), .A(n15506), .B(n14908), .ZN(
        n14897) );
  NAND3_X1 U16686 ( .A1(n14899), .A2(n14898), .A3(n14897), .ZN(P1_U3249) );
  MUX2_X1 U16687 ( .A(n12034), .B(P1_REG2_REG_7__SCAN_IN), .S(n14911), .Z(
        n14900) );
  NAND3_X1 U16688 ( .A1(n14902), .A2(n14901), .A3(n14900), .ZN(n14903) );
  NAND3_X1 U16689 ( .A1(n15513), .A2(n14904), .A3(n14903), .ZN(n14915) );
  AOI21_X1 U16690 ( .B1(n15492), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n14905), .ZN(
        n14914) );
  MUX2_X1 U16691 ( .A(n10923), .B(P1_REG1_REG_7__SCAN_IN), .S(n14911), .Z(
        n14906) );
  NAND3_X1 U16692 ( .A1(n14908), .A2(n14907), .A3(n14906), .ZN(n14909) );
  NAND3_X1 U16693 ( .A1(n15506), .A2(n14910), .A3(n14909), .ZN(n14913) );
  NAND2_X1 U16694 ( .A1(n15500), .A2(n14911), .ZN(n14912) );
  NAND4_X1 U16695 ( .A1(n14915), .A2(n14914), .A3(n14913), .A4(n14912), .ZN(
        P1_U3250) );
  OAI21_X1 U16696 ( .B1(n14919), .B2(n14918), .A(n14917), .ZN(n14920) );
  NAND3_X1 U16697 ( .A1(n6733), .A2(n15506), .A3(n14920), .ZN(n14932) );
  OAI21_X1 U16698 ( .B1(n15497), .B2(n14922), .A(n14921), .ZN(n14923) );
  AOI21_X1 U16699 ( .B1(n14924), .B2(n15500), .A(n14923), .ZN(n14931) );
  MUX2_X1 U16700 ( .A(n12330), .B(P1_REG2_REG_10__SCAN_IN), .S(n14924), .Z(
        n14925) );
  NAND3_X1 U16701 ( .A1(n14927), .A2(n14926), .A3(n14925), .ZN(n14928) );
  NAND3_X1 U16702 ( .A1(n15513), .A2(n14929), .A3(n14928), .ZN(n14930) );
  NAND3_X1 U16703 ( .A1(n14932), .A2(n14931), .A3(n14930), .ZN(P1_U3253) );
  OR2_X1 U16704 ( .A1(n14933), .A2(n14940), .ZN(n14934) );
  AND2_X1 U16705 ( .A1(n14936), .A2(n14934), .ZN(n14938) );
  XNOR2_X1 U16706 ( .A(n14951), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n14937) );
  AND2_X1 U16707 ( .A1(n14934), .A2(n14937), .ZN(n14935) );
  NAND2_X1 U16708 ( .A1(n14936), .A2(n14935), .ZN(n14953) );
  OAI211_X1 U16709 ( .C1(n14938), .C2(n14937), .A(n15513), .B(n14953), .ZN(
        n14950) );
  XNOR2_X1 U16710 ( .A(n14955), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n14944) );
  OAI22_X1 U16711 ( .A1(n14941), .A2(n14940), .B1(P1_REG1_REG_15__SCAN_IN), 
        .B2(n14939), .ZN(n14943) );
  AOI211_X1 U16712 ( .C1(n14944), .C2(n14943), .A(n14954), .B(n14942), .ZN(
        n14945) );
  INV_X1 U16713 ( .A(n14945), .ZN(n14946) );
  NAND2_X1 U16714 ( .A1(n14947), .A2(n14946), .ZN(n14948) );
  AOI21_X1 U16715 ( .B1(n15492), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n14948), 
        .ZN(n14949) );
  OAI211_X1 U16716 ( .C1(n14975), .C2(n14951), .A(n14950), .B(n14949), .ZN(
        P1_U3259) );
  NAND2_X1 U16717 ( .A1(n14955), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14952) );
  NAND2_X1 U16718 ( .A1(n14953), .A2(n14952), .ZN(n14964) );
  INV_X1 U16719 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15221) );
  XNOR2_X1 U16720 ( .A(n14965), .B(n15221), .ZN(n14963) );
  XNOR2_X1 U16721 ( .A(n14964), .B(n14963), .ZN(n14962) );
  XNOR2_X1 U16722 ( .A(n14965), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14970) );
  XOR2_X1 U16723 ( .A(n14971), .B(n14970), .Z(n14956) );
  NAND2_X1 U16724 ( .A1(n15506), .A2(n14956), .ZN(n14957) );
  NAND2_X1 U16725 ( .A1(n14958), .A2(n14957), .ZN(n14960) );
  INV_X1 U16726 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15458) );
  NOR2_X1 U16727 ( .A1(n15497), .A2(n15458), .ZN(n14959) );
  AOI211_X1 U16728 ( .C1(n15500), .C2(n14965), .A(n14960), .B(n14959), .ZN(
        n14961) );
  OAI21_X1 U16729 ( .B1(n14962), .B2(n14989), .A(n14961), .ZN(P1_U3260) );
  NAND2_X1 U16730 ( .A1(n14964), .A2(n14963), .ZN(n14967) );
  NAND2_X1 U16731 ( .A1(n14965), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14966) );
  NAND2_X1 U16732 ( .A1(n14967), .A2(n14966), .ZN(n14984) );
  XNOR2_X1 U16733 ( .A(n14984), .B(n14974), .ZN(n14982) );
  XNOR2_X1 U16734 ( .A(n14982), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n14979) );
  INV_X1 U16735 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14969) );
  XOR2_X1 U16736 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14980), .Z(n14977) );
  NAND2_X1 U16737 ( .A1(n15492), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n14972) );
  OAI211_X1 U16738 ( .C1(n14975), .C2(n14974), .A(n14973), .B(n14972), .ZN(
        n14976) );
  AOI21_X1 U16739 ( .B1(n14977), .B2(n15506), .A(n14976), .ZN(n14978) );
  OAI21_X1 U16740 ( .B1(n14979), .B2(n14989), .A(n14978), .ZN(P1_U3261) );
  INV_X1 U16741 ( .A(n14992), .ZN(n14988) );
  NAND2_X1 U16742 ( .A1(n14982), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n14986) );
  NAND2_X1 U16743 ( .A1(n14984), .A2(n14983), .ZN(n14985) );
  NAND2_X1 U16744 ( .A1(n14986), .A2(n14985), .ZN(n14987) );
  INV_X1 U16745 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n15185) );
  XNOR2_X1 U16746 ( .A(n14987), .B(n15185), .ZN(n14990) );
  AOI22_X1 U16747 ( .A1(n14988), .A2(n15506), .B1(n15513), .B2(n14990), .ZN(
        n14995) );
  NOR2_X1 U16748 ( .A1(n14990), .A2(n14989), .ZN(n14991) );
  AOI211_X1 U16749 ( .C1(n14992), .C2(n15506), .A(n14991), .B(n15500), .ZN(
        n14994) );
  OAI211_X1 U16750 ( .C1(n7068), .C2(n15497), .A(n14997), .B(n14996), .ZN(
        P1_U3262) );
  XNOR2_X1 U16751 ( .A(n15008), .B(n15376), .ZN(n14999) );
  NAND2_X1 U16752 ( .A1(n14999), .A2(n15168), .ZN(n15276) );
  NOR2_X1 U16753 ( .A1(n15220), .A2(n15000), .ZN(n15003) );
  NAND2_X1 U16754 ( .A1(n15002), .A2(n15001), .ZN(n15279) );
  NOR2_X1 U16755 ( .A1(n15533), .A2(n15279), .ZN(n15010) );
  AOI211_X1 U16756 ( .C1(n15004), .C2(n15524), .A(n15003), .B(n15010), .ZN(
        n15005) );
  OAI21_X1 U16757 ( .B1(n15276), .B2(n15174), .A(n15005), .ZN(P1_U3263) );
  AOI21_X1 U16758 ( .B1(n15006), .B2(n15012), .A(n15270), .ZN(n15007) );
  NAND2_X1 U16759 ( .A1(n15008), .A2(n15007), .ZN(n15280) );
  NOR2_X1 U16760 ( .A1(n15220), .A2(n15009), .ZN(n15011) );
  AOI211_X1 U16761 ( .C1(n15012), .C2(n15524), .A(n15011), .B(n15010), .ZN(
        n15013) );
  OAI21_X1 U16762 ( .B1(n15280), .B2(n15174), .A(n15013), .ZN(P1_U3264) );
  INV_X1 U16763 ( .A(n15284), .ZN(n15029) );
  NAND2_X1 U16764 ( .A1(n15285), .A2(n15220), .ZN(n15028) );
  INV_X1 U16765 ( .A(n15020), .ZN(n15022) );
  INV_X1 U16766 ( .A(n10032), .ZN(n15021) );
  AOI211_X2 U16767 ( .C1(n15023), .C2(n15022), .A(n15270), .B(n15021), .ZN(
        n15283) );
  AOI22_X1 U16768 ( .A1(n15024), .A2(n15526), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n15274), .ZN(n15025) );
  OAI21_X1 U16769 ( .B1(n15383), .B2(n15234), .A(n15025), .ZN(n15026) );
  AOI21_X1 U16770 ( .B1(n15283), .B2(n15522), .A(n15026), .ZN(n15027) );
  OAI211_X1 U16771 ( .C1(n15248), .C2(n15029), .A(n15028), .B(n15027), .ZN(
        P1_U3265) );
  AOI22_X1 U16772 ( .A1(n15030), .A2(n15260), .B1(n15370), .B2(n15031), .ZN(
        n15036) );
  INV_X1 U16773 ( .A(n15030), .ZN(n15033) );
  INV_X1 U16774 ( .A(n15031), .ZN(n15032) );
  AOI22_X1 U16775 ( .A1(n15033), .A2(n15260), .B1(n15370), .B2(n15032), .ZN(
        n15035) );
  AOI22_X1 U16776 ( .A1(n15038), .A2(n15258), .B1(n15257), .B2(n15037), .ZN(
        n15039) );
  INV_X1 U16777 ( .A(n15041), .ZN(n15055) );
  AOI211_X1 U16778 ( .C1(n15042), .C2(n15055), .A(n15270), .B(n15020), .ZN(
        n15289) );
  AOI22_X1 U16779 ( .A1(n15043), .A2(n15526), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n15274), .ZN(n15044) );
  OAI21_X1 U16780 ( .B1(n7759), .B2(n15234), .A(n15044), .ZN(n15045) );
  AOI21_X1 U16781 ( .B1(n15289), .B2(n15522), .A(n15045), .ZN(n15046) );
  OAI21_X1 U16782 ( .B1(n6499), .B2(n15274), .A(n15046), .ZN(P1_U3266) );
  INV_X1 U16783 ( .A(n15292), .ZN(n15051) );
  INV_X1 U16784 ( .A(n15071), .ZN(n15066) );
  NAND3_X1 U16785 ( .A1(n15091), .A2(n15066), .A3(n15070), .ZN(n15074) );
  NAND2_X1 U16786 ( .A1(n15074), .A2(n15048), .ZN(n15049) );
  AOI211_X1 U16787 ( .C1(n15052), .C2(n15526), .A(n15051), .B(n15295), .ZN(
        n15064) );
  INV_X1 U16788 ( .A(n15054), .ZN(n15056) );
  OAI211_X1 U16789 ( .C1(n7758), .C2(n15056), .A(n15055), .B(n15168), .ZN(
        n15291) );
  INV_X1 U16790 ( .A(n15291), .ZN(n15062) );
  OAI22_X1 U16791 ( .A1(n7758), .A2(n15234), .B1(n15057), .B2(n15220), .ZN(
        n15061) );
  XNOR2_X1 U16792 ( .A(n15059), .B(n15058), .ZN(n15293) );
  NOR2_X1 U16793 ( .A1(n15293), .A2(n15248), .ZN(n15060) );
  AOI211_X1 U16794 ( .C1(n15062), .C2(n15522), .A(n15061), .B(n15060), .ZN(
        n15063) );
  OAI21_X1 U16795 ( .B1(n15064), .B2(n15533), .A(n15063), .ZN(P1_U3267) );
  INV_X1 U16796 ( .A(n15065), .ZN(n15067) );
  NAND2_X1 U16797 ( .A1(n15069), .A2(n15068), .ZN(n15301) );
  INV_X1 U16798 ( .A(n15091), .ZN(n15073) );
  INV_X1 U16799 ( .A(n15070), .ZN(n15072) );
  OAI21_X1 U16800 ( .B1(n15073), .B2(n15072), .A(n15071), .ZN(n15075) );
  AOI21_X1 U16801 ( .B1(n15075), .B2(n15074), .A(n15160), .ZN(n15302) );
  INV_X1 U16802 ( .A(n15300), .ZN(n15076) );
  OAI21_X1 U16803 ( .B1(n15302), .B2(n15076), .A(n15220), .ZN(n15084) );
  INV_X1 U16804 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n15077) );
  OAI22_X1 U16805 ( .A1(n15078), .A2(n15217), .B1(n15077), .B2(n15220), .ZN(
        n15082) );
  XOR2_X1 U16806 ( .A(n15079), .B(n15298), .Z(n15080) );
  NAND2_X1 U16807 ( .A1(n15080), .A2(n15168), .ZN(n15299) );
  NOR2_X1 U16808 ( .A1(n15299), .A2(n15174), .ZN(n15081) );
  AOI211_X1 U16809 ( .C1(n15524), .C2(n15298), .A(n15082), .B(n15081), .ZN(
        n15083) );
  OAI211_X1 U16810 ( .C1(n15301), .C2(n15248), .A(n15084), .B(n15083), .ZN(
        P1_U3268) );
  INV_X1 U16811 ( .A(n15109), .ZN(n15086) );
  NAND2_X1 U16812 ( .A1(n15086), .A2(n15085), .ZN(n15088) );
  AOI21_X1 U16813 ( .B1(n15092), .B2(n15088), .A(n15087), .ZN(n15096) );
  AOI22_X1 U16814 ( .A1(n15090), .A2(n15258), .B1(n15257), .B2(n15089), .ZN(
        n15095) );
  OAI211_X1 U16815 ( .C1(n15093), .C2(n15092), .A(n15091), .B(n15260), .ZN(
        n15094) );
  INV_X1 U16816 ( .A(n15307), .ZN(n15105) );
  INV_X1 U16817 ( .A(n15112), .ZN(n15098) );
  INV_X1 U16818 ( .A(n15079), .ZN(n15097) );
  AOI211_X1 U16819 ( .C1(n15099), .C2(n15098), .A(n15270), .B(n15097), .ZN(
        n15306) );
  INV_X1 U16820 ( .A(n15100), .ZN(n15101) );
  AOI22_X1 U16821 ( .A1(n15101), .A2(n15526), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n15274), .ZN(n15102) );
  OAI21_X1 U16822 ( .B1(n15396), .B2(n15234), .A(n15102), .ZN(n15103) );
  AOI21_X1 U16823 ( .B1(n15306), .B2(n15522), .A(n15103), .ZN(n15104) );
  OAI21_X1 U16824 ( .B1(n15105), .B2(n15274), .A(n15104), .ZN(P1_U3269) );
  XOR2_X1 U16825 ( .A(n15111), .B(n15106), .Z(n15108) );
  OAI21_X1 U16826 ( .B1(n15108), .B2(n15160), .A(n15107), .ZN(n15310) );
  INV_X1 U16827 ( .A(n15310), .ZN(n15119) );
  AOI21_X1 U16828 ( .B1(n15111), .B2(n15110), .A(n15109), .ZN(n15312) );
  AOI211_X1 U16829 ( .C1(n15113), .C2(n15130), .A(n15270), .B(n15112), .ZN(
        n15311) );
  NAND2_X1 U16830 ( .A1(n15311), .A2(n15522), .ZN(n15116) );
  AOI22_X1 U16831 ( .A1(n15114), .A2(n15526), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15274), .ZN(n15115) );
  OAI211_X1 U16832 ( .C1(n15400), .C2(n15234), .A(n15116), .B(n15115), .ZN(
        n15117) );
  AOI21_X1 U16833 ( .B1(n15312), .B2(n15519), .A(n15117), .ZN(n15118) );
  OAI21_X1 U16834 ( .B1(n15119), .B2(n15533), .A(n15118), .ZN(P1_U3270) );
  NAND3_X1 U16835 ( .A1(n15120), .A2(n15158), .A3(n15159), .ZN(n15157) );
  AOI21_X1 U16836 ( .B1(n15157), .B2(n15121), .A(n10020), .ZN(n15140) );
  AOI21_X1 U16837 ( .B1(n15148), .B2(n15122), .A(n15140), .ZN(n15125) );
  OAI21_X1 U16838 ( .B1(n15129), .B2(n15128), .A(n15127), .ZN(n15317) );
  INV_X1 U16839 ( .A(n15130), .ZN(n15131) );
  AOI211_X1 U16840 ( .C1(n15132), .C2(n15146), .A(n15270), .B(n15131), .ZN(
        n15316) );
  NAND2_X1 U16841 ( .A1(n15316), .A2(n15522), .ZN(n15135) );
  AOI22_X1 U16842 ( .A1(n15133), .A2(n15526), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n15274), .ZN(n15134) );
  OAI211_X1 U16843 ( .C1(n15234), .C2(n15404), .A(n15135), .B(n15134), .ZN(
        n15136) );
  AOI21_X1 U16844 ( .B1(n15317), .B2(n15519), .A(n15136), .ZN(n15137) );
  OAI21_X1 U16845 ( .B1(n15315), .B2(n15533), .A(n15137), .ZN(P1_U3271) );
  NOR2_X1 U16846 ( .A1(n15139), .A2(n15138), .ZN(n15141) );
  AOI211_X1 U16847 ( .C1(n15141), .C2(n15157), .A(n15160), .B(n15140), .ZN(
        n15143) );
  NOR2_X1 U16848 ( .A1(n15143), .A2(n15142), .ZN(n15324) );
  OAI21_X1 U16849 ( .B1(n15145), .B2(n10020), .A(n15144), .ZN(n15320) );
  INV_X1 U16850 ( .A(n15167), .ZN(n15147) );
  OAI211_X1 U16851 ( .C1(n15148), .C2(n15147), .A(n15146), .B(n15168), .ZN(
        n15321) );
  INV_X1 U16852 ( .A(n15149), .ZN(n15150) );
  AOI22_X1 U16853 ( .A1(n15150), .A2(n15526), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n15274), .ZN(n15153) );
  NAND2_X1 U16854 ( .A1(n15151), .A2(n15524), .ZN(n15152) );
  OAI211_X1 U16855 ( .C1(n15321), .C2(n15174), .A(n15153), .B(n15152), .ZN(
        n15154) );
  AOI21_X1 U16856 ( .B1(n15320), .B2(n15519), .A(n15154), .ZN(n15155) );
  OAI21_X1 U16857 ( .B1(n15324), .B2(n15533), .A(n15155), .ZN(P1_U3272) );
  AOI21_X1 U16858 ( .B1(n15156), .B2(n15158), .A(n15354), .ZN(n15166) );
  INV_X1 U16859 ( .A(n15157), .ZN(n15162) );
  AOI21_X1 U16860 ( .B1(n15120), .B2(n15159), .A(n15158), .ZN(n15161) );
  NOR3_X1 U16861 ( .A1(n15162), .A2(n15161), .A3(n15160), .ZN(n15163) );
  AOI211_X1 U16862 ( .C1(n15166), .C2(n15165), .A(n15164), .B(n15163), .ZN(
        n15326) );
  OAI211_X1 U16863 ( .C1(n15183), .C2(n15328), .A(n15168), .B(n15167), .ZN(
        n15325) );
  INV_X1 U16864 ( .A(n15169), .ZN(n15170) );
  AOI22_X1 U16865 ( .A1(n15170), .A2(n15526), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n15274), .ZN(n15173) );
  NAND2_X1 U16866 ( .A1(n15171), .A2(n15524), .ZN(n15172) );
  OAI211_X1 U16867 ( .C1(n15325), .C2(n15174), .A(n15173), .B(n15172), .ZN(
        n15175) );
  INV_X1 U16868 ( .A(n15175), .ZN(n15176) );
  OAI21_X1 U16869 ( .B1(n15326), .B2(n15533), .A(n15176), .ZN(P1_U3273) );
  XNOR2_X1 U16870 ( .A(n15178), .B(n15177), .ZN(n15335) );
  OAI21_X1 U16871 ( .B1(n15179), .B2(n7736), .A(n15120), .ZN(n15180) );
  NAND2_X1 U16872 ( .A1(n15180), .A2(n15260), .ZN(n15334) );
  OAI211_X1 U16873 ( .C1(n15217), .C2(n15181), .A(n15334), .B(n15329), .ZN(
        n15182) );
  NAND2_X1 U16874 ( .A1(n15182), .A2(n15220), .ZN(n15189) );
  INV_X1 U16875 ( .A(n15198), .ZN(n15184) );
  AOI211_X1 U16876 ( .C1(n15332), .C2(n15184), .A(n15270), .B(n15183), .ZN(
        n15330) );
  OAI22_X1 U16877 ( .A1(n15186), .A2(n15234), .B1(n15185), .B2(n15220), .ZN(
        n15187) );
  AOI21_X1 U16878 ( .B1(n15330), .B2(n15522), .A(n15187), .ZN(n15188) );
  OAI211_X1 U16879 ( .C1(n15335), .C2(n15248), .A(n15189), .B(n15188), .ZN(
        P1_U3274) );
  XOR2_X1 U16880 ( .A(n15190), .B(n15192), .Z(n15341) );
  OAI211_X1 U16881 ( .C1(n15193), .C2(n15192), .A(n15191), .B(n15260), .ZN(
        n15195) );
  INV_X1 U16882 ( .A(n15340), .ZN(n15197) );
  INV_X1 U16883 ( .A(n15196), .ZN(n15337) );
  OAI21_X1 U16884 ( .B1(n15197), .B2(n15337), .A(n15220), .ZN(n15205) );
  AOI211_X1 U16885 ( .C1(n15199), .C2(n15219), .A(n15270), .B(n15198), .ZN(
        n15338) );
  AOI22_X1 U16886 ( .A1(n15533), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n15200), 
        .B2(n15526), .ZN(n15201) );
  OAI21_X1 U16887 ( .B1(n15202), .B2(n15234), .A(n15201), .ZN(n15203) );
  AOI21_X1 U16888 ( .B1(n15338), .B2(n15522), .A(n15203), .ZN(n15204) );
  OAI211_X1 U16889 ( .C1(n15341), .C2(n15248), .A(n15205), .B(n15204), .ZN(
        P1_U3275) );
  INV_X1 U16890 ( .A(n12763), .ZN(n15207) );
  AOI21_X1 U16891 ( .B1(n15207), .B2(n15206), .A(n6554), .ZN(n15210) );
  INV_X1 U16892 ( .A(n15208), .ZN(n15209) );
  NOR2_X1 U16893 ( .A1(n15210), .A2(n15209), .ZN(n15212) );
  OAI21_X1 U16894 ( .B1(n15212), .B2(n15213), .A(n15211), .ZN(n15348) );
  OAI211_X1 U16895 ( .C1(n15215), .C2(n9825), .A(n15260), .B(n15214), .ZN(
        n15347) );
  OAI211_X1 U16896 ( .C1(n15217), .C2(n15216), .A(n15347), .B(n15342), .ZN(
        n15218) );
  NAND2_X1 U16897 ( .A1(n15218), .A2(n15220), .ZN(n15225) );
  AOI211_X1 U16898 ( .C1(n15345), .C2(n15230), .A(n15270), .B(n7772), .ZN(
        n15343) );
  INV_X1 U16899 ( .A(n15345), .ZN(n15222) );
  OAI22_X1 U16900 ( .A1(n15222), .A2(n15234), .B1(n15221), .B2(n15220), .ZN(
        n15223) );
  AOI21_X1 U16901 ( .B1(n15343), .B2(n15522), .A(n15223), .ZN(n15224) );
  OAI211_X1 U16902 ( .C1(n15348), .C2(n15248), .A(n15225), .B(n15224), .ZN(
        P1_U3276) );
  NOR2_X1 U16903 ( .A1(n15250), .A2(n15226), .ZN(n15255) );
  INV_X1 U16904 ( .A(n15227), .ZN(n15228) );
  NOR2_X1 U16905 ( .A1(n15255), .A2(n15228), .ZN(n15229) );
  XNOR2_X1 U16906 ( .A(n15229), .B(n15236), .ZN(n15355) );
  INV_X1 U16907 ( .A(n15269), .ZN(n15232) );
  INV_X1 U16908 ( .A(n15230), .ZN(n15231) );
  AOI211_X1 U16909 ( .C1(n15351), .C2(n15232), .A(n15270), .B(n15231), .ZN(
        n15349) );
  INV_X1 U16910 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n15233) );
  OAI22_X1 U16911 ( .A1(n15235), .A2(n15234), .B1(n15233), .B2(n15220), .ZN(
        n15246) );
  OAI21_X1 U16912 ( .B1(n6584), .B2(n9812), .A(n15237), .ZN(n15238) );
  NAND2_X1 U16913 ( .A1(n15238), .A2(n15260), .ZN(n15352) );
  OAI22_X1 U16914 ( .A1(n15242), .A2(n15241), .B1(n15240), .B2(n15239), .ZN(
        n15350) );
  AOI21_X1 U16915 ( .B1(n15243), .B2(n15526), .A(n15350), .ZN(n15244) );
  AOI21_X1 U16916 ( .B1(n15352), .B2(n15244), .A(n15533), .ZN(n15245) );
  AOI211_X1 U16917 ( .C1(n15349), .C2(n15522), .A(n15246), .B(n15245), .ZN(
        n15247) );
  OAI21_X1 U16918 ( .B1(n15248), .B2(n15355), .A(n15247), .ZN(P1_U3277) );
  INV_X1 U16919 ( .A(n15249), .ZN(n15267) );
  INV_X1 U16920 ( .A(n15250), .ZN(n15253) );
  AOI21_X1 U16921 ( .B1(n15253), .B2(n15252), .A(n15251), .ZN(n15254) );
  OAI21_X1 U16922 ( .B1(n15255), .B2(n15254), .A(n15370), .ZN(n15266) );
  AOI22_X1 U16923 ( .A1(n15259), .A2(n15258), .B1(n15257), .B2(n15256), .ZN(
        n15265) );
  OAI211_X1 U16924 ( .C1(n15263), .C2(n15262), .A(n15261), .B(n15260), .ZN(
        n15264) );
  NAND3_X1 U16925 ( .A1(n15266), .A2(n15265), .A3(n15264), .ZN(n15357) );
  AOI21_X1 U16926 ( .B1(n15267), .B2(n15526), .A(n15357), .ZN(n15275) );
  AOI22_X1 U16927 ( .A1(n15271), .A2(n15524), .B1(P1_REG2_REG_15__SCAN_IN), 
        .B2(n15274), .ZN(n15273) );
  AOI211_X1 U16928 ( .C1(n15271), .C2(n7764), .A(n15270), .B(n15269), .ZN(
        n15356) );
  NAND2_X1 U16929 ( .A1(n15356), .A2(n15522), .ZN(n15272) );
  OAI211_X1 U16930 ( .C1(n15275), .C2(n15274), .A(n15273), .B(n15272), .ZN(
        P1_U3278) );
  INV_X1 U16931 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n15277) );
  AND2_X2 U16932 ( .A1(n15276), .A2(n15279), .ZN(n15373) );
  OAI21_X1 U16933 ( .B1(n15376), .B2(n10080), .A(n15278), .ZN(P1_U3559) );
  INV_X1 U16934 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n15281) );
  OAI21_X1 U16935 ( .B1(n15380), .B2(n10080), .A(n15282), .ZN(P1_U3558) );
  INV_X1 U16936 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n15286) );
  NAND2_X1 U16937 ( .A1(n15552), .A2(n15286), .ZN(n15287) );
  OAI21_X1 U16938 ( .B1(n15383), .B2(n10080), .A(n15288), .ZN(P1_U3556) );
  INV_X1 U16939 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n15290) );
  INV_X1 U16940 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n15296) );
  OAI211_X1 U16941 ( .C1(n15293), .C2(n15354), .A(n15292), .B(n15291), .ZN(
        n15294) );
  NOR2_X1 U16942 ( .A1(n15295), .A2(n15294), .ZN(n15386) );
  MUX2_X1 U16943 ( .A(n15296), .B(n15386), .S(n15554), .Z(n15297) );
  OAI21_X1 U16944 ( .B1(n7758), .B2(n10080), .A(n15297), .ZN(P1_U3554) );
  INV_X1 U16945 ( .A(n15298), .ZN(n15392) );
  INV_X1 U16946 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n15304) );
  OAI211_X1 U16947 ( .C1(n15301), .C2(n15354), .A(n15300), .B(n15299), .ZN(
        n15303) );
  NOR2_X1 U16948 ( .A1(n15303), .A2(n15302), .ZN(n15389) );
  MUX2_X1 U16949 ( .A(n15304), .B(n15389), .S(n15554), .Z(n15305) );
  INV_X1 U16950 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n15308) );
  NOR2_X1 U16951 ( .A1(n15307), .A2(n15306), .ZN(n15393) );
  MUX2_X1 U16952 ( .A(n15308), .B(n15393), .S(n15554), .Z(n15309) );
  AOI211_X1 U16953 ( .C1(n15370), .C2(n15312), .A(n15311), .B(n15310), .ZN(
        n15397) );
  MUX2_X1 U16954 ( .A(n15313), .B(n15397), .S(n15554), .Z(n15314) );
  OAI21_X1 U16955 ( .B1(n15400), .B2(n10080), .A(n15314), .ZN(P1_U3551) );
  INV_X1 U16956 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n15318) );
  MUX2_X1 U16957 ( .A(n15318), .B(n15401), .S(n15554), .Z(n15319) );
  OAI21_X1 U16958 ( .B1(n10080), .B2(n15404), .A(n15319), .ZN(P1_U3550) );
  NAND2_X1 U16959 ( .A1(n15320), .A2(n15370), .ZN(n15322) );
  NAND4_X1 U16960 ( .A1(n15324), .A2(n15323), .A3(n15322), .A4(n15321), .ZN(
        n15405) );
  MUX2_X1 U16961 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15405), .S(n15554), .Z(
        P1_U3549) );
  OAI211_X1 U16962 ( .C1(n15328), .C2(n15327), .A(n15326), .B(n15325), .ZN(
        n15406) );
  MUX2_X1 U16963 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15406), .S(n15554), .Z(
        P1_U3548) );
  INV_X1 U16964 ( .A(n15329), .ZN(n15331) );
  AOI211_X1 U16965 ( .C1(n15332), .C2(n15547), .A(n15331), .B(n15330), .ZN(
        n15333) );
  OAI211_X1 U16966 ( .C1(n15354), .C2(n15335), .A(n15334), .B(n15333), .ZN(
        n15407) );
  MUX2_X1 U16967 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15407), .S(n15554), .Z(
        P1_U3547) );
  NOR3_X1 U16968 ( .A1(n15338), .A2(n15337), .A3(n15336), .ZN(n15339) );
  OAI211_X1 U16969 ( .C1(n15354), .C2(n15341), .A(n15340), .B(n15339), .ZN(
        n15408) );
  MUX2_X1 U16970 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15408), .S(n15554), .Z(
        P1_U3546) );
  INV_X1 U16971 ( .A(n15342), .ZN(n15344) );
  AOI211_X1 U16972 ( .C1(n15345), .C2(n15547), .A(n15344), .B(n15343), .ZN(
        n15346) );
  OAI211_X1 U16973 ( .C1(n15354), .C2(n15348), .A(n15347), .B(n15346), .ZN(
        n15409) );
  MUX2_X1 U16974 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15409), .S(n15554), .Z(
        P1_U3545) );
  AOI211_X1 U16975 ( .C1(n15351), .C2(n15547), .A(n15350), .B(n15349), .ZN(
        n15353) );
  OAI211_X1 U16976 ( .C1(n15355), .C2(n15354), .A(n15353), .B(n15352), .ZN(
        n15410) );
  MUX2_X1 U16977 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15410), .S(n15554), .Z(
        P1_U3544) );
  NOR2_X1 U16978 ( .A1(n15357), .A2(n15356), .ZN(n15411) );
  MUX2_X1 U16979 ( .A(n15358), .B(n15411), .S(n15554), .Z(n15359) );
  OAI21_X1 U16980 ( .B1(n15414), .B2(n10080), .A(n15359), .ZN(P1_U3543) );
  AOI211_X1 U16981 ( .C1(n15362), .C2(n15370), .A(n15361), .B(n15360), .ZN(
        n15415) );
  MUX2_X1 U16982 ( .A(n15363), .B(n15415), .S(n15554), .Z(n15364) );
  OAI21_X1 U16983 ( .B1(n7762), .B2(n10080), .A(n15364), .ZN(P1_U3542) );
  INV_X1 U16984 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n15371) );
  NAND2_X1 U16985 ( .A1(n15366), .A2(n15365), .ZN(n15368) );
  AOI211_X1 U16986 ( .C1(n15370), .C2(n15369), .A(n15368), .B(n15367), .ZN(
        n15418) );
  MUX2_X1 U16987 ( .A(n15371), .B(n15418), .S(n15554), .Z(n15372) );
  OAI21_X1 U16988 ( .B1(n15421), .B2(n10080), .A(n15372), .ZN(P1_U3541) );
  OAI21_X1 U16989 ( .B1(n15376), .B2(n10072), .A(n15375), .ZN(P1_U3527) );
  OAI21_X1 U16990 ( .B1(n15380), .B2(n10072), .A(n15379), .ZN(P1_U3526) );
  INV_X1 U16991 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n15387) );
  MUX2_X1 U16992 ( .A(n15387), .B(n15386), .S(n15550), .Z(n15388) );
  OAI21_X1 U16993 ( .B1(n7758), .B2(n10072), .A(n15388), .ZN(P1_U3522) );
  OAI21_X1 U16994 ( .B1(n15392), .B2(n10072), .A(n15391), .ZN(P1_U3521) );
  MUX2_X1 U16995 ( .A(n15394), .B(n15393), .S(n15550), .Z(n15395) );
  OAI21_X1 U16996 ( .B1(n15396), .B2(n10072), .A(n15395), .ZN(P1_U3520) );
  INV_X1 U16997 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n15398) );
  MUX2_X1 U16998 ( .A(n15398), .B(n15397), .S(n15550), .Z(n15399) );
  OAI21_X1 U16999 ( .B1(n15400), .B2(n10072), .A(n15399), .ZN(P1_U3519) );
  MUX2_X1 U17000 ( .A(n15402), .B(n15401), .S(n15550), .Z(n15403) );
  OAI21_X1 U17001 ( .B1(n10072), .B2(n15404), .A(n15403), .ZN(P1_U3518) );
  MUX2_X1 U17002 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15405), .S(n15550), .Z(
        P1_U3517) );
  MUX2_X1 U17003 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15406), .S(n15550), .Z(
        P1_U3516) );
  MUX2_X1 U17004 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15407), .S(n15550), .Z(
        P1_U3515) );
  MUX2_X1 U17005 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15408), .S(n15550), .Z(
        P1_U3513) );
  MUX2_X1 U17006 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15409), .S(n15550), .Z(
        P1_U3510) );
  MUX2_X1 U17007 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15410), .S(n15550), .Z(
        P1_U3507) );
  MUX2_X1 U17008 ( .A(n15412), .B(n15411), .S(n15550), .Z(n15413) );
  OAI21_X1 U17009 ( .B1(n15414), .B2(n10072), .A(n15413), .ZN(P1_U3504) );
  INV_X1 U17010 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n15416) );
  MUX2_X1 U17011 ( .A(n15416), .B(n15415), .S(n15550), .Z(n15417) );
  OAI21_X1 U17012 ( .B1(n7762), .B2(n10072), .A(n15417), .ZN(P1_U3501) );
  MUX2_X1 U17013 ( .A(n15419), .B(n15418), .S(n15550), .Z(n15420) );
  OAI21_X1 U17014 ( .B1(n15421), .B2(n10072), .A(n15420), .ZN(P1_U3498) );
  NOR4_X1 U17015 ( .A1(n6630), .A2(P1_IR_REG_30__SCAN_IN), .A3(n15422), .A4(
        P1_U3086), .ZN(n15423) );
  AOI21_X1 U17016 ( .B1(n15424), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15423), 
        .ZN(n15425) );
  OAI21_X1 U17017 ( .B1(n15427), .B2(n15426), .A(n15425), .ZN(P1_U3324) );
  OAI222_X1 U17018 ( .A1(n15435), .A2(n15431), .B1(n15433), .B2(n15430), .C1(
        P1_U3086), .C2(n15428), .ZN(P1_U3326) );
  OAI222_X1 U17019 ( .A1(P1_U3086), .A2(n15436), .B1(n15435), .B2(n15434), 
        .C1(n15433), .C2(n15432), .ZN(P1_U3328) );
  MUX2_X1 U17020 ( .A(n15438), .B(n15437), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U17021 ( .A(n15439), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XOR2_X1 U17022 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15440), .Z(SUB_1596_U53) );
  INV_X1 U17023 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15443) );
  INV_X1 U17024 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15444) );
  NAND2_X1 U17025 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15444), .ZN(n15446) );
  AOI22_X1 U17026 ( .A1(n15447), .A2(n15446), .B1(P3_ADDR_REG_15__SCAN_IN), 
        .B2(n15445), .ZN(n15453) );
  XOR2_X1 U17027 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n15453), .Z(n15455) );
  XNOR2_X1 U17028 ( .A(n15455), .B(P3_ADDR_REG_16__SCAN_IN), .ZN(n15449) );
  NOR2_X1 U17029 ( .A1(n15452), .A2(n6580), .ZN(n15450) );
  XOR2_X1 U17030 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n15450), .Z(SUB_1596_U64)
         );
  INV_X1 U17031 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15451) );
  NAND2_X1 U17032 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15453), .ZN(n15457) );
  INV_X1 U17033 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15454) );
  NAND2_X1 U17034 ( .A1(n15455), .A2(n15454), .ZN(n15456) );
  NAND2_X1 U17035 ( .A1(n15457), .A2(n15456), .ZN(n15465) );
  XNOR2_X1 U17036 ( .A(n15465), .B(n15458), .ZN(n15467) );
  XNOR2_X1 U17037 ( .A(n15467), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n15459) );
  NAND2_X1 U17038 ( .A1(n7116), .A2(n15462), .ZN(n15460) );
  XNOR2_X1 U17039 ( .A(n15460), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  AND2_X1 U17040 ( .A1(n15475), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n15476) );
  NOR2_X1 U17041 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n15475), .ZN(n15464) );
  NOR2_X1 U17042 ( .A1(n15476), .A2(n15464), .ZN(n15468) );
  NOR2_X1 U17043 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n15465), .ZN(n15466) );
  AOI21_X1 U17044 ( .B1(n15467), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n15466), 
        .ZN(n15477) );
  XOR2_X1 U17045 ( .A(n15468), .B(n15477), .Z(n15470) );
  XNOR2_X1 U17046 ( .A(n15470), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(n15469) );
  XNOR2_X1 U17047 ( .A(n15471), .B(n15469), .ZN(SUB_1596_U62) );
  INV_X1 U17048 ( .A(n15471), .ZN(n15474) );
  INV_X1 U17049 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15473) );
  AOI21_X1 U17050 ( .B1(n15471), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n15470), 
        .ZN(n15472) );
  OAI22_X1 U17051 ( .A1(n15477), .A2(n15476), .B1(P1_ADDR_REG_18__SCAN_IN), 
        .B2(n15475), .ZN(n15480) );
  XNOR2_X1 U17052 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P3_ADDR_REG_19__SCAN_IN), 
        .ZN(n15478) );
  XNOR2_X1 U17053 ( .A(n15478), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n15479) );
  XNOR2_X1 U17054 ( .A(n15480), .B(n15479), .ZN(n15481) );
  XNOR2_X1 U17055 ( .A(n15482), .B(n15481), .ZN(SUB_1596_U4) );
  AOI21_X1 U17056 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15483) );
  OAI21_X1 U17057 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15483), 
        .ZN(U28) );
  AOI21_X1 U17058 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15484) );
  OAI21_X1 U17059 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15484), 
        .ZN(U29) );
  XOR2_X1 U17060 ( .A(n15486), .B(n15485), .Z(n15487) );
  XNOR2_X1 U17061 ( .A(n15487), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  OAI21_X1 U17062 ( .B1(n15489), .B2(P1_REG1_REG_0__SCAN_IN), .A(n15488), .ZN(
        n15491) );
  XNOR2_X1 U17063 ( .A(n15491), .B(n15490), .ZN(n15495) );
  AOI22_X1 U17064 ( .A1(n15492), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15493) );
  OAI21_X1 U17065 ( .B1(n15495), .B2(n15494), .A(n15493), .ZN(P1_U3243) );
  NOR2_X1 U17066 ( .A1(n15497), .A2(n15496), .ZN(n15498) );
  AOI211_X1 U17067 ( .C1(n15500), .C2(n15507), .A(n15499), .B(n15498), .ZN(
        n15516) );
  MUX2_X1 U17068 ( .A(n10918), .B(P1_REG1_REG_4__SCAN_IN), .S(n15507), .Z(
        n15501) );
  NAND3_X1 U17069 ( .A1(n15503), .A2(n15502), .A3(n15501), .ZN(n15504) );
  NAND3_X1 U17070 ( .A1(n15506), .A2(n15505), .A3(n15504), .ZN(n15515) );
  MUX2_X1 U17071 ( .A(n11563), .B(P1_REG2_REG_4__SCAN_IN), .S(n15507), .Z(
        n15508) );
  NAND3_X1 U17072 ( .A1(n15510), .A2(n15509), .A3(n15508), .ZN(n15511) );
  NAND3_X1 U17073 ( .A1(n15513), .A2(n15512), .A3(n15511), .ZN(n15514) );
  AND3_X1 U17074 ( .A1(n15516), .A2(n15515), .A3(n15514), .ZN(n15518) );
  NAND2_X1 U17075 ( .A1(n15518), .A2(n15517), .ZN(P1_U3247) );
  NAND2_X1 U17076 ( .A1(n15520), .A2(n15519), .ZN(n15530) );
  NAND2_X1 U17077 ( .A1(n15522), .A2(n15521), .ZN(n15529) );
  NAND2_X1 U17078 ( .A1(n15524), .A2(n15523), .ZN(n15528) );
  AOI22_X1 U17079 ( .A1(n15533), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n15526), 
        .B2(n15525), .ZN(n15527) );
  AND4_X1 U17080 ( .A1(n15530), .A2(n15529), .A3(n15528), .A4(n15527), .ZN(
        n15531) );
  OAI21_X1 U17081 ( .B1(n15533), .B2(n15532), .A(n15531), .ZN(P1_U3290) );
  AND2_X1 U17082 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15539), .ZN(P1_U3294) );
  INV_X1 U17083 ( .A(n15539), .ZN(n15538) );
  NOR2_X1 U17084 ( .A1(n15538), .A2(n15534), .ZN(P1_U3295) );
  AND2_X1 U17085 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15539), .ZN(P1_U3296) );
  AND2_X1 U17086 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15539), .ZN(P1_U3297) );
  AND2_X1 U17087 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15539), .ZN(P1_U3298) );
  AND2_X1 U17088 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15539), .ZN(P1_U3299) );
  AND2_X1 U17089 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15539), .ZN(P1_U3300) );
  AND2_X1 U17090 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15539), .ZN(P1_U3301) );
  AND2_X1 U17091 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15539), .ZN(P1_U3302) );
  AND2_X1 U17092 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15539), .ZN(P1_U3303) );
  AND2_X1 U17093 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15539), .ZN(P1_U3304) );
  AND2_X1 U17094 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15539), .ZN(P1_U3305) );
  AND2_X1 U17095 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15539), .ZN(P1_U3306) );
  NOR2_X1 U17096 ( .A1(n15538), .A2(n15535), .ZN(P1_U3307) );
  AND2_X1 U17097 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15539), .ZN(P1_U3308) );
  AND2_X1 U17098 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15539), .ZN(P1_U3309) );
  NOR2_X1 U17099 ( .A1(n15538), .A2(n15536), .ZN(P1_U3310) );
  AND2_X1 U17100 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15539), .ZN(P1_U3311) );
  AND2_X1 U17101 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15539), .ZN(P1_U3312) );
  AND2_X1 U17102 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15539), .ZN(P1_U3313) );
  AND2_X1 U17103 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15539), .ZN(P1_U3314) );
  AND2_X1 U17104 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15539), .ZN(P1_U3315) );
  NOR2_X1 U17105 ( .A1(n15538), .A2(n15537), .ZN(P1_U3316) );
  AND2_X1 U17106 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15539), .ZN(P1_U3317) );
  AND2_X1 U17107 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15539), .ZN(P1_U3318) );
  AND2_X1 U17108 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15539), .ZN(P1_U3319) );
  AND2_X1 U17109 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15539), .ZN(P1_U3320) );
  AND2_X1 U17110 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15539), .ZN(P1_U3321) );
  AND2_X1 U17111 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15539), .ZN(P1_U3322) );
  AND2_X1 U17112 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15539), .ZN(P1_U3323) );
  INV_X1 U17113 ( .A(n15540), .ZN(n15542) );
  AOI211_X1 U17114 ( .C1(n15543), .C2(n15547), .A(n15542), .B(n15541), .ZN(
        n15551) );
  AOI22_X1 U17115 ( .A1(n15550), .A2(n15551), .B1(n9675), .B2(n15549), .ZN(
        P1_U3477) );
  INV_X1 U17116 ( .A(n15544), .ZN(n15546) );
  AOI211_X1 U17117 ( .C1(n15548), .C2(n15547), .A(n15546), .B(n15545), .ZN(
        n15553) );
  AOI22_X1 U17118 ( .A1(n15550), .A2(n15553), .B1(n9692), .B2(n15549), .ZN(
        P1_U3480) );
  AOI22_X1 U17119 ( .A1(n15554), .A2(n15551), .B1(n14895), .B2(n15552), .ZN(
        P1_U3534) );
  AOI22_X1 U17120 ( .A1(n15554), .A2(n15553), .B1(n10923), .B2(n15552), .ZN(
        P1_U3535) );
  NOR2_X1 U17121 ( .A1(n15585), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U17122 ( .A1(n15613), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n15610), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n15558) );
  AOI22_X1 U17123 ( .A1(n15585), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n15557) );
  OAI22_X1 U17124 ( .A1(n15597), .A2(P2_REG1_REG_0__SCAN_IN), .B1(
        P2_REG2_REG_0__SCAN_IN), .B2(n15591), .ZN(n15555) );
  OAI21_X1 U17125 ( .B1(n15587), .B2(n15555), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n15556) );
  OAI211_X1 U17126 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n15558), .A(n15557), .B(
        n15556), .ZN(P2_U3214) );
  OAI22_X1 U17127 ( .A1(n15608), .A2(n15560), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15559), .ZN(n15561) );
  AOI21_X1 U17128 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n15585), .A(n15561), .ZN(
        n15570) );
  OAI211_X1 U17129 ( .C1(n15564), .C2(n15563), .A(n15613), .B(n15562), .ZN(
        n15569) );
  AOI211_X1 U17130 ( .C1(n15566), .C2(n15565), .A(n6476), .B(n15597), .ZN(
        n15567) );
  INV_X1 U17131 ( .A(n15567), .ZN(n15568) );
  NAND3_X1 U17132 ( .A1(n15570), .A2(n15569), .A3(n15568), .ZN(P2_U3217) );
  INV_X1 U17133 ( .A(n15571), .ZN(n15573) );
  NAND3_X1 U17134 ( .A1(n15574), .A2(n15573), .A3(n15572), .ZN(n15575) );
  NAND2_X1 U17135 ( .A1(n15576), .A2(n15575), .ZN(n15581) );
  XNOR2_X1 U17136 ( .A(n15578), .B(n15577), .ZN(n15579) );
  AOI222_X1 U17137 ( .A1(n15581), .A2(n15613), .B1(n15580), .B2(n15587), .C1(
        n15579), .C2(n15610), .ZN(n15583) );
  OAI211_X1 U17138 ( .C1(n15584), .C2(n15618), .A(n15583), .B(n15582), .ZN(
        P2_U3226) );
  NAND2_X1 U17139 ( .A1(n15585), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n15590) );
  NAND2_X1 U17140 ( .A1(n15587), .A2(n15586), .ZN(n15588) );
  AND3_X1 U17141 ( .A1(n15590), .A2(n15589), .A3(n15588), .ZN(n15603) );
  AOI21_X1 U17142 ( .B1(n15593), .B2(n15592), .A(n15591), .ZN(n15595) );
  NAND2_X1 U17143 ( .A1(n15595), .A2(n15594), .ZN(n15602) );
  AOI211_X1 U17144 ( .C1(n15599), .C2(n15598), .A(n15597), .B(n15596), .ZN(
        n15600) );
  INV_X1 U17145 ( .A(n15600), .ZN(n15601) );
  NAND3_X1 U17146 ( .A1(n15603), .A2(n15602), .A3(n15601), .ZN(P2_U3227) );
  INV_X1 U17147 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15617) );
  XOR2_X1 U17148 ( .A(n15605), .B(n15604), .Z(n15611) );
  OAI21_X1 U17149 ( .B1(n15608), .B2(n15607), .A(n15606), .ZN(n15609) );
  AOI21_X1 U17150 ( .B1(n15611), .B2(n15610), .A(n15609), .ZN(n15616) );
  XOR2_X1 U17151 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n15612), .Z(n15614) );
  NAND2_X1 U17152 ( .A1(n15614), .A2(n15613), .ZN(n15615) );
  OAI211_X1 U17153 ( .C1(n15618), .C2(n15617), .A(n15616), .B(n15615), .ZN(
        P2_U3228) );
  OAI22_X1 U17154 ( .A1(n15622), .A2(n15621), .B1(n15620), .B2(n15619), .ZN(
        n15623) );
  AOI21_X1 U17155 ( .B1(n15625), .B2(n15624), .A(n15623), .ZN(n15626) );
  OAI21_X1 U17156 ( .B1(n15628), .B2(n15627), .A(n15626), .ZN(n15629) );
  AOI21_X1 U17157 ( .B1(n15631), .B2(n15630), .A(n15629), .ZN(n15632) );
  OAI21_X1 U17158 ( .B1(n14312), .B2(n15633), .A(n15632), .ZN(P2_U3258) );
  NOR2_X1 U17159 ( .A1(n15642), .A2(n15634), .ZN(n15639) );
  AND2_X1 U17160 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15637), .ZN(P2_U3266) );
  AND2_X1 U17161 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15637), .ZN(P2_U3267) );
  AND2_X1 U17162 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15637), .ZN(P2_U3268) );
  AND2_X1 U17163 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15637), .ZN(P2_U3269) );
  AND2_X1 U17164 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15637), .ZN(P2_U3270) );
  AND2_X1 U17165 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15637), .ZN(P2_U3271) );
  AND2_X1 U17166 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15637), .ZN(P2_U3272) );
  AND2_X1 U17167 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15637), .ZN(P2_U3273) );
  AND2_X1 U17168 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15637), .ZN(P2_U3274) );
  AND2_X1 U17169 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15637), .ZN(P2_U3275) );
  AND2_X1 U17170 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15637), .ZN(P2_U3276) );
  AND2_X1 U17171 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15637), .ZN(P2_U3277) );
  AND2_X1 U17172 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15637), .ZN(P2_U3278) );
  AND2_X1 U17173 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15637), .ZN(P2_U3279) );
  AND2_X1 U17174 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15637), .ZN(P2_U3280) );
  AND2_X1 U17175 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15637), .ZN(P2_U3281) );
  AND2_X1 U17176 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15637), .ZN(P2_U3282) );
  AND2_X1 U17177 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15637), .ZN(P2_U3283) );
  AND2_X1 U17178 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15637), .ZN(P2_U3284) );
  AND2_X1 U17179 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15637), .ZN(P2_U3285) );
  AND2_X1 U17180 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15637), .ZN(P2_U3286) );
  NOR2_X1 U17181 ( .A1(n15639), .A2(n15635), .ZN(P2_U3287) );
  NOR2_X1 U17182 ( .A1(n15639), .A2(n15636), .ZN(P2_U3288) );
  AND2_X1 U17183 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15637), .ZN(P2_U3289) );
  AND2_X1 U17184 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15637), .ZN(P2_U3290) );
  AND2_X1 U17185 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15637), .ZN(P2_U3291) );
  AND2_X1 U17186 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15637), .ZN(P2_U3292) );
  AND2_X1 U17187 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15637), .ZN(P2_U3293) );
  AND2_X1 U17188 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15637), .ZN(P2_U3294) );
  NOR2_X1 U17189 ( .A1(n15639), .A2(n15638), .ZN(P2_U3295) );
  AOI22_X1 U17190 ( .A1(n15645), .A2(n15641), .B1(n15640), .B2(n15642), .ZN(
        P2_U3416) );
  AOI22_X1 U17191 ( .A1(n15645), .A2(n15644), .B1(n15643), .B2(n15642), .ZN(
        P2_U3417) );
  INV_X1 U17192 ( .A(n15646), .ZN(n15652) );
  OAI21_X1 U17193 ( .B1(n15649), .B2(n15648), .A(n15647), .ZN(n15651) );
  AOI211_X1 U17194 ( .C1(n15653), .C2(n15652), .A(n15651), .B(n15650), .ZN(
        n15667) );
  INV_X1 U17195 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15654) );
  AOI22_X1 U17196 ( .A1(n15666), .A2(n15667), .B1(n15654), .B2(n15664), .ZN(
        P2_U3436) );
  INV_X1 U17197 ( .A(n15655), .ZN(n15659) );
  NAND2_X1 U17198 ( .A1(n15657), .A2(n15656), .ZN(n15658) );
  OAI211_X1 U17199 ( .C1(n15661), .C2(n15660), .A(n15659), .B(n15658), .ZN(
        n15662) );
  NOR2_X1 U17200 ( .A1(n15663), .A2(n15662), .ZN(n15669) );
  INV_X1 U17201 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15665) );
  AOI22_X1 U17202 ( .A1(n15666), .A2(n15669), .B1(n15665), .B2(n15664), .ZN(
        P2_U3442) );
  AOI22_X1 U17203 ( .A1(n15670), .A2(n15667), .B1(n8971), .B2(n15668), .ZN(
        P2_U3501) );
  AOI22_X1 U17204 ( .A1(n15670), .A2(n15669), .B1(n11073), .B2(n15668), .ZN(
        P2_U3503) );
  NOR2_X1 U17205 ( .A1(P3_U3897), .A2(n15671), .ZN(P3_U3150) );
  INV_X1 U17206 ( .A(n15672), .ZN(n15676) );
  OAI22_X1 U17207 ( .A1(n15676), .A2(n15675), .B1(n15674), .B2(n15673), .ZN(
        n15677) );
  AOI211_X1 U17208 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15685), .A(n15678), .B(
        n15677), .ZN(n15679) );
  AOI22_X1 U17209 ( .A1(n15691), .A2(n15680), .B1(n15679), .B2(n9345), .ZN(
        P3_U3231) );
  INV_X1 U17210 ( .A(n15681), .ZN(n15682) );
  AOI21_X1 U17211 ( .B1(n15684), .B2(n15683), .A(n15682), .ZN(n15690) );
  AOI22_X1 U17212 ( .A1(n15687), .A2(n15686), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15685), .ZN(n15688) );
  OAI221_X1 U17213 ( .B1(n15691), .B2(n15690), .C1(n9345), .C2(n15689), .A(
        n15688), .ZN(P3_U3232) );
  AOI22_X1 U17214 ( .A1(n15722), .A2(n15692), .B1(n8105), .B2(n15721), .ZN(
        P3_U3393) );
  INV_X1 U17215 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15693) );
  AOI22_X1 U17216 ( .A1(n15722), .A2(n15694), .B1(n15693), .B2(n15721), .ZN(
        P3_U3396) );
  INV_X1 U17217 ( .A(n15695), .ZN(n15696) );
  AOI211_X1 U17218 ( .C1(n15698), .C2(n15720), .A(n15697), .B(n15696), .ZN(
        n15724) );
  AOI22_X1 U17219 ( .A1(n15722), .A2(n15724), .B1(n8139), .B2(n15721), .ZN(
        P3_U3399) );
  NOR2_X1 U17220 ( .A1(n15715), .A2(n15699), .ZN(n15701) );
  AOI211_X1 U17221 ( .C1(n15702), .C2(n15720), .A(n15701), .B(n15700), .ZN(
        n15726) );
  AOI22_X1 U17222 ( .A1(n15722), .A2(n15726), .B1(n8154), .B2(n15721), .ZN(
        P3_U3402) );
  AOI22_X1 U17223 ( .A1(n15705), .A2(n15720), .B1(n15704), .B2(n15703), .ZN(
        n15706) );
  AND2_X1 U17224 ( .A1(n15707), .A2(n15706), .ZN(n15728) );
  INV_X1 U17225 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15708) );
  AOI22_X1 U17226 ( .A1(n15722), .A2(n15728), .B1(n15708), .B2(n15721), .ZN(
        P3_U3405) );
  NAND2_X1 U17227 ( .A1(n15709), .A2(n15720), .ZN(n15711) );
  NAND2_X1 U17228 ( .A1(n15711), .A2(n15710), .ZN(n15712) );
  NOR2_X1 U17229 ( .A1(n15713), .A2(n15712), .ZN(n15730) );
  INV_X1 U17230 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15714) );
  AOI22_X1 U17231 ( .A1(n15722), .A2(n15730), .B1(n15714), .B2(n15721), .ZN(
        P3_U3408) );
  NOR2_X1 U17232 ( .A1(n15716), .A2(n15715), .ZN(n15718) );
  AOI211_X1 U17233 ( .C1(n15720), .C2(n15719), .A(n15718), .B(n15717), .ZN(
        n15733) );
  AOI22_X1 U17234 ( .A1(n15722), .A2(n15733), .B1(n8199), .B2(n15721), .ZN(
        P3_U3411) );
  AOI22_X1 U17235 ( .A1(n15734), .A2(n15724), .B1(n15723), .B2(n15731), .ZN(
        P3_U3462) );
  AOI22_X1 U17236 ( .A1(n15734), .A2(n15726), .B1(n15725), .B2(n15731), .ZN(
        P3_U3463) );
  AOI22_X1 U17237 ( .A1(n15734), .A2(n15728), .B1(n15727), .B2(n15731), .ZN(
        P3_U3464) );
  AOI22_X1 U17238 ( .A1(n15734), .A2(n15730), .B1(n15729), .B2(n15731), .ZN(
        P3_U3465) );
  AOI22_X1 U17239 ( .A1(n15734), .A2(n15733), .B1(n15732), .B2(n15731), .ZN(
        P3_U3466) );
  XNOR2_X1 U17240 ( .A(n15736), .B(n15735), .ZN(n15737) );
  XNOR2_X1 U17241 ( .A(n15737), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  AOI21_X1 U17242 ( .B1(n15740), .B2(n15739), .A(n15738), .ZN(SUB_1596_U5) );
  INV_X1 U7187 ( .A(n8984), .ZN(n8970) );
  BUF_X2 U7213 ( .A(n10292), .Z(n10191) );
  NAND2_X1 U7217 ( .A1(n7278), .A2(n10019), .ZN(n7277) );
  CLKBUF_X2 U7224 ( .A(n8970), .Z(n9465) );
  CLKBUF_X1 U7358 ( .A(n8983), .Z(n9469) );
  CLKBUF_X1 U7359 ( .A(n8926), .Z(n11815) );
  CLKBUF_X1 U10264 ( .A(n8934), .Z(n11455) );
endmodule

