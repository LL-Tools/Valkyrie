

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9566, n9567, n9568, n9569, n9570, n9572, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
         n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234,
         n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
         n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
         n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
         n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
         n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
         n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282,
         n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
         n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
         n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306,
         n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314,
         n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
         n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
         n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338,
         n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346,
         n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354,
         n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
         n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
         n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378,
         n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386,
         n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
         n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
         n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410,
         n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418,
         n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426,
         n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434,
         n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
         n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450,
         n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
         n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466,
         n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474,
         n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482,
         n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490,
         n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498,
         n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506,
         n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
         n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522,
         n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530,
         n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538,
         n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546,
         n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554,
         n21555, n21556, n21557, n21558;

  INV_X1 U11010 ( .A(n20309), .ZN(n20253) );
  NOR2_X1 U11011 ( .A1(n17524), .A2(n18985), .ZN(n18675) );
  NAND2_X1 U11012 ( .A1(n9835), .A2(n20313), .ZN(n20366) );
  CLKBUF_X1 U11013 ( .A(n10691), .Z(n14624) );
  NAND2_X1 U11014 ( .A1(n14072), .A2(n20550), .ZN(n14194) );
  INV_X1 U11015 ( .A(n18583), .ZN(n10114) );
  NAND2_X1 U11016 ( .A1(n11319), .A2(n11318), .ZN(n11772) );
  OR2_X1 U11017 ( .A1(n13121), .A2(n13120), .ZN(n18985) );
  INV_X4 U11018 ( .A(n10620), .ZN(n11113) );
  NAND2_X1 U11019 ( .A1(n12281), .A2(n10592), .ZN(n12448) );
  AND2_X2 U11022 ( .A1(n10686), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10806) );
  CLKBUF_X2 U11023 ( .A(n10710), .Z(n14435) );
  CLKBUF_X2 U11024 ( .A(n10766), .Z(n9577) );
  CLKBUF_X1 U11025 ( .A(n14481), .Z(n9585) );
  NAND2_X1 U11027 ( .A1(n11462), .A2(n11461), .ZN(n12227) );
  NAND2_X1 U11028 ( .A1(n12534), .A2(n10323), .ZN(n10078) );
  AND2_X2 U11029 ( .A1(n9580), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10823) );
  INV_X1 U11030 ( .A(n17276), .ZN(n18107) );
  AND2_X1 U11032 ( .A1(n14618), .A2(n10551), .ZN(n14472) );
  CLKBUF_X3 U11033 ( .A(n10824), .Z(n9591) );
  CLKBUF_X2 U11034 ( .A(n11367), .Z(n11789) );
  CLKBUF_X2 U11035 ( .A(n11366), .Z(n12885) );
  CLKBUF_X2 U11036 ( .A(n11424), .Z(n11511) );
  CLKBUF_X2 U11037 ( .A(n11376), .Z(n12877) );
  CLKBUF_X2 U11038 ( .A(n11369), .Z(n12852) );
  CLKBUF_X2 U11039 ( .A(n11374), .Z(n12886) );
  CLKBUF_X2 U11040 ( .A(n11375), .Z(n12878) );
  INV_X1 U11041 ( .A(n18077), .ZN(n18008) );
  NAND2_X2 U11042 ( .A1(n10514), .A2(n10513), .ZN(n10594) );
  INV_X2 U11043 ( .A(n10598), .ZN(n10585) );
  NAND2_X1 U11044 ( .A1(n17221), .A2(n13000), .ZN(n9640) );
  INV_X1 U11045 ( .A(n9843), .ZN(n20763) );
  CLKBUF_X2 U11046 ( .A(n11430), .Z(n11431) );
  CLKBUF_X3 U11047 ( .A(n10560), .Z(n14630) );
  BUF_X1 U11048 ( .A(n10576), .Z(n10851) );
  AND2_X1 U11049 ( .A1(n9812), .A2(n10698), .ZN(n9924) );
  AND2_X1 U11050 ( .A1(n14618), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10811) );
  INV_X1 U11051 ( .A(n12004), .ZN(n12080) );
  NAND2_X1 U11052 ( .A1(n9845), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10067) );
  BUF_X1 U11054 ( .A(n10823), .Z(n9587) );
  INV_X1 U11055 ( .A(n9639), .ZN(n12477) );
  AND2_X1 U11056 ( .A1(n10851), .A2(n9641), .ZN(n10052) );
  INV_X1 U11057 ( .A(n11152), .ZN(n10629) );
  AND2_X1 U11058 ( .A1(n9581), .A2(n10551), .ZN(n14474) );
  INV_X1 U11059 ( .A(n13034), .ZN(n17322) );
  NOR2_X1 U11060 ( .A1(n20715), .A2(n20763), .ZN(n10178) );
  OR2_X1 U11061 ( .A1(n10899), .A2(n10597), .ZN(n11030) );
  AND2_X1 U11062 ( .A1(n10576), .A2(n12286), .ZN(n13148) );
  OR2_X1 U11063 ( .A1(n10817), .A2(n10816), .ZN(n12291) );
  BUF_X1 U11065 ( .A(n13228), .Z(n17329) );
  NAND2_X1 U11066 ( .A1(n10179), .A2(n10178), .ZN(n11979) );
  AND4_X1 U11067 ( .A1(n11350), .A2(n11349), .A3(n11348), .A4(n11347), .ZN(
        n11351) );
  OR2_X1 U11068 ( .A1(n11014), .A2(n11015), .ZN(n11020) );
  NAND2_X1 U11070 ( .A1(n15601), .A2(n15600), .ZN(n16438) );
  OR2_X1 U11071 ( .A1(n14353), .A2(n14356), .ZN(n16057) );
  INV_X1 U11072 ( .A(n20472), .ZN(n9823) );
  INV_X1 U11073 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13452) );
  AND2_X1 U11074 ( .A1(n13379), .A2(n13421), .ZN(n18868) );
  INV_X2 U11075 ( .A(n12726), .ZN(n13625) );
  INV_X1 U11076 ( .A(n14053), .ZN(n20733) );
  AND2_X1 U11077 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11594), .ZN(
        n11606) );
  XNOR2_X1 U11078 ( .A(n15162), .B(n15161), .ZN(n15351) );
  NAND2_X1 U11079 ( .A1(n13648), .A2(n13652), .ZN(n20679) );
  XNOR2_X1 U11080 ( .A(n11584), .B(n12122), .ZN(n21155) );
  CLKBUF_X3 U11081 ( .A(n13754), .Z(n15909) );
  INV_X1 U11082 ( .A(n16151), .ZN(n19647) );
  CLKBUF_X2 U11083 ( .A(n10592), .Z(n9596) );
  OAI21_X1 U11084 ( .B1(n19927), .B2(n19926), .A(n19925), .ZN(n19951) );
  INV_X1 U11085 ( .A(n20366), .ZN(n20352) );
  NAND2_X1 U11086 ( .A1(n12999), .A2(n17220), .ZN(n10445) );
  OR2_X1 U11087 ( .A1(n13217), .A2(n13216), .ZN(n13495) );
  OR2_X1 U11088 ( .A1(n13704), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n15937) );
  OR2_X1 U11089 ( .A1(n20246), .A2(n20091), .ZN(n20111) );
  NAND2_X2 U11090 ( .A1(n17524), .A2(n13748), .ZN(n18672) );
  AND2_X1 U11091 ( .A1(n10602), .A2(n12513), .ZN(n9566) );
  INV_X2 U11092 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13810) );
  AND2_X1 U11093 ( .A1(n9830), .A2(n9899), .ZN(n9567) );
  NAND2_X2 U11094 ( .A1(n13838), .A2(n13837), .ZN(n20680) );
  NAND2_X2 U11095 ( .A1(n12140), .A2(n12139), .ZN(n13838) );
  AND2_X1 U11096 ( .A1(n12996), .A2(n17220), .ZN(n9568) );
  AND2_X2 U11097 ( .A1(n12996), .A2(n17220), .ZN(n13361) );
  NAND2_X2 U11098 ( .A1(n10225), .A2(n10222), .ZN(n9968) );
  NAND2_X2 U11099 ( .A1(n10185), .A2(n9855), .ZN(n10225) );
  NOR2_X2 U11100 ( .A1(n13165), .A2(n13488), .ZN(n13286) );
  BUF_X2 U11101 ( .A(n10559), .Z(n14605) );
  NAND2_X2 U11102 ( .A1(n9957), .A2(n9958), .ZN(n12143) );
  NAND2_X2 U11103 ( .A1(n9956), .A2(n9959), .ZN(n9957) );
  NAND2_X2 U11104 ( .A1(n10115), .A2(n10073), .ZN(n14191) );
  AND2_X1 U11105 ( .A1(n12147), .A2(n12146), .ZN(n10115) );
  OAI21_X2 U11106 ( .B1(n11476), .B2(n11465), .A(n11467), .ZN(n10068) );
  OAI21_X2 U11107 ( .B1(n11396), .B2(n12222), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11476) );
  XNOR2_X2 U11108 ( .A(n13764), .B(n13762), .ZN(n13640) );
  NAND2_X1 U11109 ( .A1(n13780), .A2(n10677), .ZN(n19749) );
  AND2_X1 U11110 ( .A1(n10477), .A2(n14307), .ZN(n9569) );
  AND2_X2 U11111 ( .A1(n10477), .A2(n14307), .ZN(n9570) );
  AND2_X2 U11112 ( .A1(n10477), .A2(n14307), .ZN(n14628) );
  AND2_X4 U11113 ( .A1(n15991), .A2(n15993), .ZN(n15976) );
  NAND2_X2 U11115 ( .A1(n10474), .A2(n9643), .ZN(n11381) );
  NOR3_X2 U11116 ( .A1(n17232), .A2(n17987), .A3(n17994), .ZN(n17993) );
  AND2_X1 U11117 ( .A1(n10186), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9572) );
  AOI21_X2 U11118 ( .B1(n11440), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10183), 
        .ZN(n10182) );
  XNOR2_X2 U11119 ( .A(n9885), .B(n16697), .ZN(n16389) );
  AOI211_X2 U11120 ( .C1(n16957), .C2(n10160), .A(n17016), .B(n17021), .ZN(
        n17001) );
  OAI21_X1 U11121 ( .B1(n12806), .B2(n10374), .A(n10373), .ZN(n10372) );
  NOR2_X1 U11122 ( .A1(n14729), .A2(n14369), .ZN(n12906) );
  AND2_X1 U11123 ( .A1(n10050), .A2(n10338), .ZN(n11200) );
  CLKBUF_X1 U11124 ( .A(n12871), .Z(n11914) );
  OAI21_X1 U11125 ( .B1(n16320), .B2(n9893), .A(n9890), .ZN(n16270) );
  AOI21_X1 U11126 ( .B1(n9602), .B2(n10404), .A(n9660), .ZN(n10403) );
  OAI21_X1 U11127 ( .B1(n19987), .B2(n19986), .A(n19985), .ZN(n20005) );
  INV_X2 U11128 ( .A(n18681), .ZN(n18667) );
  NAND2_X2 U11129 ( .A1(n18426), .A2(n18530), .ZN(n18681) );
  XOR2_X1 U11130 ( .A(n11019), .B(n11020), .Z(n15604) );
  OR2_X1 U11131 ( .A1(n11020), .A2(n11019), .ZN(n11029) );
  INV_X1 U11132 ( .A(n20313), .ZN(n20458) );
  NAND2_X1 U11133 ( .A1(n13902), .A2(n13901), .ZN(n13903) );
  CLKBUF_X1 U11134 ( .A(n21228), .Z(n9778) );
  INV_X1 U11135 ( .A(n18672), .ZN(n18658) );
  NOR2_X1 U11136 ( .A1(n18536), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18506) );
  AND2_X1 U11137 ( .A1(n9975), .A2(n9973), .ZN(n11469) );
  NAND2_X2 U11138 ( .A1(n10922), .A2(n11030), .ZN(n10919) );
  NAND2_X1 U11139 ( .A1(n10637), .A2(n10638), .ZN(n10654) );
  NAND2_X1 U11140 ( .A1(n16419), .A2(n16747), .ZN(n16429) );
  NAND2_X1 U11141 ( .A1(n10005), .A2(n9981), .ZN(n9910) );
  NAND2_X1 U11142 ( .A1(n9810), .A2(n9808), .ZN(n10618) );
  NAND2_X1 U11143 ( .A1(n10898), .A2(n10897), .ZN(n10899) );
  NOR2_X1 U11144 ( .A1(n13381), .A2(n19405), .ZN(n13440) );
  CLKBUF_X2 U11145 ( .A(n10629), .Z(n11147) );
  MUX2_X1 U11146 ( .A(n10850), .B(n12484), .S(n12482), .Z(n11052) );
  AND2_X1 U11148 ( .A1(n16838), .A2(n18996), .ZN(n13418) );
  NAND2_X1 U11150 ( .A1(n11505), .A2(n11506), .ZN(n11976) );
  NAND2_X1 U11151 ( .A1(n11355), .A2(n11391), .ZN(n12220) );
  AND2_X1 U11152 ( .A1(n9673), .A2(n9824), .ZN(n13392) );
  NAND2_X1 U11153 ( .A1(n20757), .A2(n11391), .ZN(n11390) );
  INV_X1 U11154 ( .A(n11383), .ZN(n11355) );
  CLKBUF_X2 U11155 ( .A(n12286), .Z(n19806) );
  NAND2_X1 U11156 ( .A1(n12283), .A2(n20304), .ZN(n12287) );
  OR2_X1 U11157 ( .A1(n13071), .A2(n13070), .ZN(n19001) );
  NAND2_X1 U11158 ( .A1(n9843), .A2(n11385), .ZN(n14713) );
  AND2_X1 U11159 ( .A1(n11565), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11616) );
  CLKBUF_X2 U11161 ( .A(n10805), .Z(n9579) );
  INV_X4 U11162 ( .A(n17239), .ZN(n17293) );
  AND2_X1 U11163 ( .A1(n14596), .A2(n10551), .ZN(n10804) );
  AND2_X1 U11164 ( .A1(n14596), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10805) );
  CLKBUF_X2 U11165 ( .A(n11423), .Z(n11410) );
  CLKBUF_X2 U11166 ( .A(n11368), .Z(n12876) );
  CLKBUF_X2 U11167 ( .A(n12887), .Z(n11859) );
  INV_X1 U11168 ( .A(n13361), .ZN(n13478) );
  INV_X4 U11169 ( .A(n18077), .ZN(n17278) );
  BUF_X2 U11170 ( .A(n14472), .Z(n9588) );
  BUF_X2 U11171 ( .A(n12879), .Z(n12857) );
  INV_X4 U11172 ( .A(n10445), .ZN(n17330) );
  CLKBUF_X2 U11173 ( .A(n10560), .Z(n14596) );
  CLKBUF_X2 U11174 ( .A(n11432), .Z(n12880) );
  NAND2_X1 U11175 ( .A1(n12986), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14333) );
  INV_X4 U11176 ( .A(n9640), .ZN(n14312) );
  AND2_X1 U11177 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11594) );
  NOR2_X2 U11178 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17221) );
  NOR2_X1 U11179 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13000) );
  INV_X4 U11180 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10551) );
  XNOR2_X1 U11181 ( .A(n10074), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15361) );
  OR2_X1 U11182 ( .A1(n16555), .A2(n19706), .ZN(n9928) );
  AND2_X1 U11183 ( .A1(n12809), .A2(n10325), .ZN(n9984) );
  NAND4_X1 U11184 ( .A1(n10410), .A2(n10413), .A3(n10409), .A4(n10408), .ZN(
        n12769) );
  XNOR2_X1 U11185 ( .A(n10417), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15196) );
  XNOR2_X1 U11186 ( .A(n10018), .B(n14352), .ZN(n10053) );
  OR2_X1 U11187 ( .A1(n12700), .A2(n10407), .ZN(n10410) );
  NAND2_X1 U11188 ( .A1(n11200), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16515) );
  OAI21_X1 U11189 ( .B1(n16169), .B2(n16173), .A(n9819), .ZN(n10018) );
  AOI21_X1 U11190 ( .B1(n10103), .B2(n10375), .A(n16230), .ZN(n16234) );
  NAND2_X1 U11191 ( .A1(n9688), .A2(n10039), .ZN(n16451) );
  NAND2_X1 U11192 ( .A1(n12701), .A2(n10416), .ZN(n10414) );
  AND2_X1 U11193 ( .A1(n12589), .A2(n12588), .ZN(n9937) );
  OAI21_X1 U11194 ( .B1(n9605), .B2(n10348), .A(n9645), .ZN(n10347) );
  OAI21_X1 U11195 ( .B1(n11914), .B2(n14730), .A(n14729), .ZN(n15165) );
  NAND2_X1 U11196 ( .A1(n9900), .A2(n11196), .ZN(n10050) );
  XNOR2_X1 U11197 ( .A(n9807), .B(n16302), .ZN(n16611) );
  OAI21_X1 U11198 ( .B1(n12719), .B2(n12718), .A(n15324), .ZN(n9855) );
  AND2_X1 U11199 ( .A1(n10043), .A2(n10041), .ZN(n9605) );
  AOI211_X1 U11200 ( .C1(n19609), .C2(n15604), .A(n15603), .B(n15602), .ZN(
        n15605) );
  NAND2_X1 U11201 ( .A1(n12719), .A2(n15324), .ZN(n15218) );
  NAND2_X1 U11202 ( .A1(n10071), .A2(n10069), .ZN(n12719) );
  NOR2_X1 U11203 ( .A1(n16270), .A2(n16271), .ZN(n12606) );
  NAND2_X1 U11204 ( .A1(n10029), .A2(n10026), .ZN(n11006) );
  NAND3_X1 U11205 ( .A1(n10123), .A2(n9655), .A3(n9863), .ZN(n9862) );
  AOI21_X1 U11206 ( .B1(n12786), .B2(n9919), .A(n9917), .ZN(n12788) );
  AND2_X1 U11207 ( .A1(n10049), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10048) );
  AND2_X1 U11208 ( .A1(n9638), .A2(n16366), .ZN(n10194) );
  AND2_X1 U11209 ( .A1(n10338), .A2(n10051), .ZN(n10049) );
  NAND3_X1 U11210 ( .A1(n16333), .A2(n10908), .A3(n9599), .ZN(n10055) );
  AND2_X1 U11211 ( .A1(n10394), .A2(n10393), .ZN(n10392) );
  AND2_X1 U11212 ( .A1(n10338), .A2(n9772), .ZN(n10039) );
  NAND2_X1 U11213 ( .A1(n9800), .A2(n9796), .ZN(n20297) );
  NAND2_X1 U11214 ( .A1(n10116), .A2(n10403), .ZN(n15322) );
  AND2_X1 U11215 ( .A1(n16332), .A2(n16334), .ZN(n10908) );
  AOI21_X1 U11216 ( .B1(n9925), .B2(n11196), .A(n12570), .ZN(n10338) );
  XNOR2_X1 U11217 ( .A(n12737), .B(n12736), .ZN(n14379) );
  NOR2_X1 U11218 ( .A1(n9995), .A2(n17154), .ZN(n9994) );
  AND2_X1 U11219 ( .A1(n9799), .A2(n9797), .ZN(n9796) );
  NAND2_X1 U11220 ( .A1(n9935), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11184) );
  AND2_X1 U11221 ( .A1(n11194), .A2(n11192), .ZN(n16376) );
  OAI221_X1 U11222 ( .B1(n20894), .B2(n21000), .C1(n20894), .C2(n20879), .A(
        n21197), .ZN(n20897) );
  OR2_X1 U11223 ( .A1(n12732), .A2(n12089), .ZN(n14339) );
  XNOR2_X1 U11224 ( .A(n12756), .B(n11154), .ZN(n15946) );
  AND2_X1 U11225 ( .A1(n15247), .A2(n10117), .ZN(n9848) );
  OAI21_X1 U11226 ( .B1(n12755), .B2(n12757), .A(n12756), .ZN(n14687) );
  NAND2_X1 U11227 ( .A1(n10087), .A2(n15876), .ZN(n9885) );
  NAND2_X1 U11228 ( .A1(n9936), .A2(n11189), .ZN(n16397) );
  NAND2_X1 U11229 ( .A1(n12732), .A2(n14732), .ZN(n14731) );
  AND2_X1 U11230 ( .A1(n12195), .A2(n9849), .ZN(n15247) );
  INV_X4 U11231 ( .A(n20575), .ZN(n20560) );
  AOI21_X1 U11232 ( .B1(n9960), .B2(n12156), .A(n9680), .ZN(n9961) );
  INV_X1 U11233 ( .A(n14146), .ZN(n9858) );
  NOR2_X1 U11234 ( .A1(n15645), .A2(n15629), .ZN(n15630) );
  AND2_X2 U11235 ( .A1(n14787), .A2(n9736), .ZN(n12732) );
  AND2_X1 U11236 ( .A1(n14657), .A2(n11177), .ZN(n16414) );
  AND2_X1 U11237 ( .A1(n10219), .A2(n10004), .ZN(n12195) );
  XNOR2_X1 U11238 ( .A(n12155), .B(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9960) );
  OAI211_X1 U11239 ( .C1(n20208), .C2(n20188), .A(n20187), .B(n20253), .ZN(
        n20210) );
  NAND2_X1 U11240 ( .A1(n16989), .A2(n17180), .ZN(n17181) );
  AND2_X1 U11241 ( .A1(n14787), .A2(n9723), .ZN(n14745) );
  NAND2_X1 U11242 ( .A1(n10424), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10423) );
  NAND2_X1 U11243 ( .A1(n10416), .A2(n12198), .ZN(n10424) );
  NAND2_X1 U11244 ( .A1(n9623), .A2(n9831), .ZN(n11189) );
  NAND2_X1 U11245 ( .A1(n9867), .A2(n12154), .ZN(n12155) );
  NOR3_X2 U11246 ( .A1(n11024), .A2(n11190), .A3(n21478), .ZN(n16160) );
  NAND2_X1 U11247 ( .A1(n18399), .A2(n16935), .ZN(n18464) );
  NAND2_X1 U11248 ( .A1(n9881), .A2(n10106), .ZN(n18399) );
  INV_X1 U11249 ( .A(n20166), .ZN(n20175) );
  NAND2_X1 U11250 ( .A1(n11622), .A2(n11621), .ZN(n14244) );
  AOI21_X1 U11251 ( .B1(n15604), .B2(n11025), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16159) );
  NAND2_X1 U11252 ( .A1(n20962), .A2(n21189), .ZN(n20991) );
  NAND2_X1 U11253 ( .A1(n9880), .A2(n9760), .ZN(n10106) );
  NAND2_X1 U11254 ( .A1(n20834), .A2(n21189), .ZN(n20871) );
  NOR2_X2 U11255 ( .A1(n21244), .A2(n21190), .ZN(n21293) );
  AND2_X1 U11256 ( .A1(n9939), .A2(n9898), .ZN(n9831) );
  NAND2_X1 U11257 ( .A1(n9939), .A2(n10844), .ZN(n11168) );
  NOR2_X2 U11258 ( .A1(n20246), .A2(n20219), .ZN(n20242) );
  NAND2_X1 U11259 ( .A1(n11546), .A2(n11547), .ZN(n12148) );
  INV_X1 U11260 ( .A(n19844), .ZN(n19982) );
  OR2_X1 U11261 ( .A1(n20214), .A2(n20091), .ZN(n20123) );
  AOI21_X1 U11262 ( .B1(n12143), .B2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12144) );
  OAI211_X1 U11263 ( .C1(n15550), .C2(n11751), .A(n11599), .B(n11598), .ZN(
        n13960) );
  NAND2_X1 U11264 ( .A1(n20465), .A2(n19652), .ZN(n20214) );
  NAND2_X1 U11265 ( .A1(n20465), .A2(n16799), .ZN(n20246) );
  NAND2_X1 U11266 ( .A1(n18498), .A2(n17176), .ZN(n18808) );
  OR2_X1 U11267 ( .A1(n15547), .A2(n12134), .ZN(n12140) );
  XNOR2_X1 U11268 ( .A(n12176), .B(n11615), .ZN(n12165) );
  NAND2_X1 U11269 ( .A1(n11001), .A2(n11000), .ZN(n15639) );
  AND2_X1 U11270 ( .A1(n10365), .A2(n10093), .ZN(n10092) );
  NOR2_X1 U11271 ( .A1(n16458), .A2(n12577), .ZN(n9942) );
  INV_X1 U11272 ( .A(n20091), .ZN(n20078) );
  NOR2_X1 U11273 ( .A1(n15671), .A2(n11190), .ZN(n10994) );
  AND2_X1 U11274 ( .A1(n16635), .A2(n12571), .ZN(n16509) );
  NAND2_X1 U11275 ( .A1(n9823), .A2(n19739), .ZN(n20219) );
  AND2_X1 U11276 ( .A1(n9823), .A2(n20461), .ZN(n20313) );
  NAND2_X1 U11277 ( .A1(n18506), .A2(n18489), .ZN(n18488) );
  OR2_X1 U11278 ( .A1(n15653), .A2(n10992), .ZN(n15671) );
  NAND2_X1 U11279 ( .A1(n18680), .A2(n17151), .ZN(n18586) );
  AND2_X1 U11280 ( .A1(n16688), .A2(n12569), .ZN(n16635) );
  AND2_X1 U11281 ( .A1(n13761), .A2(n13767), .ZN(n13778) );
  NAND2_X1 U11282 ( .A1(n9876), .A2(n9875), .ZN(n18536) );
  OR3_X1 U11283 ( .A1(n18708), .A2(n18702), .A3(n17169), .ZN(n17203) );
  NAND2_X1 U11284 ( .A1(n13642), .A2(n13765), .ZN(n13779) );
  INV_X1 U11285 ( .A(n11571), .ZN(n11498) );
  OR2_X1 U11286 ( .A1(n13640), .A2(n13641), .ZN(n13643) );
  NOR2_X1 U11287 ( .A1(n20216), .A2(n10790), .ZN(n10791) );
  INV_X1 U11288 ( .A(n18543), .ZN(n9876) );
  AND2_X1 U11289 ( .A1(n13718), .A2(n13639), .ZN(n13641) );
  NOR2_X1 U11290 ( .A1(n15553), .A2(n9687), .ZN(n9852) );
  AND2_X1 U11291 ( .A1(n9696), .A2(n13720), .ZN(n10676) );
  NAND2_X1 U11292 ( .A1(n9612), .A2(n10659), .ZN(n20216) );
  AND2_X1 U11293 ( .A1(n13747), .A2(n13746), .ZN(n19421) );
  NAND2_X1 U11294 ( .A1(n10001), .A2(n9695), .ZN(n11496) );
  OR2_X1 U11295 ( .A1(n18568), .A2(n9627), .ZN(n18543) );
  AND2_X1 U11296 ( .A1(n10674), .A2(n13720), .ZN(n10677) );
  NAND2_X1 U11297 ( .A1(n18603), .A2(n16930), .ZN(n18568) );
  AND2_X1 U11298 ( .A1(n10353), .A2(n10659), .ZN(n10660) );
  AND2_X1 U11299 ( .A1(n10674), .A2(n16732), .ZN(n10657) );
  AND2_X2 U11300 ( .A1(n18792), .A2(n18298), .ZN(n19404) );
  NAND2_X1 U11301 ( .A1(n18792), .A2(n13397), .ZN(n19399) );
  AND2_X1 U11302 ( .A1(n9868), .A2(n9700), .ZN(n12115) );
  NOR2_X1 U11303 ( .A1(n16983), .A2(n16982), .ZN(n18598) );
  BUF_X2 U11304 ( .A(n10653), .Z(n19727) );
  AND2_X1 U11305 ( .A1(n16732), .A2(n15938), .ZN(n10353) );
  NAND2_X1 U11306 ( .A1(n12545), .A2(n14187), .ZN(n12587) );
  OR2_X1 U11307 ( .A1(n11469), .A2(n11471), .ZN(n11472) );
  OAI21_X1 U11308 ( .B1(n15938), .B2(n13632), .A(n13174), .ZN(n16758) );
  AND2_X1 U11309 ( .A1(n10947), .A2(n10250), .ZN(n10963) );
  NAND2_X1 U11310 ( .A1(n9787), .A2(n9786), .ZN(n16983) );
  NAND2_X1 U11311 ( .A1(n10644), .A2(n10654), .ZN(n15938) );
  CLKBUF_X1 U11312 ( .A(n10643), .Z(n10655) );
  NAND2_X1 U11313 ( .A1(n10640), .A2(n10639), .ZN(n10644) );
  NAND2_X1 U11314 ( .A1(n10080), .A2(n10626), .ZN(n10239) );
  NAND2_X1 U11315 ( .A1(n11468), .A2(n9910), .ZN(n20772) );
  NAND2_X1 U11316 ( .A1(n9971), .A2(n11460), .ZN(n9977) );
  CLKBUF_X1 U11317 ( .A(n10641), .Z(n10642) );
  NAND2_X1 U11318 ( .A1(n13384), .A2(n13383), .ZN(n18958) );
  NOR2_X1 U11319 ( .A1(n14662), .A2(n15882), .ZN(n12316) );
  NAND2_X1 U11320 ( .A1(n13806), .A2(n15978), .ZN(n14151) );
  OR2_X1 U11321 ( .A1(n10618), .A2(n10617), .ZN(n10619) );
  XNOR2_X1 U11322 ( .A(n10618), .B(n10616), .ZN(n10641) );
  NAND2_X1 U11323 ( .A1(n11321), .A2(n11320), .ZN(n11854) );
  INV_X1 U11324 ( .A(n11852), .ZN(n11321) );
  OAI211_X1 U11325 ( .C1(n11150), .C2(n16715), .A(n10631), .B(n10630), .ZN(
        n13772) );
  NAND2_X1 U11326 ( .A1(n14255), .A2(n14254), .ZN(n15934) );
  NAND2_X1 U11327 ( .A1(n12305), .A2(n12304), .ZN(n14664) );
  NAND3_X2 U11328 ( .A1(n18297), .A2(n18295), .A3(n18298), .ZN(n18355) );
  OR2_X1 U11329 ( .A1(n13440), .A2(n13094), .ZN(n13180) );
  CLKBUF_X1 U11330 ( .A(n10623), .Z(n10632) );
  NAND2_X1 U11331 ( .A1(n13198), .A2(n13433), .ZN(n16808) );
  NAND2_X1 U11332 ( .A1(n13926), .A2(n13925), .ZN(n13928) );
  OR2_X1 U11333 ( .A1(n14195), .A2(n17396), .ZN(n10334) );
  NAND2_X1 U11334 ( .A1(n9649), .A2(n18978), .ZN(n13198) );
  OR2_X1 U11335 ( .A1(n10620), .A2(n10612), .ZN(n10614) );
  OAI211_X1 U11336 ( .C1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n13240), .A(
        n11997), .B(n11996), .ZN(n12000) );
  OAI21_X1 U11337 ( .B1(n9593), .B2(n10612), .A(n12288), .ZN(n12294) );
  CLKBUF_X1 U11338 ( .A(n12508), .Z(n15586) );
  AOI21_X1 U11339 ( .B1(n13073), .B2(n13072), .A(n13418), .ZN(n13194) );
  INV_X1 U11340 ( .A(n12448), .ZN(n12431) );
  NOR2_X1 U11341 ( .A1(n11441), .A2(n10072), .ZN(n12174) );
  NAND2_X1 U11342 ( .A1(n10188), .A2(n10052), .ZN(n10190) );
  NAND2_X1 U11343 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17067), .ZN(
        n18372) );
  NAND2_X1 U11344 ( .A1(n12782), .A2(n12726), .ZN(n12729) );
  INV_X2 U11345 ( .A(n12287), .ZN(n9598) );
  INV_X1 U11346 ( .A(n12554), .ZN(n12504) );
  AND2_X1 U11347 ( .A1(n10590), .A2(n12499), .ZN(n10130) );
  NAND2_X1 U11348 ( .A1(n13392), .A2(n19001), .ZN(n13073) );
  CLKBUF_X2 U11349 ( .A(n11355), .Z(n20747) );
  OR2_X1 U11351 ( .A1(n11390), .A2(n11386), .ZN(n12212) );
  AND2_X1 U11352 ( .A1(n9701), .A2(n11993), .ZN(n11961) );
  OR2_X1 U11353 ( .A1(n11422), .A2(n11421), .ZN(n12169) );
  OR2_X1 U11354 ( .A1(n10776), .A2(n10775), .ZN(n10865) );
  CLKBUF_X1 U11355 ( .A(n10589), .Z(n19777) );
  INV_X1 U11356 ( .A(n10584), .ZN(n12512) );
  NAND2_X1 U11357 ( .A1(n9575), .A2(n12124), .ZN(n11995) );
  OR2_X1 U11358 ( .A1(n10841), .A2(n10840), .ZN(n10850) );
  NAND2_X1 U11359 ( .A1(n9646), .A2(n9608), .ZN(n10352) );
  NAND2_X1 U11360 ( .A1(n20742), .A2(n9953), .ZN(n14010) );
  OR2_X1 U11361 ( .A1(n13367), .A2(n13366), .ZN(n13404) );
  OR2_X1 U11362 ( .A1(n11438), .A2(n11437), .ZN(n12123) );
  NAND2_X1 U11363 ( .A1(n10490), .A2(n10489), .ZN(n10589) );
  AND4_X1 U11364 ( .A1(n10724), .A2(n10723), .A3(n10722), .A4(n10721), .ZN(
        n10739) );
  NAND2_X2 U11365 ( .A1(n10502), .A2(n10501), .ZN(n10593) );
  NOR2_X1 U11366 ( .A1(n18518), .A2(n18520), .ZN(n17745) );
  NAND2_X1 U11367 ( .A1(n10463), .A2(n10488), .ZN(n10489) );
  NAND3_X2 U11368 ( .A1(n9676), .A2(n10475), .A3(n11300), .ZN(n9843) );
  NAND2_X1 U11369 ( .A1(n11616), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11633) );
  AND3_X1 U11370 ( .A1(n11297), .A2(n11299), .A3(n11298), .ZN(n9676) );
  CLKBUF_X3 U11371 ( .A(n10804), .Z(n9578) );
  AND4_X1 U11372 ( .A1(n11338), .A2(n11337), .A3(n11336), .A4(n11335), .ZN(
        n11354) );
  NOR2_X2 U11373 ( .A1(n20709), .A2(n20712), .ZN(n20710) );
  AND4_X1 U11374 ( .A1(n11346), .A2(n11345), .A3(n11344), .A4(n11343), .ZN(
        n11352) );
  AOI21_X1 U11375 ( .B1(n14596), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n10255), .ZN(n10254) );
  BUF_X2 U11376 ( .A(n13207), .Z(n18061) );
  NAND2_X2 U11377 ( .A1(n19531), .A2(n19466), .ZN(n19522) );
  BUF_X2 U11378 ( .A(n13207), .Z(n17323) );
  AND4_X1 U11379 ( .A1(n10481), .A2(n10480), .A3(n10479), .A4(n10478), .ZN(
        n10482) );
  AND4_X1 U11380 ( .A1(n11304), .A2(n11303), .A3(n11302), .A4(n11301), .ZN(
        n11312) );
  NAND2_X2 U11381 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20446), .ZN(n20444) );
  AND2_X2 U11382 ( .A1(n14560), .A2(n10551), .ZN(n14479) );
  INV_X1 U11383 ( .A(n13507), .ZN(n18006) );
  CLKBUF_X3 U11384 ( .A(n10811), .Z(n9592) );
  INV_X2 U11385 ( .A(n17509), .ZN(U215) );
  BUF_X2 U11386 ( .A(n11412), .Z(n11425) );
  AOI22_X1 U11387 ( .A1(n14629), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10564) );
  INV_X1 U11388 ( .A(n14088), .ZN(n14604) );
  BUF_X2 U11389 ( .A(n10559), .Z(n14629) );
  INV_X2 U11390 ( .A(n17512), .ZN(n17514) );
  NAND2_X2 U11391 ( .A1(n13809), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14088) );
  AND2_X2 U11392 ( .A1(n14104), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10560) );
  AND2_X2 U11393 ( .A1(n13994), .A2(n14013), .ZN(n12879) );
  AND2_X2 U11394 ( .A1(n14014), .A2(n13994), .ZN(n11374) );
  AND2_X1 U11395 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10477) );
  AND2_X2 U11396 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13809) );
  AND2_X2 U11397 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14013) );
  NOR2_X2 U11398 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14014) );
  AND2_X2 U11399 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13978) );
  INV_X2 U11400 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17217) );
  INV_X1 U11401 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19391) );
  NOR2_X1 U11402 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13426) );
  NAND2_X1 U11403 ( .A1(n10604), .A2(n12534), .ZN(n10620) );
  INV_X1 U11404 ( .A(n12534), .ZN(n10006) );
  OAI21_X1 U11405 ( .B1(n10795), .B2(n10742), .A(n9983), .ZN(n10743) );
  NAND2_X2 U11406 ( .A1(n11389), .A2(n11388), .ZN(n11399) );
  OR2_X1 U11407 ( .A1(n10799), .A2(n10798), .ZN(n10800) );
  INV_X2 U11408 ( .A(n11385), .ZN(n20757) );
  NAND2_X1 U11409 ( .A1(n10676), .A2(n15909), .ZN(n20183) );
  AND3_X4 U11410 ( .A1(n12909), .A2(P1_STATE2_REG_1__SCAN_IN), .A3(n20562), 
        .ZN(n20575) );
  XNOR2_X1 U11411 ( .A(n11917), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12909) );
  NOR2_X2 U11412 ( .A1(n10066), .A2(n10061), .ZN(n10065) );
  NOR3_X2 U11413 ( .A1(n18118), .A2(n13135), .A3(n17779), .ZN(n9653) );
  NAND2_X1 U11414 ( .A1(n13780), .A2(n10676), .ZN(n19919) );
  NAND2_X1 U11415 ( .A1(n13780), .A2(n10660), .ZN(n19977) );
  OAI211_X2 U11416 ( .C1(n20838), .C2(n9706), .A(n9838), .B(n11481), .ZN(
        n13307) );
  NAND2_X1 U11417 ( .A1(n10666), .A2(n9861), .ZN(n10795) );
  NAND2_X1 U11418 ( .A1(n10065), .A2(n10064), .ZN(n9575) );
  NAND2_X1 U11419 ( .A1(n10065), .A2(n10064), .ZN(n9576) );
  NOR2_X2 U11420 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17693), .ZN(n17678) );
  NAND2_X2 U11421 ( .A1(n10220), .A2(n20838), .ZN(n11475) );
  AOI21_X2 U11422 ( .B1(n11068), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10615), .ZN(n10616) );
  AND2_X4 U11423 ( .A1(n11207), .A2(n14007), .ZN(n11412) );
  NAND2_X2 U11424 ( .A1(n10550), .A2(n10549), .ZN(n10584) );
  AND2_X2 U11425 ( .A1(n14354), .A2(n14355), .ZN(n14353) );
  NOR2_X2 U11426 ( .A1(n15649), .A2(n10396), .ZN(n14354) );
  NAND2_X2 U11427 ( .A1(n9658), .A2(n11388), .ZN(n13300) );
  OR2_X2 U11428 ( .A1(n14809), .A2(n14797), .ZN(n14795) );
  NOR2_X2 U11429 ( .A1(n17064), .A2(n17710), .ZN(n18403) );
  AND2_X1 U11430 ( .A1(n10646), .A2(n13754), .ZN(n9861) );
  NOR2_X2 U11431 ( .A1(n20742), .A2(n11381), .ZN(n12117) );
  INV_X2 U11432 ( .A(n12124), .ZN(n20742) );
  OR2_X1 U11433 ( .A1(n12222), .A2(n11464), .ZN(n9845) );
  NAND2_X2 U11434 ( .A1(n11992), .A2(n20562), .ZN(n17350) );
  NOR2_X2 U11435 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17601), .ZN(n17587) );
  OR2_X1 U11436 ( .A1(n15547), .A2(n15553), .ZN(n21244) );
  NAND2_X2 U11437 ( .A1(n11572), .A2(n11593), .ZN(n15547) );
  NOR2_X2 U11438 ( .A1(n14932), .A2(n10329), .ZN(n14887) );
  NAND2_X2 U11439 ( .A1(n14968), .A2(n14952), .ZN(n14932) );
  NOR2_X2 U11440 ( .A1(n14066), .A2(n15772), .ZN(n12799) );
  AND2_X1 U11441 ( .A1(n9570), .A2(n10551), .ZN(n10766) );
  INV_X2 U11442 ( .A(n14088), .ZN(n9580) );
  INV_X1 U11443 ( .A(n14088), .ZN(n9581) );
  INV_X1 U11444 ( .A(n9581), .ZN(n9582) );
  CLKBUF_X1 U11445 ( .A(n14481), .Z(n9583) );
  AND2_X1 U11446 ( .A1(n9569), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14481) );
  AND2_X1 U11447 ( .A1(n14625), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10824) );
  NOR2_X2 U11448 ( .A1(n14194), .A2(n10332), .ZN(n14245) );
  INV_X1 U11449 ( .A(n12480), .ZN(n9593) );
  NOR2_X2 U11450 ( .A1(n14890), .A2(n14875), .ZN(n14853) );
  NOR3_X4 U11451 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17896) );
  BUF_X4 U11452 ( .A(n10592), .Z(n9595) );
  AND2_X4 U11453 ( .A1(n14560), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10699) );
  BUF_X4 U11454 ( .A(n10559), .Z(n14560) );
  INV_X1 U11455 ( .A(n12287), .ZN(n9597) );
  NAND2_X1 U11456 ( .A1(n16838), .A2(n13392), .ZN(n13072) );
  AND2_X1 U11457 ( .A1(n10027), .A2(n10054), .ZN(n9846) );
  AND2_X1 U11458 ( .A1(n10031), .A2(n16202), .ZN(n10027) );
  INV_X1 U11459 ( .A(n10423), .ZN(n10184) );
  NAND2_X1 U11460 ( .A1(n12695), .A2(n10416), .ZN(n10002) );
  INV_X1 U11461 ( .A(n11610), .ZN(n9851) );
  AOI21_X1 U11462 ( .B1(n13194), .B2(n19554), .A(n13193), .ZN(n13395) );
  INV_X1 U11463 ( .A(n13982), .ZN(n13297) );
  AOI21_X1 U11464 ( .B1(n9920), .B2(n12218), .A(n14227), .ZN(n12250) );
  INV_X1 U11465 ( .A(n10198), .ZN(n9920) );
  AOI21_X1 U11466 ( .B1(n14213), .B2(n12217), .A(n13299), .ZN(n12218) );
  OAI21_X1 U11467 ( .B1(n14213), .B2(n10200), .A(n10199), .ZN(n10198) );
  AOI22_X1 U11468 ( .A1(n13806), .A2(n12511), .B1(n12948), .B2(n12510), .ZN(
        n13825) );
  INV_X1 U11469 ( .A(n13808), .ZN(n12511) );
  INV_X1 U11470 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U11471 ( .A1(n9861), .A2(n9886), .ZN(n9982) );
  NOR2_X1 U11472 ( .A1(n10659), .A2(n9887), .ZN(n9886) );
  NAND2_X1 U11473 ( .A1(n11949), .A2(n11948), .ZN(n11957) );
  XNOR2_X1 U11474 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11956) );
  AND2_X1 U11475 ( .A1(n11498), .A2(n11600), .ZN(n9874) );
  INV_X1 U11476 ( .A(n12184), .ZN(n10405) );
  XNOR2_X1 U11477 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11050) );
  AND3_X2 U11478 ( .A1(n10868), .A2(n13810), .A3(n10169), .ZN(n10559) );
  INV_X1 U11479 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U11480 ( .A1(n11113), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10622) );
  NAND2_X1 U11481 ( .A1(n9791), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10606) );
  OR2_X1 U11482 ( .A1(n10599), .A2(n10573), .ZN(n9792) );
  INV_X1 U11483 ( .A(n9828), .ZN(n13373) );
  AND3_X2 U11484 ( .A1(n17217), .A2(n19391), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12991) );
  NOR2_X1 U11485 ( .A1(n11391), .A2(n11383), .ZN(n13243) );
  NAND2_X1 U11486 ( .A1(n14899), .A2(n10440), .ZN(n14791) );
  AND2_X1 U11487 ( .A1(n11869), .A2(n10441), .ZN(n10440) );
  AND2_X1 U11488 ( .A1(n14807), .A2(n12703), .ZN(n11869) );
  OR2_X1 U11489 ( .A1(n14911), .A2(n14912), .ZN(n14942) );
  INV_X1 U11490 ( .A(n12902), .ZN(n11910) );
  OR2_X1 U11491 ( .A1(n11385), .A2(n21239), .ZN(n11751) );
  INV_X1 U11492 ( .A(n11751), .ZN(n11727) );
  INV_X1 U11493 ( .A(n12904), .ZN(n12900) );
  NAND2_X1 U11494 ( .A1(n10420), .A2(n10416), .ZN(n15177) );
  NOR2_X1 U11495 ( .A1(n10423), .A2(n10422), .ZN(n10421) );
  INV_X1 U11496 ( .A(n15241), .ZN(n10422) );
  NOR2_X1 U11497 ( .A1(n14923), .A2(n14935), .ZN(n10330) );
  NAND2_X1 U11498 ( .A1(n12148), .A2(n13462), .ZN(n9867) );
  OR2_X1 U11499 ( .A1(n11517), .A2(n11516), .ZN(n12149) );
  AND2_X1 U11500 ( .A1(n11601), .A2(n13462), .ZN(n9956) );
  NOR2_X1 U11501 ( .A1(n11383), .A2(n10072), .ZN(n11492) );
  INV_X1 U11502 ( .A(n10067), .ZN(n9844) );
  NAND2_X1 U11503 ( .A1(n11499), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9837) );
  NAND2_X1 U11504 ( .A1(n9974), .A2(n11444), .ZN(n9973) );
  INV_X1 U11505 ( .A(n10182), .ZN(n9974) );
  INV_X1 U11506 ( .A(n14010), .ZN(n13980) );
  NAND2_X1 U11507 ( .A1(n11504), .A2(n11503), .ZN(n20872) );
  INV_X1 U11508 ( .A(n20775), .ZN(n20878) );
  OR2_X1 U11509 ( .A1(n11166), .A2(n12482), .ZN(n10863) );
  INV_X1 U11510 ( .A(n16237), .ZN(n10315) );
  NAND2_X1 U11511 ( .A1(n9617), .A2(n11085), .ZN(n10246) );
  NAND2_X1 U11512 ( .A1(n16146), .A2(n10388), .ZN(n10386) );
  NOR2_X1 U11513 ( .A1(n15593), .A2(n10233), .ZN(n10231) );
  AOI21_X1 U11514 ( .B1(n10092), .B2(n10095), .A(n9689), .ZN(n10091) );
  INV_X1 U11515 ( .A(n10092), .ZN(n9892) );
  NAND2_X1 U11516 ( .A1(n10028), .A2(n10034), .ZN(n10996) );
  NOR2_X1 U11517 ( .A1(n15635), .A2(n15650), .ZN(n10397) );
  NAND2_X1 U11518 ( .A1(n10030), .A2(n16202), .ZN(n10029) );
  NAND2_X1 U11519 ( .A1(n9846), .A2(n10055), .ZN(n10026) );
  INV_X1 U11520 ( .A(n10034), .ZN(n10030) );
  INV_X1 U11521 ( .A(n15721), .ZN(n10399) );
  NOR2_X1 U11522 ( .A1(n10367), .A2(n10097), .ZN(n10096) );
  INV_X1 U11523 ( .A(n10370), .ZN(n10097) );
  OR2_X1 U11524 ( .A1(n14267), .A2(n11190), .ZN(n10959) );
  NAND2_X1 U11525 ( .A1(n9927), .A2(n9926), .ZN(n11194) );
  AND2_X1 U11526 ( .A1(n10779), .A2(n11025), .ZN(n9926) );
  AND2_X1 U11527 ( .A1(n10844), .A2(n11166), .ZN(n9898) );
  AND2_X1 U11528 ( .A1(n10844), .A2(n9908), .ZN(n9897) );
  AND2_X1 U11529 ( .A1(n11166), .A2(n11167), .ZN(n9908) );
  NAND2_X1 U11530 ( .A1(n9678), .A2(n14120), .ZN(n10611) );
  NAND2_X1 U11531 ( .A1(n9834), .A2(n13758), .ZN(n13760) );
  NAND2_X1 U11532 ( .A1(n18616), .A2(n16925), .ZN(n17085) );
  OR2_X1 U11533 ( .A1(n16916), .A2(n16962), .ZN(n16923) );
  OAI21_X1 U11534 ( .B1(n13092), .B2(n13091), .A(n13184), .ZN(n13389) );
  INV_X1 U11535 ( .A(n13073), .ZN(n13399) );
  NAND2_X1 U11536 ( .A1(n10225), .A2(n10224), .ZN(n10076) );
  NOR2_X1 U11537 ( .A1(n10221), .A2(n9686), .ZN(n9967) );
  NOR2_X1 U11538 ( .A1(n12721), .A2(n9726), .ZN(n10222) );
  NOR3_X1 U11539 ( .A1(n15381), .A2(n12256), .A3(n12255), .ZN(n12916) );
  AND2_X1 U11540 ( .A1(n12699), .A2(n10412), .ZN(n10411) );
  AND2_X1 U11541 ( .A1(n10415), .A2(n12201), .ZN(n10412) );
  NAND2_X1 U11542 ( .A1(n10414), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10407) );
  AND2_X1 U11543 ( .A1(n14054), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13609) );
  NAND2_X1 U11544 ( .A1(n11976), .A2(n11981), .ZN(n11977) );
  NAND2_X1 U11545 ( .A1(n11975), .A2(n11974), .ZN(n11978) );
  AND2_X1 U11546 ( .A1(n14650), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14054) );
  OR2_X1 U11547 ( .A1(n10982), .A2(n10964), .ZN(n15709) );
  AND2_X1 U11548 ( .A1(n9662), .A2(n15770), .ZN(n10235) );
  AND2_X1 U11549 ( .A1(n10050), .A2(n10049), .ZN(n14346) );
  AND2_X1 U11550 ( .A1(n10979), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16232) );
  NAND2_X1 U11551 ( .A1(n12612), .A2(n16243), .ZN(n10376) );
  NAND2_X1 U11552 ( .A1(n10100), .A2(n12609), .ZN(n10103) );
  XNOR2_X1 U11553 ( .A(n16758), .B(n13637), .ZN(n13717) );
  NAND2_X1 U11554 ( .A1(n12532), .A2(n12497), .ZN(n13806) );
  OR2_X1 U11555 ( .A1(n20465), .A2(n19652), .ZN(n19844) );
  OR2_X1 U11556 ( .A1(n20465), .A2(n16799), .ZN(n20017) );
  NAND2_X1 U11557 ( .A1(n20472), .A2(n19739), .ZN(n20091) );
  INV_X1 U11558 ( .A(n20259), .ZN(n20256) );
  OR2_X1 U11559 ( .A1(n20259), .A2(n20258), .ZN(n9799) );
  INV_X1 U11560 ( .A(n20128), .ZN(n20309) );
  AND4_X1 U11561 ( .A1(n13419), .A2(n13196), .A3(n18157), .A4(n13189), .ZN(
        n13094) );
  AND3_X1 U11562 ( .A1(n13108), .A2(n9659), .A3(n13107), .ZN(n19554) );
  AND3_X1 U11563 ( .A1(n13106), .A2(n13105), .A3(n13104), .ZN(n13107) );
  AND4_X1 U11564 ( .A1(n13099), .A2(n13098), .A3(n13097), .A4(n13096), .ZN(
        n13108) );
  OR2_X1 U11565 ( .A1(n14042), .A2(n14227), .ZN(n15339) );
  NAND2_X1 U11566 ( .A1(n12533), .A2(n11056), .ZN(n19579) );
  NAND2_X1 U11567 ( .A1(n10125), .A2(n10127), .ZN(n16554) );
  NAND2_X1 U11568 ( .A1(n9648), .A2(n9567), .ZN(n10125) );
  AND2_X1 U11569 ( .A1(n16419), .A2(n14342), .ZN(n16425) );
  AND2_X1 U11570 ( .A1(n12763), .A2(n12762), .ZN(n12764) );
  OR2_X1 U11571 ( .A1(n14687), .A2(n19728), .ZN(n12763) );
  AND2_X1 U11572 ( .A1(n9567), .A2(n19721), .ZN(n9930) );
  INV_X1 U11573 ( .A(n16553), .ZN(n10126) );
  NAND2_X1 U11574 ( .A1(n19444), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n17518) );
  AND2_X1 U11575 ( .A1(n19727), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n9889) );
  NAND2_X1 U11576 ( .A1(n9612), .A2(n9989), .ZN(n9988) );
  NOR2_X1 U11577 ( .A1(n10666), .A2(n9990), .ZN(n9989) );
  INV_X1 U11578 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n9990) );
  NAND2_X1 U11579 ( .A1(n10666), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n9894) );
  AND2_X1 U11580 ( .A1(n19727), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n9888) );
  NAND2_X1 U11581 ( .A1(n20752), .A2(n11385), .ZN(n9955) );
  OR2_X1 U11582 ( .A1(n11542), .A2(n11541), .ZN(n12159) );
  NAND2_X1 U11583 ( .A1(n11961), .A2(n13462), .ZN(n11966) );
  AOI21_X1 U11584 ( .B1(n11952), .B2(n11951), .A(n11950), .ZN(n9916) );
  NAND2_X1 U11585 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n14489) );
  INV_X1 U11586 ( .A(n10607), .ZN(n10604) );
  NOR2_X1 U11587 ( .A1(n12595), .A2(n12597), .ZN(n12594) );
  AOI21_X1 U11588 ( .B1(n15584), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10624) );
  NOR2_X1 U11589 ( .A1(n10035), .A2(n9679), .ZN(n10034) );
  INV_X1 U11590 ( .A(n16203), .ZN(n10035) );
  AND2_X1 U11591 ( .A1(n10684), .A2(n10683), .ZN(n9811) );
  NAND2_X1 U11592 ( .A1(n12553), .A2(n10458), .ZN(n10342) );
  NAND2_X1 U11593 ( .A1(n9566), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10458) );
  NAND2_X1 U11594 ( .A1(n10603), .A2(n10345), .ZN(n10344) );
  NAND2_X1 U11595 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10345) );
  AOI21_X1 U11596 ( .B1(n14108), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10168), 
        .ZN(n9808) );
  AND2_X1 U11597 ( .A1(n14136), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10168) );
  AND2_X1 U11598 ( .A1(n14122), .A2(n12558), .ZN(n10131) );
  NAND2_X1 U11599 ( .A1(n10193), .A2(n10192), .ZN(n12537) );
  NAND2_X1 U11600 ( .A1(n12501), .A2(n19777), .ZN(n10192) );
  INV_X2 U11601 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10868) );
  NAND2_X1 U11602 ( .A1(n10848), .A2(n10847), .ZN(n10855) );
  AND2_X2 U11603 ( .A1(n10582), .A2(n13148), .ZN(n12534) );
  NOR2_X1 U11604 ( .A1(n10470), .A2(n11575), .ZN(n11576) );
  INV_X1 U11605 ( .A(n11390), .ZN(n13611) );
  NAND2_X1 U11606 ( .A1(n14780), .A2(n9667), .ZN(n11913) );
  INV_X1 U11607 ( .A(n14781), .ZN(n11887) );
  NOR2_X2 U11608 ( .A1(n14911), .A2(n11754), .ZN(n14899) );
  OR2_X1 U11609 ( .A1(n11753), .A2(n14913), .ZN(n11754) );
  NAND2_X1 U11610 ( .A1(n9756), .A2(n10436), .ZN(n10435) );
  INV_X1 U11611 ( .A(n15056), .ZN(n10436) );
  INV_X1 U11612 ( .A(n14746), .ZN(n10335) );
  AND2_X1 U11613 ( .A1(n12199), .A2(n10070), .ZN(n10069) );
  INV_X1 U11614 ( .A(n15242), .ZN(n10071) );
  AND2_X1 U11615 ( .A1(n12201), .A2(n12200), .ZN(n10070) );
  NOR2_X1 U11616 ( .A1(n10416), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10415) );
  NOR2_X1 U11617 ( .A1(n15332), .A2(n12192), .ZN(n10118) );
  INV_X1 U11618 ( .A(n15258), .ZN(n10004) );
  INV_X1 U11619 ( .A(n14932), .ZN(n10331) );
  INV_X1 U11620 ( .A(n17359), .ZN(n10404) );
  INV_X1 U11621 ( .A(n12085), .ZN(n12060) );
  INV_X1 U11622 ( .A(n11308), .ZN(n11309) );
  AOI22_X1 U11623 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11411), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11307) );
  NAND2_X1 U11624 ( .A1(n9859), .A2(n11397), .ZN(n10005) );
  AND3_X1 U11625 ( .A1(n11459), .A2(n11458), .A3(n11457), .ZN(n11470) );
  NOR2_X1 U11626 ( .A1(n11491), .A2(n11490), .ZN(n12135) );
  INV_X1 U11627 ( .A(n11961), .ZN(n11958) );
  INV_X1 U11628 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21123) );
  NAND2_X1 U11629 ( .A1(n20720), .A2(n10072), .ZN(n11519) );
  NOR2_X1 U11630 ( .A1(n10242), .A2(n10241), .ZN(n10240) );
  INV_X1 U11631 ( .A(n10461), .ZN(n10242) );
  NOR2_X1 U11632 ( .A1(n15745), .A2(n10294), .ZN(n10293) );
  AND2_X1 U11633 ( .A1(n10903), .A2(n10904), .ZN(n10897) );
  NAND2_X1 U11634 ( .A1(n10597), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10864) );
  NAND2_X1 U11635 ( .A1(n10853), .A2(n10852), .ZN(n10876) );
  AND2_X1 U11636 ( .A1(n15959), .A2(n14612), .ZN(n10267) );
  AND2_X1 U11637 ( .A1(n9728), .A2(n16004), .ZN(n10268) );
  AOI21_X1 U11638 ( .B1(n10385), .B2(n12325), .A(n10381), .ZN(n10380) );
  INV_X1 U11639 ( .A(n13158), .ZN(n10381) );
  AND2_X1 U11640 ( .A1(n13629), .A2(n15978), .ZN(n14571) );
  NAND2_X1 U11641 ( .A1(n12680), .A2(n10014), .ZN(n10013) );
  NAND2_X1 U11642 ( .A1(n10012), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10011) );
  NAND2_X1 U11643 ( .A1(n12583), .A2(n9670), .ZN(n10010) );
  NOR2_X1 U11644 ( .A1(n12634), .A2(n10319), .ZN(n12638) );
  NAND2_X1 U11645 ( .A1(n10320), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10319) );
  NOR2_X1 U11646 ( .A1(n10322), .A2(n10321), .ZN(n10320) );
  NAND2_X1 U11647 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10322) );
  NOR2_X1 U11648 ( .A1(n15861), .A2(n10302), .ZN(n10301) );
  NAND2_X1 U11649 ( .A1(n14351), .A2(n21531), .ZN(n10044) );
  AND2_X1 U11650 ( .A1(n10046), .A2(n16202), .ZN(n10045) );
  AND2_X1 U11651 ( .A1(n11012), .A2(n11005), .ZN(n10046) );
  AOI21_X1 U11652 ( .B1(n14350), .B2(n16173), .A(n16189), .ZN(n11012) );
  AND2_X1 U11653 ( .A1(n11005), .A2(n10245), .ZN(n10033) );
  INV_X1 U11654 ( .A(n10033), .ZN(n9815) );
  NOR2_X1 U11655 ( .A1(n14348), .A2(n14349), .ZN(n9817) );
  NAND2_X1 U11656 ( .A1(n11003), .A2(n11002), .ZN(n11017) );
  NOR2_X1 U11657 ( .A1(n11190), .A2(n16186), .ZN(n11002) );
  INV_X1 U11658 ( .A(n15734), .ZN(n10400) );
  INV_X1 U11659 ( .A(n12592), .ZN(n10230) );
  INV_X1 U11660 ( .A(n12795), .ZN(n11106) );
  INV_X1 U11661 ( .A(n16301), .ZN(n10367) );
  INV_X1 U11662 ( .A(n13884), .ZN(n10402) );
  NOR2_X1 U11663 ( .A1(n12603), .A2(n10371), .ZN(n10370) );
  INV_X1 U11664 ( .A(n13618), .ZN(n12388) );
  NOR2_X1 U11665 ( .A1(n13941), .A2(n10229), .ZN(n10228) );
  INV_X1 U11666 ( .A(n14235), .ZN(n10229) );
  INV_X1 U11667 ( .A(n13913), .ZN(n10227) );
  CLKBUF_X1 U11668 ( .A(n10842), .Z(n11188) );
  INV_X1 U11669 ( .A(n16397), .ZN(n9935) );
  NAND2_X1 U11670 ( .A1(n10738), .A2(n10737), .ZN(n10244) );
  AND4_X1 U11671 ( .A1(n10732), .A2(n10731), .A3(n10730), .A4(n10729), .ZN(
        n10738) );
  AND4_X1 U11672 ( .A1(n10736), .A2(n10735), .A3(n10734), .A4(n10733), .ZN(
        n10737) );
  NAND2_X1 U11673 ( .A1(n13928), .A2(n12297), .ZN(n12305) );
  CLKBUF_X1 U11674 ( .A(n12583), .Z(n12584) );
  NAND2_X1 U11675 ( .A1(n11042), .A2(n11041), .ZN(n12495) );
  OR2_X1 U11676 ( .A1(n11040), .A2(n11039), .ZN(n11042) );
  AND4_X1 U11677 ( .A1(n10589), .A2(n12286), .A3(n10594), .A4(n10593), .ZN(
        n9794) );
  AND2_X1 U11678 ( .A1(n11051), .A2(n11035), .ZN(n12492) );
  INV_X1 U11679 ( .A(n18992), .ZN(n13186) );
  NAND2_X1 U11680 ( .A1(n17221), .A2(n12999), .ZN(n10444) );
  NAND2_X1 U11681 ( .A1(n13000), .A2(n17220), .ZN(n18085) );
  NAND2_X1 U11682 ( .A1(n12998), .A2(n13451), .ZN(n13095) );
  AND2_X1 U11683 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12984) );
  NAND2_X1 U11684 ( .A1(n18377), .A2(n18583), .ZN(n10354) );
  NAND2_X1 U11685 ( .A1(n9991), .A2(n18583), .ZN(n10362) );
  NAND2_X1 U11686 ( .A1(n10105), .A2(n9992), .ZN(n9991) );
  AND2_X1 U11687 ( .A1(n10104), .A2(n18773), .ZN(n9992) );
  OR2_X1 U11688 ( .A1(n9999), .A2(n18601), .ZN(n9996) );
  INV_X1 U11689 ( .A(n16930), .ZN(n9999) );
  AOI21_X1 U11690 ( .B1(n16930), .B2(n9998), .A(n10350), .ZN(n9997) );
  NOR2_X1 U11691 ( .A1(n10114), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10113) );
  INV_X1 U11692 ( .A(n18568), .ZN(n10351) );
  NAND2_X1 U11693 ( .A1(n9788), .A2(n10137), .ZN(n9787) );
  INV_X1 U11694 ( .A(n16980), .ZN(n10137) );
  XNOR2_X1 U11695 ( .A(n13404), .B(n10352), .ZN(n16904) );
  AND2_X1 U11696 ( .A1(n13395), .A2(n13378), .ZN(n13421) );
  AND3_X1 U11697 ( .A1(n13023), .A2(n13022), .A3(n13021), .ZN(n13026) );
  AND2_X1 U11698 ( .A1(n12986), .A2(n13452), .ZN(n13061) );
  INV_X1 U11699 ( .A(n13229), .ZN(n17312) );
  INV_X1 U11700 ( .A(n13369), .ZN(n9827) );
  OR3_X1 U11701 ( .A1(n14213), .A2(n14227), .A3(n11979), .ZN(n12964) );
  OR2_X1 U11702 ( .A1(n12239), .A2(n12237), .ZN(n13982) );
  AOI21_X1 U11703 ( .B1(n11576), .B2(n11751), .A(n10430), .ZN(n10429) );
  INV_X1 U11704 ( .A(n11592), .ZN(n10430) );
  NAND2_X1 U11705 ( .A1(n21239), .A2(n21191), .ZN(n12902) );
  AND2_X1 U11706 ( .A1(n11609), .A2(n9626), .ZN(n9857) );
  NAND2_X1 U11707 ( .A1(n12165), .A2(n11727), .ZN(n11622) );
  INV_X1 U11708 ( .A(n11785), .ZN(n12903) );
  NOR2_X1 U11709 ( .A1(n11901), .A2(n15189), .ZN(n11909) );
  NAND2_X1 U11710 ( .A1(n11909), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11916) );
  CLKBUF_X1 U11711 ( .A(n11913), .Z(n11912) );
  AOI21_X1 U11712 ( .B1(n14942), .B2(n14914), .A(n14913), .ZN(n14945) );
  NAND2_X1 U11713 ( .A1(n13615), .A2(n13616), .ZN(n13614) );
  INV_X1 U11714 ( .A(n10076), .ZN(n9913) );
  NAND2_X1 U11715 ( .A1(n15395), .A2(n9923), .ZN(n15381) );
  NAND2_X1 U11716 ( .A1(n13650), .A2(n15394), .ZN(n9923) );
  INV_X1 U11717 ( .A(n12695), .ZN(n12697) );
  NAND2_X1 U11718 ( .A1(n12696), .A2(n15185), .ZN(n12700) );
  AND2_X1 U11719 ( .A1(n12695), .A2(n10406), .ZN(n15232) );
  NAND2_X1 U11720 ( .A1(n15324), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10406) );
  NAND2_X1 U11721 ( .A1(n10330), .A2(n14901), .ZN(n10329) );
  NOR2_X1 U11722 ( .A1(n10416), .A2(n21428), .ZN(n9872) );
  INV_X1 U11723 ( .A(n9960), .ZN(n14192) );
  NAND2_X1 U11724 ( .A1(n14191), .A2(n14192), .ZN(n14190) );
  NAND2_X1 U11725 ( .A1(n12250), .A2(n12246), .ZN(n13648) );
  NAND2_X1 U11726 ( .A1(n11460), .A2(n9980), .ZN(n9979) );
  NOR2_X1 U11727 ( .A1(n11460), .A2(n9980), .ZN(n9978) );
  NAND2_X1 U11728 ( .A1(n11481), .A2(n9706), .ZN(n10427) );
  NOR2_X1 U11729 ( .A1(n9706), .A2(n11481), .ZN(n10425) );
  OAI21_X1 U11730 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n21000), .A(
        n20878), .ZN(n20840) );
  AND2_X1 U11731 ( .A1(n15550), .A2(n15547), .ZN(n20834) );
  INV_X1 U11732 ( .A(n21122), .ZN(n20992) );
  NOR2_X1 U11733 ( .A1(n15550), .A2(n15551), .ZN(n21092) );
  INV_X1 U11734 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21157) );
  AND2_X1 U11735 ( .A1(n21054), .A2(n20878), .ZN(n21197) );
  NOR2_X1 U11736 ( .A1(n21127), .A2(n21126), .ZN(n21237) );
  INV_X2 U11737 ( .A(n11993), .ZN(n20715) );
  INV_X1 U11738 ( .A(n20840), .ZN(n21245) );
  NAND2_X1 U11739 ( .A1(n15539), .A2(n10072), .ZN(n20775) );
  NAND2_X1 U11740 ( .A1(n15573), .A2(n15538), .ZN(n15539) );
  NAND2_X1 U11741 ( .A1(n10312), .A2(n10316), .ZN(n10306) );
  AOI21_X1 U11742 ( .B1(n10299), .B2(n10293), .A(n10286), .ZN(n10285) );
  INV_X1 U11743 ( .A(n15745), .ZN(n10286) );
  INV_X1 U11744 ( .A(n10293), .ZN(n10287) );
  NOR2_X1 U11745 ( .A1(n16266), .A2(n10296), .ZN(n10295) );
  INV_X1 U11746 ( .A(n16281), .ZN(n10296) );
  NAND2_X1 U11747 ( .A1(n10298), .A2(n9609), .ZN(n10297) );
  OR2_X1 U11748 ( .A1(n12336), .A2(n12335), .ZN(n13899) );
  AND2_X1 U11749 ( .A1(n13904), .A2(n9630), .ZN(n16023) );
  INV_X1 U11750 ( .A(n12325), .ZN(n10382) );
  NAND2_X1 U11751 ( .A1(n15881), .A2(n10388), .ZN(n10387) );
  CLKBUF_X1 U11752 ( .A(n13156), .Z(n13157) );
  NAND2_X1 U11753 ( .A1(n15630), .A2(n9734), .ZN(n12756) );
  XNOR2_X1 U11754 ( .A(n11161), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12617) );
  AOI21_X1 U11755 ( .B1(n10091), .B2(n9892), .A(n9891), .ZN(n9890) );
  INV_X1 U11756 ( .A(n10091), .ZN(n9893) );
  INV_X1 U11757 ( .A(n16278), .ZN(n9891) );
  NAND2_X1 U11758 ( .A1(n11157), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12634) );
  INV_X1 U11759 ( .A(n12631), .ZN(n11157) );
  NAND2_X1 U11760 ( .A1(n10050), .A2(n9909), .ZN(n16157) );
  AND2_X1 U11761 ( .A1(n10049), .A2(n10340), .ZN(n9909) );
  AND2_X1 U11762 ( .A1(n12475), .A2(n12474), .ZN(n15635) );
  NAND2_X1 U11763 ( .A1(n16637), .A2(n12576), .ZN(n16491) );
  NAND2_X1 U11764 ( .A1(n11200), .A2(n11199), .ZN(n16211) );
  NAND2_X1 U11765 ( .A1(n10056), .A2(n9614), .ZN(n10054) );
  NAND2_X1 U11766 ( .A1(n9606), .A2(n9663), .ZN(n10056) );
  NAND2_X1 U11767 ( .A1(n10928), .A2(n10094), .ZN(n10135) );
  INV_X1 U11768 ( .A(n11200), .ZN(n16227) );
  NAND2_X1 U11769 ( .A1(n10974), .A2(n16251), .ZN(n16242) );
  NAND2_X1 U11770 ( .A1(n9934), .A2(n11196), .ZN(n9933) );
  NAND2_X1 U11771 ( .A1(n16250), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10127) );
  OR2_X1 U11772 ( .A1(n15807), .A2(n10972), .ZN(n16288) );
  NOR2_X1 U11773 ( .A1(n12604), .A2(n10369), .ZN(n10368) );
  INV_X1 U11774 ( .A(n16306), .ZN(n10369) );
  NAND2_X1 U11775 ( .A1(n12602), .A2(n10370), .ZN(n10363) );
  NAND2_X1 U11776 ( .A1(n16320), .A2(n10918), .ZN(n12602) );
  NAND2_X1 U11777 ( .A1(n9927), .A2(n10779), .ZN(n11191) );
  AND2_X1 U11778 ( .A1(n16404), .A2(n11188), .ZN(n10122) );
  NAND2_X1 U11779 ( .A1(n10083), .A2(n11185), .ZN(n10121) );
  INV_X1 U11780 ( .A(n11182), .ZN(n10083) );
  INV_X1 U11781 ( .A(n10122), .ZN(n11185) );
  NAND2_X1 U11782 ( .A1(n16414), .A2(n9901), .ZN(n10128) );
  NAND2_X1 U11783 ( .A1(n9902), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9901) );
  NAND2_X1 U11784 ( .A1(n16397), .A2(n16717), .ZN(n16402) );
  INV_X1 U11785 ( .A(n11184), .ZN(n16404) );
  NOR2_X1 U11786 ( .A1(n12587), .A2(n14119), .ZN(n12547) );
  NAND2_X1 U11787 ( .A1(n13173), .A2(n20304), .ZN(n13757) );
  OR2_X1 U11788 ( .A1(n20017), .A2(n20091), .ZN(n19846) );
  NOR2_X1 U11789 ( .A1(n20463), .A2(n9805), .ZN(n9804) );
  OR2_X1 U11790 ( .A1(n17421), .A2(n16742), .ZN(n16743) );
  NAND2_X1 U11791 ( .A1(n9861), .A2(n19727), .ZN(n16795) );
  NAND2_X1 U11792 ( .A1(n20251), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n9822) );
  NAND2_X1 U11793 ( .A1(n20352), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n9821) );
  NAND2_X1 U11794 ( .A1(n15909), .A2(n10660), .ZN(n9798) );
  AND2_X1 U11795 ( .A1(n20253), .A2(n16773), .ZN(n19803) );
  AND2_X1 U11796 ( .A1(n20253), .A2(n16771), .ZN(n19802) );
  INV_X1 U11797 ( .A(n10795), .ZN(n20303) );
  INV_X2 U11798 ( .A(n9595), .ZN(n15978) );
  NOR2_X1 U11799 ( .A1(n17712), .A2(n10159), .ZN(n10157) );
  NAND2_X1 U11800 ( .A1(n19565), .A2(n18978), .ZN(n16825) );
  NOR3_X1 U11801 ( .A1(n13543), .A2(n13542), .A3(n13541), .ZN(n16833) );
  OR2_X1 U11802 ( .A1(n13219), .A2(n21512), .ZN(n13543) );
  NAND2_X1 U11803 ( .A1(n9996), .A2(n9997), .ZN(n18581) );
  INV_X1 U11804 ( .A(n18985), .ZN(n18298) );
  XNOR2_X1 U11805 ( .A(n9781), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17120) );
  INV_X1 U11806 ( .A(n18863), .ZN(n18712) );
  NOR2_X1 U11807 ( .A1(n18583), .A2(n18760), .ZN(n10104) );
  OAI21_X1 U11808 ( .B1(n18623), .B2(n9879), .A(n9877), .ZN(n18616) );
  AOI21_X1 U11809 ( .B1(n16921), .B2(n18928), .A(n9878), .ZN(n9877) );
  INV_X1 U11810 ( .A(n18617), .ZN(n9878) );
  XNOR2_X1 U11811 ( .A(n16920), .B(n16918), .ZN(n18623) );
  NAND2_X1 U11812 ( .A1(n18623), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18625) );
  AOI21_X1 U11813 ( .B1(n13093), .B2(n10472), .A(n13389), .ZN(n13744) );
  NOR2_X1 U11814 ( .A1(n9826), .A2(n9825), .ZN(n9824) );
  INV_X1 U11815 ( .A(n19554), .ZN(n18978) );
  NOR2_X1 U11816 ( .A1(n12909), .A2(n14650), .ZN(n11992) );
  INV_X1 U11817 ( .A(n20574), .ZN(n20553) );
  NAND2_X1 U11818 ( .A1(n13610), .A2(n13609), .ZN(n15142) );
  OAI21_X1 U11819 ( .B1(n14213), .B2(n13608), .A(n13607), .ZN(n13610) );
  AND2_X1 U11820 ( .A1(n13606), .A2(n13605), .ZN(n13607) );
  OAI21_X1 U11821 ( .B1(n14743), .B2(n14744), .A(n11912), .ZN(n15181) );
  NAND2_X1 U11822 ( .A1(n15339), .A2(n12708), .ZN(n15344) );
  INV_X1 U11823 ( .A(n15344), .ZN(n20641) );
  NAND2_X1 U11824 ( .A1(n14061), .A2(n21163), .ZN(n20712) );
  INV_X1 U11825 ( .A(n15339), .ZN(n20650) );
  NAND2_X1 U11826 ( .A1(n12741), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12786) );
  OAI211_X1 U11827 ( .C1(n9968), .C2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n9965), .B(n9964), .ZN(n12779) );
  INV_X1 U11828 ( .A(n9966), .ZN(n9965) );
  OAI21_X1 U11829 ( .B1(n15365), .B2(n10204), .A(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10203) );
  NOR2_X1 U11830 ( .A1(n10205), .A2(n12723), .ZN(n10204) );
  AOI21_X1 U11831 ( .B1(n15365), .B2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12268), .ZN(n12269) );
  NAND2_X1 U11832 ( .A1(n12204), .A2(n9774), .ZN(n12203) );
  NAND2_X1 U11833 ( .A1(n9854), .A2(n10075), .ZN(n10074) );
  NAND2_X1 U11834 ( .A1(n15178), .A2(n10416), .ZN(n10075) );
  NAND2_X1 U11835 ( .A1(n10225), .A2(n9853), .ZN(n9854) );
  NOR2_X1 U11836 ( .A1(n10206), .A2(n10205), .ZN(n15365) );
  INV_X1 U11837 ( .A(n12740), .ZN(n10206) );
  NAND2_X1 U11838 ( .A1(n10419), .A2(n10418), .ZN(n10417) );
  OAI21_X1 U11839 ( .B1(n15200), .B2(n15385), .A(n10416), .ZN(n10418) );
  NAND2_X1 U11840 ( .A1(n12913), .A2(n15324), .ZN(n10419) );
  NOR2_X1 U11841 ( .A1(n15403), .A2(n12263), .ZN(n15391) );
  NOR2_X1 U11842 ( .A1(n10209), .A2(n20677), .ZN(n10208) );
  OR2_X1 U11843 ( .A1(n10210), .A2(n12253), .ZN(n10209) );
  INV_X1 U11844 ( .A(n20666), .ZN(n20699) );
  NAND2_X1 U11845 ( .A1(n20772), .A2(n11475), .ZN(n21188) );
  AOI21_X1 U11846 ( .B1(n9609), .B2(n10274), .A(n9761), .ZN(n10271) );
  NAND2_X1 U11847 ( .A1(n15617), .A2(n9609), .ZN(n10273) );
  NOR2_X1 U11848 ( .A1(n16038), .A2(n16021), .ZN(n16031) );
  OR2_X1 U11849 ( .A1(n12353), .A2(n12352), .ZN(n14080) );
  OAI21_X1 U11850 ( .B1(n13823), .B2(n9566), .A(n14187), .ZN(n13177) );
  NAND2_X1 U11851 ( .A1(n19696), .A2(n14156), .ZN(n19662) );
  NAND2_X1 U11852 ( .A1(n19579), .A2(n11155), .ZN(n16419) );
  INV_X1 U11853 ( .A(n16419), .ZN(n16354) );
  XNOR2_X1 U11854 ( .A(n9866), .B(n9938), .ZN(n12546) );
  INV_X1 U11855 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U11856 ( .A1(n14346), .A2(n9775), .ZN(n9866) );
  XNOR2_X1 U11857 ( .A(n16451), .B(n21531), .ZN(n14368) );
  INV_X1 U11858 ( .A(n10372), .ZN(n12815) );
  INV_X1 U11859 ( .A(n10103), .ZN(n12812) );
  NAND2_X1 U11860 ( .A1(n12804), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16556) );
  OR2_X1 U11861 ( .A1(n16265), .A2(n19706), .ZN(n12809) );
  AND2_X1 U11862 ( .A1(n10327), .A2(n10326), .ZN(n10325) );
  NAND2_X1 U11863 ( .A1(n16261), .A2(n19712), .ZN(n10326) );
  INV_X1 U11864 ( .A(n12805), .ZN(n10327) );
  AOI21_X1 U11865 ( .B1(n10086), .B2(n9604), .A(n10949), .ZN(n10085) );
  AND2_X1 U11866 ( .A1(n12591), .A2(n9770), .ZN(n9899) );
  INV_X1 U11867 ( .A(n16731), .ZN(n16722) );
  NAND2_X1 U11868 ( .A1(n12552), .A2(n12551), .ZN(n19728) );
  AND2_X1 U11869 ( .A1(n12547), .A2(n15978), .ZN(n19726) );
  INV_X1 U11870 ( .A(n19728), .ZN(n19712) );
  CLKBUF_X1 U11871 ( .A(n16731), .Z(n19724) );
  INV_X1 U11872 ( .A(n19726), .ZN(n19706) );
  INV_X1 U11873 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20248) );
  INV_X1 U11874 ( .A(n19652), .ZN(n16799) );
  OR2_X1 U11875 ( .A1(n13717), .A2(n13716), .ZN(n13719) );
  INV_X1 U11876 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20480) );
  INV_X1 U11877 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20471) );
  NAND2_X1 U11878 ( .A1(n13806), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16765) );
  INV_X1 U11879 ( .A(n13779), .ZN(n9836) );
  INV_X1 U11880 ( .A(n20315), .ZN(n20262) );
  INV_X1 U11881 ( .A(n20321), .ZN(n20264) );
  INV_X1 U11882 ( .A(n20339), .ZN(n20282) );
  INV_X1 U11883 ( .A(n20361), .ZN(n20295) );
  OR2_X1 U11884 ( .A1(n14134), .A2(n14133), .ZN(n17414) );
  NOR2_X1 U11885 ( .A1(n13197), .A2(n13392), .ZN(n17523) );
  INV_X1 U11886 ( .A(n13198), .ZN(n18295) );
  NAND2_X1 U11887 ( .A1(n19561), .A2(n19401), .ZN(n18293) );
  NOR2_X1 U11888 ( .A1(n19402), .A2(n18293), .ZN(n19565) );
  NOR2_X1 U11889 ( .A1(n18403), .A2(n10155), .ZN(n10154) );
  INV_X1 U11890 ( .A(n17926), .ZN(n17866) );
  NOR2_X2 U11891 ( .A1(n19539), .A2(n17929), .ZN(n17914) );
  NAND2_X1 U11892 ( .A1(n17986), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n17977) );
  NAND2_X1 U11893 ( .A1(n17977), .A2(n18148), .ZN(n17982) );
  AND2_X1 U11894 ( .A1(n17993), .A2(P3_EBX_REG_25__SCAN_IN), .ZN(n17986) );
  AND2_X1 U11895 ( .A1(n13180), .A2(n13123), .ZN(n18154) );
  AND2_X1 U11896 ( .A1(n18154), .A2(n19010), .ZN(n18151) );
  NOR2_X1 U11897 ( .A1(n18318), .A2(n18181), .ZN(n18175) );
  NAND2_X1 U11898 ( .A1(n9650), .A2(P3_EAX_REG_15__SCAN_IN), .ZN(n18231) );
  NAND2_X1 U11899 ( .A1(n17120), .A2(n18675), .ZN(n9780) );
  NOR2_X1 U11900 ( .A1(n16990), .A2(n9783), .ZN(n9782) );
  NOR2_X1 U11901 ( .A1(n17001), .A2(n10163), .ZN(n9783) );
  INV_X2 U11902 ( .A(n18432), .ZN(n18530) );
  INV_X1 U11903 ( .A(n18588), .ZN(n18556) );
  AND2_X1 U11904 ( .A1(n18680), .A2(n17153), .ZN(n18588) );
  OAI22_X1 U11905 ( .A1(n16951), .A2(n16950), .B1(n16949), .B2(n16948), .ZN(
        n17126) );
  AND2_X1 U11906 ( .A1(n18722), .A2(n18944), .ZN(n18881) );
  NAND2_X1 U11907 ( .A1(n10197), .A2(n11966), .ZN(n11922) );
  NAND2_X1 U11908 ( .A1(n11976), .A2(n11920), .ZN(n10197) );
  AND2_X1 U11909 ( .A1(n11924), .A2(n11923), .ZN(n11930) );
  AOI21_X1 U11910 ( .B1(n11961), .B2(n11982), .A(n9914), .ZN(n11924) );
  INV_X1 U11911 ( .A(n11925), .ZN(n9914) );
  INV_X1 U11912 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n9887) );
  NAND2_X1 U11913 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n9801) );
  OAI21_X1 U11914 ( .B1(n19977), .B2(n10751), .A(n9905), .ZN(n10755) );
  NOR2_X1 U11915 ( .A1(n10761), .A2(n10760), .ZN(n10762) );
  OAI22_X1 U11916 ( .A1(n20088), .A2(n10650), .B1(n10649), .B2(n10795), .ZN(
        n10651) );
  OAI21_X1 U11917 ( .B1(n20127), .B2(n10658), .A(n9906), .ZN(n10663) );
  OAI21_X1 U11918 ( .B1(n19977), .B2(n10661), .A(n9795), .ZN(n10662) );
  NAND2_X1 U11919 ( .A1(n9861), .A2(n9888), .ZN(n10009) );
  NAND2_X1 U11920 ( .A1(n9861), .A2(n9677), .ZN(n10007) );
  AOI22_X1 U11921 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n9588), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10838) );
  XNOR2_X1 U11922 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10858) );
  AOI21_X1 U11923 ( .B1(n11937), .B2(n11936), .A(n11935), .ZN(n11944) );
  AOI21_X1 U11924 ( .B1(n11957), .B2(n11956), .A(n11955), .ZN(n11967) );
  AND2_X1 U11925 ( .A1(n9727), .A2(n14873), .ZN(n10441) );
  NAND2_X1 U11926 ( .A1(n13611), .A2(n20747), .ZN(n11392) );
  NAND2_X1 U11927 ( .A1(n9972), .A2(n10182), .ZN(n12126) );
  NAND2_X1 U11928 ( .A1(n9955), .A2(n9840), .ZN(n11398) );
  AND3_X1 U11929 ( .A1(n20747), .A2(n11390), .A3(n9843), .ZN(n9840) );
  NOR2_X1 U11930 ( .A1(n9970), .A2(n11439), .ZN(n9969) );
  NOR2_X1 U11931 ( .A1(n11993), .A2(n10072), .ZN(n11493) );
  INV_X1 U11932 ( .A(n11492), .ZN(n11506) );
  CLKBUF_X1 U11933 ( .A(n10601), .Z(n12482) );
  AOI21_X1 U11934 ( .B1(n10019), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A(n9749), .ZN(n14597) );
  AOI21_X1 U11935 ( .B1(n14624), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A(n9754), .ZN(n14603) );
  NAND2_X1 U11936 ( .A1(n10020), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n14554) );
  AOI21_X1 U11937 ( .B1(n14624), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n9755), .ZN(n14565) );
  AOI21_X1 U11938 ( .B1(n10019), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A(n9716), .ZN(n14525) );
  AOI21_X1 U11939 ( .B1(n10019), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A(n9717), .ZN(n14518) );
  AOI21_X1 U11940 ( .B1(n10019), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A(n9759), .ZN(n14468) );
  AOI21_X1 U11941 ( .B1(n10019), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A(n9715), .ZN(n14461) );
  NOR2_X1 U11942 ( .A1(n10382), .A2(n10389), .ZN(n10378) );
  AND2_X1 U11943 ( .A1(n9596), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10014) );
  NAND2_X1 U11944 ( .A1(n10252), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10607) );
  NOR2_X1 U11945 ( .A1(n16180), .A2(n10282), .ZN(n10281) );
  NOR2_X1 U11946 ( .A1(n10993), .A2(n10032), .ZN(n10031) );
  INV_X1 U11947 ( .A(n16218), .ZN(n10032) );
  NAND2_X1 U11948 ( .A1(n12289), .A2(n10585), .ZN(n10591) );
  AND2_X1 U11949 ( .A1(n10595), .A2(n19806), .ZN(n10575) );
  NAND2_X1 U11950 ( .A1(n10606), .A2(n9790), .ZN(n10623) );
  NAND2_X1 U11951 ( .A1(n10605), .A2(n10604), .ZN(n9790) );
  OAI211_X1 U11952 ( .C1(n11152), .C2(n14281), .A(n10614), .B(n10613), .ZN(
        n10615) );
  INV_X1 U11953 ( .A(n9947), .ZN(n9946) );
  OAI21_X1 U11954 ( .B1(n12482), .B2(n12492), .A(n12495), .ZN(n9947) );
  INV_X1 U11955 ( .A(n12492), .ZN(n9948) );
  NAND2_X1 U11956 ( .A1(n10256), .A2(n10551), .ZN(n10255) );
  NAND2_X1 U11957 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10256) );
  AOI21_X1 U11958 ( .B1(n14596), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n10259), .ZN(n10258) );
  NAND2_X1 U11959 ( .A1(n10260), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10259) );
  NAND2_X1 U11960 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10260) );
  NOR2_X1 U11961 ( .A1(n10642), .A2(n15938), .ZN(n10664) );
  NAND2_X1 U11962 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10057) );
  NAND2_X1 U11963 ( .A1(n10560), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10134) );
  NAND2_X1 U11964 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10133) );
  AND2_X1 U11965 ( .A1(n20248), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11036) );
  XNOR2_X1 U11966 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10854) );
  INV_X1 U11967 ( .A(n13082), .ZN(n13181) );
  AND2_X1 U11968 ( .A1(n19391), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12997) );
  AND2_X1 U11969 ( .A1(n13452), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12996) );
  NAND2_X1 U11970 ( .A1(n16959), .A2(n16958), .ZN(n16967) );
  NAND2_X1 U11971 ( .A1(n13404), .A2(n10352), .ZN(n16908) );
  AOI22_X1 U11972 ( .A1(n12887), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11375), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11297) );
  INV_X1 U11973 ( .A(n11544), .ZN(n11545) );
  NAND2_X1 U11974 ( .A1(n11375), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11347) );
  NOR2_X1 U11975 ( .A1(n14758), .A2(n10438), .ZN(n10437) );
  INV_X1 U11976 ( .A(n10439), .ZN(n10438) );
  AND2_X1 U11977 ( .A1(n14770), .A2(n11887), .ZN(n10439) );
  OR2_X1 U11978 ( .A1(n14834), .A2(n14852), .ZN(n12702) );
  AND2_X1 U11979 ( .A1(n14899), .A2(n10441), .ZN(n12704) );
  INV_X1 U11980 ( .A(n12868), .ZN(n12896) );
  NOR2_X1 U11981 ( .A1(n10435), .A2(n10433), .ZN(n10432) );
  NOR2_X1 U11982 ( .A1(n10337), .A2(n14759), .ZN(n10336) );
  INV_X1 U11983 ( .A(n12915), .ZN(n10337) );
  INV_X1 U11984 ( .A(n12156), .ZN(n9962) );
  NAND2_X1 U11985 ( .A1(n10201), .A2(n9953), .ZN(n10200) );
  INV_X1 U11986 ( .A(n12210), .ZN(n10201) );
  NAND2_X1 U11987 ( .A1(n9681), .A2(n11381), .ZN(n10199) );
  INV_X1 U11988 ( .A(n11397), .ZN(n9980) );
  OR2_X1 U11989 ( .A1(n11456), .A2(n11455), .ZN(n12116) );
  INV_X1 U11990 ( .A(n11493), .ZN(n11505) );
  CLKBUF_X1 U11991 ( .A(n12206), .Z(n12207) );
  INV_X1 U11992 ( .A(n9706), .ZN(n9839) );
  AOI22_X1 U11993 ( .A1(n11376), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11375), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11378) );
  NAND2_X1 U11994 ( .A1(n9915), .A2(n11965), .ZN(n11975) );
  AND2_X1 U11995 ( .A1(n11964), .A2(n11963), .ZN(n11965) );
  OAI21_X1 U11996 ( .B1(n9916), .B2(n11954), .A(n11959), .ZN(n9915) );
  NOR2_X1 U11997 ( .A1(n10218), .A2(n10215), .ZN(n11334) );
  NAND2_X1 U11998 ( .A1(n10217), .A2(n10216), .ZN(n10215) );
  NAND2_X1 U11999 ( .A1(n9692), .A2(n11207), .ZN(n10216) );
  NAND2_X1 U12000 ( .A1(n12887), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10063) );
  NAND2_X1 U12001 ( .A1(n11376), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10062) );
  NAND2_X1 U12002 ( .A1(n10573), .A2(n12283), .ZN(n10601) );
  AND2_X1 U12003 ( .A1(n9729), .A2(n10251), .ZN(n10250) );
  INV_X1 U12004 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10251) );
  INV_X1 U12005 ( .A(n10900), .ZN(n10249) );
  INV_X1 U12006 ( .A(n10899), .ZN(n10248) );
  AOI21_X1 U12007 ( .B1(n10019), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A(n9753), .ZN(n14591) );
  AOI21_X1 U12008 ( .B1(n10019), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(n9752), .ZN(n14584) );
  AOI21_X1 U12009 ( .B1(n10019), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A(n9750), .ZN(n14543) );
  AOI21_X1 U12010 ( .B1(n10019), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A(n9751), .ZN(n14536) );
  AOI21_X1 U12011 ( .B1(n14596), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A(n9758), .ZN(n14500) );
  INV_X1 U12012 ( .A(n16009), .ZN(n10269) );
  NOR2_X1 U12013 ( .A1(n19806), .A2(n10585), .ZN(n10188) );
  NAND2_X1 U12014 ( .A1(n10323), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12494) );
  AND2_X1 U12015 ( .A1(n12594), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12649) );
  INV_X1 U12016 ( .A(n12798), .ZN(n11105) );
  INV_X1 U12017 ( .A(n14360), .ZN(n10234) );
  AND2_X1 U12018 ( .A1(n15681), .A2(n11025), .ZN(n16200) );
  AND4_X1 U12019 ( .A1(n12813), .A2(n10977), .A3(n16243), .A4(n12612), .ZN(
        n10981) );
  NOR2_X1 U12020 ( .A1(n16230), .A2(n16231), .ZN(n9606) );
  NOR2_X1 U12021 ( .A1(n12808), .A2(n10102), .ZN(n10101) );
  INV_X1 U12022 ( .A(n12607), .ZN(n10102) );
  INV_X1 U12023 ( .A(n15784), .ZN(n11099) );
  AND2_X1 U12024 ( .A1(n9620), .A2(n13789), .ZN(n10401) );
  NOR2_X1 U12025 ( .A1(n16638), .A2(n16648), .ZN(n10196) );
  INV_X1 U12026 ( .A(n16376), .ZN(n11193) );
  NOR2_X1 U12027 ( .A1(n10697), .A2(n10696), .ZN(n12319) );
  INV_X1 U12028 ( .A(n10850), .ZN(n12300) );
  AOI21_X1 U12029 ( .B1(n11113), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10344), .ZN(
        n10343) );
  NAND2_X1 U12030 ( .A1(n10342), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10341) );
  NAND2_X1 U12031 ( .A1(n11068), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10346) );
  NAND2_X1 U12032 ( .A1(n12537), .A2(n19806), .ZN(n12556) );
  INV_X1 U12033 ( .A(n12549), .ZN(n13812) );
  OR2_X1 U12034 ( .A1(n14549), .A2(n13631), .ZN(n13637) );
  NAND2_X1 U12035 ( .A1(n9944), .A2(n9943), .ZN(n12532) );
  NAND2_X1 U12036 ( .A1(n15584), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9943) );
  NAND2_X1 U12037 ( .A1(n9945), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9944) );
  OAI21_X1 U12038 ( .B1(n12493), .B2(n9948), .A(n9946), .ZN(n9945) );
  OR2_X1 U12039 ( .A1(n14549), .A2(n13630), .ZN(n13762) );
  AND2_X1 U12040 ( .A1(n14571), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13759) );
  NAND2_X1 U12041 ( .A1(n13760), .A2(n13759), .ZN(n13767) );
  CLKBUF_X1 U12042 ( .A(n11045), .Z(n11046) );
  AOI22_X1 U12043 ( .A1(n9581), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10546) );
  INV_X1 U12044 ( .A(n10593), .ZN(n10581) );
  INV_X1 U12045 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20176) );
  INV_X1 U12046 ( .A(n18996), .ZN(n13189) );
  NAND2_X1 U12047 ( .A1(n12997), .A2(n17220), .ZN(n10446) );
  AND2_X1 U12048 ( .A1(n12996), .A2(n17221), .ZN(n13228) );
  AND3_X1 U12049 ( .A1(n17223), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12986) );
  NAND2_X1 U12050 ( .A1(n10166), .A2(n16816), .ZN(n10165) );
  NOR3_X1 U12051 ( .A1(n18372), .A2(n17576), .A3(n10165), .ZN(n16956) );
  INV_X1 U12052 ( .A(n10109), .ZN(n10108) );
  INV_X1 U12053 ( .A(n16943), .ZN(n9995) );
  NAND2_X1 U12054 ( .A1(n10351), .A2(n10113), .ZN(n17096) );
  AND2_X1 U12055 ( .A1(n16971), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16972) );
  AND2_X1 U12056 ( .A1(n19554), .A2(n19010), .ZN(n13375) );
  NAND2_X1 U12057 ( .A1(n13048), .A2(n10173), .ZN(n10172) );
  NAND2_X1 U12058 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10173) );
  INV_X1 U12059 ( .A(n13054), .ZN(n9826) );
  INV_X1 U12060 ( .A(n13451), .ZN(n13427) );
  INV_X1 U12061 ( .A(n13370), .ZN(n13419) );
  NAND2_X1 U12062 ( .A1(n13396), .A2(n13418), .ZN(n13381) );
  AND2_X1 U12063 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12999) );
  AND2_X1 U12064 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13451), .ZN(
        n14328) );
  AND3_X1 U12065 ( .A1(n13037), .A2(n13036), .A3(n13035), .ZN(n13040) );
  OR2_X1 U12066 ( .A1(n11633), .A2(n15343), .ZN(n11650) );
  NAND2_X1 U12067 ( .A1(n14787), .A2(n12915), .ZN(n12914) );
  AND2_X1 U12068 ( .A1(n14854), .A2(n14837), .ZN(n14839) );
  AND2_X1 U12069 ( .A1(n12037), .A2(n12036), .ZN(n14966) );
  AND2_X1 U12070 ( .A1(n12030), .A2(n12029), .ZN(n15058) );
  INV_X1 U12071 ( .A(n20709), .ZN(n20711) );
  AND2_X1 U12072 ( .A1(n13677), .A2(n13676), .ZN(n20600) );
  NAND2_X1 U12073 ( .A1(n20639), .A2(n13675), .ZN(n13677) );
  OR3_X1 U12074 ( .A1(n14213), .A2(n14227), .A3(n13674), .ZN(n13675) );
  INV_X1 U12075 ( .A(n12108), .ZN(n12979) );
  NAND2_X1 U12076 ( .A1(n11324), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11894) );
  INV_X1 U12077 ( .A(n11879), .ZN(n11324) );
  NAND2_X1 U12078 ( .A1(n11886), .A2(n11885), .ZN(n14781) );
  NAND2_X1 U12079 ( .A1(n11323), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11875) );
  INV_X1 U12080 ( .A(n11832), .ZN(n11323) );
  INV_X1 U12081 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14800) );
  INV_X1 U12082 ( .A(n11878), .ZN(n14794) );
  OR2_X1 U12083 ( .A1(n11848), .A2(n12710), .ZN(n11832) );
  CLKBUF_X1 U12084 ( .A(n14791), .Z(n14792) );
  INV_X1 U12085 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12710) );
  NAND2_X1 U12086 ( .A1(n11322), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11848) );
  INV_X1 U12087 ( .A(n11854), .ZN(n11322) );
  OR2_X1 U12088 ( .A1(n14872), .A2(n12702), .ZN(n14836) );
  OR2_X1 U12089 ( .A1(n14872), .A2(n14852), .ZN(n14850) );
  AND2_X1 U12090 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11318) );
  INV_X1 U12091 ( .A(n11713), .ZN(n11319) );
  INV_X1 U12092 ( .A(n14899), .ZN(n14915) );
  AND2_X1 U12093 ( .A1(n11682), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11730) );
  AND2_X1 U12094 ( .A1(n11316), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11682) );
  INV_X1 U12095 ( .A(n11666), .ZN(n11316) );
  NAND2_X1 U12096 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n11315), .ZN(
        n11666) );
  INV_X1 U12097 ( .A(n11650), .ZN(n11315) );
  NOR2_X1 U12098 ( .A1(n11655), .A2(n11654), .ZN(n15056) );
  AOI21_X1 U12099 ( .B1(n12157), .B2(n11727), .A(n11569), .ZN(n15154) );
  NOR2_X1 U12100 ( .A1(n11605), .A2(n11549), .ZN(n11565) );
  NAND2_X1 U12101 ( .A1(n11606), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11605) );
  OR2_X1 U12102 ( .A1(n14213), .A2(n12969), .ZN(n14042) );
  OAI22_X1 U12103 ( .A1(n9967), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n12724), .B2(n12776), .ZN(n9966) );
  NAND2_X1 U12104 ( .A1(n15210), .A2(n15183), .ZN(n12204) );
  NOR2_X1 U12105 ( .A1(n10416), .A2(n12721), .ZN(n9853) );
  AND2_X1 U12106 ( .A1(n12083), .A2(n12082), .ZN(n14746) );
  NAND2_X1 U12107 ( .A1(n14787), .A2(n10336), .ZN(n14761) );
  AND2_X1 U12108 ( .A1(n12072), .A2(n12071), .ZN(n14797) );
  NAND2_X1 U12109 ( .A1(n14839), .A2(n12770), .ZN(n14812) );
  NAND2_X1 U12110 ( .A1(n12069), .A2(n12068), .ZN(n14809) );
  INV_X1 U12111 ( .A(n14811), .ZN(n12068) );
  INV_X1 U12112 ( .A(n14812), .ZN(n12069) );
  OR2_X1 U12113 ( .A1(n15410), .A2(n15412), .ZN(n15403) );
  OR2_X1 U12114 ( .A1(n15450), .A2(n12262), .ZN(n15410) );
  AND2_X1 U12115 ( .A1(n20702), .A2(n12262), .ZN(n10207) );
  AND2_X1 U12116 ( .A1(n12058), .A2(n12057), .ZN(n14855) );
  XNOR2_X1 U12117 ( .A(n15332), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15241) );
  NAND2_X1 U12118 ( .A1(n12194), .A2(n10118), .ZN(n10117) );
  NAND2_X1 U12119 ( .A1(n14887), .A2(n14888), .ZN(n14890) );
  NAND2_X1 U12120 ( .A1(n15482), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15450) );
  AND2_X1 U12121 ( .A1(n12048), .A2(n12047), .ZN(n14923) );
  NAND2_X1 U12122 ( .A1(n10331), .A2(n12045), .ZN(n14933) );
  AND2_X1 U12123 ( .A1(n20679), .A2(n12257), .ZN(n10210) );
  NAND2_X1 U12124 ( .A1(n12186), .A2(n15284), .ZN(n15297) );
  NAND2_X1 U12125 ( .A1(n9873), .A2(n17358), .ZN(n15342) );
  NAND2_X1 U12126 ( .A1(n17361), .A2(n17359), .ZN(n9873) );
  AND2_X1 U12127 ( .A1(n12026), .A2(n12025), .ZN(n14993) );
  CLKBUF_X1 U12128 ( .A(n14992), .Z(n15059) );
  NAND2_X1 U12129 ( .A1(n10333), .A2(n14247), .ZN(n10332) );
  INV_X1 U12130 ( .A(n10334), .ZN(n10333) );
  NAND2_X1 U12131 ( .A1(n9963), .A2(n12164), .ZN(n17361) );
  OR2_X1 U12132 ( .A1(n12109), .A2(n12108), .ZN(n9958) );
  NAND2_X1 U12133 ( .A1(n15565), .A2(n10072), .ZN(n21377) );
  OAI21_X1 U12134 ( .B1(n11979), .B2(n20733), .A(n13300), .ZN(n12222) );
  OR2_X1 U12135 ( .A1(n12221), .A2(n12220), .ZN(n12969) );
  INV_X1 U12136 ( .A(n13975), .ZN(n11462) );
  NOR2_X1 U12137 ( .A1(n11310), .A2(n11309), .ZN(n11311) );
  INV_X1 U12138 ( .A(n21155), .ZN(n20713) );
  NAND2_X1 U12139 ( .A1(n11586), .A2(n10072), .ZN(n10181) );
  INV_X1 U12140 ( .A(n20838), .ZN(n11468) );
  NAND2_X1 U12141 ( .A1(n10140), .A2(n11472), .ZN(n11571) );
  NAND2_X1 U12142 ( .A1(n11577), .A2(n12115), .ZN(n10140) );
  NOR2_X1 U12143 ( .A1(n11399), .A2(n11980), .ZN(n12972) );
  OR2_X1 U12144 ( .A1(n13304), .A2(n13303), .ZN(n14037) );
  AND2_X1 U12145 ( .A1(n11501), .A2(n21235), .ZN(n20874) );
  INV_X1 U12146 ( .A(n20902), .ZN(n20962) );
  OR2_X1 U12147 ( .A1(n15543), .A2(n20713), .ZN(n21122) );
  INV_X1 U12148 ( .A(n21244), .ZN(n20714) );
  AND2_X1 U12149 ( .A1(n15543), .A2(n20713), .ZN(n21091) );
  AND2_X1 U12150 ( .A1(n14059), .A2(n14063), .ZN(n14223) );
  CLKBUF_X1 U12151 ( .A(n12225), .Z(n14058) );
  INV_X1 U12152 ( .A(n21308), .ZN(n21379) );
  NAND2_X1 U12153 ( .A1(n10601), .A2(n10574), .ZN(n12508) );
  INV_X1 U12154 ( .A(n10998), .ZN(n11001) );
  NOR2_X2 U12155 ( .A1(n10990), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n15653) );
  AND2_X1 U12156 ( .A1(n10038), .A2(n10961), .ZN(n15735) );
  NAND2_X1 U12157 ( .A1(n10934), .A2(n9738), .ZN(n10038) );
  NAND2_X1 U12158 ( .A1(n10919), .A2(n10036), .ZN(n10942) );
  AND2_X1 U12159 ( .A1(n9621), .A2(n10938), .ZN(n10036) );
  NAND2_X1 U12160 ( .A1(n10248), .A2(n10249), .ZN(n10909) );
  INV_X1 U12161 ( .A(n10887), .ZN(n10025) );
  NAND2_X1 U12162 ( .A1(n10021), .A2(n10887), .ZN(n10024) );
  AND2_X1 U12163 ( .A1(n11043), .A2(n12495), .ZN(n12951) );
  NAND2_X1 U12164 ( .A1(n15590), .A2(n12684), .ZN(n15816) );
  AND2_X1 U12165 ( .A1(n11119), .A2(n15714), .ZN(n11120) );
  AND2_X1 U12166 ( .A1(n13966), .A2(n13905), .ZN(n10270) );
  INV_X1 U12167 ( .A(n14571), .ZN(n14549) );
  NOR2_X2 U12168 ( .A1(n15600), .A2(n12754), .ZN(n12753) );
  AOI21_X1 U12169 ( .B1(n14630), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(n9766), .ZN(n14632) );
  AOI21_X1 U12170 ( .B1(n14630), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A(n9767), .ZN(n14622) );
  NOR2_X1 U12171 ( .A1(n10264), .A2(n10263), .ZN(n10262) );
  INV_X1 U12172 ( .A(n10267), .ZN(n10263) );
  NAND2_X1 U12173 ( .A1(n15952), .A2(n14612), .ZN(n10266) );
  AND2_X1 U12174 ( .A1(n12462), .A2(n12461), .ZN(n15734) );
  AND2_X1 U12175 ( .A1(n12458), .A2(n12457), .ZN(n15749) );
  CLKBUF_X1 U12176 ( .A(n12800), .Z(n12801) );
  INV_X1 U12177 ( .A(n16772), .ZN(n12527) );
  AND2_X1 U12178 ( .A1(n12420), .A2(n12419), .ZN(n13884) );
  NAND2_X1 U12179 ( .A1(n12389), .A2(n9610), .ZN(n13885) );
  AND2_X1 U12180 ( .A1(n12341), .A2(n12340), .ZN(n13167) );
  INV_X1 U12181 ( .A(n10190), .ZN(n12513) );
  CLKBUF_X1 U12182 ( .A(n12512), .Z(n12559) );
  NOR2_X1 U12183 ( .A1(n10593), .A2(n15584), .ZN(n13629) );
  INV_X1 U12184 ( .A(n12494), .ZN(n14153) );
  NOR2_X1 U12185 ( .A1(n12941), .A2(n20381), .ZN(n13703) );
  INV_X1 U12186 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16206) );
  INV_X1 U12187 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12597) );
  AND2_X1 U12188 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11158) );
  NAND2_X1 U12189 ( .A1(n11106), .A2(n11105), .ZN(n12796) );
  INV_X1 U12190 ( .A(n12634), .ZN(n10318) );
  NOR2_X1 U12191 ( .A1(n12634), .A2(n10322), .ZN(n12637) );
  AND2_X1 U12192 ( .A1(n9693), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10300) );
  NAND2_X1 U12193 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n10280), .ZN(
        n12627) );
  AND4_X1 U12194 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10280) );
  NAND2_X1 U12195 ( .A1(n10082), .A2(n10239), .ZN(n10081) );
  NAND2_X1 U12196 ( .A1(n10239), .A2(n10238), .ZN(n10059) );
  INV_X1 U12197 ( .A(n16160), .ZN(n11028) );
  INV_X1 U12198 ( .A(n12749), .ZN(n11027) );
  NAND2_X1 U12199 ( .A1(n12748), .A2(n10349), .ZN(n10348) );
  INV_X1 U12200 ( .A(n16159), .ZN(n10349) );
  AND2_X1 U12201 ( .A1(n10451), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10340) );
  INV_X1 U12202 ( .A(n10042), .ZN(n10041) );
  OAI21_X1 U12203 ( .B1(n14351), .B2(n9771), .A(n10136), .ZN(n10042) );
  NAND2_X1 U12204 ( .A1(n9818), .A2(n10136), .ZN(n9820) );
  NAND2_X1 U12205 ( .A1(n11006), .A2(n10033), .ZN(n9818) );
  NAND2_X1 U12206 ( .A1(n10397), .A2(n15621), .ZN(n10396) );
  OAI211_X1 U12207 ( .C1(n11006), .C2(n9816), .A(n9814), .B(n9813), .ZN(n16169) );
  INV_X1 U12208 ( .A(n9817), .ZN(n9816) );
  NAND2_X1 U12209 ( .A1(n11006), .A2(n9622), .ZN(n9813) );
  INV_X1 U12210 ( .A(n10397), .ZN(n10395) );
  NOR2_X1 U12211 ( .A1(n16479), .A2(n16492), .ZN(n10051) );
  INV_X1 U12212 ( .A(n11006), .ZN(n16177) );
  AND2_X1 U12213 ( .A1(n9730), .A2(n12821), .ZN(n10398) );
  INV_X1 U12214 ( .A(n15678), .ZN(n15694) );
  OR2_X1 U12215 ( .A1(n10987), .A2(n16508), .ZN(n16219) );
  NAND2_X1 U12216 ( .A1(n10966), .A2(n10965), .ZN(n12814) );
  OR2_X1 U12217 ( .A1(n15709), .A2(n11190), .ZN(n10966) );
  INV_X1 U12218 ( .A(n10100), .ZN(n12806) );
  NAND2_X1 U12219 ( .A1(n9606), .A2(n12609), .ZN(n10374) );
  AND2_X1 U12220 ( .A1(n12464), .A2(n12463), .ZN(n15721) );
  AND2_X1 U12221 ( .A1(n12460), .A2(n9730), .ZN(n15720) );
  NAND2_X1 U12222 ( .A1(n12460), .A2(n9712), .ZN(n15732) );
  NAND2_X1 U12223 ( .A1(n12612), .A2(n12610), .ZN(n10099) );
  AND2_X1 U12224 ( .A1(n12451), .A2(n12450), .ZN(n14068) );
  AND2_X1 U12225 ( .A1(n10366), .A2(n16289), .ZN(n10365) );
  NAND2_X1 U12226 ( .A1(n10096), .A2(n10094), .ZN(n10093) );
  OR2_X1 U12227 ( .A1(n10368), .A2(n10367), .ZN(n10366) );
  INV_X1 U12228 ( .A(n10096), .ZN(n10095) );
  INV_X1 U12229 ( .A(n16286), .ZN(n16275) );
  CLKBUF_X1 U12230 ( .A(n13787), .Z(n13788) );
  AND2_X1 U12231 ( .A1(n12389), .A2(n9620), .ZN(n13887) );
  NAND2_X1 U12232 ( .A1(n13895), .A2(n11087), .ZN(n15812) );
  AND2_X1 U12233 ( .A1(n12387), .A2(n12386), .ZN(n13618) );
  INV_X1 U12234 ( .A(n10196), .ZN(n9985) );
  AND2_X1 U12235 ( .A1(n16683), .A2(n16673), .ZN(n16637) );
  INV_X1 U12236 ( .A(n14082), .ZN(n10226) );
  INV_X1 U12237 ( .A(n9830), .ZN(n16353) );
  INV_X1 U12238 ( .A(n16637), .ZN(n16662) );
  NAND2_X1 U12239 ( .A1(n9862), .A2(n9638), .ZN(n9900) );
  NOR2_X1 U12240 ( .A1(n14669), .A2(n12575), .ZN(n16683) );
  NOR2_X1 U12241 ( .A1(n9671), .A2(n10244), .ZN(n10243) );
  INV_X1 U12242 ( .A(n9924), .ZN(n10040) );
  NAND2_X1 U12243 ( .A1(n14656), .A2(n14655), .ZN(n14657) );
  XNOR2_X1 U12244 ( .A(n11168), .B(n11166), .ZN(n14656) );
  NAND2_X1 U12245 ( .A1(n12536), .A2(n12507), .ZN(n13808) );
  INV_X1 U12246 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19722) );
  NAND2_X1 U12247 ( .A1(n10006), .A2(n10588), .ZN(n10324) );
  NOR2_X1 U12248 ( .A1(n12587), .A2(n12566), .ZN(n12791) );
  AND2_X1 U12249 ( .A1(n12277), .A2(n12276), .ZN(n12278) );
  AOI21_X1 U12250 ( .B1(n16732), .B2(n13755), .A(n13636), .ZN(n13716) );
  CLKBUF_X1 U12251 ( .A(n13921), .Z(n14665) );
  INV_X1 U12252 ( .A(n12509), .ZN(n9809) );
  NOR2_X2 U12253 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14104) );
  CLKBUF_X1 U12254 ( .A(n13809), .Z(n14103) );
  NAND2_X1 U12255 ( .A1(n13640), .A2(n13641), .ZN(n13642) );
  AND2_X1 U12256 ( .A1(n10584), .A2(n10598), .ZN(n10170) );
  AND2_X1 U12257 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19873) );
  NAND2_X1 U12258 ( .A1(n20253), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19795) );
  AND2_X1 U12259 ( .A1(n19554), .A2(n18985), .ZN(n13380) );
  INV_X1 U12260 ( .A(n13744), .ZN(n19405) );
  NOR2_X1 U12261 ( .A1(n16809), .A2(n16808), .ZN(n19402) );
  NOR2_X1 U12262 ( .A1(n18403), .A2(n10159), .ZN(n10153) );
  NOR2_X1 U12263 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17845), .ZN(n17823) );
  NOR2_X1 U12264 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17879), .ZN(n17878) );
  NOR2_X1 U12265 ( .A1(n19389), .A2(n16825), .ZN(n17902) );
  INV_X1 U12266 ( .A(n17902), .ZN(n17917) );
  NAND2_X1 U12267 ( .A1(n18052), .A2(P3_EBX_REG_21__SCAN_IN), .ZN(n17231) );
  NAND2_X1 U12268 ( .A1(n18001), .A2(P3_EBX_REG_22__SCAN_IN), .ZN(n17994) );
  AND4_X1 U12269 ( .A1(n13004), .A2(n13003), .A3(n13002), .A4(n13001), .ZN(
        n13005) );
  OR2_X1 U12270 ( .A1(n13520), .A2(n13519), .ZN(n16899) );
  OR2_X1 U12271 ( .A1(n13352), .A2(n13351), .ZN(n16960) );
  NAND2_X1 U12272 ( .A1(n10171), .A2(n19561), .ZN(n13219) );
  NAND2_X1 U12273 ( .A1(n13438), .A2(n13203), .ZN(n10171) );
  NOR2_X1 U12274 ( .A1(n18293), .A2(n18256), .ZN(n18273) );
  NAND2_X1 U12275 ( .A1(n17162), .A2(n9884), .ZN(n9883) );
  NAND2_X1 U12276 ( .A1(n17049), .A2(n10114), .ZN(n9884) );
  NOR2_X1 U12277 ( .A1(n18373), .A2(n10167), .ZN(n10166) );
  AND2_X1 U12278 ( .A1(n18471), .A2(n9703), .ZN(n17067) );
  INV_X1 U12279 ( .A(n18406), .ZN(n10145) );
  NAND2_X1 U12280 ( .A1(n18471), .A2(n9616), .ZN(n18405) );
  NOR2_X1 U12281 ( .A1(n17064), .A2(n10147), .ZN(n10146) );
  INV_X1 U12282 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10147) );
  NOR2_X1 U12283 ( .A1(n17078), .A2(n17079), .ZN(n18471) );
  NAND2_X1 U12284 ( .A1(n17745), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17078) );
  NAND2_X1 U12285 ( .A1(n10144), .A2(n10143), .ZN(n18518) );
  NOR2_X1 U12286 ( .A1(n16815), .A2(n18589), .ZN(n10143) );
  NOR2_X1 U12287 ( .A1(n18630), .A2(n18629), .ZN(n18615) );
  AND2_X1 U12288 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18642) );
  NOR2_X1 U12289 ( .A1(n16970), .A2(n10139), .ZN(n16968) );
  AND2_X1 U12290 ( .A1(n13405), .A2(n13410), .ZN(n10139) );
  XNOR2_X1 U12291 ( .A(n13404), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18678) );
  AND2_X1 U12292 ( .A1(n16952), .A2(n17142), .ZN(n10110) );
  NAND2_X1 U12293 ( .A1(n9993), .A2(n9994), .ZN(n17160) );
  AND2_X1 U12294 ( .A1(n17191), .A2(n10114), .ZN(n9993) );
  INV_X1 U12295 ( .A(n10354), .ZN(n10357) );
  INV_X1 U12296 ( .A(n10356), .ZN(n10355) );
  INV_X1 U12297 ( .A(n10106), .ZN(n10361) );
  AND2_X1 U12298 ( .A1(n18418), .A2(n18716), .ZN(n18401) );
  INV_X1 U12299 ( .A(n10362), .ZN(n9881) );
  INV_X1 U12300 ( .A(n18808), .ZN(n18709) );
  INV_X1 U12301 ( .A(n18578), .ZN(n10111) );
  INV_X1 U12302 ( .A(n10113), .ZN(n10112) );
  INV_X1 U12303 ( .A(n18498), .ZN(n18866) );
  NAND2_X1 U12304 ( .A1(n10351), .A2(n10350), .ZN(n18582) );
  NAND2_X1 U12305 ( .A1(n18601), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18603) );
  AND2_X1 U12306 ( .A1(n16963), .A2(n16961), .ZN(n18609) );
  NOR2_X1 U12307 ( .A1(n18626), .A2(n16977), .ZN(n18608) );
  NOR2_X1 U12308 ( .A1(n18628), .A2(n18627), .ZN(n18626) );
  AOI21_X1 U12309 ( .B1(n16968), .B2(n10138), .A(n16970), .ZN(n18655) );
  INV_X1 U12310 ( .A(n16969), .ZN(n10138) );
  OR2_X1 U12311 ( .A1(n16972), .A2(n9785), .ZN(n18656) );
  NOR2_X1 U12312 ( .A1(n16971), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9785) );
  NOR2_X1 U12313 ( .A1(n18655), .A2(n18656), .ZN(n18654) );
  NAND2_X1 U12314 ( .A1(n16907), .A2(n16906), .ZN(n18652) );
  AOI21_X2 U12315 ( .B1(n13375), .B2(n13199), .A(n16808), .ZN(n13384) );
  AND3_X1 U12316 ( .A1(n13419), .A2(n13196), .A3(n18298), .ZN(n13199) );
  INV_X1 U12317 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19407) );
  INV_X1 U12318 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17223) );
  NOR2_X2 U12319 ( .A1(n19557), .A2(n13381), .ZN(n19406) );
  NOR2_X1 U12320 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18977), .ZN(n19263) );
  INV_X1 U12321 ( .A(n13392), .ZN(n18989) );
  OR2_X1 U12322 ( .A1(n13033), .A2(n13032), .ZN(n18992) );
  INV_X1 U12323 ( .A(n19263), .ZN(n19011) );
  OR2_X1 U12324 ( .A1(n19399), .A2(n13745), .ZN(n13746) );
  INV_X1 U12325 ( .A(n12964), .ZN(n12980) );
  AND2_X1 U12326 ( .A1(n20540), .A2(n14841), .ZN(n20505) );
  INV_X1 U12327 ( .A(n17350), .ZN(n20536) );
  NOR2_X1 U12328 ( .A1(n14950), .A2(n14840), .ZN(n20540) );
  INV_X1 U12329 ( .A(n20553), .ZN(n20541) );
  NAND2_X1 U12330 ( .A1(n10428), .A2(n10429), .ZN(n13833) );
  NAND2_X1 U12331 ( .A1(n21382), .A2(n11991), .ZN(n20562) );
  INV_X1 U12332 ( .A(n20579), .ZN(n20565) );
  NOR2_X1 U12333 ( .A1(n12095), .A2(n12094), .ZN(n20574) );
  NAND2_X1 U12334 ( .A1(n14950), .A2(n20562), .ZN(n20517) );
  NOR2_X2 U12335 ( .A1(n12095), .A2(n12090), .ZN(n20532) );
  INV_X1 U12336 ( .A(n20599), .ZN(n15062) );
  INV_X1 U12337 ( .A(n20594), .ZN(n20590) );
  AND2_X1 U12338 ( .A1(n13246), .A2(n13609), .ZN(n20599) );
  OR2_X1 U12339 ( .A1(n13604), .A2(n13625), .ZN(n13244) );
  NAND2_X1 U12340 ( .A1(n15157), .A2(n9842), .ZN(n15127) );
  INV_X1 U12341 ( .A(n15135), .ZN(n15129) );
  OR2_X1 U12342 ( .A1(n14715), .A2(n20711), .ZN(n15135) );
  AND2_X1 U12343 ( .A1(n15157), .A2(n13613), .ZN(n15143) );
  INV_X2 U12344 ( .A(n15142), .ZN(n15157) );
  INV_X1 U12345 ( .A(n15143), .ZN(n15156) );
  NOR2_X1 U12346 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14220), .ZN(n20612) );
  INV_X1 U12347 ( .A(n21378), .ZN(n20624) );
  OAI21_X1 U12348 ( .B1(n12979), .B2(n21308), .A(n12980), .ZN(n13268) );
  INV_X1 U12349 ( .A(n20639), .ZN(n13601) );
  INV_X1 U12350 ( .A(n13550), .ZN(n20637) );
  INV_X1 U12351 ( .A(n13268), .ZN(n13550) );
  NOR2_X1 U12352 ( .A1(n20712), .A2(n15112), .ZN(n12714) );
  INV_X1 U12353 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15251) );
  OAI21_X1 U12354 ( .B1(n14945), .B2(n14928), .A(n14927), .ZN(n15290) );
  INV_X1 U12355 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15343) );
  INV_X1 U12356 ( .A(n20654), .ZN(n15347) );
  NAND2_X1 U12357 ( .A1(n12777), .A2(n9912), .ZN(n12725) );
  NAND2_X1 U12358 ( .A1(n9913), .A2(n12724), .ZN(n9912) );
  NOR2_X1 U12359 ( .A1(n15406), .A2(n9675), .ZN(n15395) );
  OAI21_X1 U12360 ( .B1(n15430), .B2(n12198), .A(n10416), .ZN(n15219) );
  AOI21_X1 U12361 ( .B1(n9921), .B2(n9922), .A(n15517), .ZN(n15406) );
  NOR2_X1 U12362 ( .A1(n10207), .A2(n15412), .ZN(n9922) );
  NAND3_X1 U12363 ( .A1(n9613), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n10414), .ZN(n10408) );
  NOR2_X1 U12364 ( .A1(n15481), .A2(n10207), .ZN(n15424) );
  NAND2_X1 U12365 ( .A1(n9871), .A2(n9870), .ZN(n9869) );
  NAND2_X1 U12366 ( .A1(n15325), .A2(n10416), .ZN(n9870) );
  NAND2_X1 U12367 ( .A1(n15323), .A2(n9872), .ZN(n9871) );
  NAND2_X1 U12368 ( .A1(n14190), .A2(n12156), .ZN(n17368) );
  AND2_X1 U12369 ( .A1(n20679), .A2(n20701), .ZN(n20675) );
  NAND2_X1 U12370 ( .A1(n12252), .A2(n12251), .ZN(n20677) );
  OR2_X1 U12371 ( .A1(n20679), .A2(n13650), .ZN(n20702) );
  NAND2_X1 U12372 ( .A1(n12250), .A2(n14649), .ZN(n13652) );
  NAND2_X1 U12373 ( .A1(n9690), .A2(n10426), .ZN(n21127) );
  INV_X1 U12374 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20708) );
  NOR2_X1 U12375 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15565) );
  INV_X1 U12376 ( .A(n20833), .ZN(n20799) );
  OAI211_X1 U12377 ( .C1(n21163), .C2(n20777), .A(n20776), .B(n21245), .ZN(
        n20794) );
  OAI22_X1 U12378 ( .A1(n20845), .A2(n20844), .B1(n21239), .B2(n20843), .ZN(
        n20867) );
  AND2_X1 U12379 ( .A1(n20834), .A2(n21091), .ZN(n20896) );
  NAND2_X1 U12380 ( .A1(n20962), .A2(n10452), .ZN(n20956) );
  OAI211_X1 U12381 ( .C1(n20930), .C2(n21000), .A(n21197), .B(n20929), .ZN(
        n20959) );
  OAI211_X1 U12382 ( .C1(n21015), .C2(n21000), .A(n21050), .B(n20999), .ZN(
        n21018) );
  OAI211_X1 U12383 ( .C1(n21163), .C2(n21024), .A(n21023), .B(n21245), .ZN(
        n21042) );
  INV_X1 U12384 ( .A(n20764), .ZN(n9954) );
  OAI22_X1 U12385 ( .A1(n21056), .A2(n21055), .B1(n21054), .B2(n21053), .ZN(
        n21087) );
  OAI211_X1 U12386 ( .C1(n21163), .C2(n21099), .A(n21098), .B(n21245), .ZN(
        n21119) );
  INV_X1 U12387 ( .A(n21115), .ZN(n21118) );
  OAI211_X1 U12388 ( .C1(n21130), .C2(n21239), .A(n21197), .B(n21129), .ZN(
        n21151) );
  OAI211_X1 U12389 ( .C1(n21163), .C2(n21162), .A(n21161), .B(n21245), .ZN(
        n21181) );
  INV_X1 U12390 ( .A(n21059), .ZN(n21252) );
  INV_X1 U12391 ( .A(n21079), .ZN(n21282) );
  OAI211_X1 U12392 ( .C1(n21247), .C2(n21163), .A(n21246), .B(n21245), .ZN(
        n21294) );
  INV_X1 U12393 ( .A(n13609), .ZN(n14227) );
  OR2_X1 U12394 ( .A1(n14213), .A2(n21000), .ZN(n15573) );
  INV_X1 U12395 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n14650) );
  OR2_X1 U12396 ( .A1(n12950), .A2(n17428), .ZN(n15590) );
  OAI21_X1 U12397 ( .B1(n16057), .B2(n19611), .A(n10392), .ZN(n10391) );
  AOI21_X1 U12398 ( .B1(n15612), .B2(n19609), .A(n15611), .ZN(n10393) );
  NOR2_X1 U12399 ( .A1(n10279), .A2(n10277), .ZN(n10276) );
  NAND2_X1 U12400 ( .A1(n15647), .A2(n9609), .ZN(n10278) );
  AOI21_X1 U12401 ( .B1(n9611), .B2(n10306), .A(n9765), .ZN(n10305) );
  NAND2_X1 U12402 ( .A1(n10309), .A2(n10308), .ZN(n10307) );
  NAND2_X1 U12403 ( .A1(n15715), .A2(n9609), .ZN(n10311) );
  INV_X1 U12404 ( .A(n10284), .ZN(n10283) );
  NAND2_X1 U12405 ( .A1(n10297), .A2(n9737), .ZN(n10292) );
  NAND2_X1 U12406 ( .A1(n10290), .A2(n10288), .ZN(n15759) );
  INV_X1 U12407 ( .A(n10289), .ZN(n10288) );
  OR2_X1 U12408 ( .A1(n10297), .A2(n10291), .ZN(n10290) );
  OAI21_X1 U12409 ( .B1(n10291), .B2(n10295), .A(n16259), .ZN(n10289) );
  AOI21_X1 U12410 ( .B1(n15774), .B2(n9609), .A(n16266), .ZN(n15758) );
  AND2_X1 U12411 ( .A1(n12677), .A2(n12676), .ZN(n15791) );
  NAND2_X1 U12412 ( .A1(n12617), .A2(n15584), .ZN(n12619) );
  INV_X1 U12413 ( .A(n15933), .ZN(n19611) );
  NAND2_X1 U12414 ( .A1(n14277), .A2(n15791), .ZN(n15912) );
  INV_X1 U12415 ( .A(n19625), .ZN(n15930) );
  NAND2_X1 U12416 ( .A1(n9609), .A2(n15791), .ZN(n15944) );
  INV_X1 U12417 ( .A(n15912), .ZN(n15931) );
  OR2_X1 U12418 ( .A1(n12444), .A2(n12443), .ZN(n16027) );
  OR2_X1 U12419 ( .A1(n12430), .A2(n12429), .ZN(n16033) );
  OR2_X1 U12420 ( .A1(n12414), .A2(n12413), .ZN(n16039) );
  OR2_X1 U12421 ( .A1(n12399), .A2(n12398), .ZN(n14391) );
  NAND2_X1 U12422 ( .A1(n13904), .A2(n10270), .ZN(n14393) );
  INV_X1 U12423 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14281) );
  NAND2_X1 U12424 ( .A1(n15960), .A2(n15959), .ZN(n15958) );
  AND2_X1 U12425 ( .A1(n16151), .A2(n13148), .ZN(n16137) );
  INV_X1 U12426 ( .A(n10379), .ZN(n13159) );
  AOI21_X1 U12427 ( .B1(n10387), .B2(n10384), .A(n10382), .ZN(n10379) );
  OR2_X1 U12428 ( .A1(n15881), .A2(n16146), .ZN(n10383) );
  AND2_X1 U12429 ( .A1(n16056), .A2(n16144), .ZN(n16156) );
  AND2_X1 U12430 ( .A1(n16151), .A2(n10596), .ZN(n19648) );
  INV_X1 U12431 ( .A(n16144), .ZN(n19649) );
  NOR2_X1 U12432 ( .A1(n14151), .A2(n14150), .ZN(n14152) );
  INV_X2 U12433 ( .A(n19662), .ZN(n19693) );
  INV_X1 U12434 ( .A(n13805), .ZN(n19700) );
  CLKBUF_X2 U12435 ( .A(n13795), .Z(n19701) );
  INV_X1 U12436 ( .A(n13704), .ZN(n19698) );
  NAND2_X1 U12437 ( .A1(n9567), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16262) );
  NAND2_X1 U12438 ( .A1(n16275), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10015) );
  INV_X1 U12439 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15861) );
  INV_X1 U12440 ( .A(n16429), .ZN(n16409) );
  INV_X1 U12441 ( .A(n16732), .ZN(n13720) );
  INV_X1 U12442 ( .A(n16425), .ZN(n16406) );
  NAND2_X1 U12443 ( .A1(n14357), .A2(n9940), .ZN(n16435) );
  NAND2_X1 U12444 ( .A1(n9942), .A2(n9941), .ZN(n9940) );
  INV_X1 U12445 ( .A(n9942), .ZN(n16446) );
  INV_X1 U12446 ( .A(n16458), .ZN(n16469) );
  NAND2_X1 U12447 ( .A1(n9907), .A2(n16198), .ZN(n16490) );
  NAND2_X1 U12448 ( .A1(n16211), .A2(n16479), .ZN(n9907) );
  INV_X1 U12449 ( .A(n16515), .ZN(n16226) );
  INV_X1 U12450 ( .A(n10376), .ZN(n10375) );
  NAND2_X1 U12451 ( .A1(n10364), .A2(n16301), .ZN(n16291) );
  NAND2_X1 U12452 ( .A1(n10363), .A2(n10368), .ZN(n10364) );
  NAND2_X1 U12453 ( .A1(n10363), .A2(n16306), .ZN(n9807) );
  CLKBUF_X1 U12454 ( .A(n16367), .Z(n16669) );
  NAND2_X1 U12455 ( .A1(n9900), .A2(n9925), .ZN(n16670) );
  OAI211_X1 U12456 ( .C1(n11183), .C2(n10122), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n10121), .ZN(n10129) );
  NOR2_X1 U12457 ( .A1(n12587), .A2(n13808), .ZN(n19719) );
  INV_X1 U12458 ( .A(n14155), .ZN(n16742) );
  INV_X1 U12459 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14307) );
  INV_X1 U12460 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17343) );
  NAND2_X1 U12461 ( .A1(n13828), .A2(n13827), .ZN(n17344) );
  NAND2_X1 U12462 ( .A1(n9903), .A2(n9768), .ZN(n19850) );
  OAI21_X1 U12463 ( .B1(n19848), .B2(n20120), .A(n19845), .ZN(n19868) );
  OAI211_X1 U12464 ( .C1(n16781), .C2(n16780), .A(n20253), .B(n16779), .ZN(
        n19972) );
  NOR2_X1 U12465 ( .A1(n20463), .A2(n10120), .ZN(n10119) );
  NAND2_X1 U12466 ( .A1(n9806), .A2(n9804), .ZN(n20011) );
  INV_X1 U12467 ( .A(n19988), .ZN(n20036) );
  INV_X1 U12468 ( .A(n20030), .ZN(n20037) );
  INV_X1 U12469 ( .A(n20095), .ZN(n20114) );
  INV_X1 U12470 ( .A(n20088), .ZN(n10648) );
  AND2_X1 U12471 ( .A1(n16802), .A2(n16801), .ZN(n20171) );
  NAND2_X1 U12472 ( .A1(n16777), .A2(n16776), .ZN(n20189) );
  NAND2_X1 U12473 ( .A1(n19774), .A2(n19773), .ZN(n20199) );
  NAND2_X1 U12474 ( .A1(n19783), .A2(n19782), .ZN(n20202) );
  NAND2_X1 U12475 ( .A1(n19791), .A2(n19790), .ZN(n20205) );
  INV_X1 U12476 ( .A(n20184), .ZN(n20213) );
  NAND2_X1 U12477 ( .A1(n16786), .A2(n16785), .ZN(n20226) );
  NAND2_X1 U12478 ( .A1(n19768), .A2(n19767), .ZN(n20231) );
  NAND2_X1 U12479 ( .A1(n19805), .A2(n19804), .ZN(n20241) );
  INV_X1 U12480 ( .A(n20337), .ZN(n20278) );
  INV_X1 U12481 ( .A(n20345), .ZN(n20284) );
  INV_X1 U12482 ( .A(n20343), .ZN(n20283) );
  INV_X1 U12483 ( .A(n20349), .ZN(n20288) );
  OR2_X1 U12484 ( .A1(n20257), .A2(n20294), .ZN(n9800) );
  OR2_X1 U12485 ( .A1(n20259), .A2(n20255), .ZN(n9833) );
  NAND2_X1 U12486 ( .A1(n16775), .A2(n16774), .ZN(n20315) );
  INV_X1 U12487 ( .A(n20249), .ZN(n20306) );
  INV_X1 U12488 ( .A(n19747), .ZN(n20307) );
  INV_X1 U12489 ( .A(n20226), .ZN(n20324) );
  NAND2_X1 U12490 ( .A1(n16788), .A2(n16787), .ZN(n20321) );
  NOR2_X1 U12491 ( .A1(n19795), .A2(n9596), .ZN(n20319) );
  INV_X1 U12492 ( .A(n16803), .ZN(n20320) );
  INV_X1 U12493 ( .A(n20268), .ZN(n20325) );
  AND2_X1 U12494 ( .A1(n20253), .A2(n19762), .ZN(n20326) );
  INV_X1 U12495 ( .A(n20194), .ZN(n20330) );
  INV_X1 U12496 ( .A(n20231), .ZN(n20336) );
  NAND2_X1 U12497 ( .A1(n19766), .A2(n19765), .ZN(n20333) );
  INV_X1 U12498 ( .A(n20273), .ZN(n20331) );
  AND2_X1 U12499 ( .A1(n20253), .A2(n19770), .ZN(n20332) );
  NAND2_X1 U12500 ( .A1(n19776), .A2(n19775), .ZN(n20339) );
  NOR2_X1 U12501 ( .A1(n19795), .A2(n19777), .ZN(n20337) );
  AND2_X1 U12502 ( .A1(n20253), .A2(n19779), .ZN(n20338) );
  INV_X1 U12503 ( .A(n20199), .ZN(n20342) );
  NOR2_X1 U12504 ( .A1(n19795), .A2(n10597), .ZN(n20343) );
  AND2_X1 U12505 ( .A1(n20253), .A2(n19787), .ZN(n20344) );
  NOR2_X1 U12506 ( .A1(n19795), .A2(n10581), .ZN(n20349) );
  NAND2_X1 U12507 ( .A1(n19793), .A2(n19792), .ZN(n20351) );
  AND2_X1 U12508 ( .A1(n20253), .A2(n19797), .ZN(n20350) );
  INV_X1 U12509 ( .A(n20205), .ZN(n20356) );
  INV_X1 U12510 ( .A(n20241), .ZN(n20367) );
  INV_X1 U12511 ( .A(n20246), .ZN(n9835) );
  NAND2_X1 U12512 ( .A1(n19801), .A2(n19800), .ZN(n20361) );
  NOR2_X1 U12513 ( .A1(n20308), .A2(n20305), .ZN(n20360) );
  AND2_X1 U12514 ( .A1(n20253), .A2(n19810), .ZN(n20359) );
  NAND3_X1 U12515 ( .A1(n16757), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n17428) );
  AND2_X1 U12516 ( .A1(n14139), .A2(n14138), .ZN(n17425) );
  INV_X1 U12517 ( .A(n19571), .ZN(n19557) );
  NAND2_X1 U12518 ( .A1(n17000), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16999) );
  NAND2_X1 U12519 ( .A1(n17580), .A2(n17744), .ZN(n17568) );
  NOR2_X1 U12520 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17611), .ZN(n17610) );
  NAND2_X1 U12521 ( .A1(n17681), .A2(n17744), .ZN(n17665) );
  NAND2_X1 U12522 ( .A1(n10150), .A2(n10149), .ZN(n17726) );
  NOR2_X1 U12523 ( .A1(n17712), .A2(n10155), .ZN(n10158) );
  NOR2_X1 U12524 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17791), .ZN(n17772) );
  OR2_X1 U12525 ( .A1(n16825), .A2(n16824), .ZN(n17926) );
  AOI21_X1 U12526 ( .B1(n19440), .B2(n19385), .A(n16810), .ZN(n17929) );
  NAND2_X1 U12527 ( .A1(n17899), .A2(n17917), .ZN(n17933) );
  NOR2_X1 U12528 ( .A1(n17231), .A2(n19010), .ZN(n18001) );
  NOR2_X1 U12529 ( .A1(n18021), .A2(n17676), .ZN(n18052) );
  NOR2_X1 U12530 ( .A1(n21491), .A2(n18056), .ZN(n13469) );
  AND2_X1 U12531 ( .A1(n13658), .A2(n13657), .ZN(n14326) );
  NAND2_X1 U12532 ( .A1(n18131), .A2(n9757), .ZN(n18118) );
  AND2_X1 U12533 ( .A1(n18154), .A2(n9829), .ZN(n18131) );
  INV_X1 U12534 ( .A(n13134), .ZN(n9829) );
  NOR2_X1 U12535 ( .A1(n13134), .A2(n17233), .ZN(n18137) );
  INV_X2 U12536 ( .A(n18151), .ZN(n18148) );
  INV_X1 U12537 ( .A(n18171), .ZN(n18166) );
  NAND2_X1 U12538 ( .A1(n18194), .A2(n9635), .ZN(n18181) );
  NAND2_X1 U12539 ( .A1(n18194), .A2(n18157), .ZN(n18189) );
  NAND2_X1 U12540 ( .A1(n18194), .A2(n9633), .ZN(n18190) );
  NAND2_X1 U12541 ( .A1(n16835), .A2(P3_EAX_REG_17__SCAN_IN), .ZN(n18225) );
  INV_X1 U12542 ( .A(n18221), .ZN(n18223) );
  NOR2_X1 U12543 ( .A1(n18231), .A2(n18300), .ZN(n18156) );
  INV_X1 U12544 ( .A(n18229), .ZN(n18214) );
  NOR2_X1 U12545 ( .A1(n16834), .A2(n10176), .ZN(n10175) );
  INV_X1 U12546 ( .A(n18251), .ZN(n18241) );
  INV_X1 U12547 ( .A(n17153), .ZN(n17151) );
  OR2_X1 U12548 ( .A1(n16893), .A2(n16892), .ZN(n16979) );
  INV_X1 U12549 ( .A(n16899), .ZN(n16964) );
  INV_X1 U12550 ( .A(n10352), .ZN(n16958) );
  INV_X1 U12551 ( .A(n19010), .ZN(n18157) );
  AND3_X1 U12552 ( .A1(n18157), .A2(P3_EAX_REG_2__SCAN_IN), .A3(n13339), .ZN(
        n13353) );
  INV_X1 U12553 ( .A(n13543), .ZN(n13540) );
  OR2_X1 U12554 ( .A1(n18251), .A2(n13372), .ZN(n18255) );
  AND2_X1 U12555 ( .A1(n18295), .A2(n18294), .ZN(n18296) );
  INV_X1 U12556 ( .A(n9883), .ZN(n17027) );
  NOR2_X1 U12557 ( .A1(n18372), .A2(n10164), .ZN(n17055) );
  INV_X1 U12558 ( .A(n10166), .ZN(n10164) );
  NOR2_X1 U12559 ( .A1(n18372), .A2(n18373), .ZN(n18357) );
  NAND2_X1 U12560 ( .A1(n18471), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18454) );
  INV_X1 U12561 ( .A(n17077), .ZN(n18519) );
  INV_X1 U12562 ( .A(n19015), .ZN(n19336) );
  NAND2_X1 U12563 ( .A1(n18642), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18630) );
  INV_X1 U12564 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18629) );
  INV_X1 U12565 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18657) );
  INV_X1 U12566 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18673) );
  OR2_X1 U12567 ( .A1(n19011), .A2(n19085), .ZN(n19015) );
  INV_X1 U12568 ( .A(n18675), .ZN(n18612) );
  AOI21_X1 U12569 ( .B1(n17181), .B2(n19404), .A(n10141), .ZN(n17193) );
  INV_X1 U12570 ( .A(n10142), .ZN(n10141) );
  AOI21_X1 U12571 ( .B1(n17182), .B2(n18712), .A(n9732), .ZN(n10142) );
  NAND2_X1 U12572 ( .A1(n10105), .A2(n10104), .ZN(n16933) );
  OR2_X1 U12573 ( .A1(n18906), .A2(n17151), .ZN(n18873) );
  INV_X1 U12574 ( .A(n18873), .ZN(n18894) );
  NAND2_X1 U12575 ( .A1(n18625), .A2(n16921), .ZN(n18618) );
  INV_X1 U12576 ( .A(n18855), .ZN(n18955) );
  AND2_X1 U12577 ( .A1(n13403), .A2(n19561), .ZN(n18944) );
  NOR2_X1 U12578 ( .A1(n19555), .A2(n17518), .ZN(n19561) );
  INV_X1 U12579 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19555) );
  INV_X1 U12580 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19444) );
  INV_X1 U12581 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19539) );
  AND2_X2 U12582 ( .A1(n12934), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20709)
         );
  NAND2_X1 U12584 ( .A1(n15361), .A2(n20650), .ZN(n15179) );
  NOR2_X1 U12585 ( .A1(n10205), .A2(n12778), .ZN(n9919) );
  NAND2_X1 U12586 ( .A1(n12787), .A2(n9918), .ZN(n9917) );
  AND2_X1 U12587 ( .A1(n10203), .A2(n10202), .ZN(n15357) );
  AOI21_X1 U12588 ( .B1(n15356), .B2(n15355), .A(n15354), .ZN(n10202) );
  NOR2_X1 U12589 ( .A1(n12271), .A2(n12270), .ZN(n12272) );
  INV_X1 U12590 ( .A(n12269), .ZN(n12270) );
  AND2_X1 U12591 ( .A1(n12920), .A2(n12919), .ZN(n12921) );
  OAI21_X1 U12592 ( .B1(n12546), .B2(n16396), .A(n11202), .ZN(P2_U2983) );
  NAND2_X1 U12593 ( .A1(n9637), .A2(n16415), .ZN(n12839) );
  INV_X1 U12594 ( .A(n14367), .ZN(n10016) );
  NAND2_X1 U12595 ( .A1(n12614), .A2(n16394), .ZN(n12615) );
  OAI211_X1 U12596 ( .C1(n16710), .C2(n12546), .A(n9937), .B(n12590), .ZN(
        P2_U3015) );
  NAND2_X1 U12597 ( .A1(n9637), .A2(n19721), .ZN(n12767) );
  OAI211_X1 U12598 ( .C1(n14368), .C2(n16710), .A(n9951), .B(n9950), .ZN(
        P2_U3018) );
  NOR2_X1 U12599 ( .A1(n14363), .A2(n14362), .ZN(n9951) );
  NAND2_X1 U12600 ( .A1(n10053), .A2(n19726), .ZN(n9950) );
  OAI21_X1 U12601 ( .B1(n12846), .B2(n16710), .A(n12828), .ZN(n12829) );
  INV_X1 U12602 ( .A(n9932), .ZN(n9931) );
  NAND2_X1 U12603 ( .A1(n9648), .A2(n9930), .ZN(n9929) );
  OAI211_X1 U12604 ( .C1(n10328), .C2(n16556), .A(n9984), .B(n12810), .ZN(
        P2_U3029) );
  NAND2_X1 U12605 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n10949), .ZN(
        n10328) );
  NAND2_X1 U12606 ( .A1(n10084), .A2(n10085), .ZN(n12810) );
  INV_X1 U12607 ( .A(n17986), .ZN(n17981) );
  INV_X1 U12608 ( .A(n18154), .ZN(n18145) );
  INV_X1 U12609 ( .A(n16991), .ZN(n9784) );
  INV_X2 U12610 ( .A(n11409), .ZN(n11808) );
  NAND3_X2 U12611 ( .A1(n10013), .A2(n10011), .A3(n10010), .ZN(n11068) );
  AND2_X1 U12612 ( .A1(n9614), .A2(n10928), .ZN(n9599) );
  INV_X1 U12613 ( .A(n14348), .ZN(n10136) );
  NAND2_X1 U12614 ( .A1(n10434), .A2(n9756), .ZN(n14991) );
  NOR2_X1 U12615 ( .A1(n13915), .A2(n13783), .ZN(n9600) );
  AND2_X2 U12616 ( .A1(n14007), .A2(n13994), .ZN(n11430) );
  AND2_X1 U12617 ( .A1(n9629), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9601) );
  NAND2_X1 U12618 ( .A1(n20733), .A2(n11993), .ZN(n12108) );
  AND2_X1 U12619 ( .A1(n10405), .A2(n17358), .ZN(n9602) );
  AND3_X1 U12620 ( .A1(n10851), .A2(n9641), .A3(n10596), .ZN(n9603) );
  AND2_X1 U12621 ( .A1(n16710), .A2(n12789), .ZN(n9604) );
  INV_X2 U12622 ( .A(n15324), .ZN(n10416) );
  INV_X1 U12623 ( .A(n15332), .ZN(n15324) );
  AND2_X1 U12624 ( .A1(n10691), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10710) );
  CLKBUF_X3 U12625 ( .A(n13228), .Z(n18098) );
  NAND2_X1 U12626 ( .A1(n14780), .A2(n10439), .ZN(n14757) );
  AND2_X1 U12627 ( .A1(n14899), .A2(n9727), .ZN(n14871) );
  AND2_X1 U12628 ( .A1(n14899), .A2(n11771), .ZN(n14884) );
  NAND2_X1 U12629 ( .A1(n15630), .A2(n10232), .ZN(n9607) );
  AND4_X1 U12630 ( .A1(n13334), .A2(n13333), .A3(n13332), .A4(n13331), .ZN(
        n9608) );
  INV_X1 U12632 ( .A(n10223), .ZN(n10221) );
  AND2_X1 U12633 ( .A1(n12388), .A2(n9762), .ZN(n9610) );
  NOR2_X1 U12634 ( .A1(n15688), .A2(n15687), .ZN(n15675) );
  AND2_X1 U12635 ( .A1(n10310), .A2(n9609), .ZN(n9611) );
  NAND2_X1 U12636 ( .A1(n14414), .A2(n16014), .ZN(n16008) );
  OR3_X1 U12637 ( .A1(n10881), .A2(n10883), .A3(n10025), .ZN(n10886) );
  AND2_X1 U12638 ( .A1(n13754), .A2(n10664), .ZN(n9612) );
  NAND2_X1 U12639 ( .A1(n12699), .A2(n10415), .ZN(n9613) );
  OAI21_X1 U12640 ( .B1(n15449), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n10208), .ZN(n15481) );
  INV_X1 U12641 ( .A(n15481), .ZN(n9921) );
  AND2_X1 U12642 ( .A1(n10129), .A2(n9655), .ZN(n16375) );
  AND2_X1 U12643 ( .A1(n10981), .A2(n10980), .ZN(n9614) );
  INV_X1 U12644 ( .A(n15352), .ZN(n10205) );
  AND2_X1 U12645 ( .A1(n10920), .A2(n10465), .ZN(n9615) );
  AND2_X1 U12646 ( .A1(n10146), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9616) );
  AND2_X1 U12647 ( .A1(n10249), .A2(n10247), .ZN(n9617) );
  AND2_X1 U12648 ( .A1(n14414), .A2(n9728), .ZN(n16003) );
  XNOR2_X1 U12649 ( .A(n11194), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16366) );
  INV_X1 U12650 ( .A(n16366), .ZN(n9925) );
  AND2_X1 U12651 ( .A1(n10427), .A2(n10072), .ZN(n9618) );
  AND2_X1 U12652 ( .A1(n9883), .A2(n9882), .ZN(n9619) );
  AND2_X1 U12653 ( .A1(n9610), .A2(n10402), .ZN(n9620) );
  AND2_X1 U12654 ( .A1(n9615), .A2(n9739), .ZN(n9621) );
  INV_X1 U12655 ( .A(n14243), .ZN(n10434) );
  AND2_X1 U12656 ( .A1(n10033), .A2(n14349), .ZN(n9622) );
  AND2_X1 U12657 ( .A1(n9812), .A2(n9745), .ZN(n9623) );
  AND2_X1 U12658 ( .A1(n9684), .A2(n11087), .ZN(n9624) );
  OAI21_X1 U12659 ( .B1(n9609), .B2(n10314), .A(n9609), .ZN(n10312) );
  AND2_X1 U12660 ( .A1(n12031), .A2(n12034), .ZN(n9625) );
  NOR2_X1 U12661 ( .A1(n15064), .A2(n15154), .ZN(n9626) );
  NOR2_X1 U12662 ( .A1(n12794), .A2(n9733), .ZN(n10086) );
  OR2_X1 U12663 ( .A1(n10112), .A2(n10111), .ZN(n9627) );
  NOR2_X1 U12664 ( .A1(n13913), .A2(n13941), .ZN(n13940) );
  NAND2_X1 U12665 ( .A1(n13904), .A2(n13905), .ZN(n13965) );
  NAND2_X1 U12666 ( .A1(n12389), .A2(n12388), .ZN(n13617) );
  INV_X1 U12667 ( .A(n15800), .ZN(n10298) );
  AND2_X1 U12668 ( .A1(n10237), .A2(n15676), .ZN(n9628) );
  AND2_X1 U12669 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n9629) );
  OAI21_X1 U12670 ( .B1(n15740), .B2(n14277), .A(n16252), .ZN(n15715) );
  INV_X1 U12671 ( .A(n18488), .ZN(n9880) );
  AND2_X1 U12672 ( .A1(n9725), .A2(n10270), .ZN(n9630) );
  AND2_X1 U12673 ( .A1(n9628), .A2(n10236), .ZN(n9631) );
  AND2_X1 U12674 ( .A1(n9601), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9632) );
  AND2_X1 U12675 ( .A1(n12660), .A2(n9763), .ZN(n12669) );
  AND2_X1 U12676 ( .A1(n18157), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n9633) );
  AND2_X1 U12677 ( .A1(n9633), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n9634) );
  INV_X1 U12678 ( .A(n16194), .ZN(n10279) );
  NOR2_X1 U12679 ( .A1(n12658), .A2(n16206), .ZN(n12660) );
  INV_X1 U12680 ( .A(n15618), .ZN(n10274) );
  AND2_X1 U12681 ( .A1(n9634), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n9635) );
  NOR2_X2 U12682 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20463) );
  AND2_X1 U12683 ( .A1(n10196), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9636) );
  INV_X1 U12684 ( .A(n11025), .ZN(n11190) );
  OR2_X1 U12685 ( .A1(n10709), .A2(n10708), .ZN(n11166) );
  INV_X1 U12686 ( .A(n15332), .ZN(n15185) );
  NAND2_X1 U12687 ( .A1(n9959), .A2(n11601), .ZN(n15550) );
  NAND2_X1 U12688 ( .A1(n10181), .A2(n11440), .ZN(n11584) );
  XOR2_X1 U12689 ( .A(n16157), .B(n12766), .Z(n9637) );
  AND2_X1 U12690 ( .A1(n10023), .A2(n10022), .ZN(n10898) );
  NAND2_X1 U12691 ( .A1(n11193), .A2(n16687), .ZN(n9638) );
  OR2_X1 U12692 ( .A1(n12286), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n9639) );
  AND2_X1 U12693 ( .A1(n14780), .A2(n10437), .ZN(n14743) );
  NAND2_X1 U12694 ( .A1(n10919), .A2(n10920), .ZN(n10929) );
  NOR2_X1 U12695 ( .A1(n14243), .A2(n10435), .ZN(n15048) );
  NAND2_X1 U12696 ( .A1(n12460), .A2(n12459), .ZN(n15731) );
  NOR2_X1 U12697 ( .A1(n15649), .A2(n10395), .ZN(n15620) );
  NAND2_X1 U12698 ( .A1(n15675), .A2(n9628), .ZN(n15643) );
  NAND2_X1 U12699 ( .A1(n10273), .A2(n15618), .ZN(n15607) );
  AND2_X1 U12700 ( .A1(n14780), .A2(n11887), .ZN(n14769) );
  AND2_X1 U12701 ( .A1(n10589), .A2(n10593), .ZN(n9641) );
  NAND2_X1 U12702 ( .A1(n10919), .A2(n9615), .ZN(n10951) );
  NOR2_X1 U12703 ( .A1(n15326), .A2(n9869), .ZN(n9642) );
  AND4_X1 U12704 ( .A1(n11380), .A2(n11379), .A3(n11378), .A4(n11377), .ZN(
        n9643) );
  AND2_X1 U12705 ( .A1(n18194), .A2(n9634), .ZN(n9644) );
  OAI21_X1 U12706 ( .B1(n14277), .B2(n10315), .A(n15703), .ZN(n10314) );
  INV_X1 U12707 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14025) );
  AND2_X1 U12708 ( .A1(n11028), .A2(n11027), .ZN(n9645) );
  AND4_X1 U12709 ( .A1(n13338), .A2(n13337), .A3(n13336), .A4(n13335), .ZN(
        n9646) );
  AND4_X1 U12710 ( .A1(n11278), .A2(n11277), .A3(n11276), .A4(n11275), .ZN(
        n9647) );
  INV_X1 U12711 ( .A(n12480), .ZN(n12479) );
  AND2_X1 U12712 ( .A1(n16250), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9648) );
  AND2_X1 U12713 ( .A1(n13396), .A2(n13185), .ZN(n9649) );
  AND2_X1 U12714 ( .A1(n16833), .A2(n10175), .ZN(n9650) );
  NAND2_X1 U12715 ( .A1(n10919), .A2(n9621), .ZN(n9651) );
  AND4_X1 U12716 ( .A1(n10794), .A2(n10786), .A3(n10007), .A4(n10793), .ZN(
        n9652) );
  NOR2_X1 U12717 ( .A1(n16944), .A2(n10109), .ZN(n9654) );
  NAND2_X1 U12718 ( .A1(n10128), .A2(n11178), .ZN(n16401) );
  NAND2_X1 U12719 ( .A1(n11187), .A2(n11180), .ZN(n9655) );
  OAI211_X1 U12720 ( .C1(n11958), .C2(n11443), .A(n11442), .B(n11441), .ZN(
        n12122) );
  INV_X1 U12721 ( .A(n12122), .ZN(n10183) );
  MUX2_X1 U12722 ( .A(n11052), .B(n13644), .S(n10597), .Z(n10866) );
  XNOR2_X1 U12723 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11032), .ZN(
        n9656) );
  OR2_X1 U12724 ( .A1(n15649), .A2(n15650), .ZN(n9657) );
  NOR2_X1 U12725 ( .A1(n12323), .A2(n12448), .ZN(n10389) );
  INV_X1 U12726 ( .A(n10601), .ZN(n10252) );
  NAND2_X1 U12727 ( .A1(n10050), .A2(n10048), .ZN(n16184) );
  AND4_X1 U12728 ( .A1(n12232), .A2(n20715), .A3(n20733), .A4(n11381), .ZN(
        n9658) );
  AND4_X1 U12729 ( .A1(n13103), .A2(n13102), .A3(n13101), .A4(n13100), .ZN(
        n9659) );
  AND2_X1 U12730 ( .A1(n15332), .A2(n12183), .ZN(n9660) );
  AND2_X1 U12731 ( .A1(n13507), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n9661) );
  AND2_X1 U12732 ( .A1(n9857), .A2(n9858), .ZN(n14242) );
  AND2_X1 U12733 ( .A1(n9624), .A2(n11099), .ZN(n9662) );
  AND2_X1 U12734 ( .A1(n12017), .A2(n12016), .ZN(n14195) );
  AND3_X1 U12735 ( .A1(n10967), .A2(n10135), .A3(n12814), .ZN(n9663) );
  INV_X1 U12736 ( .A(n10918), .ZN(n10094) );
  AND2_X1 U12737 ( .A1(n16733), .A2(n12575), .ZN(n9664) );
  NOR2_X1 U12738 ( .A1(n10883), .A2(n10881), .ZN(n9665) );
  NOR2_X1 U12739 ( .A1(n10899), .A2(n10246), .ZN(n10910) );
  INV_X1 U12740 ( .A(n14935), .ZN(n12045) );
  AND2_X1 U12741 ( .A1(n11401), .A2(n11392), .ZN(n9666) );
  AND2_X1 U12742 ( .A1(n10437), .A2(n14744), .ZN(n9667) );
  AND2_X1 U12743 ( .A1(n14966), .A2(n14979), .ZN(n9668) );
  AND2_X1 U12744 ( .A1(n10054), .A2(n10055), .ZN(n9669) );
  AND2_X1 U12745 ( .A1(n12554), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9670) );
  AND2_X1 U12746 ( .A1(n15678), .A2(n12470), .ZN(n15666) );
  NAND4_X1 U12747 ( .A1(n10728), .A2(n10727), .A3(n10726), .A4(n10725), .ZN(
        n9671) );
  AND2_X1 U12748 ( .A1(n10248), .A2(n9617), .ZN(n9672) );
  AND4_X1 U12749 ( .A1(n13052), .A2(n13051), .A3(n13050), .A4(n13049), .ZN(
        n9673) );
  AND3_X1 U12750 ( .A1(n10047), .A2(n9988), .A3(n9987), .ZN(n9674) );
  AND2_X1 U12751 ( .A1(n20702), .A2(n12263), .ZN(n9675) );
  AND3_X1 U12752 ( .A1(n11408), .A2(n11407), .A3(n11406), .ZN(n11460) );
  INV_X1 U12753 ( .A(n11460), .ZN(n9981) );
  AND2_X1 U12754 ( .A1(n10666), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n9677) );
  AND3_X1 U12755 ( .A1(n12554), .A2(n10593), .A3(n13148), .ZN(n9678) );
  INV_X1 U12756 ( .A(n14350), .ZN(n14349) );
  OR2_X1 U12757 ( .A1(n15625), .A2(n11190), .ZN(n14350) );
  AND2_X1 U12758 ( .A1(n10988), .A2(n16200), .ZN(n9679) );
  NOR2_X1 U12759 ( .A1(n17366), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9680) );
  AND2_X1 U12760 ( .A1(n13301), .A2(n12211), .ZN(n9681) );
  AND3_X1 U12761 ( .A1(n13357), .A2(n13356), .A3(n13355), .ZN(n9682) );
  AND2_X1 U12762 ( .A1(n10863), .A2(n10862), .ZN(n9683) );
  AND2_X1 U12763 ( .A1(n12051), .A2(n12050), .ZN(n14901) );
  NAND2_X1 U12764 ( .A1(n10257), .A2(n10253), .ZN(n10583) );
  INV_X1 U12765 ( .A(n10583), .ZN(n10573) );
  INV_X1 U12766 ( .A(n12558), .ZN(n10323) );
  NOR2_X1 U12767 ( .A1(n15797), .A2(n15811), .ZN(n9684) );
  AND2_X1 U12768 ( .A1(n9833), .A2(n9832), .ZN(n9685) );
  INV_X1 U12769 ( .A(n9841), .ZN(n11401) );
  OR2_X1 U12770 ( .A1(n10416), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9686) );
  NAND2_X1 U12771 ( .A1(n11600), .A2(n11543), .ZN(n9687) );
  AND2_X1 U12772 ( .A1(n10050), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9688) );
  NAND2_X1 U12773 ( .A1(n16288), .A2(n16277), .ZN(n9689) );
  AND2_X1 U12774 ( .A1(n9856), .A2(n10427), .ZN(n9690) );
  NAND2_X1 U12775 ( .A1(n15675), .A2(n15676), .ZN(n15660) );
  AND2_X1 U12776 ( .A1(n14348), .A2(n14349), .ZN(n9691) );
  NAND2_X1 U12777 ( .A1(n10272), .A2(n10271), .ZN(n15594) );
  INV_X1 U12778 ( .A(n10385), .ZN(n10384) );
  NAND2_X1 U12779 ( .A1(n10386), .A2(n13146), .ZN(n10385) );
  AND2_X1 U12780 ( .A1(n14013), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n9692) );
  INV_X1 U12781 ( .A(n10314), .ZN(n10313) );
  INV_X1 U12782 ( .A(n10310), .ZN(n10308) );
  NAND2_X1 U12783 ( .A1(n10313), .A2(n10316), .ZN(n10310) );
  INV_X1 U12784 ( .A(n13095), .ZN(n13053) );
  INV_X1 U12785 ( .A(n20461), .ZN(n19739) );
  NAND2_X1 U12786 ( .A1(n11195), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11196) );
  INV_X1 U12787 ( .A(n11196), .ZN(n10339) );
  NAND2_X1 U12788 ( .A1(n15242), .A2(n15241), .ZN(n12695) );
  NAND2_X1 U12789 ( .A1(n10537), .A2(n10538), .ZN(n10598) );
  NOR2_X1 U12790 ( .A1(n12820), .A2(n15692), .ZN(n15678) );
  AND2_X1 U12791 ( .A1(n10301), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9693) );
  AND2_X1 U12792 ( .A1(n10228), .A2(n10226), .ZN(n9694) );
  OR2_X1 U12793 ( .A1(n12135), .A2(n11506), .ZN(n9695) );
  AND2_X1 U12794 ( .A1(n10659), .A2(n15938), .ZN(n9696) );
  AND2_X1 U12795 ( .A1(n10306), .A2(n9609), .ZN(n9697) );
  AND2_X1 U12796 ( .A1(n10416), .A2(n12201), .ZN(n9698) );
  AND2_X1 U12797 ( .A1(n10360), .A2(n10358), .ZN(n9699) );
  NAND2_X1 U12798 ( .A1(n11492), .A2(n12116), .ZN(n9700) );
  AND2_X1 U12799 ( .A1(n11383), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9701) );
  AND2_X1 U12800 ( .A1(n12612), .A2(n10101), .ZN(n9702) );
  AND2_X1 U12801 ( .A1(n9616), .A2(n10145), .ZN(n9703) );
  AND2_X1 U12802 ( .A1(n9625), .A2(n9668), .ZN(n9704) );
  NAND2_X1 U12803 ( .A1(n9837), .A2(n11480), .ZN(n11481) );
  AND2_X1 U12804 ( .A1(n12191), .A2(n12194), .ZN(n9705) );
  AND2_X1 U12805 ( .A1(n15630), .A2(n10231), .ZN(n12755) );
  AND2_X2 U12806 ( .A1(n9844), .A2(n11474), .ZN(n9706) );
  INV_X1 U12807 ( .A(n10219), .ZN(n15261) );
  AND2_X1 U12808 ( .A1(n11326), .A2(n11328), .ZN(n9707) );
  AND2_X1 U12809 ( .A1(n11440), .A2(n9979), .ZN(n9708) );
  INV_X1 U12810 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10302) );
  OAI21_X1 U12811 ( .B1(n16266), .B2(n9609), .A(n9609), .ZN(n10291) );
  NOR2_X1 U12812 ( .A1(n14194), .A2(n10334), .ZN(n14246) );
  NAND2_X1 U12813 ( .A1(n10297), .A2(n16281), .ZN(n15774) );
  NAND2_X1 U12814 ( .A1(n10292), .A2(n10283), .ZN(n15740) );
  NAND2_X1 U12815 ( .A1(n12662), .A2(n15664), .ZN(n15647) );
  NAND2_X1 U12816 ( .A1(n10278), .A2(n16194), .ZN(n15632) );
  NAND2_X1 U12817 ( .A1(n10311), .A2(n10313), .ZN(n15690) );
  INV_X1 U12818 ( .A(n15947), .ZN(n10264) );
  AND2_X1 U12819 ( .A1(n12638), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12641) );
  NAND2_X1 U12820 ( .A1(n10227), .A2(n10228), .ZN(n14081) );
  AND2_X1 U12821 ( .A1(n10307), .A2(n10306), .ZN(n9709) );
  AOI21_X1 U12822 ( .B1(n15715), .B2(n9609), .A(n16237), .ZN(n15702) );
  NAND2_X1 U12823 ( .A1(n12649), .A2(n9629), .ZN(n12654) );
  NAND2_X1 U12824 ( .A1(n12032), .A2(n12031), .ZN(n15051) );
  OR2_X1 U12825 ( .A1(n12634), .A2(n14292), .ZN(n9710) );
  NAND2_X1 U12826 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n9711) );
  AND2_X1 U12827 ( .A1(n12459), .A2(n10400), .ZN(n9712) );
  AND2_X1 U12828 ( .A1(n11105), .A2(n10230), .ZN(n9713) );
  AND2_X1 U12829 ( .A1(n11106), .A2(n9713), .ZN(n9714) );
  AND2_X1 U12830 ( .A1(n14414), .A2(n10268), .ZN(n15996) );
  NAND2_X1 U12831 ( .A1(n11156), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12626) );
  OR2_X1 U12832 ( .A1(n14194), .A2(n14195), .ZN(n14193) );
  AND2_X1 U12833 ( .A1(n10020), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n9715) );
  AND2_X1 U12834 ( .A1(n10020), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n9716) );
  AND2_X1 U12835 ( .A1(n10020), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n9717) );
  OR2_X1 U12836 ( .A1(n18509), .A2(n18811), .ZN(n18708) );
  INV_X1 U12837 ( .A(n18708), .ZN(n10105) );
  OR2_X1 U12838 ( .A1(n12621), .A2(n16418), .ZN(n9718) );
  NAND2_X1 U12839 ( .A1(n12649), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9719) );
  NAND2_X1 U12840 ( .A1(n13895), .A2(n9624), .ZN(n9720) );
  OR2_X1 U12841 ( .A1(n10303), .A2(n16368), .ZN(n9721) );
  NAND2_X1 U12842 ( .A1(n12649), .A2(n9601), .ZN(n9722) );
  NAND2_X1 U12843 ( .A1(n12250), .A2(n13297), .ZN(n20676) );
  NAND2_X1 U12844 ( .A1(n13832), .A2(n11592), .ZN(n13959) );
  NAND2_X1 U12845 ( .A1(n10383), .A2(n10388), .ZN(n13145) );
  AND2_X1 U12846 ( .A1(n10336), .A2(n10335), .ZN(n9723) );
  AND2_X1 U12847 ( .A1(n14073), .A2(n14074), .ZN(n14072) );
  AND2_X1 U12848 ( .A1(n9713), .A2(n15729), .ZN(n9724) );
  AND2_X1 U12849 ( .A1(n13895), .A2(n9662), .ZN(n15769) );
  OR2_X1 U12850 ( .A1(n10830), .A2(n10829), .ZN(n10870) );
  NAND2_X1 U12851 ( .A1(n12032), .A2(n9625), .ZN(n14965) );
  AND4_X1 U12852 ( .A1(n14392), .A2(n16033), .A3(n16039), .A4(n14391), .ZN(
        n9725) );
  AND2_X1 U12853 ( .A1(n15332), .A2(n15353), .ZN(n9726) );
  AND2_X1 U12854 ( .A1(n14886), .A2(n11771), .ZN(n9727) );
  NOR2_X1 U12855 ( .A1(n14084), .A2(n13894), .ZN(n13895) );
  INV_X1 U12856 ( .A(n9609), .ZN(n14277) );
  AND2_X1 U12857 ( .A1(n16014), .A2(n10269), .ZN(n9728) );
  AND2_X1 U12858 ( .A1(n11106), .A2(n9724), .ZN(n12817) );
  AND2_X1 U12859 ( .A1(n10946), .A2(n10455), .ZN(n9729) );
  AND2_X1 U12860 ( .A1(n12547), .A2(n9595), .ZN(n19721) );
  INV_X1 U12861 ( .A(n10983), .ZN(n10241) );
  AND2_X1 U12862 ( .A1(n9712), .A2(n10399), .ZN(n9730) );
  AND2_X1 U12863 ( .A1(n13780), .A2(n10657), .ZN(n9731) );
  OR3_X1 U12864 ( .A1(n18690), .A2(n17184), .A3(n17183), .ZN(n9732) );
  NAND2_X1 U12865 ( .A1(n15909), .A2(n10657), .ZN(n20127) );
  NAND2_X1 U12866 ( .A1(n11156), .A2(n10301), .ZN(n10303) );
  AND2_X1 U12867 ( .A1(n16733), .A2(n16567), .ZN(n9733) );
  AND2_X1 U12868 ( .A1(n10231), .A2(n12757), .ZN(n9734) );
  OR2_X1 U12869 ( .A1(n18372), .A2(n10165), .ZN(n9735) );
  INV_X1 U12870 ( .A(n11381), .ZN(n9953) );
  AND2_X1 U12871 ( .A1(n9723), .A2(n12088), .ZN(n9736) );
  AND2_X1 U12872 ( .A1(n10295), .A2(n10293), .ZN(n9737) );
  AND2_X1 U12873 ( .A1(n10597), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n9738) );
  OR2_X1 U12874 ( .A1(n11022), .A2(n10930), .ZN(n9739) );
  INV_X1 U12875 ( .A(n16225), .ZN(n10316) );
  INV_X1 U12876 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13979) );
  INV_X1 U12877 ( .A(n12721), .ZN(n10224) );
  AND2_X1 U12878 ( .A1(n15332), .A2(n12720), .ZN(n12721) );
  INV_X1 U12879 ( .A(n10233), .ZN(n10232) );
  NAND2_X1 U12880 ( .A1(n10234), .A2(n15614), .ZN(n10233) );
  INV_X1 U12881 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21239) );
  OR2_X1 U12882 ( .A1(n10720), .A2(n10719), .ZN(n11167) );
  NAND2_X1 U12883 ( .A1(n16242), .A2(n12611), .ZN(n16230) );
  OR2_X1 U12884 ( .A1(n10264), .A2(n15953), .ZN(n9740) );
  INV_X1 U12885 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16418) );
  NOR2_X1 U12886 ( .A1(n18508), .A2(n16932), .ZN(n18814) );
  NAND4_X1 U12887 ( .A1(n10428), .A2(n13615), .A3(n13616), .A4(n10429), .ZN(
        n13832) );
  AND2_X1 U12888 ( .A1(n10946), .A2(n10037), .ZN(n9741) );
  AND2_X1 U12889 ( .A1(n10331), .A2(n10330), .ZN(n9742) );
  AND2_X1 U12890 ( .A1(n10597), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n9743) );
  AND2_X1 U12891 ( .A1(n10356), .A2(n18361), .ZN(n9744) );
  AND2_X1 U12892 ( .A1(n10698), .A2(n11167), .ZN(n9745) );
  AND2_X1 U12893 ( .A1(n10268), .A2(n15998), .ZN(n9746) );
  NAND2_X1 U12894 ( .A1(n11532), .A2(n11531), .ZN(n11600) );
  AND2_X1 U12895 ( .A1(n9630), .A2(n16017), .ZN(n9747) );
  AND2_X1 U12896 ( .A1(n9724), .A2(n11120), .ZN(n9748) );
  INV_X1 U12897 ( .A(n13966), .ZN(n13964) );
  OR2_X1 U12898 ( .A1(n12382), .A2(n12381), .ZN(n13966) );
  NAND2_X1 U12899 ( .A1(n12997), .A2(n17221), .ZN(n13229) );
  INV_X1 U12900 ( .A(n17744), .ZN(n17862) );
  NAND2_X1 U12901 ( .A1(n10318), .A2(n10320), .ZN(n12636) );
  NAND2_X1 U12902 ( .A1(n12660), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12663) );
  NAND2_X1 U12903 ( .A1(n12660), .A2(n10281), .ZN(n12666) );
  INV_X1 U12904 ( .A(n17161), .ZN(n9882) );
  INV_X1 U12905 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10247) );
  AND2_X1 U12906 ( .A1(n10020), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n9749) );
  AND2_X1 U12907 ( .A1(n10020), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n9750) );
  AND2_X1 U12908 ( .A1(n10020), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n9751) );
  AND2_X1 U12909 ( .A1(n10020), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n9752) );
  AND2_X1 U12910 ( .A1(n10020), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n9753) );
  AND2_X1 U12911 ( .A1(n10020), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n9754) );
  AND2_X1 U12912 ( .A1(n10020), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n9755) );
  INV_X1 U12913 ( .A(n15644), .ZN(n10236) );
  INV_X1 U12914 ( .A(n15661), .ZN(n10237) );
  INV_X1 U12915 ( .A(n15047), .ZN(n10433) );
  OR2_X1 U12916 ( .A1(n11639), .A2(n11638), .ZN(n9756) );
  NOR2_X1 U12917 ( .A1(n13891), .A2(n13890), .ZN(n14073) );
  NAND2_X1 U12918 ( .A1(n12649), .A2(n9632), .ZN(n12658) );
  INV_X1 U12919 ( .A(n15664), .ZN(n10277) );
  AND3_X1 U12920 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(P3_EBX_REG_6__SCAN_IN), .ZN(n9757) );
  INV_X1 U12921 ( .A(n16189), .ZN(n10245) );
  INV_X1 U12922 ( .A(n10574), .ZN(n14120) );
  INV_X1 U12923 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n9998) );
  AND2_X1 U12924 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n9758) );
  AND2_X1 U12925 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n9759) );
  INV_X1 U12926 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n10072) );
  NOR2_X1 U12927 ( .A1(n16934), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9760) );
  AND2_X1 U12928 ( .A1(n10163), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10161) );
  INV_X1 U12929 ( .A(n10161), .ZN(n10155) );
  AND2_X1 U12930 ( .A1(n10467), .A2(n12672), .ZN(n9761) );
  INV_X1 U12931 ( .A(n10159), .ZN(n10156) );
  NAND2_X1 U12932 ( .A1(n10160), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10159) );
  NAND2_X1 U12933 ( .A1(n12404), .A2(n12403), .ZN(n9762) );
  AND2_X1 U12934 ( .A1(n12816), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12576) );
  INV_X1 U12935 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n10037) );
  INV_X1 U12936 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10350) );
  AND2_X1 U12937 ( .A1(n10281), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9763) );
  OR2_X1 U12938 ( .A1(n12206), .A2(n20715), .ZN(n9764) );
  INV_X1 U12939 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10160) );
  INV_X1 U12940 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10317) );
  INV_X1 U12941 ( .A(n19978), .ZN(n10120) );
  NAND2_X1 U12942 ( .A1(n18615), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18594) );
  INV_X1 U12943 ( .A(n18594), .ZN(n10144) );
  INV_X1 U12944 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10167) );
  AND2_X1 U12945 ( .A1(n12658), .A2(n12659), .ZN(n9765) );
  AND2_X1 U12946 ( .A1(n10020), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n9766) );
  AND2_X1 U12947 ( .A1(n10020), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n9767) );
  INV_X1 U12948 ( .A(n16259), .ZN(n10294) );
  INV_X1 U12949 ( .A(n20044), .ZN(n9805) );
  AND2_X1 U12950 ( .A1(n19849), .A2(n20252), .ZN(n9768) );
  AND2_X1 U12951 ( .A1(n18471), .A2(n10146), .ZN(n9769) );
  NOR2_X1 U12952 ( .A1(n16567), .A2(n12792), .ZN(n9770) );
  INV_X1 U12953 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10282) );
  INV_X1 U12954 ( .A(n16266), .ZN(n10299) );
  NOR2_X1 U12955 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9771) );
  AND3_X1 U12956 ( .A1(n11199), .A2(n14347), .A3(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n9772) );
  AND2_X1 U12957 ( .A1(n10108), .A2(n10110), .ZN(n9773) );
  INV_X1 U12958 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10359) );
  INV_X1 U12959 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10163) );
  INV_X1 U12960 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n10174) );
  INV_X1 U12961 ( .A(n16432), .ZN(n9941) );
  OR2_X1 U12962 ( .A1(n15182), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9774) );
  AND2_X1 U12963 ( .A1(n10340), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9775) );
  INV_X1 U12964 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n9875) );
  INV_X1 U12965 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17154) );
  INV_X1 U12966 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10321) );
  AND2_X1 U12967 ( .A1(n15385), .A2(n15394), .ZN(n9776) );
  AND2_X1 U12968 ( .A1(n9636), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9777) );
  AOI22_X2 U12969 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20762), .B1(DATAI_17_), 
        .B2(n20710), .ZN(n21257) );
  AOI22_X2 U12970 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20762), .B1(DATAI_28_), 
        .B2(n20710), .ZN(n21218) );
  AOI22_X2 U12971 ( .A1(DATAI_21_), .A2(n20710), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20762), .ZN(n21281) );
  AOI22_X2 U12972 ( .A1(DATAI_31_), .A2(n20710), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20762), .ZN(n21234) );
  AOI22_X2 U12973 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20762), .B1(DATAI_30_), 
        .B2(n20710), .ZN(n21226) );
  AOI22_X2 U12974 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20762), .B1(DATAI_26_), 
        .B2(n20710), .ZN(n21210) );
  NOR2_X2 U12975 ( .A1(n20712), .A2(n20711), .ZN(n20762) );
  OR3_X1 U12976 ( .A1(n16491), .A2(n16479), .A3(n16492), .ZN(n16458) );
  NAND2_X1 U12977 ( .A1(n17154), .A2(n17030), .ZN(n10109) );
  NOR2_X4 U12978 ( .A1(n21315), .A2(n21389), .ZN(n21355) );
  AOI22_X2 U12979 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20762), .B1(DATAI_27_), 
        .B2(n20710), .ZN(n21214) );
  CLKBUF_X1 U12980 ( .A(n20895), .Z(n9779) );
  NAND3_X1 U12981 ( .A1(n9784), .A2(n9782), .A3(n9780), .ZN(n16992) );
  NAND2_X1 U12982 ( .A1(n17132), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9781) );
  NAND2_X1 U12983 ( .A1(n17200), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18370) );
  NOR2_X2 U12984 ( .A1(n18808), .A2(n16988), .ZN(n17200) );
  NAND2_X2 U12985 ( .A1(n18584), .A2(n16987), .ZN(n18498) );
  OR2_X2 U12986 ( .A1(n18608), .A2(n17102), .ZN(n9786) );
  NAND2_X1 U12987 ( .A1(n18608), .A2(n17102), .ZN(n9788) );
  AND2_X2 U12988 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17220) );
  INV_X1 U12989 ( .A(n9789), .ZN(n10605) );
  OAI211_X1 U12990 ( .C1(n10193), .C2(n10191), .A(n10189), .B(n10190), .ZN(
        n9789) );
  NAND3_X1 U12991 ( .A1(n10077), .A2(n9793), .A3(n9792), .ZN(n9791) );
  NAND3_X1 U12992 ( .A1(n10006), .A2(n10588), .A3(n10323), .ZN(n9793) );
  NAND2_X1 U12993 ( .A1(n10131), .A2(n10132), .ZN(n10077) );
  NAND2_X1 U12994 ( .A1(n9794), .A2(n10170), .ZN(n14122) );
  NAND2_X1 U12995 ( .A1(n10586), .A2(n9794), .ZN(n11049) );
  NAND3_X1 U12996 ( .A1(n15909), .A2(n10660), .A3(
        P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n9795) );
  AOI21_X1 U12997 ( .B1(n9798), .B2(n20252), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n9832) );
  OAI22_X1 U12998 ( .A1(n9798), .A2(n10752), .B1(n10753), .B2(n20127), .ZN(
        n10754) );
  OR2_X1 U12999 ( .A1(n9798), .A2(n20302), .ZN(n9797) );
  NAND2_X1 U13000 ( .A1(n9803), .A2(n9801), .ZN(n10673) );
  INV_X1 U13001 ( .A(n9896), .ZN(n9802) );
  NAND2_X1 U13002 ( .A1(n20014), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n9803) );
  NAND2_X1 U13003 ( .A1(n20014), .A2(n20304), .ZN(n9806) );
  NAND2_X2 U13004 ( .A1(n9809), .A2(n10611), .ZN(n14108) );
  NAND2_X2 U13005 ( .A1(n10078), .A2(n12498), .ZN(n12509) );
  NAND2_X1 U13006 ( .A1(n10623), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9810) );
  NAND3_X1 U13007 ( .A1(n9811), .A2(n10685), .A3(n10682), .ZN(n9812) );
  AOI21_X1 U13008 ( .B1(n9817), .B2(n9815), .A(n9691), .ZN(n9814) );
  NAND2_X1 U13009 ( .A1(n9820), .A2(n14349), .ZN(n9819) );
  NAND2_X2 U13010 ( .A1(n16389), .A2(n16388), .ZN(n16333) );
  NAND3_X1 U13011 ( .A1(n9822), .A2(n9821), .A3(n20463), .ZN(n20259) );
  NAND2_X1 U13012 ( .A1(n12583), .A2(n12554), .ZN(n12549) );
  NOR2_X2 U13013 ( .A1(n10579), .A2(n10580), .ZN(n12583) );
  NAND3_X1 U13014 ( .A1(n13057), .A2(n13055), .A3(n13056), .ZN(n9825) );
  INV_X2 U13015 ( .A(n18085), .ZN(n18028) );
  AND2_X2 U13016 ( .A1(n9828), .A2(n9827), .ZN(n13396) );
  OR2_X2 U13017 ( .A1(n13194), .A2(n13399), .ZN(n9828) );
  NAND2_X2 U13018 ( .A1(n16367), .A2(n11196), .ZN(n9830) );
  NAND2_X2 U13019 ( .A1(n9830), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9986) );
  NAND2_X1 U13020 ( .A1(n9830), .A2(n12591), .ZN(n16286) );
  NAND2_X1 U13021 ( .A1(n9830), .A2(n16522), .ZN(n16248) );
  OAI21_X2 U13022 ( .B1(n9831), .B2(n11167), .A(n11179), .ZN(n16412) );
  AOI22_X1 U13023 ( .A1(n10122), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n16376), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n9863) );
  NAND2_X1 U13024 ( .A1(n13754), .A2(n13755), .ZN(n9834) );
  XNOR2_X2 U13025 ( .A(n13778), .B(n9836), .ZN(n20465) );
  XNOR2_X2 U13026 ( .A(n13307), .B(n20872), .ZN(n20720) );
  NAND2_X1 U13027 ( .A1(n9910), .A2(n9839), .ZN(n9838) );
  AND2_X4 U13028 ( .A1(n9911), .A2(n13978), .ZN(n11759) );
  AND2_X4 U13029 ( .A1(n14025), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9911) );
  AND2_X1 U13030 ( .A1(n20763), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12904) );
  NAND2_X1 U13031 ( .A1(n11383), .A2(n9843), .ZN(n11386) );
  OAI211_X1 U13032 ( .C1(n11385), .C2(n9953), .A(n14010), .B(n9843), .ZN(
        n12234) );
  NAND2_X1 U13033 ( .A1(n9955), .A2(n9843), .ZN(n9841) );
  AND2_X1 U13034 ( .A1(n20599), .A2(n9843), .ZN(n20596) );
  NAND2_X1 U13035 ( .A1(n12975), .A2(n9843), .ZN(n14043) );
  AND2_X1 U13036 ( .A1(n20752), .A2(n9843), .ZN(n9842) );
  OR2_X2 U13037 ( .A1(n15332), .A2(n12185), .ZN(n15284) );
  NAND2_X1 U13038 ( .A1(n12189), .A2(n15282), .ZN(n15257) );
  NOR2_X2 U13039 ( .A1(n15297), .A2(n12188), .ZN(n15282) );
  NAND2_X2 U13040 ( .A1(n9848), .A2(n9847), .ZN(n15242) );
  NAND4_X1 U13041 ( .A1(n10116), .A2(n9705), .A3(n10403), .A4(n10003), .ZN(
        n9847) );
  NAND2_X1 U13042 ( .A1(n10003), .A2(n12191), .ZN(n15246) );
  NAND2_X2 U13043 ( .A1(n9850), .A2(n9602), .ZN(n10116) );
  INV_X1 U13044 ( .A(n15283), .ZN(n9849) );
  AND2_X2 U13045 ( .A1(n9963), .A2(n12164), .ZN(n9850) );
  INV_X2 U13046 ( .A(n15553), .ZN(n11520) );
  NAND2_X2 U13047 ( .A1(n9851), .A2(n11612), .ZN(n12176) );
  NAND3_X1 U13048 ( .A1(n9852), .A2(n11498), .A3(n11497), .ZN(n11610) );
  XNOR2_X2 U13049 ( .A(n11496), .B(n9860), .ZN(n11497) );
  NAND2_X2 U13050 ( .A1(n10002), .A2(n10184), .ZN(n10185) );
  NAND3_X1 U13051 ( .A1(n13780), .A2(n10657), .A3(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n9905) );
  NAND3_X1 U13052 ( .A1(n9856), .A2(n10426), .A3(n9618), .ZN(n10001) );
  NAND2_X1 U13053 ( .A1(n10000), .A2(n11481), .ZN(n9856) );
  NAND3_X1 U13054 ( .A1(n9857), .A2(n9858), .A3(n14244), .ZN(n14243) );
  NAND2_X1 U13055 ( .A1(n9858), .A2(n11609), .ZN(n14144) );
  NOR2_X4 U13056 ( .A1(n14791), .A2(n14794), .ZN(n14780) );
  INV_X1 U13057 ( .A(n9859), .ZN(n9971) );
  NAND2_X2 U13058 ( .A1(n11499), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9859) );
  NAND2_X1 U13059 ( .A1(n9859), .A2(n9978), .ZN(n9976) );
  INV_X1 U13060 ( .A(n11497), .ZN(n11570) );
  NAND2_X1 U13061 ( .A1(n11497), .A2(n11498), .ZN(n11593) );
  INV_X1 U13062 ( .A(n11495), .ZN(n9860) );
  NAND2_X1 U13063 ( .A1(n9862), .A2(n10194), .ZN(n16367) );
  OAI211_X1 U13064 ( .C1(n10339), .C2(n9862), .A(n9933), .B(n16523), .ZN(
        n16250) );
  NAND3_X2 U13065 ( .A1(n9652), .A2(n21558), .A3(n9864), .ZN(n9939) );
  NOR2_X2 U13066 ( .A1(n10803), .A2(n10802), .ZN(n9864) );
  NAND3_X1 U13068 ( .A1(n11475), .A2(n10072), .A3(n20772), .ZN(n9868) );
  NAND2_X1 U13069 ( .A1(n15334), .A2(n15331), .ZN(n15323) );
  NAND3_X1 U13070 ( .A1(n9874), .A2(n11497), .A3(n11520), .ZN(n11544) );
  INV_X1 U13071 ( .A(n16921), .ZN(n9879) );
  OR2_X2 U13072 ( .A1(n16944), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17162) );
  NAND2_X1 U13073 ( .A1(n9885), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16332) );
  NAND2_X1 U13074 ( .A1(n9861), .A2(n9889), .ZN(n9983) );
  NAND2_X1 U13075 ( .A1(n10669), .A2(n10666), .ZN(n9896) );
  OAI22_X1 U13076 ( .A1(n19879), .A2(n10782), .B1(n9895), .B2(n9894), .ZN(
        n10783) );
  INV_X1 U13077 ( .A(n10669), .ZN(n9895) );
  OAI22_X1 U13078 ( .A1(n10799), .A2(n10758), .B1(n10759), .B2(n9896), .ZN(
        n10760) );
  OAI21_X1 U13079 ( .B1(n9896), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n10119), 
        .ZN(n16779) );
  INV_X1 U13080 ( .A(n16412), .ZN(n9902) );
  NAND2_X1 U13081 ( .A1(n9939), .A2(n9897), .ZN(n11179) );
  NAND3_X1 U13082 ( .A1(n13780), .A2(n10657), .A3(
        P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n9906) );
  NAND3_X1 U13083 ( .A1(n13780), .A2(n10657), .A3(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n9904) );
  NAND2_X1 U13084 ( .A1(n9731), .A2(n20304), .ZN(n9903) );
  OAI21_X1 U13085 ( .B1(n19816), .B2(n10784), .A(n9904), .ZN(n10785) );
  INV_X1 U13086 ( .A(n9910), .ZN(n10220) );
  AND2_X2 U13087 ( .A1(n9911), .A2(n13994), .ZN(n11369) );
  AND2_X2 U13088 ( .A1(n11208), .A2(n9911), .ZN(n11367) );
  AND2_X2 U13089 ( .A1(n11207), .A2(n9911), .ZN(n11366) );
  NAND3_X1 U13090 ( .A1(n11207), .A2(n9911), .A3(
        P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10217) );
  NAND3_X1 U13091 ( .A1(n11208), .A2(n9911), .A3(
        P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10212) );
  NAND3_X1 U13092 ( .A1(n9911), .A2(n13994), .A3(
        P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10213) );
  NOR2_X4 U13093 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13994) );
  AOI21_X1 U13094 ( .B1(n15022), .B2(n20696), .A(n12907), .ZN(n9918) );
  NAND3_X1 U13095 ( .A1(n10846), .A2(n10779), .A3(n9924), .ZN(n10088) );
  NAND2_X1 U13096 ( .A1(n9924), .A2(n10462), .ZN(n10781) );
  INV_X1 U13097 ( .A(n11189), .ZN(n9927) );
  NAND3_X1 U13098 ( .A1(n9931), .A2(n9929), .A3(n9928), .ZN(P2_U3028) );
  OAI21_X1 U13099 ( .B1(n10127), .B2(n16710), .A(n10126), .ZN(n9932) );
  INV_X1 U13100 ( .A(n10194), .ZN(n9934) );
  NAND2_X1 U13101 ( .A1(n11179), .A2(n10040), .ZN(n9936) );
  AND2_X1 U13102 ( .A1(n9939), .A2(n10845), .ZN(n10846) );
  AND2_X1 U13103 ( .A1(n9949), .A2(n12793), .ZN(n16568) );
  OR2_X1 U13104 ( .A1(n9567), .A2(n9604), .ZN(n9949) );
  AND2_X4 U13105 ( .A1(n14014), .A2(n11208), .ZN(n12887) );
  AND2_X2 U13106 ( .A1(n9952), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11208) );
  MUX2_X1 U13107 ( .A(n12232), .B(n11384), .S(n9953), .Z(n11389) );
  NAND2_X1 U13108 ( .A1(n9954), .A2(n11381), .ZN(n21063) );
  INV_X1 U13109 ( .A(n11391), .ZN(n20752) );
  NAND2_X1 U13110 ( .A1(n11593), .A2(n15553), .ZN(n9959) );
  OAI21_X2 U13111 ( .B1(n14191), .B2(n9962), .A(n9961), .ZN(n9963) );
  NAND2_X1 U13112 ( .A1(n10076), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9964) );
  NAND2_X1 U13113 ( .A1(n9968), .A2(n9967), .ZN(n12777) );
  AND2_X2 U13114 ( .A1(n9968), .A2(n10223), .ZN(n15162) );
  NAND2_X1 U13115 ( .A1(n9979), .A2(n11444), .ZN(n9970) );
  NAND3_X1 U13116 ( .A1(n9977), .A2(n9969), .A3(n9976), .ZN(n9975) );
  NAND3_X1 U13117 ( .A1(n9708), .A2(n9977), .A3(n9976), .ZN(n9972) );
  NAND3_X1 U13118 ( .A1(n9977), .A2(n9979), .A3(n9976), .ZN(n11586) );
  OAI21_X1 U13119 ( .B1(n20216), .B2(n10647), .A(n9982), .ZN(n10652) );
  INV_X2 U13120 ( .A(n9986), .ZN(n16352) );
  AOI21_X2 U13121 ( .B1(n16331), .B2(n16638), .A(n16325), .ZN(n16629) );
  NOR2_X2 U13122 ( .A1(n9986), .A2(n9985), .ZN(n16325) );
  NAND3_X1 U13123 ( .A1(n13780), .A2(n10677), .A3(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n9987) );
  INV_X2 U13124 ( .A(n13754), .ZN(n13780) );
  XNOR2_X2 U13125 ( .A(n11061), .B(n10636), .ZN(n13754) );
  AND2_X1 U13126 ( .A1(n17191), .A2(n16943), .ZN(n16944) );
  NAND2_X1 U13127 ( .A1(n9994), .A2(n17191), .ZN(n17049) );
  NAND3_X1 U13128 ( .A1(n9996), .A2(n9997), .A3(n18814), .ZN(n18509) );
  INV_X1 U13129 ( .A(n11475), .ZN(n10000) );
  AND2_X2 U13130 ( .A1(n11387), .A2(n11400), .ZN(n11388) );
  NAND2_X1 U13131 ( .A1(n15257), .A2(n12195), .ZN(n10003) );
  NAND2_X1 U13133 ( .A1(n10611), .A2(n12498), .ZN(n10012) );
  OAI21_X1 U13134 ( .B1(n16275), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10015), .ZN(n16580) );
  XNOR2_X1 U13135 ( .A(n10015), .B(n16567), .ZN(n16274) );
  INV_X1 U13136 ( .A(n10078), .ZN(n12680) );
  OAI211_X1 U13137 ( .C1(n14368), .C2(n16396), .A(n10017), .B(n10016), .ZN(
        P2_U2986) );
  NAND2_X1 U13138 ( .A1(n10053), .A2(n16394), .ZN(n10017) );
  CLKBUF_X1 U13139 ( .A(n14596), .Z(n10019) );
  CLKBUF_X1 U13140 ( .A(n10686), .Z(n10020) );
  AND2_X2 U13141 ( .A1(n10686), .A2(n10551), .ZN(n10818) );
  INV_X1 U13142 ( .A(n10891), .ZN(n10021) );
  INV_X1 U13143 ( .A(n10883), .ZN(n10022) );
  NOR2_X1 U13144 ( .A1(n10024), .A2(n10881), .ZN(n10023) );
  NAND3_X1 U13145 ( .A1(n10054), .A2(n10055), .A3(n10031), .ZN(n10028) );
  NAND3_X1 U13146 ( .A1(n10054), .A2(n10055), .A3(n16218), .ZN(n16199) );
  NAND2_X1 U13147 ( .A1(n10947), .A2(n10946), .ZN(n10935) );
  NAND2_X1 U13148 ( .A1(n10947), .A2(n9741), .ZN(n10934) );
  AND2_X1 U13149 ( .A1(n10050), .A2(n10039), .ZN(n16185) );
  NAND3_X1 U13150 ( .A1(n10996), .A2(n10045), .A3(n10044), .ZN(n10043) );
  NAND3_X1 U13151 ( .A1(n15909), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A3(
        n10660), .ZN(n10047) );
  NAND2_X1 U13152 ( .A1(n9612), .A2(n19727), .ZN(n20088) );
  NAND2_X2 U13153 ( .A1(n16333), .A2(n10908), .ZN(n16320) );
  NAND2_X1 U13154 ( .A1(n10058), .A2(n10057), .ZN(n10532) );
  AND3_X4 U13155 ( .A1(n10868), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n13810), .ZN(n10686) );
  NAND2_X1 U13156 ( .A1(n10560), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10058) );
  XNOR2_X2 U13157 ( .A(n10060), .B(n10059), .ZN(n10653) );
  NAND2_X1 U13158 ( .A1(n10643), .A2(n10619), .ZN(n10060) );
  NAND2_X1 U13159 ( .A1(n10641), .A2(n10654), .ZN(n10643) );
  NAND3_X1 U13160 ( .A1(n11330), .A2(n10063), .A3(n10062), .ZN(n10061) );
  NAND2_X4 U13161 ( .A1(n10065), .A2(n10064), .ZN(n14053) );
  NAND3_X1 U13162 ( .A1(n11333), .A2(n11327), .A3(n11329), .ZN(n10066) );
  AND4_X2 U13163 ( .A1(n9707), .A2(n11331), .A3(n11332), .A4(n11334), .ZN(
        n10064) );
  XNOR2_X2 U13164 ( .A(n10068), .B(n10067), .ZN(n20838) );
  NAND3_X1 U13165 ( .A1(n20642), .A2(n10180), .A3(n10466), .ZN(n10073) );
  NAND2_X1 U13166 ( .A1(n12561), .A2(n10077), .ZN(n12562) );
  NAND2_X1 U13167 ( .A1(n10081), .A2(n10079), .ZN(n11061) );
  NAND3_X1 U13168 ( .A1(n10643), .A2(n10619), .A3(n10239), .ZN(n10079) );
  INV_X1 U13169 ( .A(n10627), .ZN(n10080) );
  INV_X1 U13170 ( .A(n10238), .ZN(n10082) );
  NAND2_X1 U13171 ( .A1(n10627), .A2(n10628), .ZN(n10238) );
  NAND2_X1 U13172 ( .A1(n9567), .A2(n10086), .ZN(n10084) );
  AND2_X2 U13173 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11045) );
  NAND3_X1 U13174 ( .A1(n10090), .A2(n10089), .A3(n10088), .ZN(n10087) );
  NAND2_X1 U13175 ( .A1(n10842), .A2(n11168), .ZN(n10089) );
  NAND2_X1 U13176 ( .A1(n10781), .A2(n10780), .ZN(n10090) );
  OAI21_X1 U13177 ( .B1(n16320), .B2(n10095), .A(n10092), .ZN(n16276) );
  NAND2_X1 U13178 ( .A1(n16558), .A2(n9702), .ZN(n10098) );
  NAND2_X1 U13179 ( .A1(n10098), .A2(n10099), .ZN(n16245) );
  NAND2_X1 U13180 ( .A1(n16558), .A2(n10101), .ZN(n10100) );
  NAND2_X1 U13181 ( .A1(n16558), .A2(n12607), .ZN(n12807) );
  INV_X1 U13182 ( .A(n16944), .ZN(n10107) );
  NAND2_X1 U13183 ( .A1(n10107), .A2(n9773), .ZN(n16947) );
  NAND2_X2 U13184 ( .A1(n14328), .A2(n17217), .ZN(n17239) );
  NAND2_X2 U13185 ( .A1(n20680), .A2(n12142), .ZN(n20642) );
  NAND2_X2 U13186 ( .A1(n10185), .A2(n15218), .ZN(n15210) );
  NAND3_X1 U13187 ( .A1(n11182), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n11183), .ZN(n10123) );
  NAND2_X1 U13188 ( .A1(n10124), .A2(n11185), .ZN(n16387) );
  NAND2_X1 U13189 ( .A1(n11183), .A2(n11182), .ZN(n10124) );
  NAND3_X1 U13190 ( .A1(n10128), .A2(n11178), .A3(n16402), .ZN(n11181) );
  OAI211_X1 U13191 ( .C1(n10595), .C2(n10593), .A(n10130), .B(n10591), .ZN(
        n10132) );
  NAND2_X1 U13192 ( .A1(n10587), .A2(n11049), .ZN(n10588) );
  NAND2_X1 U13193 ( .A1(n10134), .A2(n10133), .ZN(n10527) );
  NOR2_X1 U13194 ( .A1(n9605), .A2(n16159), .ZN(n12747) );
  AND2_X2 U13195 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13451) );
  OR2_X1 U13196 ( .A1(n17000), .A2(n10163), .ZN(n10162) );
  OR3_X1 U13197 ( .A1(n17000), .A2(n10163), .A3(n17712), .ZN(n10150) );
  AOI21_X1 U13198 ( .B1(n17000), .B2(n10161), .A(n10156), .ZN(n10151) );
  NOR2_X1 U13199 ( .A1(n17726), .A2(n10148), .ZN(n17682) );
  OAI21_X1 U13200 ( .B1(n10162), .B2(n18403), .A(n10152), .ZN(n10148) );
  AOI21_X1 U13201 ( .B1(n17000), .B2(n10158), .A(n10157), .ZN(n10149) );
  NAND2_X2 U13202 ( .A1(n10162), .A2(n10151), .ZN(n17744) );
  AOI21_X1 U13203 ( .B1(n17000), .B2(n10154), .A(n10153), .ZN(n10152) );
  NAND2_X2 U13204 ( .A1(n10558), .A2(n12558), .ZN(n12498) );
  NOR2_X2 U13205 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10186) );
  NAND2_X2 U13206 ( .A1(n10526), .A2(n10525), .ZN(n12286) );
  INV_X1 U13207 ( .A(n18057), .ZN(n18112) );
  NOR2_X1 U13208 ( .A1(n9661), .A2(n10172), .ZN(n13050) );
  AND2_X4 U13209 ( .A1(n12991), .A2(n13452), .ZN(n18057) );
  NAND3_X1 U13210 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(P3_EAX_REG_13__SCAN_IN), .ZN(n10176) );
  INV_X1 U13211 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10177) );
  AND2_X4 U13212 ( .A1(n10177), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11207) );
  INV_X1 U13213 ( .A(n12206), .ZN(n10179) );
  OR2_X1 U13214 ( .A1(n20645), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10180) );
  NAND3_X1 U13215 ( .A1(n10185), .A2(n15218), .A3(n9776), .ZN(n12913) );
  OAI22_X1 U13217 ( .A1(n14090), .A2(n14092), .B1(n14089), .B2(n10186), .ZN(
        n14091) );
  NAND2_X1 U13218 ( .A1(n19806), .A2(n10585), .ZN(n10191) );
  INV_X1 U13219 ( .A(n10191), .ZN(n10187) );
  NAND3_X1 U13220 ( .A1(n10187), .A2(n19777), .A3(n12501), .ZN(n10189) );
  NAND2_X1 U13221 ( .A1(n12282), .A2(n10595), .ZN(n10193) );
  NAND2_X1 U13222 ( .A1(n16352), .A2(n9777), .ZN(n10195) );
  NAND2_X1 U13223 ( .A1(n16352), .A2(n9636), .ZN(n16615) );
  NAND2_X1 U13224 ( .A1(n16352), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16331) );
  NAND2_X1 U13225 ( .A1(n10195), .A2(n16590), .ZN(n16287) );
  NAND2_X2 U13226 ( .A1(n11978), .A2(n11977), .ZN(n14213) );
  AND2_X2 U13227 ( .A1(n11207), .A2(n14013), .ZN(n11424) );
  AND2_X2 U13228 ( .A1(n14014), .A2(n13978), .ZN(n11432) );
  NAND4_X1 U13229 ( .A1(n10214), .A2(n10213), .A3(n10212), .A4(n10211), .ZN(
        n10218) );
  NAND3_X1 U13230 ( .A1(n14014), .A2(n13978), .A3(
        P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10211) );
  NAND3_X1 U13231 ( .A1(n11207), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A3(
        n14007), .ZN(n10214) );
  NAND2_X1 U13232 ( .A1(n15185), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10219) );
  NAND3_X1 U13233 ( .A1(n11498), .A2(n11520), .A3(n11497), .ZN(n11601) );
  NAND2_X1 U13234 ( .A1(n15324), .A2(n12722), .ZN(n10223) );
  NAND2_X1 U13235 ( .A1(n10227), .A2(n9694), .ZN(n14084) );
  NAND2_X1 U13236 ( .A1(n11106), .A2(n9748), .ZN(n15688) );
  NAND2_X1 U13237 ( .A1(n15630), .A2(n15614), .ZN(n15616) );
  NAND2_X1 U13238 ( .A1(n13895), .A2(n10235), .ZN(n12795) );
  NAND2_X1 U13239 ( .A1(n15675), .A2(n9631), .ZN(n15645) );
  NAND2_X1 U13240 ( .A1(n10982), .A2(n10240), .ZN(n10990) );
  NAND2_X1 U13241 ( .A1(n10982), .A2(n10983), .ZN(n10989) );
  NAND2_X1 U13242 ( .A1(n10990), .A2(n9743), .ZN(n10991) );
  NAND2_X2 U13243 ( .A1(n10739), .A2(n10243), .ZN(n11025) );
  NAND2_X1 U13244 ( .A1(n10947), .A2(n9729), .ZN(n10961) );
  NAND2_X4 U13245 ( .A1(n10608), .A2(n9603), .ZN(n11152) );
  NOR2_X2 U13246 ( .A1(n10607), .A2(n12504), .ZN(n10608) );
  AND2_X2 U13247 ( .A1(n12512), .A2(n10598), .ZN(n12554) );
  NAND4_X1 U13248 ( .A1(n10552), .A2(n10554), .A3(n10553), .A4(n10254), .ZN(
        n10253) );
  NAND4_X1 U13249 ( .A1(n10555), .A2(n10556), .A3(n10557), .A4(n10258), .ZN(
        n10257) );
  NAND2_X1 U13250 ( .A1(n15960), .A2(n10267), .ZN(n10265) );
  OAI211_X1 U13251 ( .C1(n14595), .C2(n9740), .A(n10261), .B(n14617), .ZN(
        n14640) );
  NAND2_X1 U13252 ( .A1(n15960), .A2(n10262), .ZN(n10261) );
  NAND2_X1 U13253 ( .A1(n15948), .A2(n15947), .ZN(n16045) );
  NAND2_X1 U13254 ( .A1(n10265), .A2(n10266), .ZN(n15948) );
  AND2_X2 U13255 ( .A1(n14414), .A2(n9746), .ZN(n15991) );
  NAND2_X1 U13256 ( .A1(n13904), .A2(n9747), .ZN(n16013) );
  NAND2_X1 U13257 ( .A1(n15617), .A2(n9609), .ZN(n10272) );
  NAND2_X1 U13258 ( .A1(n10275), .A2(n9609), .ZN(n12668) );
  NAND2_X1 U13259 ( .A1(n12662), .A2(n10276), .ZN(n10275) );
  NAND3_X1 U13260 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12621) );
  OAI22_X1 U13261 ( .A1(n9609), .A2(n10287), .B1(n9609), .B2(n10285), .ZN(
        n10284) );
  NAND2_X1 U13262 ( .A1(n11156), .A2(n10300), .ZN(n12631) );
  NAND2_X1 U13263 ( .A1(n15715), .A2(n9697), .ZN(n10304) );
  NAND2_X1 U13264 ( .A1(n10304), .A2(n10305), .ZN(n15663) );
  INV_X1 U13265 ( .A(n15715), .ZN(n10309) );
  NAND2_X1 U13266 ( .A1(n12584), .A2(n10324), .ZN(n13807) );
  AND2_X2 U13267 ( .A1(n12032), .A2(n9704), .ZN(n14968) );
  NAND4_X1 U13268 ( .A1(n10346), .A2(n10606), .A3(n10343), .A4(n10341), .ZN(
        n10637) );
  XNOR2_X1 U13269 ( .A(n9656), .B(n10347), .ZN(n12548) );
  XNOR2_X1 U13270 ( .A(n16959), .B(n10352), .ZN(n13405) );
  NAND2_X1 U13271 ( .A1(n18378), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10360) );
  NAND3_X1 U13272 ( .A1(n10360), .A2(n10354), .A3(n9744), .ZN(n17191) );
  NOR2_X1 U13273 ( .A1(n10357), .A2(n10355), .ZN(n10358) );
  NAND2_X1 U13274 ( .A1(n10114), .A2(n10359), .ZN(n10356) );
  OAI21_X1 U13275 ( .B1(n10362), .B2(n10361), .A(n16940), .ZN(n17198) );
  OAI21_X1 U13276 ( .B1(n18488), .B2(n16934), .A(n16933), .ZN(n18476) );
  NAND2_X1 U13277 ( .A1(n12602), .A2(n12601), .ZN(n16309) );
  INV_X1 U13278 ( .A(n12601), .ZN(n10371) );
  AOI21_X1 U13279 ( .B1(n10376), .B2(n9606), .A(n16232), .ZN(n10373) );
  NAND2_X1 U13280 ( .A1(n15881), .A2(n10378), .ZN(n10377) );
  NAND2_X1 U13281 ( .A1(n10377), .A2(n10380), .ZN(n13156) );
  INV_X1 U13282 ( .A(n10389), .ZN(n10388) );
  NAND2_X1 U13283 ( .A1(n15613), .A2(n10390), .ZN(P2_U2827) );
  INV_X1 U13284 ( .A(n10391), .ZN(n10390) );
  OR2_X1 U13285 ( .A1(n15955), .A2(n15937), .ZN(n10394) );
  NAND2_X1 U13286 ( .A1(n12460), .A2(n10398), .ZN(n12820) );
  NAND2_X1 U13287 ( .A1(n12389), .A2(n10401), .ZN(n13787) );
  NAND2_X1 U13288 ( .A1(n12700), .A2(n10411), .ZN(n10409) );
  NAND2_X1 U13289 ( .A1(n12700), .A2(n12699), .ZN(n15224) );
  NAND2_X1 U13290 ( .A1(n12701), .A2(n9698), .ZN(n10413) );
  NAND2_X1 U13291 ( .A1(n15242), .A2(n10421), .ZN(n10420) );
  NAND2_X1 U13292 ( .A1(n11475), .A2(n10425), .ZN(n10426) );
  NAND2_X1 U13293 ( .A1(n15547), .A2(n11576), .ZN(n10428) );
  INV_X1 U13294 ( .A(n14243), .ZN(n10431) );
  NAND2_X1 U13295 ( .A1(n10431), .A2(n10432), .ZN(n14911) );
  INV_X1 U13296 ( .A(n16402), .ZN(n16403) );
  INV_X1 U13297 ( .A(n12627), .ZN(n11156) );
  NAND2_X1 U13298 ( .A1(n11007), .A2(n11008), .ZN(n11014) );
  NAND2_X1 U13299 ( .A1(n12343), .A2(n12342), .ZN(n13165) );
  INV_X1 U13300 ( .A(n13156), .ZN(n12343) );
  NAND2_X1 U13301 ( .A1(n10593), .A2(n10594), .ZN(n10590) );
  INV_X1 U13302 ( .A(n10594), .ZN(n10597) );
  NAND2_X1 U13303 ( .A1(n12279), .A2(n12278), .ZN(n13929) );
  AND2_X1 U13304 ( .A1(n12289), .A2(n9595), .ZN(n10599) );
  BUF_X1 U13305 ( .A(n12695), .Z(n15430) );
  INV_X1 U13306 ( .A(n12115), .ZN(n11578) );
  NAND2_X1 U13307 ( .A1(n12453), .A2(n12452), .ZN(n14066) );
  NAND2_X1 U13308 ( .A1(n11181), .A2(n11186), .ZN(n11182) );
  INV_X1 U13309 ( .A(n13787), .ZN(n12453) );
  XNOR2_X1 U13310 ( .A(n12753), .B(n12481), .ZN(n12692) );
  NAND2_X1 U13311 ( .A1(n14690), .A2(n19724), .ZN(n12765) );
  XNOR2_X2 U13312 ( .A(n14548), .B(n14547), .ZN(n15973) );
  AOI21_X2 U13313 ( .B1(n15976), .B2(n14510), .A(n14509), .ZN(n14548) );
  AOI22_X1 U13314 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9572), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10542) );
  AOI22_X1 U13315 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10506) );
  NAND2_X1 U13316 ( .A1(n10691), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10486) );
  NAND2_X1 U13317 ( .A1(n10581), .A2(n10594), .ZN(n12289) );
  INV_X1 U13318 ( .A(n10594), .ZN(n10576) );
  INV_X1 U13319 ( .A(n14710), .ZN(n15071) );
  XOR2_X1 U13320 ( .A(n14369), .B(n14729), .Z(n14710) );
  AND2_X1 U13321 ( .A1(n10653), .A2(n15938), .ZN(n10674) );
  NAND2_X1 U13322 ( .A1(n12548), .A2(n19726), .ZN(n12590) );
  INV_X1 U13323 ( .A(n11979), .ZN(n12225) );
  NAND2_X1 U13324 ( .A1(n12871), .A2(n14730), .ZN(n14729) );
  NOR2_X2 U13325 ( .A1(n11913), .A2(n11915), .ZN(n12871) );
  INV_X1 U13326 ( .A(n14145), .ZN(n11609) );
  NAND2_X1 U13327 ( .A1(n10668), .A2(n19727), .ZN(n19879) );
  NAND2_X1 U13328 ( .A1(n10668), .A2(n10659), .ZN(n10799) );
  OR2_X1 U13330 ( .A1(n12220), .A2(n11995), .ZN(n12243) );
  XNOR2_X1 U13331 ( .A(n12906), .B(n12905), .ZN(n14721) );
  INV_X1 U13332 ( .A(n14575), .ZN(n14574) );
  INV_X1 U13333 ( .A(n12286), .ZN(n10596) );
  OR2_X1 U13334 ( .A1(n15929), .A2(n15928), .ZN(P2_U2853) );
  OR2_X1 U13335 ( .A1(n15880), .A2(n15879), .ZN(P2_U2849) );
  INV_X1 U13336 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n15584) );
  NOR2_X4 U13337 ( .A1(n18353), .A2(n18298), .ZN(n10447) );
  AND2_X1 U13338 ( .A1(n12814), .A2(n12813), .ZN(n10448) );
  NOR2_X1 U13339 ( .A1(n17397), .A2(n14246), .ZN(n10449) );
  NAND2_X2 U13340 ( .A1(n15157), .A2(n13612), .ZN(n15158) );
  OR2_X1 U13341 ( .A1(n14144), .A2(n15064), .ZN(n10450) );
  NOR2_X1 U13342 ( .A1(n12759), .A2(n16186), .ZN(n10451) );
  NOR2_X1 U13343 ( .A1(n15543), .A2(n21155), .ZN(n10452) );
  NOR2_X1 U13344 ( .A1(n14354), .A2(n15622), .ZN(n10453) );
  AND3_X1 U13345 ( .A1(n13343), .A2(n13342), .A3(n13341), .ZN(n10454) );
  OR2_X1 U13346 ( .A1(n11022), .A2(n10936), .ZN(n10455) );
  AND4_X1 U13347 ( .A1(n13695), .A2(n13694), .A3(n13693), .A4(n13692), .ZN(
        n10456) );
  INV_X1 U13348 ( .A(n19524), .ZN(n19568) );
  NOR2_X1 U13349 ( .A1(n15636), .A2(n15620), .ZN(n10457) );
  INV_X1 U13350 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18882) );
  INV_X1 U13351 ( .A(n15412), .ZN(n12197) );
  NAND2_X1 U13352 ( .A1(n12641), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10459) );
  INV_X1 U13353 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11465) );
  INV_X1 U13354 ( .A(n16396), .ZN(n16415) );
  INV_X1 U13355 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12778) );
  INV_X1 U13356 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15834) );
  INV_X1 U13357 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13074) );
  OR2_X1 U13358 ( .A1(n14413), .A2(n14412), .ZN(n16014) );
  OR2_X1 U13359 ( .A1(n12369), .A2(n12368), .ZN(n13905) );
  AND2_X1 U13360 ( .A1(n19531), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19468) );
  AND2_X1 U13361 ( .A1(n10701), .A2(n10700), .ZN(n10460) );
  OR2_X1 U13362 ( .A1(n11022), .A2(n10986), .ZN(n10461) );
  INV_X1 U13363 ( .A(n16029), .ZN(n16037) );
  NAND2_X1 U13364 ( .A1(n15999), .A2(n19806), .ZN(n16029) );
  INV_X1 U13365 ( .A(n14713), .ZN(n11461) );
  AND2_X1 U13366 ( .A1(n10843), .A2(n11190), .ZN(n10462) );
  AND4_X1 U13367 ( .A1(n10485), .A2(n10484), .A3(n10483), .A4(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10463) );
  INV_X1 U13368 ( .A(n10653), .ZN(n10659) );
  INV_X1 U13369 ( .A(n19727), .ZN(n10666) );
  AND2_X1 U13370 ( .A1(n12774), .A2(n12773), .ZN(n10464) );
  INV_X1 U13371 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16311) );
  INV_X1 U13372 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15739) );
  OR2_X1 U13373 ( .A1(n11022), .A2(n11093), .ZN(n10465) );
  OR2_X1 U13374 ( .A1(n12143), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10466) );
  INV_X1 U13375 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13077) );
  NAND2_X1 U13376 ( .A1(n12669), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10467) );
  INV_X1 U13377 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17886) );
  INV_X1 U13378 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21000) );
  INV_X1 U13379 ( .A(n21163), .ZN(n21376) );
  OR2_X1 U13380 ( .A1(n15867), .A2(n15866), .ZN(P2_U2848) );
  OR2_X1 U13381 ( .A1(n15853), .A2(n15852), .ZN(P2_U2846) );
  AND2_X1 U13382 ( .A1(n11597), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10470) );
  OR2_X1 U13383 ( .A1(n15972), .A2(n15964), .ZN(n10471) );
  AND2_X1 U13384 ( .A1(n17930), .A2(n13414), .ZN(n13496) );
  AND2_X1 U13385 ( .A1(n13182), .A2(n13386), .ZN(n10472) );
  AND2_X1 U13386 ( .A1(n12765), .A2(n12764), .ZN(n10473) );
  INV_X1 U13387 ( .A(n11759), .ZN(n11409) );
  AND2_X2 U13388 ( .A1(n13978), .A2(n14013), .ZN(n11375) );
  AND4_X1 U13389 ( .A1(n11373), .A2(n11372), .A3(n11371), .A4(n11370), .ZN(
        n10474) );
  AND4_X1 U13390 ( .A1(n11296), .A2(n11295), .A3(n11294), .A4(n11293), .ZN(
        n10475) );
  XNOR2_X1 U13391 ( .A(n11469), .B(n11470), .ZN(n11577) );
  AND4_X1 U13392 ( .A1(n11282), .A2(n11281), .A3(n11280), .A4(n11279), .ZN(
        n10476) );
  NAND2_X1 U13393 ( .A1(n13717), .A2(n13716), .ZN(n13718) );
  INV_X1 U13394 ( .A(n19604), .ZN(n19705) );
  INV_X1 U13395 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13998) );
  AND2_X1 U13396 ( .A1(n21157), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11936) );
  AOI22_X1 U13397 ( .A1(n11411), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11424), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11377) );
  NAND2_X1 U13398 ( .A1(n12225), .A2(n12091), .ZN(n11463) );
  NAND2_X1 U13399 ( .A1(n12482), .A2(n10861), .ZN(n10862) );
  INV_X1 U13400 ( .A(n10589), .ZN(n10595) );
  AOI22_X1 U13401 ( .A1(n10691), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10547) );
  OR2_X1 U13402 ( .A1(n11530), .A2(n11529), .ZN(n12150) );
  NOR2_X1 U13403 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20708), .ZN(
        n11970) );
  NOR2_X1 U13404 ( .A1(n9596), .A2(n10584), .ZN(n10587) );
  OR2_X1 U13405 ( .A1(n11274), .A2(n11273), .ZN(n11898) );
  AND2_X1 U13406 ( .A1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11320) );
  OR2_X1 U13407 ( .A1(n11564), .A2(n11563), .ZN(n12167) );
  OR2_X1 U13408 ( .A1(n11969), .A2(n11968), .ZN(n11972) );
  INV_X1 U13409 ( .A(n11439), .ZN(n11440) );
  INV_X1 U13410 ( .A(n14068), .ZN(n12452) );
  INV_X1 U13411 ( .A(n13167), .ZN(n12342) );
  NAND2_X1 U13412 ( .A1(n14664), .A2(n12309), .ZN(n14662) );
  NAND2_X1 U13413 ( .A1(n12508), .A2(n10575), .ZN(n10580) );
  AND2_X1 U13414 ( .A1(n10594), .A2(n20304), .ZN(n12281) );
  AND2_X1 U13415 ( .A1(n10487), .A2(n10486), .ZN(n10488) );
  AND2_X1 U13416 ( .A1(n19395), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13088) );
  MUX2_X1 U13417 ( .A(n12085), .B(n11995), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n11997) );
  NAND2_X1 U13418 ( .A1(n11374), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11339) );
  AND2_X1 U13419 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11317) );
  NAND2_X1 U13420 ( .A1(n12197), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12198) );
  AND2_X1 U13421 ( .A1(n11972), .A2(n11971), .ZN(n11981) );
  INV_X1 U13422 ( .A(n12220), .ZN(n12232) );
  XNOR2_X1 U13423 ( .A(n10855), .B(n10849), .ZN(n12484) );
  OR2_X1 U13424 ( .A1(n14552), .A2(n15964), .ZN(n14570) );
  INV_X1 U13425 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16292) );
  AND2_X1 U13426 ( .A1(n16770), .A2(n20459), .ZN(n16771) );
  AOI21_X1 U13427 ( .B1(n13090), .B2(n13089), .A(n13088), .ZN(n13184) );
  AND2_X1 U13428 ( .A1(n13394), .A2(n13377), .ZN(n13378) );
  INV_X1 U13429 ( .A(n14950), .ZN(n20555) );
  INV_X1 U13430 ( .A(n15052), .ZN(n12034) );
  INV_X1 U13431 ( .A(n15058), .ZN(n12031) );
  AND4_X1 U13432 ( .A1(n11342), .A2(n11341), .A3(n11340), .A4(n11339), .ZN(
        n11353) );
  NAND2_X1 U13433 ( .A1(n13995), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12868) );
  NAND2_X1 U13434 ( .A1(n11730), .A2(n11317), .ZN(n11713) );
  AOI21_X1 U13435 ( .B1(n12110), .B2(n11727), .A(n11608), .ZN(n14145) );
  AND2_X1 U13436 ( .A1(n11461), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11597) );
  OR2_X1 U13437 ( .A1(n12173), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17359) );
  AND2_X1 U13438 ( .A1(n12216), .A2(n12215), .ZN(n13299) );
  AND2_X1 U13439 ( .A1(n14053), .A2(n11391), .ZN(n13462) );
  INV_X1 U13440 ( .A(n12212), .ZN(n13995) );
  NOR2_X1 U13441 ( .A1(n20994), .A2(n20993), .ZN(n21094) );
  NAND2_X1 U13442 ( .A1(n20747), .A2(n12169), .ZN(n11441) );
  AND2_X2 U13443 ( .A1(n11519), .A2(n11518), .ZN(n15553) );
  AOI21_X1 U13444 ( .B1(n9609), .B2(n15799), .A(n16294), .ZN(n15800) );
  XNOR2_X1 U13445 ( .A(n13772), .B(n10635), .ZN(n10636) );
  NAND2_X1 U13446 ( .A1(n13769), .A2(n13768), .ZN(n13902) );
  OR2_X1 U13447 ( .A1(n14570), .A2(n14578), .ZN(n14611) );
  NAND2_X1 U13448 ( .A1(n15666), .A2(n15667), .ZN(n15649) );
  AND2_X1 U13449 ( .A1(n12455), .A2(n12454), .ZN(n15772) );
  AND2_X1 U13450 ( .A1(n12359), .A2(n12358), .ZN(n13488) );
  OR2_X1 U13451 ( .A1(n14353), .A2(n15599), .ZN(n15601) );
  AND2_X1 U13452 ( .A1(n12467), .A2(n12466), .ZN(n15692) );
  OR2_X1 U13453 ( .A1(n15754), .A2(n10976), .ZN(n12612) );
  OR2_X1 U13454 ( .A1(n10971), .A2(n16602), .ZN(n16301) );
  NAND2_X1 U13455 ( .A1(n13923), .A2(n13922), .ZN(n13921) );
  NAND2_X1 U13456 ( .A1(n14153), .A2(n12496), .ZN(n12497) );
  INV_X1 U13457 ( .A(n19795), .ZN(n19807) );
  AND2_X1 U13458 ( .A1(n18583), .A2(n21475), .ZN(n18462) );
  INV_X1 U13459 ( .A(n18868), .ZN(n18861) );
  NOR2_X1 U13460 ( .A1(n16965), .A2(n16964), .ZN(n16963) );
  NOR2_X1 U13461 ( .A1(n13197), .A2(n13195), .ZN(n13382) );
  AND3_X1 U13462 ( .A1(n13060), .A2(n13059), .A3(n13058), .ZN(n13065) );
  AND2_X1 U13463 ( .A1(n14733), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n12103) );
  NAND2_X1 U13464 ( .A1(n12097), .A2(n12096), .ZN(n14950) );
  AND2_X1 U13465 ( .A1(n12063), .A2(n12062), .ZN(n14837) );
  INV_X1 U13466 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15267) );
  INV_X1 U13467 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11549) );
  NAND2_X1 U13468 ( .A1(n12698), .A2(n10416), .ZN(n12699) );
  INV_X1 U13469 ( .A(n20702), .ZN(n15449) );
  INV_X1 U13470 ( .A(n21188), .ZN(n21194) );
  OR2_X1 U13471 ( .A1(n15547), .A2(n11520), .ZN(n20902) );
  NOR2_X1 U13472 ( .A1(n20873), .A2(n20775), .ZN(n21050) );
  INV_X1 U13473 ( .A(n15547), .ZN(n15551) );
  INV_X1 U13474 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21186) );
  OR2_X1 U13475 ( .A1(n20775), .A2(n21000), .ZN(n20764) );
  INV_X1 U13476 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15790) );
  INV_X1 U13477 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n14292) );
  NAND2_X1 U13478 ( .A1(n14253), .A2(n12682), .ZN(n15875) );
  NAND2_X1 U13479 ( .A1(n13149), .A2(n12527), .ZN(n16140) );
  AND2_X1 U13480 ( .A1(n16151), .A2(n12515), .ZN(n13149) );
  NAND2_X1 U13481 ( .A1(n12525), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n16772)
         );
  INV_X1 U13482 ( .A(n12941), .ZN(n12685) );
  INV_X1 U13483 ( .A(n12612), .ZN(n12811) );
  OR2_X1 U13484 ( .A1(n10959), .A2(n16604), .ZN(n16307) );
  AND2_X1 U13485 ( .A1(n10896), .A2(n10895), .ZN(n16388) );
  AOI22_X1 U13486 ( .A1(n13757), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20463), .B2(n20248), .ZN(n13174) );
  INV_X1 U13487 ( .A(n20463), .ZN(n20252) );
  NAND2_X1 U13488 ( .A1(n13389), .A2(n13387), .ZN(n19401) );
  NAND2_X1 U13489 ( .A1(n17665), .A2(n18413), .ZN(n17664) );
  INV_X1 U13490 ( .A(n17933), .ZN(n17699) );
  INV_X1 U13491 ( .A(n17929), .ZN(n17899) );
  OR2_X1 U13492 ( .A1(n18586), .A2(n18581), .ZN(n16997) );
  INV_X1 U13493 ( .A(n18759), .ZN(n18766) );
  AND2_X2 U13494 ( .A1(n18868), .A2(n18839), .ZN(n18792) );
  INV_X1 U13495 ( .A(n14332), .ZN(n17227) );
  AOI221_X1 U13496 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n19555), .C1(n19444), 
        .C2(P3_STATE2_REG_2__SCAN_IN), .A(n17227), .ZN(n18977) );
  INV_X1 U13497 ( .A(n19438), .ZN(n19385) );
  OR2_X1 U13498 ( .A1(n12960), .A2(n14227), .ZN(n12965) );
  OR2_X1 U13499 ( .A1(n12104), .A2(n12103), .ZN(n12105) );
  AND2_X1 U13500 ( .A1(n20545), .A2(n14948), .ZN(n20511) );
  AND2_X1 U13501 ( .A1(n20562), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20579) );
  AND2_X1 U13502 ( .A1(n15157), .A2(n20763), .ZN(n14714) );
  NOR2_X2 U13503 ( .A1(n14715), .A2(n20709), .ZN(n15137) );
  INV_X1 U13504 ( .A(n20633), .ZN(n13587) );
  NAND2_X1 U13505 ( .A1(n11583), .A2(n11582), .ZN(n13616) );
  OR2_X1 U13506 ( .A1(n15029), .A2(n20668), .ZN(n12920) );
  AND2_X1 U13507 ( .A1(n12250), .A2(n12228), .ZN(n20696) );
  OAI22_X1 U13508 ( .A1(n20730), .A2(n20729), .B1(n20728), .B2(n21054), .ZN(
        n20768) );
  OAI21_X1 U13509 ( .B1(n20730), .B2(n20726), .A(n20724), .ZN(n20769) );
  OAI22_X1 U13510 ( .A1(n20806), .A2(n20805), .B1(n21054), .B2(n20932), .ZN(
        n20829) );
  OAI211_X1 U13511 ( .C1(n20806), .C2(n20804), .A(n21050), .B(n20803), .ZN(
        n20830) );
  OAI21_X1 U13512 ( .B1(n20844), .B2(n20842), .A(n20841), .ZN(n20868) );
  INV_X1 U13513 ( .A(n20956), .ZN(n20921) );
  OAI22_X1 U13514 ( .A1(n20934), .A2(n20933), .B1(n20932), .B2(n21185), .ZN(
        n20958) );
  OAI211_X1 U13515 ( .C1(n21163), .C2(n11500), .A(n20969), .B(n21245), .ZN(
        n20988) );
  INV_X1 U13516 ( .A(n20983), .ZN(n21017) );
  INV_X1 U13517 ( .A(n21085), .ZN(n21041) );
  AND2_X1 U13518 ( .A1(n15543), .A2(n21155), .ZN(n21189) );
  OAI22_X1 U13519 ( .A1(n21134), .A2(n21133), .B1(n21185), .B2(n21132), .ZN(
        n21150) );
  NOR2_X2 U13520 ( .A1(n21244), .A2(n21122), .ZN(n21180) );
  OAI211_X1 U13521 ( .C1(n21227), .C2(n21198), .A(n21197), .B(n21196), .ZN(
        n21230) );
  INV_X1 U13522 ( .A(n21063), .ZN(n21258) );
  INV_X1 U13523 ( .A(n21075), .ZN(n21276) );
  INV_X1 U13524 ( .A(n14223), .ZN(n14214) );
  INV_X1 U13525 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21315) );
  CLKBUF_X1 U13526 ( .A(n21342), .Z(n21351) );
  AND2_X1 U13527 ( .A1(n19700), .A2(n12691), .ZN(n15933) );
  INV_X1 U13528 ( .A(n15875), .ZN(n19609) );
  NAND2_X1 U13529 ( .A1(n13719), .A2(n13718), .ZN(n20461) );
  AND2_X1 U13530 ( .A1(n13149), .A2(n16770), .ZN(n16136) );
  INV_X1 U13531 ( .A(n19648), .ZN(n16056) );
  NOR2_X1 U13532 ( .A1(n16758), .A2(n13176), .ZN(n19652) );
  NOR2_X1 U13533 ( .A1(n19700), .A2(n13703), .ZN(n13795) );
  AND2_X1 U13534 ( .A1(n12685), .A2(n9595), .ZN(n13877) );
  OAI21_X1 U13535 ( .B1(n12846), .B2(n16396), .A(n12845), .ZN(n12847) );
  INV_X1 U13536 ( .A(n16555), .ZN(n12614) );
  AND2_X1 U13537 ( .A1(n15814), .A2(n15813), .ZN(n16608) );
  NOR2_X2 U13538 ( .A1(n19579), .A2(n9595), .ZN(n16394) );
  INV_X1 U13539 ( .A(n12793), .ZN(n12794) );
  INV_X1 U13540 ( .A(n16342), .ZN(n16652) );
  INV_X1 U13541 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16715) );
  CLKBUF_X1 U13542 ( .A(n14657), .Z(n14675) );
  NOR2_X1 U13543 ( .A1(n12587), .A2(n12586), .ZN(n16731) );
  OAI21_X1 U13544 ( .B1(n16765), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16743), 
        .ZN(n20128) );
  AND2_X1 U13545 ( .A1(n19822), .A2(n19818), .ZN(n19839) );
  INV_X1 U13546 ( .A(n19846), .ZN(n19869) );
  OAI21_X1 U13547 ( .B1(n19884), .B2(n19883), .A(n19882), .ZN(n19907) );
  NAND2_X1 U13548 ( .A1(n20472), .A2(n20461), .ZN(n19875) );
  INV_X1 U13549 ( .A(n19975), .ZN(n19915) );
  OAI21_X1 U13550 ( .B1(n16781), .B2(n19912), .A(n16768), .ZN(n19971) );
  NOR2_X1 U13551 ( .A1(n19980), .A2(n19979), .ZN(n20004) );
  OAI21_X1 U13552 ( .B1(n20016), .B2(n20252), .A(n20015), .ZN(n20035) );
  NAND2_X1 U13553 ( .A1(n20050), .A2(n20049), .ZN(n20074) );
  NAND2_X1 U13554 ( .A1(n20090), .A2(n20089), .ZN(n20113) );
  INV_X1 U13555 ( .A(n20123), .ZN(n20147) );
  NAND2_X1 U13556 ( .A1(n16798), .A2(n16797), .ZN(n20172) );
  NOR2_X1 U13557 ( .A1(n20214), .A2(n19875), .ZN(n20184) );
  AND2_X1 U13558 ( .A1(n20222), .A2(n20217), .ZN(n20240) );
  NAND2_X1 U13559 ( .A1(n19760), .A2(n19759), .ZN(n20327) );
  NAND2_X1 U13560 ( .A1(n19785), .A2(n19784), .ZN(n20345) );
  INV_X1 U13561 ( .A(n20293), .ZN(n20357) );
  INV_X1 U13562 ( .A(n17428), .ZN(n14187) );
  INV_X1 U13563 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20391) );
  INV_X1 U13564 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20370) );
  XNOR2_X1 U13565 ( .A(n17568), .B(n17004), .ZN(n17572) );
  NOR2_X1 U13566 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17647), .ZN(n17627) );
  NOR2_X1 U13567 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17666), .ZN(n17654) );
  NOR2_X1 U13568 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17716), .ZN(n17696) );
  AND3_X1 U13569 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n17749), .ZN(n17623) );
  NOR2_X1 U13570 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17815), .ZN(n17802) );
  NOR2_X1 U13571 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17865), .ZN(n17852) );
  INV_X1 U13572 ( .A(n17927), .ZN(n17884) );
  NAND2_X1 U13573 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n13469), .ZN(n18021) );
  AND2_X1 U13574 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n13537), .ZN(n13657) );
  AND2_X1 U13575 ( .A1(n18154), .A2(n18157), .ZN(n18150) );
  NOR2_X1 U13576 ( .A1(n18303), .A2(n18225), .ZN(n18224) );
  NOR2_X1 U13577 ( .A1(n18344), .A2(n18242), .ZN(n18240) );
  OR2_X1 U13578 ( .A1(n16877), .A2(n16876), .ZN(n17153) );
  NAND2_X2 U13579 ( .A1(n18297), .A2(n18296), .ZN(n18353) );
  OR2_X1 U13580 ( .A1(n18481), .A2(n17169), .ZN(n18359) );
  AND2_X1 U13581 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18685), .ZN(n18432) );
  NAND2_X1 U13582 ( .A1(n16998), .A2(n16997), .ZN(n18554) );
  AND2_X1 U13583 ( .A1(n18814), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17176) );
  AND2_X1 U13584 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18869), .ZN(
        n18831) );
  AND2_X1 U13585 ( .A1(n19404), .A2(n18944), .ZN(n18952) );
  AND2_X1 U13586 ( .A1(n13442), .A2(n13441), .ZN(n19426) );
  INV_X1 U13587 ( .A(n19330), .ZN(n19035) );
  INV_X1 U13588 ( .A(n19384), .ZN(n19057) );
  INV_X1 U13589 ( .A(n19063), .ZN(n19103) );
  INV_X1 U13590 ( .A(n21552), .ZN(n19141) );
  INV_X1 U13591 ( .A(n21550), .ZN(n19184) );
  INV_X1 U13592 ( .A(n19190), .ZN(n19231) );
  INV_X1 U13593 ( .A(n19238), .ZN(n19279) );
  INV_X1 U13594 ( .A(n19284), .ZN(n19326) );
  AND2_X1 U13595 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19336), .ZN(n19341) );
  NOR3_X1 U13596 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19468), .A3(n19450), 
        .ZN(n19553) );
  INV_X1 U13597 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n19452) );
  INV_X1 U13598 ( .A(n12527), .ZN(n16770) );
  INV_X1 U13599 ( .A(U212), .ZN(n17470) );
  AND2_X1 U13600 ( .A1(n12964), .A2(n12965), .ZN(n21382) );
  INV_X1 U13601 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21191) );
  NOR2_X1 U13602 ( .A1(n12106), .A2(n12105), .ZN(n12107) );
  AND2_X1 U13603 ( .A1(n20511), .A2(n14949), .ZN(n17357) );
  INV_X1 U13604 ( .A(n20532), .ZN(n20589) );
  NAND2_X1 U13605 ( .A1(n20599), .A2(n20763), .ZN(n20594) );
  INV_X1 U13606 ( .A(n12706), .ZN(n15112) );
  INV_X1 U13607 ( .A(n15320), .ZN(n15148) );
  AND2_X1 U13608 ( .A1(n13548), .A2(n13547), .ZN(n20744) );
  INV_X1 U13609 ( .A(n20600), .ZN(n20626) );
  NAND2_X1 U13610 ( .A1(n12980), .A2(n13294), .ZN(n20633) );
  NOR2_X1 U13611 ( .A1(n12714), .A2(n12713), .ZN(n12715) );
  NAND2_X1 U13612 ( .A1(n15344), .A2(n13465), .ZN(n20654) );
  NAND2_X1 U13613 ( .A1(n12738), .A2(n20696), .ZN(n12746) );
  INV_X1 U13614 ( .A(n20696), .ZN(n20668) );
  NAND2_X1 U13615 ( .A1(n12250), .A2(n12224), .ZN(n20666) );
  AND3_X1 U13616 ( .A1(n15516), .A2(n15515), .A3(n20685), .ZN(n20672) );
  OAI21_X1 U13617 ( .B1(n15541), .B2(n15540), .A(n20775), .ZN(n20707) );
  AND2_X1 U13618 ( .A1(n13309), .A2(n13306), .ZN(n15577) );
  NAND2_X1 U13619 ( .A1(n20834), .A2(n20992), .ZN(n20797) );
  NAND2_X1 U13620 ( .A1(n20834), .A2(n10452), .ZN(n20833) );
  INV_X1 U13621 ( .A(n20896), .ZN(n20865) );
  NAND2_X1 U13622 ( .A1(n20962), .A2(n20992), .ZN(n20925) );
  NAND2_X1 U13623 ( .A1(n20962), .A2(n21091), .ZN(n20983) );
  NAND2_X1 U13624 ( .A1(n21092), .A2(n20992), .ZN(n21045) );
  NAND2_X1 U13625 ( .A1(n21092), .A2(n10452), .ZN(n21085) );
  NAND2_X1 U13626 ( .A1(n21092), .A2(n21189), .ZN(n21115) );
  NAND2_X1 U13627 ( .A1(n21092), .A2(n21091), .ZN(n21154) );
  OR2_X1 U13628 ( .A1(n21156), .A2(n21155), .ZN(n21233) );
  NAND2_X1 U13629 ( .A1(n20714), .A2(n21091), .ZN(n21297) );
  INV_X1 U13630 ( .A(n14054), .ZN(n15580) );
  INV_X1 U13631 ( .A(n21363), .ZN(n21299) );
  INV_X1 U13632 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21312) );
  NAND3_X1 U13633 ( .A1(n12680), .A2(n12951), .A3(n14187), .ZN(n12941) );
  INV_X1 U13634 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20122) );
  NAND2_X1 U13635 ( .A1(n12692), .A2(n15933), .ZN(n12693) );
  NAND2_X1 U13636 ( .A1(n15816), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19625) );
  INV_X1 U13637 ( .A(n16608), .ZN(n16044) );
  INV_X1 U13638 ( .A(n13177), .ZN(n15999) );
  NAND2_X1 U13639 ( .A1(n13643), .A2(n13642), .ZN(n20472) );
  NAND2_X1 U13640 ( .A1(n12282), .A2(n16151), .ZN(n16144) );
  AOI21_X2 U13641 ( .B1(n13825), .B2(n12514), .A(n17428), .ZN(n16151) );
  AND2_X1 U13642 ( .A1(n13151), .A2(n13150), .ZN(n19655) );
  NAND2_X1 U13643 ( .A1(n14154), .A2(n14153), .ZN(n19658) );
  OAI21_X2 U13644 ( .B1(n14152), .B2(n19700), .A(n15582), .ZN(n19696) );
  INV_X1 U13645 ( .A(n13877), .ZN(n13805) );
  INV_X1 U13646 ( .A(n12847), .ZN(n12848) );
  NAND2_X1 U13647 ( .A1(n11201), .A2(n9596), .ZN(n16396) );
  INV_X1 U13648 ( .A(n16394), .ZN(n16422) );
  INV_X1 U13649 ( .A(n12829), .ZN(n12830) );
  INV_X1 U13650 ( .A(n19721), .ZN(n16710) );
  INV_X1 U13651 ( .A(n16733), .ZN(n17413) );
  INV_X1 U13652 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17345) );
  NAND2_X2 U13653 ( .A1(n19982), .A2(n20078), .ZN(n19843) );
  OR2_X1 U13654 ( .A1(n19844), .A2(n19875), .ZN(n19911) );
  OR2_X1 U13655 ( .A1(n20017), .A2(n20219), .ZN(n20008) );
  AND2_X1 U13656 ( .A1(n20013), .A2(n20012), .ZN(n20030) );
  OR2_X1 U13657 ( .A1(n20017), .A2(n20458), .ZN(n20072) );
  AND2_X1 U13658 ( .A1(n20084), .A2(n20083), .ZN(n20095) );
  INV_X1 U13659 ( .A(n20351), .ZN(n20289) );
  INV_X1 U13660 ( .A(n20333), .ZN(n20274) );
  INV_X1 U13661 ( .A(n20327), .ZN(n20272) );
  INV_X1 U13662 ( .A(n20189), .ZN(n20318) );
  INV_X1 U13663 ( .A(n20202), .ZN(n20348) );
  INV_X1 U13664 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16757) );
  INV_X1 U13665 ( .A(n20456), .ZN(n20368) );
  OR2_X1 U13666 ( .A1(n20370), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n20483) );
  INV_X1 U13667 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n17521) );
  INV_X1 U13668 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18441) );
  INV_X1 U13669 ( .A(n17914), .ZN(n17880) );
  OR2_X1 U13670 ( .A1(n16825), .A2(n16819), .ZN(n17927) );
  INV_X1 U13671 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18127) );
  INV_X1 U13672 ( .A(n18150), .ZN(n17233) );
  OR2_X1 U13673 ( .A1(n18251), .A2(n16838), .ZN(n18221) );
  NOR2_X1 U13674 ( .A1(n18348), .A2(n16856), .ZN(n16859) );
  AND2_X1 U13675 ( .A1(n13696), .A2(n10456), .ZN(n16962) );
  INV_X1 U13676 ( .A(n18249), .ZN(n18197) );
  INV_X1 U13677 ( .A(n18273), .ZN(n18292) );
  INV_X1 U13678 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n21512) );
  NAND2_X1 U13679 ( .A1(n18554), .A2(n17176), .ZN(n18481) );
  INV_X1 U13680 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18684) );
  INV_X1 U13681 ( .A(n18944), .ZN(n18899) );
  NAND2_X1 U13682 ( .A1(n18881), .A2(n17176), .ZN(n18797) );
  OR2_X1 U13683 ( .A1(n18944), .A2(n18953), .ZN(n18855) );
  OR2_X1 U13684 ( .A1(n19399), .A2(n18899), .ZN(n18906) );
  INV_X1 U13685 ( .A(n18952), .ZN(n18923) );
  INV_X1 U13686 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19395) );
  INV_X1 U13687 ( .A(n19164), .ZN(n19124) );
  INV_X1 U13688 ( .A(n19209), .ZN(n19145) );
  INV_X1 U13689 ( .A(n19254), .ZN(n19188) );
  INV_X1 U13690 ( .A(n19302), .ZN(n19235) );
  INV_X1 U13691 ( .A(n19378), .ZN(n19283) );
  INV_X1 U13692 ( .A(n17909), .ZN(n19443) );
  INV_X1 U13693 ( .A(n19536), .ZN(n19449) );
  INV_X1 U13694 ( .A(n19568), .ZN(n19531) );
  NOR2_X1 U13695 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12937), .ZN(n17497)
         );
  INV_X1 U13696 ( .A(n17475), .ZN(n17472) );
  OAI21_X1 U13697 ( .B1(n15081), .B2(n17350), .A(n12107), .ZN(P1_U2812) );
  OAI21_X1 U13698 ( .B1(n15173), .B2(n20666), .A(n12272), .ZN(P1_U3003) );
  OAI211_X1 U13699 ( .C1(n15596), .C2(n14693), .A(n12694), .B(n12693), .ZN(
        P2_U2824) );
  AND2_X4 U13700 ( .A1(n13809), .A2(n13810), .ZN(n14618) );
  AOI22_X1 U13701 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10481) );
  AND2_X4 U13702 ( .A1(n11045), .A2(n10868), .ZN(n14625) );
  AOI22_X1 U13703 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10480) );
  AOI22_X1 U13704 ( .A1(n14605), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9570), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U13705 ( .A1(n10560), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10478) );
  NAND2_X1 U13706 ( .A1(n10482), .A2(n10551), .ZN(n10490) );
  AOI22_X1 U13707 ( .A1(n9581), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13708 ( .A1(n10560), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U13709 ( .A1(n14560), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9569), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10483) );
  NAND2_X1 U13710 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10487) );
  AOI22_X1 U13711 ( .A1(n9581), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10494) );
  AOI22_X1 U13712 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10493) );
  AOI22_X1 U13713 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13714 ( .A1(n14605), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14628), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10491) );
  NAND4_X1 U13715 ( .A1(n10494), .A2(n10493), .A3(n10492), .A4(n10491), .ZN(
        n10495) );
  NAND2_X1 U13716 ( .A1(n10495), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10502) );
  AOI22_X1 U13717 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13718 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13719 ( .A1(n14605), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9570), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U13720 ( .A1(n10560), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10496) );
  NAND4_X1 U13721 ( .A1(n10499), .A2(n10498), .A3(n10497), .A4(n10496), .ZN(
        n10500) );
  NAND2_X1 U13722 ( .A1(n10500), .A2(n10551), .ZN(n10501) );
  AOI22_X1 U13723 ( .A1(n9581), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10505) );
  AOI22_X1 U13724 ( .A1(n14560), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9570), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10504) );
  AOI22_X1 U13725 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10503) );
  NAND4_X1 U13726 ( .A1(n10506), .A2(n10505), .A3(n10504), .A4(n10503), .ZN(
        n10507) );
  NAND2_X1 U13727 ( .A1(n10507), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10514) );
  AOI22_X1 U13728 ( .A1(n10691), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U13729 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U13730 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9569), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13731 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10508) );
  NAND4_X1 U13732 ( .A1(n10511), .A2(n10510), .A3(n10509), .A4(n10508), .ZN(
        n10512) );
  NAND2_X1 U13733 ( .A1(n10512), .A2(n10551), .ZN(n10513) );
  AOI22_X1 U13734 ( .A1(n10691), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U13735 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U13736 ( .A1(n14560), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14628), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U13737 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10515) );
  NAND4_X1 U13738 ( .A1(n10518), .A2(n10517), .A3(n10516), .A4(n10515), .ZN(
        n10519) );
  NAND2_X1 U13739 ( .A1(n10519), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10526) );
  AOI22_X1 U13740 ( .A1(n10691), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10523) );
  AOI22_X1 U13741 ( .A1(n14560), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9570), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10522) );
  AOI22_X1 U13742 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10521) );
  AOI22_X1 U13743 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10520) );
  NAND4_X1 U13744 ( .A1(n10523), .A2(n10522), .A3(n10521), .A4(n10520), .ZN(
        n10524) );
  NAND2_X1 U13745 ( .A1(n10524), .A2(n10551), .ZN(n10525) );
  NOR2_X1 U13746 ( .A1(n10527), .A2(n10551), .ZN(n10531) );
  AOI22_X1 U13747 ( .A1(n14605), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14628), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U13748 ( .A1(n10691), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10529) );
  AOI22_X1 U13749 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10528) );
  NAND4_X1 U13750 ( .A1(n10531), .A2(n10530), .A3(n10529), .A4(n10528), .ZN(
        n10538) );
  NOR2_X1 U13751 ( .A1(n10532), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10536) );
  AOI22_X1 U13752 ( .A1(n14605), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9569), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13753 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U13754 ( .A1(n10691), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10533) );
  NAND4_X1 U13755 ( .A1(n10536), .A2(n10535), .A3(n10534), .A4(n10533), .ZN(
        n10537) );
  AOI22_X1 U13756 ( .A1(n9581), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13757 ( .A1(n14605), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14628), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10540) );
  AOI22_X1 U13758 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10539) );
  NAND4_X1 U13759 ( .A1(n10542), .A2(n10541), .A3(n10540), .A4(n10539), .ZN(
        n10543) );
  NAND2_X1 U13760 ( .A1(n10543), .A2(n10551), .ZN(n10550) );
  AOI22_X1 U13761 ( .A1(n14605), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14628), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10545) );
  AOI22_X1 U13762 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10544) );
  NAND4_X1 U13763 ( .A1(n10547), .A2(n10546), .A3(n10545), .A4(n10544), .ZN(
        n10548) );
  NAND2_X1 U13764 ( .A1(n10548), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10549) );
  INV_X1 U13765 ( .A(n14122), .ZN(n10558) );
  AOI22_X1 U13766 ( .A1(n10691), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9570), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U13767 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U13768 ( .A1(n14560), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10552) );
  AOI22_X1 U13769 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10557) );
  AOI22_X1 U13770 ( .A1(n14560), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14628), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13771 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10555) );
  BUF_X1 U13772 ( .A(n10583), .Z(n12558) );
  AOI22_X1 U13773 ( .A1(n9581), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10563) );
  AOI22_X1 U13774 ( .A1(n10691), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9570), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10562) );
  AOI22_X1 U13775 ( .A1(n14596), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10561) );
  NAND4_X1 U13776 ( .A1(n10564), .A2(n10563), .A3(n10562), .A4(n10561), .ZN(
        n10565) );
  NAND2_X1 U13777 ( .A1(n10565), .A2(n10551), .ZN(n10572) );
  AOI22_X1 U13778 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13779 ( .A1(n10691), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14604), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13780 ( .A1(n14560), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14628), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U13781 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10566) );
  NAND4_X1 U13782 ( .A1(n10569), .A2(n10568), .A3(n10567), .A4(n10566), .ZN(
        n10570) );
  NAND2_X1 U13783 ( .A1(n10570), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10571) );
  NAND2_X2 U13784 ( .A1(n10572), .A2(n10571), .ZN(n12283) );
  INV_X2 U13785 ( .A(n12283), .ZN(n10592) );
  NAND2_X1 U13786 ( .A1(n9595), .A2(n10583), .ZN(n10574) );
  NAND3_X1 U13787 ( .A1(n10851), .A2(n9596), .A3(n10581), .ZN(n10577) );
  NAND2_X1 U13788 ( .A1(n10577), .A2(n10598), .ZN(n10578) );
  NAND2_X1 U13789 ( .A1(n10578), .A2(n10591), .ZN(n10579) );
  INV_X1 U13791 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14300) );
  AND2_X1 U13792 ( .A1(n12512), .A2(n10585), .ZN(n10586) );
  AND2_X1 U13793 ( .A1(n12512), .A2(n12286), .ZN(n12499) );
  INV_X1 U13794 ( .A(n12289), .ZN(n12282) );
  XNOR2_X1 U13795 ( .A(n10594), .B(n10593), .ZN(n12501) );
  INV_X1 U13796 ( .A(n10599), .ZN(n10600) );
  NAND2_X1 U13797 ( .A1(n10605), .A2(n10600), .ZN(n12553) );
  NOR2_X1 U13798 ( .A1(n12482), .A2(n10584), .ZN(n10602) );
  NOR2_X1 U13799 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14136) );
  INV_X1 U13800 ( .A(n14136), .ZN(n10603) );
  OAI22_X1 U13801 ( .A1(n10623), .A2(n10608), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10629), .ZN(n10610) );
  AOI22_X1 U13802 ( .A1(n13812), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n14136), .ZN(n10609) );
  NAND2_X1 U13803 ( .A1(n10610), .A2(n10609), .ZN(n10638) );
  INV_X1 U13804 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10612) );
  NAND2_X1 U13805 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10613) );
  INV_X1 U13806 ( .A(n10616), .ZN(n10617) );
  INV_X1 U13807 ( .A(n11068), .ZN(n11112) );
  NAND2_X1 U13808 ( .A1(n10629), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10621) );
  OAI211_X2 U13809 ( .C1(n11112), .C2(n19722), .A(n10622), .B(n10621), .ZN(
        n10627) );
  NAND2_X1 U13810 ( .A1(n10632), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10625) );
  NAND2_X1 U13811 ( .A1(n10625), .A2(n10624), .ZN(n10628) );
  INV_X1 U13812 ( .A(n10628), .ZN(n10626) );
  INV_X2 U13813 ( .A(n11068), .ZN(n11150) );
  AOI22_X1 U13814 ( .A1(n11113), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10631) );
  NAND2_X1 U13815 ( .A1(n11147), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10630) );
  NAND2_X1 U13816 ( .A1(n10632), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10634) );
  NAND2_X1 U13817 ( .A1(n14136), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10633) );
  NAND2_X1 U13818 ( .A1(n10634), .A2(n10633), .ZN(n10635) );
  INV_X1 U13819 ( .A(n10637), .ZN(n10640) );
  INV_X1 U13820 ( .A(n10638), .ZN(n10639) );
  INV_X1 U13821 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10647) );
  INV_X1 U13822 ( .A(n10644), .ZN(n10645) );
  OR2_X1 U13823 ( .A1(n10655), .A2(n10645), .ZN(n10667) );
  INV_X1 U13824 ( .A(n10667), .ZN(n10646) );
  INV_X1 U13825 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10650) );
  INV_X1 U13826 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10649) );
  NOR2_X1 U13827 ( .A1(n10652), .A2(n10651), .ZN(n10685) );
  OR2_X1 U13828 ( .A1(n10654), .A2(n10642), .ZN(n10656) );
  NAND2_X2 U13829 ( .A1(n10656), .A2(n10655), .ZN(n16732) );
  INV_X1 U13830 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10658) );
  INV_X1 U13831 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10661) );
  NOR2_X1 U13832 ( .A1(n10663), .A2(n10662), .ZN(n10684) );
  INV_X1 U13833 ( .A(n10664), .ZN(n10665) );
  NOR2_X1 U13834 ( .A1(n13754), .A2(n10665), .ZN(n10669) );
  NOR2_X1 U13835 ( .A1(n13754), .A2(n10667), .ZN(n10668) );
  INV_X1 U13836 ( .A(n10799), .ZN(n20014) );
  INV_X1 U13837 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10671) );
  NAND2_X1 U13838 ( .A1(n10669), .A2(n19727), .ZN(n19816) );
  INV_X1 U13839 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10670) );
  OAI22_X1 U13840 ( .A1(n10671), .A2(n19879), .B1(n19816), .B2(n10670), .ZN(
        n10672) );
  NOR2_X1 U13841 ( .A1(n10673), .A2(n10672), .ZN(n10683) );
  INV_X1 U13842 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13908) );
  INV_X1 U13843 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10675) );
  OAI22_X1 U13844 ( .A1(n13908), .A2(n19749), .B1(n20183), .B2(n10675), .ZN(
        n10681) );
  INV_X1 U13845 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10679) );
  NAND2_X1 U13846 ( .A1(n10677), .A2(n15909), .ZN(n20042) );
  INV_X1 U13847 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10678) );
  OAI22_X1 U13848 ( .A1(n10679), .A2(n19919), .B1(n20042), .B2(n10678), .ZN(
        n10680) );
  NOR2_X1 U13849 ( .A1(n10681), .A2(n10680), .ZN(n10682) );
  AOI22_X1 U13850 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n14479), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U13851 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n10818), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U13852 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U13853 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9584), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10687) );
  NAND4_X1 U13854 ( .A1(n10690), .A2(n10689), .A3(n10688), .A4(n10687), .ZN(
        n10697) );
  AND2_X2 U13855 ( .A1(n9572), .A2(n10551), .ZN(n10835) );
  AOI22_X1 U13856 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n10835), .B1(
        n14435), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10695) );
  AOI22_X1 U13857 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n9588), .B1(n9590), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U13858 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n9587), .B1(n9591), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U13859 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n14473), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10692) );
  NAND4_X1 U13860 ( .A1(n10695), .A2(n10694), .A3(n10693), .A4(n10692), .ZN(
        n10696) );
  NAND2_X1 U13861 ( .A1(n12319), .A2(n9596), .ZN(n10698) );
  AOI22_X1 U13862 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n14473), .B1(
        n9591), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U13863 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n9588), .B1(n9590), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U13864 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n10710), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U13865 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10823), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10700) );
  NAND3_X1 U13866 ( .A1(n10703), .A2(n10702), .A3(n10460), .ZN(n10709) );
  AOI22_X1 U13867 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10835), .B1(
        n14479), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10707) );
  AOI22_X1 U13868 ( .A1(n10805), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10706) );
  AOI22_X1 U13869 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10818), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10705) );
  AOI22_X1 U13870 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n9585), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10704) );
  NAND4_X1 U13871 ( .A1(n10707), .A2(n10706), .A3(n10705), .A4(n10704), .ZN(
        n10708) );
  AOI22_X1 U13872 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n14435), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10714) );
  AOI22_X1 U13873 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n9578), .B1(n9579), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U13874 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10806), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13875 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10818), .B1(
        n9585), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10711) );
  NAND4_X1 U13876 ( .A1(n10714), .A2(n10713), .A3(n10712), .A4(n10711), .ZN(
        n10720) );
  AOI22_X1 U13877 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10835), .B1(
        n14479), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10718) );
  AOI22_X1 U13878 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n9590), .B1(n9591), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13879 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n9588), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13880 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n9587), .B1(n9592), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10715) );
  NAND4_X1 U13881 ( .A1(n10718), .A2(n10717), .A3(n10716), .A4(n10715), .ZN(
        n10719) );
  AND2_X1 U13882 ( .A1(n11166), .A2(n11167), .ZN(n10843) );
  NAND2_X1 U13883 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10724) );
  NAND2_X1 U13884 ( .A1(n10699), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10723) );
  NAND2_X1 U13885 ( .A1(n14435), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10722) );
  NAND2_X1 U13886 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10721) );
  NAND2_X1 U13887 ( .A1(n14479), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10728) );
  NAND2_X1 U13888 ( .A1(n10835), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10727) );
  NAND2_X1 U13889 ( .A1(n9589), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10726) );
  NAND2_X1 U13890 ( .A1(n9591), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10725) );
  NAND2_X1 U13891 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10732) );
  NAND2_X1 U13892 ( .A1(n10818), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10731) );
  NAND2_X1 U13893 ( .A1(n9577), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10730) );
  NAND2_X1 U13894 ( .A1(n9585), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10729) );
  NAND2_X1 U13895 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10736) );
  NAND2_X1 U13896 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10735) );
  NAND2_X1 U13897 ( .A1(n10823), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10734) );
  NAND2_X1 U13898 ( .A1(n9592), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10733) );
  INV_X1 U13899 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10741) );
  INV_X1 U13900 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10740) );
  OAI22_X1 U13901 ( .A1(n10741), .A2(n20216), .B1(n20088), .B2(n10740), .ZN(
        n10744) );
  INV_X1 U13902 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10742) );
  NOR2_X1 U13903 ( .A1(n10744), .A2(n10743), .ZN(n10765) );
  INV_X1 U13904 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10746) );
  INV_X1 U13905 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10745) );
  OAI22_X1 U13906 ( .A1(n10746), .A2(n19749), .B1(n20042), .B2(n10745), .ZN(
        n10750) );
  INV_X1 U13907 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10748) );
  INV_X1 U13908 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10747) );
  OAI22_X1 U13909 ( .A1(n10748), .A2(n19919), .B1(n20183), .B2(n10747), .ZN(
        n10749) );
  NOR2_X1 U13910 ( .A1(n10750), .A2(n10749), .ZN(n10764) );
  INV_X1 U13911 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10751) );
  INV_X1 U13912 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10753) );
  INV_X1 U13913 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10752) );
  NOR2_X1 U13914 ( .A1(n10755), .A2(n10754), .ZN(n10763) );
  INV_X1 U13915 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10757) );
  INV_X1 U13916 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10756) );
  OAI22_X1 U13917 ( .A1(n10757), .A2(n19879), .B1(n19816), .B2(n10756), .ZN(
        n10761) );
  INV_X1 U13918 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10759) );
  INV_X1 U13919 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10758) );
  NAND4_X1 U13920 ( .A1(n10765), .A2(n10764), .A3(n10763), .A4(n10762), .ZN(
        n10778) );
  AOI22_X1 U13921 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n14435), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10770) );
  AOI22_X1 U13922 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n9578), .B1(n9579), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10769) );
  AOI22_X1 U13923 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10806), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10768) );
  AOI22_X1 U13924 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10818), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10767) );
  NAND4_X1 U13925 ( .A1(n10770), .A2(n10769), .A3(n10768), .A4(n10767), .ZN(
        n10776) );
  AOI22_X1 U13926 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10835), .B1(
        n14479), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13927 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n9589), .B1(n9591), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U13928 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n9588), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13929 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n9587), .B1(n9592), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10771) );
  NAND4_X1 U13930 ( .A1(n10774), .A2(n10773), .A3(n10772), .A4(n10771), .ZN(
        n10775) );
  INV_X1 U13931 ( .A(n10865), .ZN(n12323) );
  NAND2_X1 U13932 ( .A1(n12323), .A2(n9595), .ZN(n10777) );
  NAND2_X1 U13933 ( .A1(n10778), .A2(n10777), .ZN(n10842) );
  INV_X1 U13934 ( .A(n10842), .ZN(n10779) );
  NAND2_X1 U13935 ( .A1(n10779), .A2(n11190), .ZN(n10780) );
  INV_X1 U13936 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10782) );
  INV_X1 U13937 ( .A(n10783), .ZN(n10787) );
  INV_X1 U13938 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10784) );
  INV_X1 U13939 ( .A(n10785), .ZN(n10786) );
  INV_X1 U13940 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10788) );
  OR2_X1 U13941 ( .A1(n19977), .A2(n10788), .ZN(n10794) );
  INV_X1 U13942 ( .A(n20127), .ZN(n10789) );
  NAND2_X1 U13943 ( .A1(n10789), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10793) );
  INV_X1 U13944 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10790) );
  INV_X1 U13945 ( .A(n10791), .ZN(n10792) );
  INV_X1 U13946 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10797) );
  INV_X1 U13947 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10796) );
  OAI22_X1 U13948 ( .A1(n10797), .A2(n20183), .B1(n20042), .B2(n10796), .ZN(
        n10803) );
  INV_X1 U13949 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10801) );
  INV_X1 U13950 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10798) );
  OAI211_X1 U13951 ( .C1(n19919), .C2(n10801), .A(n15978), .B(n10800), .ZN(
        n10802) );
  AOI22_X1 U13952 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n14435), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U13953 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n9578), .B1(n9579), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U13954 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10806), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U13955 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10818), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10807) );
  NAND4_X1 U13956 ( .A1(n10810), .A2(n10809), .A3(n10808), .A4(n10807), .ZN(
        n10817) );
  AOI22_X1 U13957 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10835), .B1(
        n14479), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10815) );
  AOI22_X1 U13958 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n9590), .B1(n9591), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13959 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n9588), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U13960 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n9587), .B1(n9592), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10812) );
  NAND4_X1 U13961 ( .A1(n10815), .A2(n10814), .A3(n10813), .A4(n10812), .ZN(
        n10816) );
  AOI22_X1 U13962 ( .A1(n14479), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10835), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U13963 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U13964 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10766), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10820) );
  AOI22_X1 U13965 ( .A1(n10818), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9583), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10819) );
  NAND4_X1 U13966 ( .A1(n10822), .A2(n10821), .A3(n10820), .A4(n10819), .ZN(
        n10830) );
  AOI22_X1 U13967 ( .A1(n10710), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U13968 ( .A1(n14472), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U13969 ( .A1(n10823), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10811), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U13970 ( .A1(n14474), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9591), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10825) );
  NAND4_X1 U13971 ( .A1(n10828), .A2(n10827), .A3(n10826), .A4(n10825), .ZN(
        n10829) );
  NAND3_X1 U13972 ( .A1(n9596), .A2(n12291), .A3(n10870), .ZN(n11173) );
  AOI22_X1 U13973 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n14479), .B1(
        n14435), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10834) );
  AOI22_X1 U13974 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10833) );
  AOI22_X1 U13975 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n9577), .B1(n9585), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10832) );
  AOI22_X1 U13976 ( .A1(n10805), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10818), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10831) );
  NAND4_X1 U13977 ( .A1(n10834), .A2(n10833), .A3(n10832), .A4(n10831), .ZN(
        n10841) );
  AOI22_X1 U13978 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10835), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U13979 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n14473), .B1(
        n9589), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10837) );
  AOI22_X1 U13980 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n9592), .B1(
        n9591), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10836) );
  NAND4_X1 U13981 ( .A1(n10839), .A2(n10838), .A3(n10837), .A4(n10836), .ZN(
        n10840) );
  NAND2_X1 U13982 ( .A1(n11173), .A2(n12300), .ZN(n10844) );
  AND2_X1 U13983 ( .A1(n10844), .A2(n10843), .ZN(n10845) );
  NAND2_X1 U13984 ( .A1(n11050), .A2(n11036), .ZN(n10848) );
  NAND2_X1 U13985 ( .A1(n20176), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10847) );
  INV_X1 U13986 ( .A(n10854), .ZN(n10849) );
  INV_X1 U13987 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13644) );
  NOR2_X1 U13988 ( .A1(n11022), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10872) );
  NAND2_X1 U13989 ( .A1(n10872), .A2(n14281), .ZN(n10853) );
  NAND2_X1 U13990 ( .A1(n12291), .A2(n11022), .ZN(n10852) );
  NAND2_X1 U13991 ( .A1(n10866), .A2(n10876), .ZN(n10883) );
  NAND2_X1 U13992 ( .A1(n10855), .A2(n10854), .ZN(n10857) );
  NAND2_X1 U13993 ( .A1(n20480), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10856) );
  NAND2_X1 U13994 ( .A1(n10857), .A2(n10856), .ZN(n10859) );
  NAND2_X1 U13995 ( .A1(n10859), .A2(n10858), .ZN(n11034) );
  OR2_X1 U13996 ( .A1(n10859), .A2(n10858), .ZN(n10860) );
  AND2_X1 U13997 ( .A1(n11034), .A2(n10860), .ZN(n11035) );
  INV_X1 U13998 ( .A(n11035), .ZN(n10861) );
  OAI21_X1 U13999 ( .B1(n9683), .B2(n10597), .A(n10864), .ZN(n10881) );
  INV_X1 U14000 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n13776) );
  MUX2_X1 U14001 ( .A(n11167), .B(n13776), .S(n10851), .Z(n10887) );
  MUX2_X1 U14002 ( .A(n12319), .B(P2_EBX_REG_5__SCAN_IN), .S(n10851), .Z(
        n10891) );
  INV_X1 U14003 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13918) );
  MUX2_X1 U14004 ( .A(n10865), .B(n13918), .S(n10597), .Z(n10903) );
  XNOR2_X1 U14005 ( .A(n10898), .B(n10903), .ZN(n15876) );
  INV_X1 U14006 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16697) );
  INV_X1 U14007 ( .A(n10876), .ZN(n10867) );
  XNOR2_X1 U14008 ( .A(n10866), .B(n10867), .ZN(n15919) );
  NAND2_X1 U14009 ( .A1(n15919), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10878) );
  INV_X1 U14010 ( .A(n10878), .ZN(n10880) );
  AND2_X1 U14011 ( .A1(n10868), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10869) );
  NOR2_X1 U14012 ( .A1(n11036), .A2(n10869), .ZN(n12486) );
  INV_X1 U14013 ( .A(n12486), .ZN(n10871) );
  INV_X1 U14014 ( .A(n10870), .ZN(n12285) );
  MUX2_X1 U14015 ( .A(n10871), .B(n12285), .S(n10252), .Z(n10873) );
  AOI21_X1 U14016 ( .B1(n10873), .B2(n11022), .A(n10872), .ZN(n15932) );
  NAND2_X1 U14017 ( .A1(n15932), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14341) );
  NAND2_X1 U14018 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n10874) );
  NOR2_X1 U14019 ( .A1(n11022), .A2(n10874), .ZN(n10875) );
  NOR2_X1 U14020 ( .A1(n10876), .A2(n10875), .ZN(n14278) );
  INV_X1 U14021 ( .A(n14278), .ZN(n10877) );
  NOR2_X1 U14022 ( .A1(n14341), .A2(n10877), .ZN(n13138) );
  NAND2_X1 U14023 ( .A1(n14341), .A2(n10877), .ZN(n13139) );
  OAI21_X1 U14024 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13138), .A(
        n13139), .ZN(n14695) );
  OAI21_X1 U14025 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n15919), .A(
        n10878), .ZN(n14697) );
  NOR2_X1 U14026 ( .A1(n14695), .A2(n14697), .ZN(n10879) );
  NOR2_X1 U14027 ( .A1(n10880), .A2(n10879), .ZN(n14660) );
  INV_X1 U14028 ( .A(n10881), .ZN(n10882) );
  XNOR2_X1 U14029 ( .A(n10883), .B(n10882), .ZN(n15900) );
  NAND2_X1 U14030 ( .A1(n15900), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14659) );
  NAND2_X1 U14031 ( .A1(n14660), .A2(n14659), .ZN(n10885) );
  INV_X1 U14032 ( .A(n15900), .ZN(n10884) );
  NAND2_X1 U14033 ( .A1(n10884), .A2(n16715), .ZN(n14658) );
  NAND2_X1 U14034 ( .A1(n10885), .A2(n14658), .ZN(n16421) );
  OAI21_X1 U14035 ( .B1(n9665), .B2(n10887), .A(n10886), .ZN(n10888) );
  INV_X1 U14036 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19717) );
  XNOR2_X1 U14037 ( .A(n10888), .B(n19717), .ZN(n16420) );
  OR2_X1 U14038 ( .A1(n16421), .A2(n16420), .ZN(n10890) );
  INV_X1 U14039 ( .A(n10888), .ZN(n15888) );
  NAND2_X1 U14040 ( .A1(n15888), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10889) );
  NAND2_X1 U14041 ( .A1(n10890), .A2(n10889), .ZN(n16398) );
  NAND2_X1 U14042 ( .A1(n16398), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10893) );
  AND2_X1 U14043 ( .A1(n10886), .A2(n10891), .ZN(n10892) );
  OR2_X1 U14044 ( .A1(n10892), .A2(n10898), .ZN(n19603) );
  NAND2_X1 U14045 ( .A1(n10893), .A2(n19603), .ZN(n10896) );
  INV_X1 U14046 ( .A(n16398), .ZN(n10894) );
  INV_X1 U14047 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16717) );
  NAND2_X1 U14048 ( .A1(n10894), .A2(n16717), .ZN(n10895) );
  INV_X1 U14049 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n11076) );
  MUX2_X1 U14050 ( .A(n11076), .B(n11025), .S(n11022), .Z(n10904) );
  INV_X1 U14051 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n14257) );
  NOR2_X1 U14052 ( .A1(n11022), .A2(n14257), .ZN(n10900) );
  NAND2_X1 U14053 ( .A1(n10899), .A2(n10900), .ZN(n10901) );
  NAND2_X1 U14054 ( .A1(n10909), .A2(n10901), .ZN(n14261) );
  NAND2_X1 U14055 ( .A1(n11025), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10902) );
  OR2_X1 U14056 ( .A1(n14261), .A2(n10902), .ZN(n16362) );
  NAND2_X1 U14057 ( .A1(n10898), .A2(n10903), .ZN(n10906) );
  INV_X1 U14058 ( .A(n10904), .ZN(n10905) );
  NAND2_X1 U14059 ( .A1(n10906), .A2(n10905), .ZN(n10907) );
  NAND2_X1 U14060 ( .A1(n10907), .A2(n10899), .ZN(n15858) );
  INV_X1 U14061 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16687) );
  OR2_X1 U14062 ( .A1(n15858), .A2(n16687), .ZN(n16381) );
  AND2_X1 U14063 ( .A1(n16362), .A2(n16381), .ZN(n16334) );
  INV_X1 U14064 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n11085) );
  INV_X1 U14065 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13970) );
  NAND2_X1 U14066 ( .A1(n10910), .A2(n13970), .ZN(n10922) );
  NAND2_X1 U14067 ( .A1(n10597), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10911) );
  NOR2_X1 U14068 ( .A1(n10910), .A2(n10911), .ZN(n10912) );
  OR2_X1 U14069 ( .A1(n10919), .A2(n10912), .ZN(n14289) );
  OR2_X1 U14070 ( .A1(n14289), .A2(n11190), .ZN(n10913) );
  INV_X1 U14071 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16638) );
  NAND2_X1 U14072 ( .A1(n10913), .A2(n16638), .ZN(n16318) );
  NAND2_X1 U14073 ( .A1(n10597), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10914) );
  OAI21_X1 U14074 ( .B1(n9672), .B2(n10914), .A(n11030), .ZN(n10915) );
  OR2_X1 U14075 ( .A1(n10915), .A2(n10910), .ZN(n10924) );
  INV_X1 U14076 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16648) );
  OAI21_X1 U14077 ( .B1(n10924), .B2(n11190), .A(n16648), .ZN(n16339) );
  INV_X1 U14078 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16677) );
  OAI21_X1 U14079 ( .B1(n14261), .B2(n11190), .A(n16677), .ZN(n16363) );
  NAND2_X1 U14080 ( .A1(n15858), .A2(n16687), .ZN(n16380) );
  AND2_X1 U14081 ( .A1(n16363), .A2(n16380), .ZN(n16335) );
  NAND2_X1 U14082 ( .A1(n10597), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10916) );
  XNOR2_X1 U14083 ( .A(n10909), .B(n10916), .ZN(n15849) );
  NAND2_X1 U14084 ( .A1(n15849), .A2(n11025), .ZN(n10917) );
  INV_X1 U14085 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16636) );
  NAND2_X1 U14086 ( .A1(n10917), .A2(n16636), .ZN(n16349) );
  AND3_X1 U14087 ( .A1(n16339), .A2(n16335), .A3(n16349), .ZN(n16319) );
  AND2_X1 U14088 ( .A1(n16318), .A2(n16319), .ZN(n10918) );
  NAND2_X1 U14089 ( .A1(n10597), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10920) );
  INV_X1 U14090 ( .A(n10920), .ZN(n10921) );
  NAND2_X1 U14091 ( .A1(n10922), .A2(n10921), .ZN(n10923) );
  NAND2_X1 U14092 ( .A1(n10929), .A2(n10923), .ZN(n14267) );
  INV_X1 U14093 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16604) );
  INV_X1 U14094 ( .A(n10924), .ZN(n15836) );
  AND2_X1 U14095 ( .A1(n11025), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10925) );
  NAND2_X1 U14096 ( .A1(n15836), .A2(n10925), .ZN(n16338) );
  AND2_X1 U14097 ( .A1(n11025), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10926) );
  NAND2_X1 U14098 ( .A1(n15849), .A2(n10926), .ZN(n16348) );
  AND2_X1 U14099 ( .A1(n16338), .A2(n16348), .ZN(n16321) );
  NAND2_X1 U14100 ( .A1(n11025), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10927) );
  OR2_X1 U14101 ( .A1(n14289), .A2(n10927), .ZN(n16317) );
  AND2_X1 U14102 ( .A1(n16321), .A2(n16317), .ZN(n12601) );
  AND2_X1 U14103 ( .A1(n16307), .A2(n12601), .ZN(n10928) );
  NAND2_X1 U14104 ( .A1(n10597), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10931) );
  INV_X1 U14105 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11093) );
  NOR2_X1 U14106 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(P2_EBX_REG_14__SCAN_IN), 
        .ZN(n10930) );
  INV_X1 U14107 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n10938) );
  NAND2_X1 U14108 ( .A1(n10942), .A2(n11030), .ZN(n10947) );
  NAND2_X1 U14109 ( .A1(n10597), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10946) );
  MUX2_X1 U14110 ( .A(n10597), .B(n10931), .S(n10935), .Z(n10932) );
  NAND2_X1 U14111 ( .A1(n10932), .A2(n10934), .ZN(n15754) );
  OR2_X1 U14112 ( .A1(n15754), .A2(n11190), .ZN(n10933) );
  INV_X1 U14113 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16543) );
  NAND2_X1 U14114 ( .A1(n10933), .A2(n16543), .ZN(n12611) );
  NOR2_X1 U14115 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(P2_EBX_REG_18__SCAN_IN), 
        .ZN(n10936) );
  NAND2_X1 U14116 ( .A1(n15735), .A2(n11025), .ZN(n10974) );
  INV_X1 U14117 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16251) );
  NAND2_X1 U14118 ( .A1(n10597), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10937) );
  XNOR2_X1 U14119 ( .A(n10961), .B(n10937), .ZN(n15726) );
  NAND2_X1 U14120 ( .A1(n15726), .A2(n11025), .ZN(n10978) );
  INV_X1 U14121 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21522) );
  AND2_X1 U14122 ( .A1(n10978), .A2(n21522), .ZN(n16231) );
  NOR2_X1 U14123 ( .A1(n11022), .A2(n10938), .ZN(n10940) );
  INV_X1 U14124 ( .A(n11030), .ZN(n10939) );
  AOI21_X1 U14125 ( .B1(n9651), .B2(n10940), .A(n10939), .ZN(n10941) );
  NAND2_X1 U14126 ( .A1(n10942), .A2(n10941), .ZN(n15781) );
  NOR2_X1 U14127 ( .A1(n15781), .A2(n11190), .ZN(n10943) );
  NAND2_X1 U14128 ( .A1(n10943), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12607) );
  INV_X1 U14129 ( .A(n10943), .ZN(n10944) );
  INV_X1 U14130 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16567) );
  NAND2_X1 U14131 ( .A1(n10944), .A2(n16567), .ZN(n10945) );
  AND2_X1 U14132 ( .A1(n12607), .A2(n10945), .ZN(n12605) );
  OR2_X1 U14133 ( .A1(n10947), .A2(n10946), .ZN(n10948) );
  AND2_X1 U14134 ( .A1(n10935), .A2(n10948), .ZN(n15766) );
  NAND2_X1 U14135 ( .A1(n15766), .A2(n11025), .ZN(n10950) );
  INV_X1 U14136 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10949) );
  NAND2_X1 U14137 ( .A1(n10950), .A2(n10949), .ZN(n12609) );
  NAND2_X1 U14138 ( .A1(n10597), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10952) );
  MUX2_X1 U14139 ( .A(n10597), .B(n10952), .S(n10951), .Z(n10953) );
  OR2_X1 U14140 ( .A1(n10951), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10956) );
  NAND2_X1 U14141 ( .A1(n10953), .A2(n10956), .ZN(n15807) );
  OR2_X1 U14142 ( .A1(n15807), .A2(n11190), .ZN(n10954) );
  INV_X1 U14143 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16590) );
  NAND2_X1 U14144 ( .A1(n10954), .A2(n16590), .ZN(n16289) );
  INV_X1 U14145 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11097) );
  NOR2_X1 U14146 ( .A1(n11022), .A2(n11097), .ZN(n10955) );
  NAND2_X1 U14147 ( .A1(n10956), .A2(n10955), .ZN(n10957) );
  AND2_X1 U14148 ( .A1(n10957), .A2(n9651), .ZN(n15786) );
  NAND2_X1 U14149 ( .A1(n15786), .A2(n11025), .ZN(n10958) );
  INV_X1 U14150 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12792) );
  NAND2_X1 U14151 ( .A1(n10958), .A2(n12792), .ZN(n16278) );
  XNOR2_X1 U14152 ( .A(n10929), .B(n10465), .ZN(n15815) );
  NAND2_X1 U14153 ( .A1(n15815), .A2(n11025), .ZN(n10971) );
  INV_X1 U14154 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16602) );
  NAND2_X1 U14155 ( .A1(n10971), .A2(n16602), .ZN(n16300) );
  NAND2_X1 U14156 ( .A1(n10959), .A2(n16604), .ZN(n16306) );
  AND4_X1 U14157 ( .A1(n16289), .A2(n16278), .A3(n16300), .A4(n16306), .ZN(
        n10960) );
  AND3_X1 U14158 ( .A1(n12605), .A2(n12609), .A3(n10960), .ZN(n10967) );
  INV_X1 U14159 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n16001) );
  NAND2_X1 U14160 ( .A1(n10963), .A2(n16001), .ZN(n10984) );
  NAND2_X1 U14161 ( .A1(n10984), .A2(n11030), .ZN(n10982) );
  NAND2_X1 U14162 ( .A1(n10597), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10962) );
  NOR2_X1 U14163 ( .A1(n10963), .A2(n10962), .ZN(n10964) );
  INV_X1 U14164 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10965) );
  NAND2_X1 U14165 ( .A1(n11025), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10968) );
  OR2_X1 U14166 ( .A1(n15709), .A2(n10968), .ZN(n12813) );
  AND2_X1 U14167 ( .A1(n11025), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10969) );
  NAND2_X1 U14168 ( .A1(n15766), .A2(n10969), .ZN(n12608) );
  AND2_X1 U14169 ( .A1(n11025), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10970) );
  NAND2_X1 U14170 ( .A1(n15786), .A2(n10970), .ZN(n16277) );
  AND2_X1 U14171 ( .A1(n16277), .A2(n16301), .ZN(n10973) );
  NAND2_X1 U14172 ( .A1(n11025), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10972) );
  AND4_X1 U14173 ( .A1(n12608), .A2(n10973), .A3(n12607), .A4(n16288), .ZN(
        n10977) );
  INV_X1 U14174 ( .A(n10974), .ZN(n10975) );
  NAND2_X1 U14175 ( .A1(n10975), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16243) );
  NAND2_X1 U14176 ( .A1(n11025), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10976) );
  INV_X1 U14177 ( .A(n10978), .ZN(n10979) );
  INV_X1 U14178 ( .A(n16232), .ZN(n10980) );
  NAND2_X1 U14179 ( .A1(n10597), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10983) );
  NAND2_X1 U14180 ( .A1(n10984), .A2(n10241), .ZN(n10985) );
  NAND2_X1 U14181 ( .A1(n10989), .A2(n10985), .ZN(n15697) );
  OR2_X1 U14182 ( .A1(n15697), .A2(n11190), .ZN(n10987) );
  INV_X1 U14183 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16508) );
  NAND2_X1 U14184 ( .A1(n10987), .A2(n16508), .ZN(n16218) );
  INV_X1 U14185 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10986) );
  XNOR2_X1 U14186 ( .A(n10989), .B(n10461), .ZN(n15681) );
  INV_X1 U14187 ( .A(n16200), .ZN(n16201) );
  INV_X1 U14188 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16495) );
  AND2_X1 U14189 ( .A1(n16201), .A2(n16495), .ZN(n10993) );
  NAND2_X1 U14190 ( .A1(n16219), .A2(n16495), .ZN(n10988) );
  NAND2_X1 U14191 ( .A1(n10991), .A2(n11030), .ZN(n10992) );
  NAND2_X1 U14192 ( .A1(n10994), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16203) );
  INV_X1 U14193 ( .A(n10994), .ZN(n10995) );
  INV_X1 U14194 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16479) );
  NAND2_X1 U14195 ( .A1(n10995), .A2(n16479), .ZN(n16202) );
  INV_X1 U14196 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15652) );
  NAND2_X1 U14197 ( .A1(n10597), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10997) );
  AOI21_X1 U14198 ( .B1(n15653), .B2(n15652), .A(n10997), .ZN(n10998) );
  NOR2_X1 U14199 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(P2_EBX_REG_25__SCAN_IN), 
        .ZN(n10999) );
  NAND2_X1 U14200 ( .A1(n15653), .A2(n10999), .ZN(n11010) );
  NAND2_X1 U14201 ( .A1(n11010), .A2(n11030), .ZN(n11007) );
  INV_X1 U14202 ( .A(n11007), .ZN(n11000) );
  INV_X1 U14203 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16186) );
  OAI21_X1 U14204 ( .B1(n15639), .B2(n11190), .A(n16186), .ZN(n11004) );
  INV_X1 U14205 ( .A(n15639), .ZN(n11003) );
  NAND2_X1 U14206 ( .A1(n11004), .A2(n11017), .ZN(n16179) );
  INV_X1 U14207 ( .A(n16179), .ZN(n11005) );
  NAND2_X1 U14208 ( .A1(n10597), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11008) );
  INV_X1 U14209 ( .A(n11008), .ZN(n11009) );
  NAND2_X1 U14210 ( .A1(n11010), .A2(n11009), .ZN(n11011) );
  NAND2_X1 U14211 ( .A1(n11014), .A2(n11011), .ZN(n15625) );
  INV_X1 U14212 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16173) );
  NAND2_X1 U14213 ( .A1(n11030), .A2(n11025), .ZN(n11016) );
  INV_X1 U14214 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16468) );
  AND2_X1 U14215 ( .A1(n11016), .A2(n16468), .ZN(n16189) );
  INV_X1 U14216 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11142) );
  NOR2_X1 U14217 ( .A1(n11022), .A2(n11142), .ZN(n11015) );
  INV_X1 U14218 ( .A(n11020), .ZN(n11013) );
  AOI21_X1 U14219 ( .B1(n11015), .B2(n11014), .A(n11013), .ZN(n15612) );
  NAND2_X1 U14220 ( .A1(n15612), .A2(n11025), .ZN(n14351) );
  OR2_X1 U14221 ( .A1(n11016), .A2(n16468), .ZN(n16190) );
  NAND2_X1 U14222 ( .A1(n11017), .A2(n16190), .ZN(n14348) );
  INV_X1 U14223 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n11018) );
  NOR2_X1 U14224 ( .A1(n11022), .A2(n11018), .ZN(n11019) );
  INV_X1 U14225 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n11021) );
  NOR2_X1 U14226 ( .A1(n11022), .A2(n11021), .ZN(n11023) );
  XNOR2_X1 U14227 ( .A(n11029), .B(n11023), .ZN(n14686) );
  INV_X1 U14228 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12766) );
  OAI21_X1 U14229 ( .B1(n14686), .B2(n11190), .A(n12766), .ZN(n12748) );
  INV_X1 U14230 ( .A(n15604), .ZN(n11024) );
  INV_X1 U14231 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21478) );
  NAND2_X1 U14232 ( .A1(n11025), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11026) );
  NOR2_X1 U14233 ( .A1(n14686), .A2(n11026), .ZN(n12749) );
  OAI21_X1 U14234 ( .B1(n11029), .B2(P2_EBX_REG_30__SCAN_IN), .A(n10597), .ZN(
        n11031) );
  NAND2_X1 U14235 ( .A1(n11031), .A2(n11030), .ZN(n12688) );
  NOR2_X1 U14236 ( .A1(n12688), .A2(n11190), .ZN(n11032) );
  NAND2_X1 U14237 ( .A1(n20471), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11033) );
  NAND2_X1 U14238 ( .A1(n11034), .A2(n11033), .ZN(n11040) );
  NAND2_X1 U14239 ( .A1(n17343), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11041) );
  OR2_X1 U14240 ( .A1(n11040), .A2(n11041), .ZN(n11051) );
  INV_X1 U14241 ( .A(n11036), .ZN(n11037) );
  XNOR2_X1 U14242 ( .A(n11050), .B(n11037), .ZN(n12485) );
  AND2_X1 U14243 ( .A1(n12484), .A2(n12485), .ZN(n11038) );
  NAND2_X1 U14244 ( .A1(n12492), .A2(n11038), .ZN(n11043) );
  NOR2_X1 U14245 ( .A1(n17343), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11039) );
  NAND3_X1 U14246 ( .A1(n12492), .A2(n12484), .A3(n12486), .ZN(n11044) );
  NAND2_X1 U14247 ( .A1(n12951), .A2(n11044), .ZN(n11048) );
  INV_X1 U14248 ( .A(n9584), .ZN(n11047) );
  AOI21_X1 U14249 ( .B1(n11046), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14121) );
  AOI21_X1 U14250 ( .B1(n11047), .B2(n14121), .A(P2_FLUSH_REG_SCAN_IN), .ZN(
        n16738) );
  MUX2_X1 U14251 ( .A(n11048), .B(n16738), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n17415) );
  NOR2_X1 U14252 ( .A1(n17415), .A2(n11049), .ZN(n11055) );
  AND2_X1 U14253 ( .A1(n12486), .A2(n11050), .ZN(n12489) );
  OAI211_X1 U14254 ( .C1(n12489), .C2(n11052), .A(n9683), .B(n11051), .ZN(
        n11053) );
  NAND2_X1 U14255 ( .A1(n11053), .A2(n12495), .ZN(n12955) );
  OR2_X1 U14256 ( .A1(n11049), .A2(n12558), .ZN(n14119) );
  NOR2_X1 U14257 ( .A1(n12955), .A2(n14119), .ZN(n11054) );
  MUX2_X1 U14258 ( .A(n11055), .B(n11054), .S(n9596), .Z(n12533) );
  NOR2_X1 U14259 ( .A1(n12558), .A2(n17428), .ZN(n11056) );
  AOI22_X1 U14260 ( .A1(n11113), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11058) );
  NAND2_X1 U14261 ( .A1(n11147), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11057) );
  OAI211_X1 U14262 ( .C1(n11150), .C2(n16604), .A(n11058), .B(n11057), .ZN(
        n14205) );
  AOI22_X1 U14263 ( .A1(n11113), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11060) );
  NAND2_X1 U14264 ( .A1(n11147), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11059) );
  OAI211_X1 U14265 ( .C1(n11150), .C2(n16638), .A(n11060), .B(n11059), .ZN(
        n13961) );
  AND2_X1 U14266 ( .A1(n14205), .A2(n13961), .ZN(n11087) );
  AOI22_X1 U14267 ( .A1(n11113), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11063) );
  NAND2_X1 U14268 ( .A1(n11147), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11062) );
  OAI211_X1 U14269 ( .C1(n11150), .C2(n19717), .A(n11063), .B(n11062), .ZN(
        n13774) );
  AND2_X1 U14270 ( .A1(n13774), .A2(n13772), .ZN(n11064) );
  NAND2_X1 U14271 ( .A1(n11061), .A2(n11064), .ZN(n13773) );
  INV_X1 U14272 ( .A(n13773), .ZN(n11073) );
  NAND2_X1 U14273 ( .A1(n11113), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11066) );
  NAND2_X1 U14274 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11065) );
  OAI211_X1 U14275 ( .C1(n11152), .C2(n13918), .A(n11066), .B(n11065), .ZN(
        n11067) );
  AOI21_X1 U14276 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n11067), .ZN(n13915) );
  INV_X1 U14277 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n11071) );
  NAND2_X1 U14278 ( .A1(n11113), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11070) );
  NAND2_X1 U14279 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11069) );
  OAI211_X1 U14280 ( .C1(n11152), .C2(n11071), .A(n11070), .B(n11069), .ZN(
        n11072) );
  AOI21_X1 U14281 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11072), .ZN(n13783) );
  NAND2_X1 U14282 ( .A1(n11073), .A2(n9600), .ZN(n13913) );
  NAND2_X1 U14283 ( .A1(n11113), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11075) );
  NAND2_X1 U14284 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11074) );
  OAI211_X1 U14285 ( .C1(n11152), .C2(n11076), .A(n11075), .B(n11074), .ZN(
        n11077) );
  AOI21_X1 U14286 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n11077), .ZN(n13941) );
  AOI22_X1 U14287 ( .A1(n11113), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11079) );
  NAND2_X1 U14288 ( .A1(n11147), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11078) );
  OAI211_X1 U14289 ( .C1(n11150), .C2(n16677), .A(n11079), .B(n11078), .ZN(
        n14235) );
  NAND2_X1 U14290 ( .A1(n11113), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11081) );
  NAND2_X1 U14291 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11080) );
  OAI211_X1 U14292 ( .C1(n11152), .C2(n10247), .A(n11081), .B(n11080), .ZN(
        n11082) );
  AOI21_X1 U14293 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11082), .ZN(n14082) );
  NAND2_X1 U14294 ( .A1(n11113), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11084) );
  NAND2_X1 U14295 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11083) );
  OAI211_X1 U14296 ( .C1(n11152), .C2(n11085), .A(n11084), .B(n11083), .ZN(
        n11086) );
  AOI21_X1 U14297 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n11086), .ZN(n13894) );
  INV_X1 U14298 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n15803) );
  NAND2_X1 U14299 ( .A1(n11113), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11089) );
  NAND2_X1 U14300 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11088) );
  OAI211_X1 U14301 ( .C1(n11152), .C2(n15803), .A(n11089), .B(n11088), .ZN(
        n11090) );
  AOI21_X1 U14302 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11090), .ZN(n15797) );
  NAND2_X1 U14303 ( .A1(n11113), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11092) );
  NAND2_X1 U14304 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11091) );
  OAI211_X1 U14305 ( .C1(n11152), .C2(n11093), .A(n11092), .B(n11091), .ZN(
        n11094) );
  AOI21_X1 U14306 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11094), .ZN(n15811) );
  NAND2_X1 U14307 ( .A1(n11113), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11096) );
  NAND2_X1 U14308 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11095) );
  OAI211_X1 U14309 ( .C1(n11152), .C2(n11097), .A(n11096), .B(n11095), .ZN(
        n11098) );
  AOI21_X1 U14310 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11098), .ZN(n15784) );
  AOI22_X1 U14311 ( .A1(n11113), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11101) );
  NAND2_X1 U14312 ( .A1(n11147), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11100) );
  OAI211_X1 U14313 ( .C1(n11150), .C2(n16567), .A(n11101), .B(n11100), .ZN(
        n15770) );
  INV_X1 U14314 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n15763) );
  NAND2_X1 U14315 ( .A1(n11113), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11103) );
  NAND2_X1 U14316 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11102) );
  OAI211_X1 U14317 ( .C1(n11152), .C2(n15763), .A(n11103), .B(n11102), .ZN(
        n11104) );
  AOI21_X1 U14318 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11104), .ZN(n12798) );
  NAND2_X1 U14319 ( .A1(n11113), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11108) );
  NAND2_X1 U14320 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11107) );
  OAI211_X1 U14321 ( .C1(n11152), .C2(n10037), .A(n11108), .B(n11107), .ZN(
        n11109) );
  AOI21_X1 U14322 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n11109), .ZN(n12592) );
  AOI22_X1 U14323 ( .A1(n11113), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11111) );
  NAND2_X1 U14324 ( .A1(n11147), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11110) );
  OAI211_X1 U14325 ( .C1(n11112), .C2(n16251), .A(n11111), .B(n11110), .ZN(
        n15729) );
  NAND2_X1 U14326 ( .A1(n11113), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11115) );
  NAND2_X1 U14327 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11114) );
  OAI211_X1 U14328 ( .C1(n11152), .C2(n16001), .A(n11115), .B(n11114), .ZN(
        n11116) );
  AOI21_X1 U14329 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11116), .ZN(n12819) );
  INV_X1 U14330 ( .A(n12819), .ZN(n11119) );
  AOI22_X1 U14331 ( .A1(n11113), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11118) );
  NAND2_X1 U14332 ( .A1(n11147), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11117) );
  OAI211_X1 U14333 ( .C1(n11150), .C2(n21522), .A(n11118), .B(n11117), .ZN(
        n15714) );
  INV_X1 U14334 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n11123) );
  NAND2_X1 U14335 ( .A1(n11113), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11122) );
  NAND2_X1 U14336 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11121) );
  OAI211_X1 U14337 ( .C1(n11152), .C2(n11123), .A(n11122), .B(n11121), .ZN(
        n11124) );
  AOI21_X1 U14338 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11124), .ZN(n15687) );
  AOI22_X1 U14339 ( .A1(n11113), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11126) );
  NAND2_X1 U14340 ( .A1(n11147), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11125) );
  OAI211_X1 U14341 ( .C1(n11150), .C2(n16495), .A(n11126), .B(n11125), .ZN(
        n15676) );
  INV_X1 U14342 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n11129) );
  NAND2_X1 U14343 ( .A1(n11113), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11128) );
  NAND2_X1 U14344 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11127) );
  OAI211_X1 U14345 ( .C1(n11152), .C2(n11129), .A(n11128), .B(n11127), .ZN(
        n11130) );
  AOI21_X1 U14346 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11130), .ZN(n15661) );
  NAND2_X1 U14347 ( .A1(n11113), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11132) );
  NAND2_X1 U14348 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11131) );
  OAI211_X1 U14349 ( .C1(n11152), .C2(n15652), .A(n11132), .B(n11131), .ZN(
        n11133) );
  AOI21_X1 U14350 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n11133), .ZN(n15644) );
  INV_X1 U14351 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U14352 ( .A1(n11113), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11135) );
  NAND2_X1 U14353 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11134) );
  OAI211_X1 U14354 ( .C1(n11152), .C2(n11136), .A(n11135), .B(n11134), .ZN(
        n11137) );
  AOI21_X1 U14355 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11137), .ZN(n15629) );
  AOI22_X1 U14356 ( .A1(n11113), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11139) );
  NAND2_X1 U14357 ( .A1(n11147), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11138) );
  OAI211_X1 U14358 ( .C1(n11150), .C2(n16173), .A(n11139), .B(n11138), .ZN(
        n15614) );
  NAND2_X1 U14359 ( .A1(n11113), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11141) );
  NAND2_X1 U14360 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11140) );
  OAI211_X1 U14361 ( .C1(n11152), .C2(n11142), .A(n11141), .B(n11140), .ZN(
        n11143) );
  AOI21_X1 U14362 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11143), .ZN(n14360) );
  INV_X1 U14363 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20441) );
  INV_X1 U14364 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16162) );
  OAI22_X1 U14365 ( .A1(n10620), .A2(n20441), .B1(n16757), .B2(n16162), .ZN(
        n11146) );
  NOR2_X1 U14366 ( .A1(n11150), .A2(n21478), .ZN(n11145) );
  AOI211_X1 U14367 ( .C1(P2_EBX_REG_29__SCAN_IN), .C2(n11147), .A(n11146), .B(
        n11145), .ZN(n15593) );
  AOI22_X1 U14368 ( .A1(n11113), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11149) );
  NAND2_X1 U14369 ( .A1(n11147), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11148) );
  OAI211_X1 U14370 ( .C1(n11150), .C2(n12766), .A(n11149), .B(n11148), .ZN(
        n12757) );
  INV_X1 U14371 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14252) );
  AOI22_X1 U14372 ( .A1(n11113), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11151) );
  OAI21_X1 U14373 ( .B1(n11152), .B2(n14252), .A(n11151), .ZN(n11153) );
  AOI21_X1 U14374 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n11153), .ZN(n11154) );
  NOR2_X1 U14375 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20462) );
  OR2_X1 U14376 ( .A1(n20462), .A2(n20463), .ZN(n16749) );
  NAND2_X1 U14377 ( .A1(n16749), .A2(n15584), .ZN(n11155) );
  AND2_X1 U14378 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n16747) );
  NOR2_X1 U14379 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12676) );
  AND2_X2 U14380 ( .A1(n20462), .A2(n12676), .ZN(n19604) );
  INV_X1 U14381 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20448) );
  NOR2_X1 U14382 ( .A1(n19705), .A2(n20448), .ZN(n12579) );
  AOI21_X1 U14383 ( .B1(n16354), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n12579), .ZN(n11164) );
  NAND2_X1 U14384 ( .A1(n12641), .A2(n11158), .ZN(n12595) );
  INV_X1 U14385 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16222) );
  INV_X1 U14386 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16180) );
  INV_X1 U14387 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16170) );
  AND2_X1 U14388 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11159) );
  NAND2_X1 U14389 ( .A1(n12669), .A2(n11159), .ZN(n12673) );
  INV_X1 U14390 ( .A(n12673), .ZN(n11160) );
  NAND2_X1 U14391 ( .A1(n11160), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11161) );
  AND2_X1 U14392 ( .A1(n20122), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12677) );
  INV_X1 U14393 ( .A(n12677), .ZN(n11162) );
  NAND2_X1 U14394 ( .A1(n15584), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13632) );
  NAND2_X1 U14395 ( .A1(n11162), .A2(n13632), .ZN(n14342) );
  NAND2_X1 U14396 ( .A1(n12617), .A2(n16425), .ZN(n11163) );
  OAI211_X1 U14397 ( .C1(n15946), .C2(n16429), .A(n11164), .B(n11163), .ZN(
        n11165) );
  AOI21_X1 U14398 ( .B1(n12548), .B2(n16394), .A(n11165), .ZN(n11202) );
  INV_X1 U14399 ( .A(n11167), .ZN(n12312) );
  INV_X1 U14400 ( .A(n12291), .ZN(n11169) );
  NOR3_X1 U14401 ( .A1(n11169), .A2(n10870), .A3(n14300), .ZN(n11172) );
  NAND2_X1 U14402 ( .A1(n12285), .A2(n14300), .ZN(n11170) );
  XNOR2_X1 U14403 ( .A(n11170), .B(n12291), .ZN(n13137) );
  INV_X1 U14404 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14302) );
  NOR2_X1 U14405 ( .A1(n13137), .A2(n14302), .ZN(n11171) );
  NOR2_X1 U14406 ( .A1(n11172), .A2(n11171), .ZN(n11174) );
  XNOR2_X1 U14407 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11174), .ZN(
        n14700) );
  XNOR2_X1 U14408 ( .A(n11173), .B(n12300), .ZN(n14699) );
  NAND2_X1 U14409 ( .A1(n14700), .A2(n14699), .ZN(n14698) );
  OR2_X1 U14410 ( .A1(n11174), .A2(n19722), .ZN(n11175) );
  NAND2_X1 U14411 ( .A1(n14698), .A2(n11175), .ZN(n11176) );
  XNOR2_X1 U14412 ( .A(n11176), .B(n16715), .ZN(n14655) );
  NAND2_X1 U14413 ( .A1(n11176), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11177) );
  NAND2_X1 U14414 ( .A1(n16412), .A2(n19717), .ZN(n11178) );
  NAND2_X1 U14415 ( .A1(n11181), .A2(n11184), .ZN(n11187) );
  XNOR2_X1 U14416 ( .A(n11188), .B(n11189), .ZN(n11186) );
  INV_X1 U14417 ( .A(n11186), .ZN(n11180) );
  NAND2_X1 U14418 ( .A1(n11187), .A2(n11180), .ZN(n11183) );
  NAND2_X1 U14419 ( .A1(n11191), .A2(n11190), .ZN(n11192) );
  INV_X1 U14420 ( .A(n11194), .ZN(n11195) );
  AND2_X1 U14421 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16631) );
  NAND2_X1 U14422 ( .A1(n16631), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16589) );
  NAND2_X1 U14423 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11197) );
  NOR2_X1 U14424 ( .A1(n16589), .A2(n11197), .ZN(n16582) );
  NAND2_X1 U14425 ( .A1(n16582), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12803) );
  AND2_X1 U14426 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16544) );
  NAND3_X1 U14427 ( .A1(n16544), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11198) );
  OR2_X1 U14428 ( .A1(n12803), .A2(n11198), .ZN(n16524) );
  NOR2_X1 U14429 ( .A1(n16524), .A2(n16251), .ZN(n16522) );
  AND2_X1 U14430 ( .A1(n16522), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12816) );
  NAND2_X1 U14431 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16492) );
  INV_X1 U14432 ( .A(n16492), .ZN(n11199) );
  AND2_X1 U14433 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16432) );
  NAND2_X1 U14434 ( .A1(n16432), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12759) );
  INV_X1 U14435 ( .A(n19579), .ZN(n11201) );
  AOI22_X1 U14436 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11206) );
  AND2_X2 U14437 ( .A1(n13979), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14007) );
  AND2_X2 U14438 ( .A1(n11208), .A2(n14007), .ZN(n11376) );
  AND2_X2 U14439 ( .A1(n11207), .A2(n14014), .ZN(n11368) );
  AOI22_X1 U14440 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12876), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11205) );
  AOI22_X1 U14441 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11204) );
  AOI22_X1 U14442 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11203) );
  NAND4_X1 U14443 ( .A1(n11206), .A2(n11205), .A3(n11204), .A4(n11203), .ZN(
        n11214) );
  AND2_X4 U14444 ( .A1(n14007), .A2(n13978), .ZN(n11423) );
  AOI22_X1 U14445 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11212) );
  AND2_X4 U14446 ( .A1(n11208), .A2(n14013), .ZN(n11411) );
  AOI22_X1 U14447 ( .A1(n11411), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U14448 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11210) );
  AOI22_X1 U14449 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11209) );
  NAND4_X1 U14450 ( .A1(n11212), .A2(n11211), .A3(n11210), .A4(n11209), .ZN(
        n11213) );
  OR2_X1 U14451 ( .A1(n11214), .A2(n11213), .ZN(n12864) );
  AOI22_X1 U14452 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11218) );
  AOI22_X1 U14453 ( .A1(n11411), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U14454 ( .A1(n12887), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12876), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14455 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11215) );
  NAND4_X1 U14456 ( .A1(n11218), .A2(n11217), .A3(n11216), .A4(n11215), .ZN(
        n11224) );
  AOI22_X1 U14457 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11222) );
  AOI22_X1 U14458 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U14459 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11220) );
  AOI22_X1 U14460 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11219) );
  NAND4_X1 U14461 ( .A1(n11222), .A2(n11221), .A3(n11220), .A4(n11219), .ZN(
        n11223) );
  NOR2_X1 U14462 ( .A1(n11224), .A2(n11223), .ZN(n11905) );
  AOI22_X1 U14463 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11228) );
  AOI22_X1 U14464 ( .A1(n11431), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11227) );
  AOI22_X1 U14465 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12876), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11226) );
  AOI22_X1 U14466 ( .A1(n12857), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11225) );
  NAND4_X1 U14467 ( .A1(n11228), .A2(n11227), .A3(n11226), .A4(n11225), .ZN(
        n11234) );
  AOI22_X1 U14468 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11859), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11232) );
  AOI22_X1 U14469 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11231) );
  AOI22_X1 U14470 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14471 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11229) );
  NAND4_X1 U14472 ( .A1(n11232), .A2(n11231), .A3(n11230), .A4(n11229), .ZN(
        n11233) );
  NOR2_X1 U14473 ( .A1(n11234), .A2(n11233), .ZN(n11889) );
  AOI22_X1 U14474 ( .A1(n11431), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11238) );
  AOI22_X1 U14475 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11425), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11237) );
  AOI22_X1 U14476 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12852), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U14477 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12857), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11235) );
  NAND4_X1 U14478 ( .A1(n11238), .A2(n11237), .A3(n11236), .A4(n11235), .ZN(
        n11244) );
  AOI22_X1 U14479 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11450), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11242) );
  AOI22_X1 U14480 ( .A1(n12887), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11241) );
  AOI22_X1 U14481 ( .A1(n12886), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11240) );
  AOI22_X1 U14482 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11239) );
  NAND4_X1 U14483 ( .A1(n11242), .A2(n11241), .A3(n11240), .A4(n11239), .ZN(
        n11243) );
  NOR2_X1 U14484 ( .A1(n11244), .A2(n11243), .ZN(n11870) );
  AOI22_X1 U14485 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11248) );
  AOI22_X1 U14486 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11247) );
  AOI22_X1 U14487 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11246) );
  AOI22_X1 U14488 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11245) );
  NAND4_X1 U14489 ( .A1(n11248), .A2(n11247), .A3(n11246), .A4(n11245), .ZN(
        n11254) );
  AOI22_X1 U14490 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11252) );
  AOI22_X1 U14491 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12876), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11251) );
  AOI22_X1 U14492 ( .A1(n12857), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11250) );
  AOI22_X1 U14493 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11249) );
  NAND4_X1 U14494 ( .A1(n11252), .A2(n11251), .A3(n11250), .A4(n11249), .ZN(
        n11253) );
  NOR2_X1 U14495 ( .A1(n11254), .A2(n11253), .ZN(n11871) );
  NOR2_X1 U14496 ( .A1(n11870), .A2(n11871), .ZN(n11881) );
  AOI22_X1 U14497 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11258) );
  AOI22_X1 U14498 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11257) );
  AOI22_X1 U14499 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11256) );
  AOI22_X1 U14500 ( .A1(n12887), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11255) );
  NAND4_X1 U14501 ( .A1(n11258), .A2(n11257), .A3(n11256), .A4(n11255), .ZN(
        n11264) );
  AOI22_X1 U14502 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11789), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11262) );
  AOI22_X1 U14503 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n12877), .B1(
        n12876), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11261) );
  AOI22_X1 U14504 ( .A1(n12857), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11260) );
  AOI22_X1 U14505 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12852), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11259) );
  NAND4_X1 U14506 ( .A1(n11262), .A2(n11261), .A3(n11260), .A4(n11259), .ZN(
        n11263) );
  OR2_X1 U14507 ( .A1(n11264), .A2(n11263), .ZN(n11880) );
  NAND2_X1 U14508 ( .A1(n11881), .A2(n11880), .ZN(n11888) );
  NOR2_X1 U14509 ( .A1(n11889), .A2(n11888), .ZN(n11897) );
  AOI22_X1 U14510 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U14511 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11267) );
  AOI22_X1 U14512 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U14513 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11265) );
  NAND4_X1 U14514 ( .A1(n11268), .A2(n11267), .A3(n11266), .A4(n11265), .ZN(
        n11274) );
  AOI22_X1 U14515 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11272) );
  AOI22_X1 U14516 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12876), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11271) );
  AOI22_X1 U14517 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11270) );
  AOI22_X1 U14518 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11269) );
  NAND4_X1 U14519 ( .A1(n11272), .A2(n11271), .A3(n11270), .A4(n11269), .ZN(
        n11273) );
  NAND2_X1 U14520 ( .A1(n11897), .A2(n11898), .ZN(n11904) );
  NOR2_X1 U14521 ( .A1(n11905), .A2(n11904), .ZN(n12865) );
  XOR2_X1 U14522 ( .A(n12864), .B(n12865), .Z(n11314) );
  AOI22_X1 U14523 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11759), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11278) );
  AOI22_X1 U14524 ( .A1(n11411), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11430), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11277) );
  AOI22_X1 U14525 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11424), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11276) );
  AOI22_X1 U14526 ( .A1(n12887), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11374), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11275) );
  AOI22_X1 U14527 ( .A1(n11367), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11366), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U14528 ( .A1(n11376), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11281) );
  AOI22_X1 U14529 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11375), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U14530 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11432), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11279) );
  NAND2_X2 U14531 ( .A1(n9647), .A2(n10476), .ZN(n11385) );
  AOI22_X1 U14532 ( .A1(n11411), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11430), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14533 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11424), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U14534 ( .A1(n11376), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11284) );
  AOI22_X1 U14535 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11432), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11283) );
  NAND4_X1 U14536 ( .A1(n11286), .A2(n11285), .A3(n11284), .A4(n11283), .ZN(
        n11292) );
  AOI22_X1 U14537 ( .A1(n11367), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11366), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11290) );
  AOI22_X1 U14538 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11759), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11289) );
  AOI22_X1 U14539 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11375), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11288) );
  AOI22_X1 U14540 ( .A1(n12887), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11374), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11287) );
  NAND4_X1 U14541 ( .A1(n11290), .A2(n11289), .A3(n11288), .A4(n11287), .ZN(
        n11291) );
  OR2_X2 U14542 ( .A1(n11292), .A2(n11291), .ZN(n11391) );
  AOI22_X1 U14543 ( .A1(n11411), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11424), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11296) );
  AOI22_X1 U14544 ( .A1(n11376), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11374), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U14545 ( .A1(n11368), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12879), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11294) );
  AOI22_X1 U14546 ( .A1(n11367), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11432), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11293) );
  AOI22_X1 U14547 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11759), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11300) );
  AOI22_X1 U14548 ( .A1(n11430), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11299) );
  AOI22_X1 U14549 ( .A1(n11366), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11298) );
  AOI22_X1 U14550 ( .A1(n11430), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11759), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11304) );
  AOI22_X1 U14551 ( .A1(n12887), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11424), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11303) );
  AOI22_X1 U14552 ( .A1(n11376), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11375), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11302) );
  AOI22_X1 U14553 ( .A1(n11366), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12879), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14554 ( .A1(n11368), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11432), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11306) );
  AOI22_X1 U14555 ( .A1(n11367), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11305) );
  NAND3_X1 U14556 ( .A1(n11307), .A2(n11306), .A3(n11305), .ZN(n11310) );
  AOI22_X1 U14557 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11374), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11308) );
  NAND2_X2 U14558 ( .A1(n11312), .A2(n11311), .ZN(n11383) );
  INV_X1 U14559 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n15077) );
  INV_X1 U14560 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15169) );
  OAI22_X1 U14561 ( .A1(n12900), .A2(n15077), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15169), .ZN(n11313) );
  AOI21_X1 U14562 ( .B1(n11314), .B2(n12896), .A(n11313), .ZN(n11325) );
  OR3_X4 U14563 ( .A1(n11772), .A2(n15267), .A3(n15251), .ZN(n11852) );
  OR2_X2 U14564 ( .A1(n11875), .A2(n14800), .ZN(n11879) );
  INV_X1 U14565 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11893) );
  OR2_X2 U14566 ( .A1(n11894), .A2(n11893), .ZN(n11901) );
  INV_X1 U14567 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15189) );
  XNOR2_X1 U14568 ( .A(n11916), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15166) );
  MUX2_X1 U14569 ( .A(n11325), .B(n15166), .S(n11910), .Z(n11915) );
  NAND2_X1 U14570 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11329) );
  NAND2_X1 U14571 ( .A1(n11411), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11328) );
  NAND2_X1 U14572 ( .A1(n11430), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11327) );
  NAND2_X1 U14573 ( .A1(n11759), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11326) );
  NAND2_X1 U14574 ( .A1(n11368), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11332) );
  NAND2_X1 U14575 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11331) );
  NAND2_X1 U14576 ( .A1(n11375), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11330) );
  NAND2_X1 U14577 ( .A1(n11374), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11333) );
  NAND2_X1 U14578 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11338) );
  NAND2_X1 U14579 ( .A1(n11411), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11337) );
  NAND2_X1 U14580 ( .A1(n11430), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11336) );
  NAND2_X1 U14581 ( .A1(n11759), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11335) );
  NAND2_X1 U14582 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11342) );
  NAND2_X1 U14583 ( .A1(n12887), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11341) );
  NAND2_X1 U14584 ( .A1(n11424), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11340) );
  NAND2_X1 U14585 ( .A1(n11367), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11346) );
  NAND2_X1 U14586 ( .A1(n11366), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11345) );
  NAND2_X1 U14587 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11344) );
  NAND2_X1 U14588 ( .A1(n11432), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11343) );
  NAND2_X1 U14589 ( .A1(n11376), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11350) );
  NAND2_X1 U14590 ( .A1(n11368), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11349) );
  NAND2_X1 U14591 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11348) );
  NAND4_X4 U14592 ( .A1(n11354), .A2(n11353), .A3(n11352), .A4(n11351), .ZN(
        n11993) );
  AOI22_X1 U14593 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11759), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U14594 ( .A1(n11411), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11430), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14595 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11424), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14596 ( .A1(n12887), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11374), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11356) );
  NAND4_X1 U14597 ( .A1(n11359), .A2(n11358), .A3(n11357), .A4(n11356), .ZN(
        n11365) );
  AOI22_X1 U14598 ( .A1(n11367), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11366), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14599 ( .A1(n11376), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14600 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11375), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11361) );
  AOI22_X1 U14601 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11432), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11360) );
  NAND4_X1 U14602 ( .A1(n11363), .A2(n11362), .A3(n11361), .A4(n11360), .ZN(
        n11364) );
  OR2_X2 U14603 ( .A1(n11365), .A2(n11364), .ZN(n12124) );
  AOI22_X1 U14604 ( .A1(n12887), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11759), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14605 ( .A1(n11367), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11366), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U14606 ( .A1(n11368), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12879), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14607 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11432), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11370) );
  AOI22_X1 U14608 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11430), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11380) );
  AOI22_X1 U14609 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11374), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11379) );
  NAND2_X1 U14610 ( .A1(n11381), .A2(n11993), .ZN(n12230) );
  OAI211_X1 U14611 ( .C1(n20747), .C2(n12108), .A(n12243), .B(n12230), .ZN(
        n11405) );
  NAND2_X1 U14612 ( .A1(n20715), .A2(n14053), .ZN(n15004) );
  NAND2_X1 U14613 ( .A1(n14010), .A2(n15004), .ZN(n11382) );
  NOR2_X1 U14614 ( .A1(n11405), .A2(n11382), .ZN(n11395) );
  NAND3_X1 U14615 ( .A1(n12117), .A2(n13243), .A3(n20757), .ZN(n12206) );
  XNOR2_X1 U14616 ( .A(n21315), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n12091) );
  NAND2_X1 U14617 ( .A1(n11391), .A2(n11385), .ZN(n11384) );
  NAND2_X1 U14618 ( .A1(n11390), .A2(n12124), .ZN(n11400) );
  NAND2_X1 U14619 ( .A1(n11386), .A2(n14713), .ZN(n11387) );
  NAND2_X1 U14620 ( .A1(n11399), .A2(n20715), .ZN(n11394) );
  NAND2_X1 U14621 ( .A1(n11398), .A2(n12212), .ZN(n11393) );
  NAND4_X1 U14622 ( .A1(n11395), .A2(n11463), .A3(n11394), .A4(n11393), .ZN(
        n11396) );
  INV_X1 U14623 ( .A(n11476), .ZN(n11499) );
  MUX2_X1 U14624 ( .A(n14054), .B(n21377), .S(n21157), .Z(n11397) );
  NAND3_X1 U14625 ( .A1(n11398), .A2(n14053), .A3(n12212), .ZN(n11408) );
  NOR2_X1 U14626 ( .A1(n14053), .A2(n11993), .ZN(n12238) );
  OAI21_X1 U14627 ( .B1(n12238), .B2(n11400), .A(n11399), .ZN(n11407) );
  NAND2_X1 U14628 ( .A1(n13980), .A2(n20757), .ZN(n12244) );
  NAND2_X1 U14629 ( .A1(n9841), .A2(n12979), .ZN(n11403) );
  AND2_X1 U14630 ( .A1(n15565), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11402) );
  NAND4_X1 U14631 ( .A1(n12244), .A2(n11403), .A3(n11402), .A4(n15004), .ZN(
        n11404) );
  NOR2_X1 U14632 ( .A1(n11405), .A2(n11404), .ZN(n11406) );
  AOI22_X1 U14633 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11416) );
  BUF_X1 U14634 ( .A(n11411), .Z(n11450) );
  AOI22_X1 U14635 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14636 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14637 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11413) );
  NAND4_X1 U14638 ( .A1(n11416), .A2(n11415), .A3(n11414), .A4(n11413), .ZN(
        n11422) );
  AOI22_X1 U14639 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11420) );
  AOI22_X1 U14640 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14641 ( .A1(n12857), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U14642 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11432), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11417) );
  NAND4_X1 U14643 ( .A1(n11420), .A2(n11419), .A3(n11418), .A4(n11417), .ZN(
        n11421) );
  INV_X1 U14644 ( .A(n12169), .ZN(n12177) );
  AND2_X1 U14645 ( .A1(n11492), .A2(n12177), .ZN(n11445) );
  AOI22_X1 U14646 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U14647 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U14648 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14649 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11426) );
  NAND4_X1 U14650 ( .A1(n11429), .A2(n11428), .A3(n11427), .A4(n11426), .ZN(
        n11438) );
  AOI22_X1 U14651 ( .A1(n11431), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11859), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U14652 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14653 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14654 ( .A1(n12857), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11432), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11433) );
  NAND4_X1 U14655 ( .A1(n11436), .A2(n11435), .A3(n11434), .A4(n11433), .ZN(
        n11437) );
  MUX2_X1 U14656 ( .A(n12174), .B(n11445), .S(n12123), .Z(n11439) );
  INV_X1 U14657 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11443) );
  AOI21_X1 U14658 ( .B1(n20715), .B2(n12123), .A(n10072), .ZN(n11442) );
  INV_X1 U14659 ( .A(n12174), .ZN(n11444) );
  INV_X1 U14660 ( .A(n11445), .ZN(n11459) );
  NAND2_X1 U14661 ( .A1(n11961), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11458) );
  AOI22_X1 U14662 ( .A1(n11431), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14663 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11448) );
  AOI22_X1 U14664 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11447) );
  AOI22_X1 U14665 ( .A1(n12886), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11446) );
  NAND4_X1 U14666 ( .A1(n11449), .A2(n11448), .A3(n11447), .A4(n11446), .ZN(
        n11456) );
  AOI22_X1 U14667 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11450), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U14668 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n12877), .B1(
        n11425), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14669 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12857), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U14670 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11432), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11451) );
  NAND4_X1 U14671 ( .A1(n11454), .A2(n11453), .A3(n11452), .A4(n11451), .ZN(
        n11455) );
  NAND2_X1 U14672 ( .A1(n11493), .A2(n12116), .ZN(n11457) );
  NAND3_X1 U14673 ( .A1(n13980), .A2(n12238), .A3(n20752), .ZN(n13975) );
  NAND2_X1 U14674 ( .A1(n11463), .A2(n12227), .ZN(n11464) );
  NAND2_X1 U14675 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11478) );
  OAI21_X1 U14676 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11478), .ZN(n21184) );
  NAND2_X1 U14677 ( .A1(n15580), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11473) );
  OAI21_X1 U14678 ( .B1(n21377), .B2(n21184), .A(n11473), .ZN(n11466) );
  INV_X1 U14679 ( .A(n11466), .ZN(n11467) );
  INV_X1 U14680 ( .A(n11470), .ZN(n11471) );
  NAND2_X1 U14681 ( .A1(n11473), .A2(n11465), .ZN(n11474) );
  INV_X1 U14682 ( .A(n11478), .ZN(n11477) );
  NAND2_X1 U14683 ( .A1(n11477), .A2(n21123), .ZN(n21093) );
  NAND2_X1 U14684 ( .A1(n11478), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11479) );
  NAND2_X1 U14685 ( .A1(n21093), .A2(n11479), .ZN(n20727) );
  INV_X1 U14686 ( .A(n21377), .ZN(n11502) );
  AOI22_X1 U14687 ( .A1(n20727), .A2(n11502), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15580), .ZN(n11480) );
  AOI22_X1 U14688 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14689 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14690 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U14691 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11482) );
  NAND4_X1 U14692 ( .A1(n11485), .A2(n11484), .A3(n11483), .A4(n11482), .ZN(
        n11491) );
  AOI22_X1 U14693 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11489) );
  INV_X1 U14694 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n21521) );
  AOI22_X1 U14695 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12876), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U14696 ( .A1(n12857), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U14697 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11486) );
  NAND4_X1 U14698 ( .A1(n11489), .A2(n11488), .A3(n11487), .A4(n11486), .ZN(
        n11490) );
  INV_X1 U14699 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11494) );
  OAI22_X1 U14700 ( .A1(n12135), .A2(n11505), .B1(n11958), .B2(n11494), .ZN(
        n11495) );
  NAND2_X1 U14701 ( .A1(n11499), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11504) );
  NAND3_X1 U14702 ( .A1(n21186), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20965) );
  INV_X1 U14703 ( .A(n20965), .ZN(n11500) );
  NAND2_X1 U14704 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11500), .ZN(
        n20963) );
  NAND2_X1 U14705 ( .A1(n21186), .A2(n20963), .ZN(n11501) );
  NOR3_X1 U14706 ( .A1(n21186), .A2(n21123), .A3(n13998), .ZN(n21247) );
  NAND2_X1 U14707 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21247), .ZN(
        n21235) );
  AOI22_X1 U14708 ( .A1(n11502), .A2(n20874), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15580), .ZN(n11503) );
  AOI22_X1 U14709 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12887), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14710 ( .A1(n11431), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11509) );
  AOI22_X1 U14711 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12857), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U14712 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11507) );
  NAND4_X1 U14713 ( .A1(n11510), .A2(n11509), .A3(n11508), .A4(n11507), .ZN(
        n11517) );
  AOI22_X1 U14714 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U14715 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12852), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U14716 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U14717 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11512) );
  NAND4_X1 U14718 ( .A1(n11515), .A2(n11514), .A3(n11513), .A4(n11512), .ZN(
        n11516) );
  AOI22_X1 U14719 ( .A1(n11976), .A2(n12149), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n11961), .ZN(n11518) );
  AOI22_X1 U14720 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14721 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14722 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U14723 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11521) );
  NAND4_X1 U14724 ( .A1(n11524), .A2(n11523), .A3(n11522), .A4(n11521), .ZN(
        n11530) );
  AOI22_X1 U14725 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11528) );
  AOI22_X1 U14726 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12876), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14727 ( .A1(n12857), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14728 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11525) );
  NAND4_X1 U14729 ( .A1(n11528), .A2(n11527), .A3(n11526), .A4(n11525), .ZN(
        n11529) );
  NAND2_X1 U14730 ( .A1(n11976), .A2(n12150), .ZN(n11532) );
  NAND2_X1 U14731 ( .A1(n11961), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11531) );
  AOI22_X1 U14732 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14733 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14734 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11534) );
  AOI22_X1 U14735 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11533) );
  NAND4_X1 U14736 ( .A1(n11536), .A2(n11535), .A3(n11534), .A4(n11533), .ZN(
        n11542) );
  AOI22_X1 U14737 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12852), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11540) );
  AOI22_X1 U14738 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U14739 ( .A1(n12857), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14740 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11537) );
  NAND4_X1 U14741 ( .A1(n11540), .A2(n11539), .A3(n11538), .A4(n11537), .ZN(
        n11541) );
  AOI22_X1 U14742 ( .A1(n11976), .A2(n12159), .B1(n11961), .B2(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11554) );
  INV_X1 U14743 ( .A(n11554), .ZN(n11543) );
  NAND2_X1 U14744 ( .A1(n11544), .A2(n11543), .ZN(n11547) );
  NAND2_X1 U14745 ( .A1(n11545), .A2(n11554), .ZN(n11546) );
  INV_X1 U14746 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11552) );
  AND2_X1 U14747 ( .A1(n11605), .A2(n11549), .ZN(n11548) );
  OR2_X1 U14748 ( .A1(n11548), .A2(n11565), .ZN(n20543) );
  NAND2_X1 U14749 ( .A1(n21239), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11785) );
  NOR2_X1 U14750 ( .A1(n11785), .A2(n11549), .ZN(n11550) );
  AOI21_X1 U14751 ( .B1(n20543), .B2(n11910), .A(n11550), .ZN(n11551) );
  OAI21_X1 U14752 ( .B1(n12900), .B2(n11552), .A(n11551), .ZN(n11553) );
  AOI21_X1 U14753 ( .B1(n12148), .B2(n11727), .A(n11553), .ZN(n15064) );
  AOI22_X1 U14754 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U14755 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14756 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14757 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11555) );
  NAND4_X1 U14758 ( .A1(n11558), .A2(n11557), .A3(n11556), .A4(n11555), .ZN(
        n11564) );
  AOI22_X1 U14759 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U14760 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12876), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14761 ( .A1(n12857), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11560) );
  AOI22_X1 U14762 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11559) );
  NAND4_X1 U14763 ( .A1(n11562), .A2(n11561), .A3(n11560), .A4(n11559), .ZN(
        n11563) );
  AOI22_X1 U14764 ( .A1(n11976), .A2(n12167), .B1(n11961), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11611) );
  NAND2_X1 U14765 ( .A1(n11610), .A2(n11611), .ZN(n12157) );
  INV_X1 U14766 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11568) );
  NOR2_X1 U14767 ( .A1(n11565), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11566) );
  OR2_X1 U14768 ( .A1(n11616), .A2(n11566), .ZN(n20534) );
  AOI22_X1 U14769 ( .A1(n20534), .A2(n11910), .B1(n12903), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11567) );
  OAI21_X1 U14770 ( .B1(n12900), .B2(n11568), .A(n11567), .ZN(n11569) );
  NAND2_X1 U14771 ( .A1(n11571), .A2(n11570), .ZN(n11572) );
  INV_X1 U14772 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15008) );
  XNOR2_X1 U14773 ( .A(n15008), .B(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n20576) );
  OAI21_X1 U14774 ( .B1(n20576), .B2(n12902), .A(n11785), .ZN(n11573) );
  AOI21_X1 U14775 ( .B1(n12904), .B2(P1_EAX_REG_2__SCAN_IN), .A(n11573), .ZN(
        n11574) );
  INV_X1 U14776 ( .A(n11574), .ZN(n11575) );
  NAND2_X1 U14777 ( .A1(n12903), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11592) );
  INV_X1 U14778 ( .A(n11577), .ZN(n11579) );
  XNOR2_X2 U14779 ( .A(n11579), .B(n11578), .ZN(n15543) );
  NAND2_X1 U14780 ( .A1(n15543), .A2(n11727), .ZN(n11583) );
  INV_X1 U14781 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n11580) );
  OAI22_X1 U14782 ( .A1(n12900), .A2(n11580), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15008), .ZN(n11581) );
  AOI21_X1 U14783 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11597), .A(
        n11581), .ZN(n11582) );
  NAND2_X1 U14784 ( .A1(n21155), .A2(n20757), .ZN(n11585) );
  NAND2_X1 U14785 ( .A1(n11585), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13247) );
  INV_X1 U14786 ( .A(n11597), .ZN(n11604) );
  NAND2_X1 U14787 ( .A1(n12904), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11588) );
  NAND2_X1 U14788 ( .A1(n21239), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11587) );
  OAI211_X1 U14789 ( .C1(n11604), .C2(n10177), .A(n11588), .B(n11587), .ZN(
        n11589) );
  AOI21_X1 U14790 ( .B1(n11586), .B2(n11727), .A(n11589), .ZN(n11590) );
  OR2_X1 U14791 ( .A1(n13247), .A2(n11590), .ZN(n13248) );
  INV_X1 U14792 ( .A(n11590), .ZN(n13249) );
  OR2_X1 U14793 ( .A1(n13249), .A2(n12902), .ZN(n11591) );
  NAND2_X1 U14794 ( .A1(n13248), .A2(n11591), .ZN(n13615) );
  NOR2_X1 U14795 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11594), .ZN(
        n11595) );
  NOR2_X1 U14796 ( .A1(n11606), .A2(n11595), .ZN(n20561) );
  INV_X1 U14797 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20566) );
  OAI22_X1 U14798 ( .A1(n20561), .A2(n12902), .B1(n11785), .B2(n20566), .ZN(
        n11596) );
  AOI21_X1 U14799 ( .B1(n12904), .B2(P1_EAX_REG_3__SCAN_IN), .A(n11596), .ZN(
        n11599) );
  NAND2_X1 U14800 ( .A1(n11597), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11598) );
  NAND2_X1 U14801 ( .A1(n13959), .A2(n13960), .ZN(n14146) );
  XNOR2_X1 U14802 ( .A(n11601), .B(n11600), .ZN(n12110) );
  INV_X1 U14803 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14039) );
  NAND2_X1 U14804 ( .A1(n21239), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11603) );
  NAND2_X1 U14805 ( .A1(n12904), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11602) );
  OAI211_X1 U14806 ( .C1(n11604), .C2(n14039), .A(n11603), .B(n11602), .ZN(
        n11607) );
  OAI21_X1 U14807 ( .B1(n11606), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11605), .ZN(n20653) );
  MUX2_X1 U14808 ( .A(n11607), .B(n20653), .S(n11910), .Z(n11608) );
  INV_X1 U14809 ( .A(n11611), .ZN(n11612) );
  INV_X1 U14810 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11614) );
  NAND2_X1 U14811 ( .A1(n11976), .A2(n12169), .ZN(n11613) );
  OAI21_X1 U14812 ( .B1(n11614), .B2(n11958), .A(n11613), .ZN(n11615) );
  INV_X1 U14813 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11619) );
  OR2_X1 U14814 ( .A1(n11616), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11617) );
  NAND2_X1 U14815 ( .A1(n11617), .A2(n11633), .ZN(n20521) );
  AOI22_X1 U14816 ( .A1(n20521), .A2(n11910), .B1(n12903), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11618) );
  OAI21_X1 U14817 ( .B1(n12900), .B2(n11619), .A(n11618), .ZN(n11620) );
  INV_X1 U14818 ( .A(n11620), .ZN(n11621) );
  AOI22_X1 U14819 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U14820 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11425), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U14821 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12852), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14822 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11623) );
  NAND4_X1 U14823 ( .A1(n11626), .A2(n11625), .A3(n11624), .A4(n11623), .ZN(
        n11632) );
  AOI22_X1 U14824 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U14825 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14826 ( .A1(n12886), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11628) );
  AOI22_X1 U14827 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12857), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11627) );
  NAND4_X1 U14828 ( .A1(n11630), .A2(n11629), .A3(n11628), .A4(n11627), .ZN(
        n11631) );
  NOR2_X1 U14829 ( .A1(n11632), .A2(n11631), .ZN(n11636) );
  XNOR2_X1 U14830 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11633), .ZN(
        n15346) );
  OAI22_X1 U14831 ( .A1(n15346), .A2(n12902), .B1(n11785), .B2(n15343), .ZN(
        n11634) );
  INV_X1 U14832 ( .A(n11634), .ZN(n11635) );
  OAI21_X1 U14833 ( .B1(n11751), .B2(n11636), .A(n11635), .ZN(n11639) );
  INV_X1 U14834 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n11637) );
  NOR2_X1 U14835 ( .A1(n12900), .A2(n11637), .ZN(n11638) );
  AOI22_X1 U14836 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U14837 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11642) );
  AOI22_X1 U14838 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n12877), .B1(
        n12876), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U14839 ( .A1(n12880), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11640) );
  NAND4_X1 U14840 ( .A1(n11643), .A2(n11642), .A3(n11641), .A4(n11640), .ZN(
        n11649) );
  AOI22_X1 U14841 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11789), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14842 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14843 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14844 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12857), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11644) );
  NAND4_X1 U14845 ( .A1(n11647), .A2(n11646), .A3(n11645), .A4(n11644), .ZN(
        n11648) );
  NOR2_X1 U14846 ( .A1(n11649), .A2(n11648), .ZN(n11652) );
  INV_X1 U14847 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20508) );
  XOR2_X1 U14848 ( .A(n20508), .B(n11650), .Z(n20506) );
  INV_X1 U14849 ( .A(n20506), .ZN(n15336) );
  AOI22_X1 U14850 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n12903), .B1(
        n11910), .B2(n15336), .ZN(n11651) );
  OAI21_X1 U14851 ( .B1(n11751), .B2(n11652), .A(n11651), .ZN(n11655) );
  INV_X1 U14852 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n11653) );
  NOR2_X1 U14853 ( .A1(n12900), .A2(n11653), .ZN(n11654) );
  AOI22_X1 U14854 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14855 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14856 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14857 ( .A1(n12886), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11656) );
  NAND4_X1 U14858 ( .A1(n11659), .A2(n11658), .A3(n11657), .A4(n11656), .ZN(
        n11665) );
  AOI22_X1 U14859 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12887), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U14860 ( .A1(n11411), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11662) );
  AOI22_X1 U14861 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U14862 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12857), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11660) );
  NAND4_X1 U14863 ( .A1(n11663), .A2(n11662), .A3(n11661), .A4(n11660), .ZN(
        n11664) );
  NOR2_X1 U14864 ( .A1(n11665), .A2(n11664), .ZN(n11670) );
  NAND2_X1 U14865 ( .A1(n12904), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11669) );
  XNOR2_X1 U14866 ( .A(n11666), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17354) );
  OAI22_X1 U14867 ( .A1(n17354), .A2(n12902), .B1(n17348), .B2(n11785), .ZN(
        n11667) );
  INV_X1 U14868 ( .A(n11667), .ZN(n11668) );
  OAI211_X1 U14869 ( .C1(n11670), .C2(n11751), .A(n11669), .B(n11668), .ZN(
        n15047) );
  AOI22_X1 U14870 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U14871 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U14872 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14873 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11671) );
  NAND4_X1 U14874 ( .A1(n11674), .A2(n11673), .A3(n11672), .A4(n11671), .ZN(
        n11680) );
  AOI22_X1 U14875 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14876 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12852), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U14877 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14878 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12857), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11675) );
  NAND4_X1 U14879 ( .A1(n11678), .A2(n11677), .A3(n11676), .A4(n11675), .ZN(
        n11679) );
  NOR2_X1 U14880 ( .A1(n11680), .A2(n11679), .ZN(n11681) );
  NOR2_X1 U14881 ( .A1(n11751), .A2(n11681), .ZN(n14977) );
  INV_X1 U14882 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n11687) );
  INV_X1 U14883 ( .A(n11730), .ZN(n11748) );
  INV_X1 U14884 ( .A(n11682), .ZN(n11684) );
  INV_X1 U14885 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11683) );
  NAND2_X1 U14886 ( .A1(n11684), .A2(n11683), .ZN(n11685) );
  NAND2_X1 U14887 ( .A1(n11748), .A2(n11685), .ZN(n15318) );
  AOI22_X1 U14888 ( .A1(n15318), .A2(n11910), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12903), .ZN(n11686) );
  OAI21_X1 U14889 ( .B1(n12900), .B2(n11687), .A(n11686), .ZN(n14941) );
  AOI22_X1 U14890 ( .A1(n11431), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14891 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12852), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14892 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U14893 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11688) );
  NAND4_X1 U14894 ( .A1(n11691), .A2(n11690), .A3(n11689), .A4(n11688), .ZN(
        n11697) );
  AOI22_X1 U14895 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11450), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14896 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14897 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12857), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14898 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11692) );
  NAND4_X1 U14899 ( .A1(n11695), .A2(n11694), .A3(n11693), .A4(n11692), .ZN(
        n11696) );
  OAI21_X1 U14900 ( .B1(n11697), .B2(n11696), .A(n11727), .ZN(n11701) );
  NAND2_X1 U14901 ( .A1(n12904), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11700) );
  INV_X1 U14902 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11712) );
  XNOR2_X1 U14903 ( .A(n11713), .B(n11712), .ZN(n15280) );
  NAND2_X1 U14904 ( .A1(n15280), .A2(n11910), .ZN(n11699) );
  NAND2_X1 U14905 ( .A1(n12903), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11698) );
  NAND4_X1 U14906 ( .A1(n11701), .A2(n11700), .A3(n11699), .A4(n11698), .ZN(
        n14928) );
  AOI22_X1 U14907 ( .A1(n11431), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14908 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U14909 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12852), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11703) );
  AOI22_X1 U14910 ( .A1(n12857), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11702) );
  NAND4_X1 U14911 ( .A1(n11705), .A2(n11704), .A3(n11703), .A4(n11702), .ZN(
        n11711) );
  AOI22_X1 U14912 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11450), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14913 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12887), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14914 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11707) );
  AOI22_X1 U14915 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11706) );
  NAND4_X1 U14916 ( .A1(n11709), .A2(n11708), .A3(n11707), .A4(n11706), .ZN(
        n11710) );
  NOR2_X1 U14917 ( .A1(n11711), .A2(n11710), .ZN(n11718) );
  NAND2_X1 U14918 ( .A1(n12904), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11717) );
  INV_X1 U14919 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n21496) );
  OAI21_X1 U14920 ( .B1(n11713), .B2(n11712), .A(n21496), .ZN(n11714) );
  NAND2_X1 U14921 ( .A1(n11714), .A2(n11772), .ZN(n15272) );
  NOR2_X1 U14922 ( .A1(n11785), .A2(n21496), .ZN(n11715) );
  AOI21_X1 U14923 ( .B1(n15272), .B2(n11910), .A(n11715), .ZN(n11716) );
  OAI211_X1 U14924 ( .C1(n11718), .C2(n11751), .A(n11717), .B(n11716), .ZN(
        n14916) );
  OAI211_X1 U14925 ( .C1(n14977), .C2(n14941), .A(n14928), .B(n14916), .ZN(
        n11753) );
  AOI22_X1 U14926 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11722) );
  AOI22_X1 U14927 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12887), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11721) );
  AOI22_X1 U14928 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12852), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14929 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12857), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11719) );
  NAND4_X1 U14930 ( .A1(n11722), .A2(n11721), .A3(n11720), .A4(n11719), .ZN(
        n11729) );
  AOI22_X1 U14931 ( .A1(n11411), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U14932 ( .A1(n11511), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U14933 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11724) );
  AOI22_X1 U14934 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11723) );
  NAND4_X1 U14935 ( .A1(n11726), .A2(n11725), .A3(n11724), .A4(n11723), .ZN(
        n11728) );
  OAI21_X1 U14936 ( .B1(n11729), .B2(n11728), .A(n11727), .ZN(n11736) );
  NAND2_X1 U14937 ( .A1(n12904), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11735) );
  NAND2_X1 U14938 ( .A1(n12903), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11734) );
  NAND2_X1 U14939 ( .A1(n11730), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11732) );
  INV_X1 U14940 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11731) );
  XNOR2_X1 U14941 ( .A(n11732), .B(n11731), .ZN(n15300) );
  NAND2_X1 U14942 ( .A1(n15300), .A2(n11910), .ZN(n11733) );
  NAND4_X1 U14943 ( .A1(n11736), .A2(n11735), .A3(n11734), .A4(n11733), .ZN(
        n14944) );
  AOI22_X1 U14944 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11740) );
  AOI22_X1 U14945 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U14946 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12852), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U14947 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11737) );
  NAND4_X1 U14948 ( .A1(n11740), .A2(n11739), .A3(n11738), .A4(n11737), .ZN(
        n11746) );
  AOI22_X1 U14949 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11744) );
  AOI22_X1 U14950 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12876), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U14951 ( .A1(n12857), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11742) );
  AOI22_X1 U14952 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11741) );
  NAND4_X1 U14953 ( .A1(n11744), .A2(n11743), .A3(n11742), .A4(n11741), .ZN(
        n11745) );
  NOR2_X1 U14954 ( .A1(n11746), .A2(n11745), .ZN(n11752) );
  NAND2_X1 U14955 ( .A1(n12904), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11750) );
  INV_X1 U14956 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11747) );
  XNOR2_X1 U14957 ( .A(n11748), .B(n11747), .ZN(n15304) );
  AOI22_X1 U14958 ( .A1(n15304), .A2(n11910), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12903), .ZN(n11749) );
  OAI211_X1 U14959 ( .C1(n11752), .C2(n11751), .A(n11750), .B(n11749), .ZN(
        n14962) );
  NAND2_X1 U14960 ( .A1(n14944), .A2(n14962), .ZN(n14913) );
  AOI22_X1 U14961 ( .A1(n11411), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14962 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U14963 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U14964 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12852), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11755) );
  NAND4_X1 U14965 ( .A1(n11758), .A2(n11757), .A3(n11756), .A4(n11755), .ZN(
        n11765) );
  AOI22_X1 U14966 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11759), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U14967 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U14968 ( .A1(n12857), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11761) );
  AOI22_X1 U14969 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11760) );
  NAND4_X1 U14970 ( .A1(n11763), .A2(n11762), .A3(n11761), .A4(n11760), .ZN(
        n11764) );
  NOR2_X1 U14971 ( .A1(n11765), .A2(n11764), .ZN(n11768) );
  AOI21_X1 U14972 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15267), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11766) );
  AOI21_X1 U14973 ( .B1(n12904), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11766), .ZN(
        n11767) );
  OAI21_X1 U14974 ( .B1(n12868), .B2(n11768), .A(n11767), .ZN(n11770) );
  XNOR2_X1 U14975 ( .A(n11772), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15265) );
  NAND2_X1 U14976 ( .A1(n15265), .A2(n11910), .ZN(n11769) );
  NAND2_X1 U14977 ( .A1(n11770), .A2(n11769), .ZN(n14900) );
  INV_X1 U14978 ( .A(n14900), .ZN(n11771) );
  OR2_X1 U14979 ( .A1(n11772), .A2(n15267), .ZN(n11773) );
  XNOR2_X1 U14980 ( .A(n11773), .B(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15255) );
  AOI22_X1 U14981 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11450), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U14982 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U14983 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11789), .B1(
        n12852), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U14984 ( .A1(n12880), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11774) );
  NAND4_X1 U14985 ( .A1(n11777), .A2(n11776), .A3(n11775), .A4(n11774), .ZN(
        n11783) );
  AOI22_X1 U14986 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n11425), .B1(
        n11859), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14987 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11431), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U14988 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U14989 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12885), .B1(
        n12857), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11778) );
  NAND4_X1 U14990 ( .A1(n11781), .A2(n11780), .A3(n11779), .A4(n11778), .ZN(
        n11782) );
  OR2_X1 U14991 ( .A1(n11783), .A2(n11782), .ZN(n11784) );
  NAND2_X1 U14992 ( .A1(n12896), .A2(n11784), .ZN(n11788) );
  INV_X1 U14993 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n15126) );
  OAI22_X1 U14994 ( .A1(n12900), .A2(n15126), .B1(n15251), .B2(n11785), .ZN(
        n11786) );
  INV_X1 U14995 ( .A(n11786), .ZN(n11787) );
  OAI211_X1 U14996 ( .C1(n15255), .C2(n12902), .A(n11788), .B(n11787), .ZN(
        n14886) );
  INV_X1 U14997 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11851) );
  XNOR2_X1 U14998 ( .A(n11852), .B(n11851), .ZN(n15239) );
  AOI22_X1 U14999 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11859), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U15000 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U15001 ( .A1(n11808), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U15002 ( .A1(n12857), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11790) );
  NAND4_X1 U15003 ( .A1(n11793), .A2(n11792), .A3(n11791), .A4(n11790), .ZN(
        n11799) );
  AOI22_X1 U15004 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U15005 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12876), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11796) );
  AOI22_X1 U15006 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11795) );
  AOI22_X1 U15007 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11794) );
  NAND4_X1 U15008 ( .A1(n11797), .A2(n11796), .A3(n11795), .A4(n11794), .ZN(
        n11798) );
  NOR2_X1 U15009 ( .A1(n11799), .A2(n11798), .ZN(n11802) );
  INV_X1 U15010 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13559) );
  OAI22_X1 U15011 ( .A1(n12900), .A2(n13559), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n11851), .ZN(n11800) );
  INV_X1 U15012 ( .A(n11800), .ZN(n11801) );
  OAI21_X1 U15013 ( .B1(n12868), .B2(n11802), .A(n11801), .ZN(n11803) );
  MUX2_X1 U15014 ( .A(n15239), .B(n11803), .S(n12902), .Z(n14873) );
  INV_X1 U15015 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14817) );
  XNOR2_X1 U15016 ( .A(n11832), .B(n14817), .ZN(n15216) );
  AOI22_X1 U15017 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12887), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U15018 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11806) );
  AOI22_X1 U15019 ( .A1(n11411), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11805) );
  AOI22_X1 U15020 ( .A1(n12886), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12857), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11804) );
  NAND4_X1 U15021 ( .A1(n11807), .A2(n11806), .A3(n11805), .A4(n11804), .ZN(
        n11814) );
  AOI22_X1 U15022 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U15023 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U15024 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U15025 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11809) );
  NAND4_X1 U15026 ( .A1(n11812), .A2(n11811), .A3(n11810), .A4(n11809), .ZN(
        n11813) );
  NOR2_X1 U15027 ( .A1(n11814), .A2(n11813), .ZN(n11817) );
  INV_X1 U15028 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n15104) );
  OAI22_X1 U15029 ( .A1(n12900), .A2(n15104), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14817), .ZN(n11815) );
  INV_X1 U15030 ( .A(n11815), .ZN(n11816) );
  OAI21_X1 U15031 ( .B1(n12868), .B2(n11817), .A(n11816), .ZN(n11818) );
  MUX2_X1 U15032 ( .A(n15216), .B(n11818), .S(n12902), .Z(n14807) );
  AOI22_X1 U15033 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11822) );
  AOI22_X1 U15034 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U15035 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12876), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11820) );
  AOI22_X1 U15036 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12857), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11819) );
  NAND4_X1 U15037 ( .A1(n11822), .A2(n11821), .A3(n11820), .A4(n11819), .ZN(
        n11828) );
  AOI22_X1 U15038 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11759), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U15039 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12852), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U15040 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U15041 ( .A1(n12880), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11823) );
  NAND4_X1 U15042 ( .A1(n11826), .A2(n11825), .A3(n11824), .A4(n11823), .ZN(
        n11827) );
  OR2_X1 U15043 ( .A1(n11828), .A2(n11827), .ZN(n11830) );
  INV_X1 U15044 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n15108) );
  OAI22_X1 U15045 ( .A1(n12900), .A2(n15108), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12710), .ZN(n11829) );
  AOI21_X1 U15046 ( .B1(n12896), .B2(n11830), .A(n11829), .ZN(n11833) );
  NAND2_X1 U15047 ( .A1(n11848), .A2(n12710), .ZN(n11831) );
  AND2_X1 U15048 ( .A1(n11832), .A2(n11831), .ZN(n14825) );
  MUX2_X1 U15049 ( .A(n11833), .B(n14825), .S(n11910), .Z(n12705) );
  AOI22_X1 U15050 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U15051 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U15052 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U15053 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12852), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11834) );
  NAND4_X1 U15054 ( .A1(n11837), .A2(n11836), .A3(n11835), .A4(n11834), .ZN(
        n11843) );
  AOI22_X1 U15055 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11841) );
  AOI22_X1 U15056 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U15057 ( .A1(n12857), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U15058 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11838) );
  NAND4_X1 U15059 ( .A1(n11841), .A2(n11840), .A3(n11839), .A4(n11838), .ZN(
        n11842) );
  NOR2_X1 U15060 ( .A1(n11843), .A2(n11842), .ZN(n11846) );
  INV_X1 U15061 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n21510) );
  AOI21_X1 U15062 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n21510), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11844) );
  AOI21_X1 U15063 ( .B1(n12904), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11844), .ZN(
        n11845) );
  OAI21_X1 U15064 ( .B1(n12868), .B2(n11846), .A(n11845), .ZN(n11850) );
  NAND2_X1 U15065 ( .A1(n11854), .A2(n21510), .ZN(n11847) );
  NAND2_X1 U15066 ( .A1(n11848), .A2(n11847), .ZN(n15227) );
  OR2_X1 U15067 ( .A1(n15227), .A2(n12902), .ZN(n11849) );
  NAND2_X1 U15068 ( .A1(n11850), .A2(n11849), .ZN(n14834) );
  INV_X1 U15069 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15235) );
  OAI21_X1 U15070 ( .B1(n11852), .B2(n11851), .A(n15235), .ZN(n11853) );
  AND2_X1 U15071 ( .A1(n11854), .A2(n11853), .ZN(n15233) );
  AOI22_X1 U15072 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11858) );
  AOI22_X1 U15073 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11857) );
  AOI22_X1 U15074 ( .A1(n11425), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U15075 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12857), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11855) );
  NAND4_X1 U15076 ( .A1(n11858), .A2(n11857), .A3(n11856), .A4(n11855), .ZN(
        n11865) );
  AOI22_X1 U15077 ( .A1(n11450), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11863) );
  AOI22_X1 U15078 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11862) );
  AOI22_X1 U15079 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U15080 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11860) );
  NAND4_X1 U15081 ( .A1(n11863), .A2(n11862), .A3(n11861), .A4(n11860), .ZN(
        n11864) );
  OR2_X1 U15082 ( .A1(n11865), .A2(n11864), .ZN(n11867) );
  INV_X1 U15083 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n15117) );
  OAI22_X1 U15084 ( .A1(n12900), .A2(n15117), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15235), .ZN(n11866) );
  AOI21_X1 U15085 ( .B1(n12896), .B2(n11867), .A(n11866), .ZN(n11868) );
  MUX2_X1 U15086 ( .A(n15233), .B(n11868), .S(n12902), .Z(n14852) );
  NOR2_X1 U15087 ( .A1(n12705), .A2(n12702), .ZN(n12703) );
  XNOR2_X1 U15088 ( .A(n11871), .B(n11870), .ZN(n11874) );
  INV_X1 U15089 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n15099) );
  OAI22_X1 U15090 ( .A1(n12900), .A2(n15099), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14800), .ZN(n11872) );
  INV_X1 U15091 ( .A(n11872), .ZN(n11873) );
  OAI21_X1 U15092 ( .B1(n12868), .B2(n11874), .A(n11873), .ZN(n11877) );
  NAND2_X1 U15093 ( .A1(n11875), .A2(n14800), .ZN(n11876) );
  NAND2_X1 U15094 ( .A1(n11879), .A2(n11876), .ZN(n15212) );
  MUX2_X1 U15095 ( .A(n11877), .B(n15212), .S(n11910), .Z(n11878) );
  XNOR2_X1 U15096 ( .A(n11879), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15203) );
  NAND2_X1 U15097 ( .A1(n15203), .A2(n11910), .ZN(n11886) );
  XNOR2_X1 U15098 ( .A(n11881), .B(n11880), .ZN(n11884) );
  NAND2_X1 U15099 ( .A1(n12904), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n11883) );
  OAI21_X1 U15100 ( .B1(n21191), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n21239), .ZN(n11882) );
  OAI211_X1 U15101 ( .C1(n11884), .C2(n12868), .A(n11883), .B(n11882), .ZN(
        n11885) );
  XNOR2_X1 U15102 ( .A(n11889), .B(n11888), .ZN(n11892) );
  INV_X1 U15103 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n15091) );
  OAI22_X1 U15104 ( .A1(n12900), .A2(n15091), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n11893), .ZN(n11890) );
  INV_X1 U15105 ( .A(n11890), .ZN(n11891) );
  OAI21_X1 U15106 ( .B1(n11892), .B2(n12868), .A(n11891), .ZN(n11896) );
  NAND2_X1 U15107 ( .A1(n11894), .A2(n11893), .ZN(n11895) );
  NAND2_X1 U15108 ( .A1(n11901), .A2(n11895), .ZN(n15193) );
  MUX2_X1 U15109 ( .A(n11896), .B(n15193), .S(n11910), .Z(n14770) );
  XOR2_X1 U15110 ( .A(n11898), .B(n11897), .Z(n11900) );
  INV_X1 U15111 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n15086) );
  OAI22_X1 U15112 ( .A1(n12900), .A2(n15086), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15189), .ZN(n11899) );
  AOI21_X1 U15113 ( .B1(n11900), .B2(n12896), .A(n11899), .ZN(n11903) );
  INV_X1 U15114 ( .A(n11901), .ZN(n11902) );
  XOR2_X1 U15115 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B(n11902), .Z(
        n15187) );
  MUX2_X1 U15116 ( .A(n11903), .B(n15187), .S(n11910), .Z(n14758) );
  XNOR2_X1 U15117 ( .A(n11905), .B(n11904), .ZN(n11908) );
  INV_X1 U15118 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n15082) );
  INV_X1 U15119 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14749) );
  OAI22_X1 U15120 ( .A1(n12900), .A2(n15082), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14749), .ZN(n11906) );
  INV_X1 U15121 ( .A(n11906), .ZN(n11907) );
  OAI21_X1 U15122 ( .B1(n11908), .B2(n12868), .A(n11907), .ZN(n11911) );
  OAI21_X1 U15123 ( .B1(n11909), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n11916), .ZN(n15174) );
  MUX2_X1 U15124 ( .A(n11911), .B(n15174), .S(n11910), .Z(n14744) );
  AOI21_X1 U15125 ( .B1(n11915), .B2(n11912), .A(n11914), .ZN(n15171) );
  INV_X1 U15126 ( .A(n15171), .ZN(n15081) );
  OR2_X2 U15127 ( .A1(n11916), .A2(n15169), .ZN(n12850) );
  INV_X1 U15128 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14734) );
  OR2_X2 U15129 ( .A1(n12850), .A2(n14734), .ZN(n12872) );
  INV_X1 U15130 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14370) );
  NOR2_X2 U15131 ( .A1(n12872), .A2(n14370), .ZN(n11917) );
  AND2_X1 U15132 ( .A1(n10177), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11918) );
  NOR2_X1 U15133 ( .A1(n11936), .A2(n11918), .ZN(n11920) );
  NAND2_X1 U15134 ( .A1(n20752), .A2(n11993), .ZN(n11919) );
  NAND2_X1 U15135 ( .A1(n11919), .A2(n20733), .ZN(n11941) );
  OAI211_X1 U15136 ( .C1(n12220), .C2(n20715), .A(n11941), .B(n11920), .ZN(
        n11921) );
  NAND2_X1 U15137 ( .A1(n11922), .A2(n11921), .ZN(n11929) );
  MUX2_X1 U15138 ( .A(n13998), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11937) );
  XNOR2_X1 U15139 ( .A(n11937), .B(n11936), .ZN(n11982) );
  NAND2_X1 U15140 ( .A1(n20752), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11925) );
  NAND2_X1 U15141 ( .A1(n11976), .A2(n14053), .ZN(n11923) );
  NAND2_X1 U15142 ( .A1(n11929), .A2(n11930), .ZN(n11928) );
  INV_X1 U15143 ( .A(n11976), .ZN(n11926) );
  NAND3_X1 U15144 ( .A1(n11926), .A2(n14053), .A3(n11925), .ZN(n11960) );
  NAND2_X1 U15145 ( .A1(n11960), .A2(n11982), .ZN(n11927) );
  NAND2_X1 U15146 ( .A1(n11928), .A2(n11927), .ZN(n11934) );
  INV_X1 U15147 ( .A(n11929), .ZN(n11932) );
  INV_X1 U15148 ( .A(n11930), .ZN(n11931) );
  NAND2_X1 U15149 ( .A1(n11932), .A2(n11931), .ZN(n11933) );
  NAND2_X1 U15150 ( .A1(n11934), .A2(n11933), .ZN(n11940) );
  NOR2_X1 U15151 ( .A1(n11465), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11935) );
  XNOR2_X1 U15152 ( .A(n13979), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11945) );
  XNOR2_X1 U15153 ( .A(n11944), .B(n11945), .ZN(n11983) );
  INV_X1 U15154 ( .A(n11983), .ZN(n11942) );
  NAND2_X1 U15155 ( .A1(n11976), .A2(n11942), .ZN(n11938) );
  OAI211_X1 U15156 ( .C1(n11942), .C2(n11958), .A(n11938), .B(n11941), .ZN(
        n11939) );
  NAND2_X1 U15157 ( .A1(n11940), .A2(n11939), .ZN(n11952) );
  INV_X1 U15158 ( .A(n11941), .ZN(n11943) );
  NAND3_X1 U15159 ( .A1(n11943), .A2(n11976), .A3(n11942), .ZN(n11951) );
  INV_X1 U15160 ( .A(n11944), .ZN(n11947) );
  INV_X1 U15161 ( .A(n11945), .ZN(n11946) );
  NAND2_X1 U15162 ( .A1(n11947), .A2(n11946), .ZN(n11949) );
  NAND2_X1 U15163 ( .A1(n21123), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11948) );
  XNOR2_X1 U15164 ( .A(n11957), .B(n11956), .ZN(n11984) );
  AND2_X1 U15165 ( .A1(n11958), .A2(n11984), .ZN(n11950) );
  INV_X1 U15166 ( .A(n11984), .ZN(n11953) );
  NOR2_X1 U15167 ( .A1(n11966), .A2(n11953), .ZN(n11954) );
  NOR2_X1 U15168 ( .A1(n14025), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11955) );
  AND2_X1 U15169 ( .A1(n11967), .A2(n11970), .ZN(n11985) );
  NAND2_X1 U15170 ( .A1(n11985), .A2(n11958), .ZN(n11959) );
  INV_X1 U15171 ( .A(n11960), .ZN(n11962) );
  NAND3_X1 U15172 ( .A1(n11962), .A2(n11961), .A3(n11985), .ZN(n11964) );
  NAND2_X1 U15173 ( .A1(n10072), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11963) );
  INV_X1 U15174 ( .A(n11966), .ZN(n11973) );
  INV_X1 U15175 ( .A(n11967), .ZN(n11969) );
  NOR2_X1 U15176 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n14039), .ZN(
        n11968) );
  INV_X1 U15177 ( .A(n11970), .ZN(n11971) );
  NAND2_X1 U15178 ( .A1(n11973), .A2(n11981), .ZN(n11974) );
  NAND2_X1 U15179 ( .A1(n12232), .A2(n20715), .ZN(n11980) );
  INV_X1 U15180 ( .A(n11981), .ZN(n11987) );
  OR4_X1 U15181 ( .A1(n11985), .A2(n11984), .A3(n11983), .A4(n11982), .ZN(
        n11986) );
  NAND2_X1 U15182 ( .A1(n11987), .A2(n11986), .ZN(n12971) );
  INV_X1 U15183 ( .A(n12971), .ZN(n11988) );
  NAND2_X1 U15184 ( .A1(n12972), .A2(n11988), .ZN(n12960) );
  OR2_X2 U15185 ( .A1(n21377), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20667) );
  INV_X2 U15186 ( .A(n20667), .ZN(n20683) );
  NOR2_X1 U15187 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21384) );
  AND2_X1 U15188 ( .A1(n21384), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14222) );
  NOR2_X1 U15189 ( .A1(n12902), .A2(n14650), .ZN(n11989) );
  MUX2_X1 U15190 ( .A(n14222), .B(n11989), .S(n10072), .Z(n11990) );
  NOR2_X1 U15191 ( .A1(n20683), .A2(n11990), .ZN(n11991) );
  NAND2_X1 U15192 ( .A1(n20742), .A2(n11993), .ZN(n12012) );
  AND2_X4 U15193 ( .A1(n9576), .A2(n11993), .ZN(n12726) );
  NAND2_X2 U15194 ( .A1(n11995), .A2(n12726), .ZN(n12085) );
  NAND2_X1 U15195 ( .A1(n12782), .A2(n13625), .ZN(n11996) );
  INV_X1 U15196 ( .A(n12012), .ZN(n12004) );
  NAND2_X1 U15197 ( .A1(n12004), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11999) );
  INV_X1 U15198 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n21464) );
  NAND2_X1 U15199 ( .A1(n12782), .A2(n21464), .ZN(n11998) );
  NAND2_X1 U15200 ( .A1(n11999), .A2(n11998), .ZN(n13242) );
  XNOR2_X1 U15201 ( .A(n12000), .B(n13242), .ZN(n13624) );
  NAND2_X1 U15202 ( .A1(n13624), .A2(n12726), .ZN(n12002) );
  INV_X1 U15203 ( .A(n12000), .ZN(n12001) );
  NAND2_X1 U15204 ( .A1(n12002), .A2(n12001), .ZN(n13891) );
  INV_X1 U15205 ( .A(n12782), .ZN(n12013) );
  MUX2_X1 U15206 ( .A(n12085), .B(n12013), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n12003) );
  OAI21_X1 U15207 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n13240), .A(
        n12003), .ZN(n13890) );
  OR2_X1 U15208 ( .A1(n12729), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n12008) );
  INV_X1 U15209 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20673) );
  NAND2_X1 U15210 ( .A1(n12080), .A2(n20673), .ZN(n12006) );
  INV_X1 U15211 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n14076) );
  NAND2_X1 U15212 ( .A1(n12726), .A2(n14076), .ZN(n12005) );
  NAND3_X1 U15213 ( .A1(n12006), .A2(n12013), .A3(n12005), .ZN(n12007) );
  NAND2_X1 U15214 ( .A1(n12008), .A2(n12007), .ZN(n14074) );
  INV_X1 U15215 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n20598) );
  NAND2_X1 U15216 ( .A1(n12060), .A2(n20598), .ZN(n12011) );
  NAND2_X1 U15217 ( .A1(n12013), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12009) );
  OAI211_X1 U15218 ( .C1(n13625), .C2(P1_EBX_REG_4__SCAN_IN), .A(n12080), .B(
        n12009), .ZN(n12010) );
  AND2_X1 U15219 ( .A1(n12011), .A2(n12010), .ZN(n20550) );
  OR2_X1 U15220 ( .A1(n12729), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n12017) );
  NAND2_X1 U15221 ( .A1(n12013), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12014) );
  NAND2_X1 U15222 ( .A1(n12080), .A2(n12014), .ZN(n12015) );
  OAI21_X1 U15223 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(n13625), .A(n12015), .ZN(
        n12016) );
  INV_X1 U15224 ( .A(n12782), .ZN(n12084) );
  NAND2_X1 U15225 ( .A1(n12084), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12018) );
  OAI211_X1 U15226 ( .C1(n13625), .C2(P1_EBX_REG_6__SCAN_IN), .A(n12080), .B(
        n12018), .ZN(n12019) );
  OAI21_X1 U15227 ( .B1(n12085), .B2(P1_EBX_REG_6__SCAN_IN), .A(n12019), .ZN(
        n17396) );
  OR2_X1 U15228 ( .A1(n12729), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n12023) );
  NAND2_X1 U15229 ( .A1(n12084), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12020) );
  NAND2_X1 U15230 ( .A1(n12080), .A2(n12020), .ZN(n12021) );
  OAI21_X1 U15231 ( .B1(P1_EBX_REG_7__SCAN_IN), .B2(n13625), .A(n12021), .ZN(
        n12022) );
  NAND2_X1 U15232 ( .A1(n12023), .A2(n12022), .ZN(n14247) );
  INV_X1 U15233 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14996) );
  NAND2_X1 U15234 ( .A1(n12060), .A2(n14996), .ZN(n12026) );
  NAND2_X1 U15235 ( .A1(n12013), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12024) );
  OAI211_X1 U15236 ( .C1(n13625), .C2(P1_EBX_REG_8__SCAN_IN), .A(n12080), .B(
        n12024), .ZN(n12025) );
  NAND2_X1 U15237 ( .A1(n14245), .A2(n14993), .ZN(n14992) );
  INV_X2 U15238 ( .A(n14992), .ZN(n12032) );
  OR2_X1 U15239 ( .A1(n12729), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n12030) );
  NAND2_X1 U15240 ( .A1(n12084), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12027) );
  NAND2_X1 U15241 ( .A1(n12080), .A2(n12027), .ZN(n12028) );
  OAI21_X1 U15242 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(n13625), .A(n12028), .ZN(
        n12029) );
  MUX2_X1 U15243 ( .A(n12085), .B(n12013), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n12033) );
  OAI21_X1 U15244 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n13240), .A(
        n12033), .ZN(n15052) );
  INV_X1 U15245 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15045) );
  NAND2_X1 U15246 ( .A1(n12060), .A2(n15045), .ZN(n12037) );
  NAND2_X1 U15247 ( .A1(n12084), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12035) );
  OAI211_X1 U15248 ( .C1(n13625), .C2(P1_EBX_REG_12__SCAN_IN), .A(n12080), .B(
        n12035), .ZN(n12036) );
  OR2_X1 U15249 ( .A1(n12729), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n12040) );
  INV_X1 U15250 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21437) );
  NAND2_X1 U15251 ( .A1(n12080), .A2(n21437), .ZN(n12038) );
  OAI211_X1 U15252 ( .C1(P1_EBX_REG_11__SCAN_IN), .C2(n13625), .A(n12038), .B(
        n12084), .ZN(n12039) );
  NAND2_X1 U15253 ( .A1(n12040), .A2(n12039), .ZN(n14979) );
  OR2_X1 U15254 ( .A1(n12729), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n12043) );
  INV_X1 U15255 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12185) );
  NAND2_X1 U15256 ( .A1(n12080), .A2(n12185), .ZN(n12041) );
  OAI211_X1 U15257 ( .C1(P1_EBX_REG_13__SCAN_IN), .C2(n13625), .A(n12041), .B(
        n12013), .ZN(n12042) );
  NAND2_X1 U15258 ( .A1(n12043), .A2(n12042), .ZN(n14952) );
  MUX2_X1 U15259 ( .A(n12085), .B(n12013), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12044) );
  OAI21_X1 U15260 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n13240), .A(
        n12044), .ZN(n14935) );
  OR2_X1 U15261 ( .A1(n12729), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n12048) );
  INV_X1 U15262 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21481) );
  NAND2_X1 U15263 ( .A1(n12080), .A2(n21481), .ZN(n12046) );
  OAI211_X1 U15264 ( .C1(P1_EBX_REG_15__SCAN_IN), .C2(n13625), .A(n12046), .B(
        n12084), .ZN(n12047) );
  INV_X1 U15265 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15041) );
  NAND2_X1 U15266 ( .A1(n12060), .A2(n15041), .ZN(n12051) );
  NAND2_X1 U15267 ( .A1(n12084), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12049) );
  OAI211_X1 U15268 ( .C1(n13625), .C2(P1_EBX_REG_16__SCAN_IN), .A(n12080), .B(
        n12049), .ZN(n12050) );
  OR2_X1 U15269 ( .A1(n12729), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n12054) );
  INV_X1 U15270 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12193) );
  NAND2_X1 U15271 ( .A1(n12080), .A2(n12193), .ZN(n12052) );
  OAI211_X1 U15272 ( .C1(P1_EBX_REG_17__SCAN_IN), .C2(n13625), .A(n12052), .B(
        n12084), .ZN(n12053) );
  NAND2_X1 U15273 ( .A1(n12054), .A2(n12053), .ZN(n14888) );
  MUX2_X1 U15274 ( .A(n12085), .B(n12013), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n12055) );
  OAI21_X1 U15275 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n13240), .A(
        n12055), .ZN(n14875) );
  OR2_X1 U15276 ( .A1(n12729), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n12058) );
  INV_X1 U15277 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15423) );
  NAND2_X1 U15278 ( .A1(n12080), .A2(n15423), .ZN(n12056) );
  OAI211_X1 U15279 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n13625), .A(n12056), .B(
        n12013), .ZN(n12057) );
  INV_X1 U15280 ( .A(n14855), .ZN(n12059) );
  AND2_X2 U15281 ( .A1(n14853), .A2(n12059), .ZN(n14854) );
  INV_X1 U15282 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15036) );
  NAND2_X1 U15283 ( .A1(n12060), .A2(n15036), .ZN(n12063) );
  NAND2_X1 U15284 ( .A1(n12084), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12061) );
  OAI211_X1 U15285 ( .C1(n13625), .C2(P1_EBX_REG_20__SCAN_IN), .A(n12080), .B(
        n12061), .ZN(n12062) );
  OR2_X1 U15286 ( .A1(n12729), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n12066) );
  NAND2_X1 U15287 ( .A1(n12080), .A2(n12201), .ZN(n12064) );
  OAI211_X1 U15288 ( .C1(P1_EBX_REG_21__SCAN_IN), .C2(n13625), .A(n12064), .B(
        n12013), .ZN(n12065) );
  NAND2_X1 U15289 ( .A1(n12066), .A2(n12065), .ZN(n12770) );
  MUX2_X1 U15290 ( .A(n12085), .B(n12013), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n12067) );
  OAI21_X1 U15291 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n13240), .A(
        n12067), .ZN(n14811) );
  OR2_X1 U15292 ( .A1(n12729), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n12072) );
  INV_X1 U15293 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15394) );
  NAND2_X1 U15294 ( .A1(n12080), .A2(n15394), .ZN(n12070) );
  OAI211_X1 U15295 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n13625), .A(n12070), .B(
        n12084), .ZN(n12071) );
  MUX2_X1 U15296 ( .A(n12085), .B(n12084), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n12073) );
  OAI21_X1 U15297 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n13240), .A(
        n12073), .ZN(n14788) );
  NOR2_X4 U15298 ( .A1(n14795), .A2(n14788), .ZN(n14787) );
  OR2_X1 U15299 ( .A1(n12729), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n12077) );
  NAND2_X1 U15300 ( .A1(n12084), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12074) );
  NAND2_X1 U15301 ( .A1(n12080), .A2(n12074), .ZN(n12075) );
  OAI21_X1 U15302 ( .B1(P1_EBX_REG_25__SCAN_IN), .B2(n13625), .A(n12075), .ZN(
        n12076) );
  NAND2_X1 U15303 ( .A1(n12077), .A2(n12076), .ZN(n12915) );
  NAND2_X1 U15304 ( .A1(n12084), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12078) );
  OAI211_X1 U15305 ( .C1(n13625), .C2(P1_EBX_REG_26__SCAN_IN), .A(n12080), .B(
        n12078), .ZN(n12079) );
  OAI21_X1 U15306 ( .B1(n12085), .B2(P1_EBX_REG_26__SCAN_IN), .A(n12079), .ZN(
        n14759) );
  OR2_X1 U15307 ( .A1(n12729), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n12083) );
  INV_X1 U15308 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12266) );
  NAND2_X1 U15309 ( .A1(n12080), .A2(n12266), .ZN(n12081) );
  OAI211_X1 U15310 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n13625), .A(n12081), .B(
        n12084), .ZN(n12082) );
  MUX2_X1 U15311 ( .A(n12085), .B(n12084), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n12087) );
  OR2_X1 U15312 ( .A1(n13240), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12086) );
  AND2_X1 U15313 ( .A1(n12087), .A2(n12086), .ZN(n12088) );
  NOR2_X1 U15314 ( .A1(n14745), .A2(n12088), .ZN(n12089) );
  OR2_X1 U15315 ( .A1(n21382), .A2(n20715), .ZN(n12095) );
  AND2_X1 U15316 ( .A1(n9576), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12093) );
  NAND2_X1 U15317 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21308) );
  NAND2_X1 U15318 ( .A1(n21308), .A2(n21191), .ZN(n14050) );
  NAND2_X1 U15319 ( .A1(n12093), .A2(n14050), .ZN(n12090) );
  NOR2_X1 U15320 ( .A1(n14339), .A2(n20589), .ZN(n12106) );
  AND2_X1 U15321 ( .A1(n14053), .A2(n21308), .ZN(n13294) );
  INV_X1 U15322 ( .A(n13294), .ZN(n12092) );
  NAND2_X1 U15323 ( .A1(n12091), .A2(n21312), .ZN(n14051) );
  OR2_X1 U15324 ( .A1(n14051), .A2(n21379), .ZN(n13295) );
  NAND2_X1 U15325 ( .A1(n12092), .A2(n13295), .ZN(n12209) );
  AND2_X1 U15326 ( .A1(n12209), .A2(n21191), .ZN(n12096) );
  OR2_X1 U15327 ( .A1(n12096), .A2(n12093), .ZN(n12094) );
  INV_X1 U15328 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14340) );
  AOI22_X1 U15329 ( .A1(n20575), .A2(n15166), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20579), .ZN(n12101) );
  INV_X1 U15330 ( .A(n12095), .ZN(n12097) );
  INV_X1 U15331 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21344) );
  INV_X1 U15332 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21340) );
  INV_X1 U15333 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21330) );
  NAND4_X1 U15334 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n14947)
         );
  INV_X1 U15335 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n14988) );
  NAND2_X1 U15336 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14980) );
  INV_X1 U15337 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21328) );
  NOR3_X1 U15338 ( .A1(n14988), .A2(n14980), .A3(n21328), .ZN(n14956) );
  NAND2_X1 U15339 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n14956), .ZN(n14842) );
  NOR3_X1 U15340 ( .A1(n21330), .A2(n14947), .A3(n14842), .ZN(n14858) );
  AND2_X1 U15341 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14862) );
  AND2_X1 U15342 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n14857) );
  AND2_X1 U15343 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n12098) );
  AND3_X1 U15344 ( .A1(n14862), .A2(n14857), .A3(n12098), .ZN(n14814) );
  NAND4_X1 U15345 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_4__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n14840)
         );
  INV_X1 U15346 ( .A(n14840), .ZN(n14813) );
  AND3_X1 U15347 ( .A1(n14858), .A2(n14814), .A3(n14813), .ZN(n14827) );
  NAND2_X1 U15348 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n14827), .ZN(n14819) );
  NOR2_X1 U15349 ( .A1(n21340), .A2(n14819), .ZN(n14799) );
  NAND2_X1 U15350 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n14799), .ZN(n14771) );
  NOR2_X1 U15351 ( .A1(n21344), .A2(n14771), .ZN(n14774) );
  AND2_X1 U15352 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n14774), .ZN(n14762) );
  AND2_X1 U15353 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n14762), .ZN(n14747) );
  NAND2_X1 U15354 ( .A1(n14747), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n12102) );
  NOR2_X1 U15355 ( .A1(n12102), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n12099) );
  NAND2_X1 U15356 ( .A1(n20555), .A2(n12099), .ZN(n12100) );
  OAI211_X1 U15357 ( .C1(n20553), .C2(n14340), .A(n12101), .B(n12100), .ZN(
        n12104) );
  INV_X1 U15358 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21349) );
  NOR2_X1 U15359 ( .A1(n21349), .A2(n12102), .ZN(n14371) );
  INV_X1 U15360 ( .A(n20517), .ZN(n14856) );
  AOI21_X1 U15361 ( .B1(n14371), .B2(n20562), .A(n14856), .ZN(n14733) );
  INV_X1 U15362 ( .A(n13462), .ZN(n12134) );
  NAND2_X1 U15363 ( .A1(n12116), .A2(n12123), .ZN(n12136) );
  NAND2_X1 U15364 ( .A1(n12136), .A2(n12135), .ZN(n12152) );
  XNOR2_X1 U15365 ( .A(n12152), .B(n12149), .ZN(n12109) );
  NAND3_X1 U15366 ( .A1(n12143), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12147) );
  NAND2_X1 U15367 ( .A1(n12110), .A2(n13462), .ZN(n12114) );
  NAND2_X1 U15368 ( .A1(n12152), .A2(n12149), .ZN(n12111) );
  XNOR2_X1 U15369 ( .A(n12111), .B(n12150), .ZN(n12112) );
  NAND2_X1 U15370 ( .A1(n12112), .A2(n12979), .ZN(n12113) );
  NAND2_X1 U15371 ( .A1(n12114), .A2(n12113), .ZN(n20645) );
  NAND2_X1 U15372 ( .A1(n12115), .A2(n14053), .ZN(n12121) );
  XNOR2_X1 U15373 ( .A(n12116), .B(n12123), .ZN(n12118) );
  INV_X1 U15374 ( .A(n12117), .ZN(n12229) );
  OAI211_X1 U15375 ( .C1(n12118), .C2(n12108), .A(n12117), .B(n11391), .ZN(
        n12119) );
  INV_X1 U15376 ( .A(n12119), .ZN(n12120) );
  NAND2_X1 U15377 ( .A1(n12121), .A2(n12120), .ZN(n12132) );
  OR2_X1 U15378 ( .A1(n12108), .A2(n12123), .ZN(n13460) );
  NAND2_X1 U15379 ( .A1(n20715), .A2(n12124), .ZN(n13459) );
  NAND2_X1 U15380 ( .A1(n13460), .A2(n13459), .ZN(n12125) );
  INV_X1 U15381 ( .A(n12125), .ZN(n12127) );
  NAND2_X1 U15382 ( .A1(n10183), .A2(n12127), .ZN(n12130) );
  OR2_X1 U15383 ( .A1(n12126), .A2(n12125), .ZN(n12129) );
  INV_X1 U15384 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13458) );
  AOI21_X1 U15385 ( .B1(n12127), .B2(n12134), .A(n13458), .ZN(n12128) );
  OAI211_X1 U15386 ( .C1(n11584), .C2(n12130), .A(n12129), .B(n12128), .ZN(
        n12131) );
  XNOR2_X1 U15387 ( .A(n12132), .B(n12131), .ZN(n13722) );
  NAND2_X1 U15388 ( .A1(n13722), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13723) );
  INV_X1 U15389 ( .A(n12131), .ZN(n13463) );
  NAND2_X1 U15390 ( .A1(n12132), .A2(n13463), .ZN(n12133) );
  NAND2_X1 U15391 ( .A1(n13723), .A2(n12133), .ZN(n12141) );
  INV_X1 U15392 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20690) );
  XNOR2_X1 U15393 ( .A(n12141), .B(n20690), .ZN(n13837) );
  XNOR2_X1 U15394 ( .A(n12136), .B(n12135), .ZN(n12138) );
  INV_X1 U15395 ( .A(n13459), .ZN(n12137) );
  AOI21_X1 U15396 ( .B1(n12138), .B2(n12979), .A(n12137), .ZN(n12139) );
  NAND2_X1 U15397 ( .A1(n12141), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12142) );
  INV_X1 U15398 ( .A(n12144), .ZN(n12145) );
  NAND2_X1 U15399 ( .A1(n12145), .A2(n20645), .ZN(n12146) );
  AND2_X1 U15400 ( .A1(n12150), .A2(n12149), .ZN(n12151) );
  NAND2_X1 U15401 ( .A1(n12152), .A2(n12151), .ZN(n12158) );
  XNOR2_X1 U15402 ( .A(n12158), .B(n12159), .ZN(n12153) );
  NAND2_X1 U15403 ( .A1(n12153), .A2(n12979), .ZN(n12154) );
  INV_X1 U15404 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14201) );
  NAND2_X1 U15405 ( .A1(n12155), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12156) );
  NAND3_X1 U15406 ( .A1(n12176), .A2(n12157), .A3(n13462), .ZN(n12163) );
  INV_X1 U15407 ( .A(n12158), .ZN(n12160) );
  NAND2_X1 U15408 ( .A1(n12160), .A2(n12159), .ZN(n12166) );
  XNOR2_X1 U15409 ( .A(n12166), .B(n12167), .ZN(n12161) );
  NAND2_X1 U15410 ( .A1(n12161), .A2(n12979), .ZN(n12162) );
  NAND2_X1 U15411 ( .A1(n12163), .A2(n12162), .ZN(n17366) );
  NAND2_X1 U15412 ( .A1(n17366), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12164) );
  NAND2_X1 U15413 ( .A1(n12165), .A2(n13462), .ZN(n12172) );
  INV_X1 U15414 ( .A(n12166), .ZN(n12168) );
  NAND2_X1 U15415 ( .A1(n12168), .A2(n12167), .ZN(n12178) );
  XNOR2_X1 U15416 ( .A(n12178), .B(n12169), .ZN(n12170) );
  NAND2_X1 U15417 ( .A1(n12170), .A2(n12979), .ZN(n12171) );
  NAND2_X1 U15418 ( .A1(n12172), .A2(n12171), .ZN(n12173) );
  NAND2_X1 U15419 ( .A1(n12173), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17358) );
  AND2_X1 U15420 ( .A1(n12174), .A2(n13462), .ZN(n12175) );
  NAND2_X4 U15421 ( .A1(n12176), .A2(n12175), .ZN(n15332) );
  OR3_X1 U15422 ( .A1(n12178), .A2(n12177), .A3(n12108), .ZN(n12181) );
  INV_X1 U15423 ( .A(n12181), .ZN(n15312) );
  NAND2_X1 U15424 ( .A1(n15312), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12180) );
  NOR2_X1 U15425 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12179) );
  AOI21_X1 U15426 ( .B1(n15332), .B2(n12180), .A(n12179), .ZN(n12184) );
  INV_X1 U15427 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17388) );
  NAND2_X1 U15428 ( .A1(n12181), .A2(n17388), .ZN(n12182) );
  NAND2_X1 U15429 ( .A1(n12182), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12183) );
  NAND2_X1 U15430 ( .A1(n15332), .A2(n12185), .ZN(n12186) );
  INV_X1 U15431 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15499) );
  NAND2_X1 U15432 ( .A1(n15332), .A2(n15499), .ZN(n15296) );
  NAND2_X1 U15433 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12187) );
  NAND2_X1 U15434 ( .A1(n15332), .A2(n12187), .ZN(n15293) );
  NAND2_X1 U15435 ( .A1(n15296), .A2(n15293), .ZN(n12188) );
  INV_X1 U15436 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21509) );
  NAND2_X1 U15437 ( .A1(n15332), .A2(n21509), .ZN(n12189) );
  OR2_X1 U15438 ( .A1(n15332), .A2(n21509), .ZN(n12190) );
  NAND2_X1 U15439 ( .A1(n15284), .A2(n12190), .ZN(n15258) );
  XNOR2_X1 U15440 ( .A(n15332), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15264) );
  NAND2_X1 U15441 ( .A1(n15332), .A2(n21481), .ZN(n15262) );
  AND2_X1 U15442 ( .A1(n15264), .A2(n15262), .ZN(n12191) );
  NOR2_X1 U15443 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12192) );
  NAND2_X1 U15444 ( .A1(n15332), .A2(n12193), .ZN(n12194) );
  OR2_X1 U15445 ( .A1(n15332), .A2(n15499), .ZN(n15295) );
  NOR2_X1 U15446 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12196) );
  OR2_X1 U15447 ( .A1(n15332), .A2(n12196), .ZN(n15291) );
  NAND2_X1 U15448 ( .A1(n15295), .A2(n15291), .ZN(n15283) );
  NAND2_X1 U15449 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15412) );
  INV_X1 U15450 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12201) );
  INV_X1 U15451 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12200) );
  INV_X1 U15452 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15415) );
  NAND2_X1 U15453 ( .A1(n15423), .A2(n15415), .ZN(n15411) );
  INV_X1 U15454 ( .A(n15411), .ZN(n12199) );
  AND2_X1 U15455 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12264) );
  NAND2_X1 U15456 ( .A1(n12264), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12254) );
  NAND2_X1 U15457 ( .A1(n15332), .A2(n12254), .ZN(n15183) );
  NOR2_X1 U15458 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12717) );
  NAND2_X1 U15459 ( .A1(n12717), .A2(n15394), .ZN(n15182) );
  MUX2_X1 U15460 ( .A(n12266), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15332), .Z(n12202) );
  OAI211_X1 U15461 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n12204), .A(
        n12203), .B(n12202), .ZN(n12205) );
  INV_X1 U15462 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12265) );
  XNOR2_X1 U15463 ( .A(n12205), .B(n12265), .ZN(n15173) );
  INV_X1 U15464 ( .A(n12207), .ZN(n13292) );
  NAND2_X1 U15465 ( .A1(n14713), .A2(n11993), .ZN(n12208) );
  AOI21_X1 U15466 ( .B1(n13292), .B2(n12209), .A(n12208), .ZN(n12210) );
  NOR2_X1 U15467 ( .A1(n12971), .A2(n21379), .ZN(n13301) );
  NAND2_X1 U15468 ( .A1(n14053), .A2(n14051), .ZN(n12211) );
  NOR2_X1 U15469 ( .A1(n12212), .A2(n20733), .ZN(n12217) );
  INV_X1 U15470 ( .A(n12972), .ZN(n12216) );
  AOI21_X1 U15471 ( .B1(n12212), .B2(n20715), .A(n12229), .ZN(n12219) );
  NAND2_X1 U15472 ( .A1(n12219), .A2(n9666), .ZN(n12221) );
  INV_X1 U15473 ( .A(n12221), .ZN(n12214) );
  NAND2_X1 U15474 ( .A1(n13611), .A2(n9576), .ZN(n12237) );
  AND2_X1 U15475 ( .A1(n12237), .A2(n11993), .ZN(n12213) );
  NAND2_X1 U15476 ( .A1(n11398), .A2(n12213), .ZN(n12240) );
  NAND2_X1 U15477 ( .A1(n12214), .A2(n12240), .ZN(n12215) );
  AND2_X1 U15478 ( .A1(n12219), .A2(n12238), .ZN(n13293) );
  INV_X1 U15479 ( .A(n13293), .ZN(n13981) );
  OAI211_X1 U15480 ( .C1(n20747), .C2(n12227), .A(n13981), .B(n12969), .ZN(
        n12223) );
  OR2_X1 U15481 ( .A1(n12223), .A2(n12222), .ZN(n12224) );
  NAND2_X1 U15482 ( .A1(n14058), .A2(n20733), .ZN(n12226) );
  OAI21_X1 U15483 ( .B1(n12227), .B2(n11383), .A(n12226), .ZN(n12228) );
  NOR2_X1 U15484 ( .A1(n14339), .A2(n20668), .ZN(n12271) );
  NAND2_X1 U15485 ( .A1(n12229), .A2(n13240), .ZN(n12231) );
  OAI211_X1 U15486 ( .C1(n12232), .C2(n15004), .A(n12231), .B(n12230), .ZN(
        n12233) );
  INV_X1 U15487 ( .A(n12233), .ZN(n12236) );
  NAND2_X1 U15488 ( .A1(n12234), .A2(n14053), .ZN(n12235) );
  OAI211_X1 U15489 ( .C1(n9666), .C2(n12013), .A(n12236), .B(n12235), .ZN(
        n12239) );
  AND2_X1 U15490 ( .A1(n12972), .A2(n9576), .ZN(n14649) );
  INV_X1 U15491 ( .A(n11399), .ZN(n12242) );
  INV_X1 U15492 ( .A(n12238), .ZN(n15002) );
  INV_X1 U15493 ( .A(n12239), .ZN(n12241) );
  OAI211_X1 U15494 ( .C1(n12242), .C2(n15002), .A(n12241), .B(n12240), .ZN(
        n13977) );
  OAI21_X1 U15495 ( .B1(n12243), .B2(n11993), .A(n12244), .ZN(n12245) );
  OR2_X1 U15496 ( .A1(n13977), .A2(n12245), .ZN(n12246) );
  INV_X1 U15497 ( .A(n20676), .ZN(n13650) );
  NAND2_X1 U15498 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12263) );
  NAND2_X1 U15499 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15440) );
  NAND2_X1 U15500 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12247) );
  NOR2_X1 U15501 ( .A1(n15440), .A2(n12247), .ZN(n15432) );
  NAND2_X1 U15502 ( .A1(n15432), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12262) );
  NAND2_X1 U15503 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15513) );
  INV_X1 U15504 ( .A(n15513), .ZN(n14200) );
  INV_X1 U15505 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20664) );
  NOR2_X1 U15506 ( .A1(n20664), .A2(n20673), .ZN(n20658) );
  NAND2_X1 U15507 ( .A1(n14200), .A2(n20658), .ZN(n14199) );
  OR2_X1 U15508 ( .A1(n14201), .A2(n14199), .ZN(n15488) );
  NAND2_X1 U15509 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15519) );
  NOR2_X1 U15510 ( .A1(n15519), .A2(n21437), .ZN(n12248) );
  AND3_X1 U15511 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15466) );
  AND2_X1 U15512 ( .A1(n12248), .A2(n15466), .ZN(n15500) );
  NAND2_X1 U15513 ( .A1(n15500), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12249) );
  OR2_X1 U15514 ( .A1(n15488), .A2(n12249), .ZN(n12257) );
  INV_X1 U15515 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20703) );
  OAI21_X1 U15516 ( .B1(n13458), .B2(n20703), .A(n20690), .ZN(n15514) );
  NAND3_X1 U15517 ( .A1(n20658), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n15514), .ZN(n15467) );
  NOR2_X1 U15518 ( .A1(n15467), .A2(n12249), .ZN(n12259) );
  NOR2_X1 U15519 ( .A1(n20676), .A2(n12259), .ZN(n12253) );
  OR2_X1 U15520 ( .A1(n13648), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12252) );
  OR2_X1 U15521 ( .A1(n12250), .A2(n20683), .ZN(n12251) );
  NOR2_X1 U15522 ( .A1(n20702), .A2(n20677), .ZN(n15517) );
  AOI21_X1 U15523 ( .B1(n20676), .B2(n13648), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12256) );
  INV_X1 U15524 ( .A(n12254), .ZN(n15372) );
  OAI22_X1 U15525 ( .A1(n15372), .A2(n13652), .B1(n13648), .B2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12255) );
  NAND3_X1 U15526 ( .A1(n12916), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12740) );
  NAND2_X1 U15527 ( .A1(n12916), .A2(n15449), .ZN(n15352) );
  NAND2_X1 U15528 ( .A1(n13458), .A2(n13652), .ZN(n20701) );
  INV_X1 U15529 ( .A(n12257), .ZN(n12258) );
  NAND2_X1 U15530 ( .A1(n20675), .A2(n12258), .ZN(n15380) );
  INV_X1 U15531 ( .A(n12259), .ZN(n12260) );
  OR2_X1 U15532 ( .A1(n20676), .A2(n12260), .ZN(n12261) );
  NAND2_X1 U15533 ( .A1(n15380), .A2(n12261), .ZN(n15482) );
  NAND3_X1 U15534 ( .A1(n12264), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12720) );
  INV_X1 U15535 ( .A(n12720), .ZN(n15176) );
  NAND2_X1 U15536 ( .A1(n15391), .A2(n15176), .ZN(n15362) );
  NAND2_X1 U15537 ( .A1(n12266), .A2(n12265), .ZN(n12722) );
  NAND2_X1 U15538 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15353) );
  NAND2_X1 U15539 ( .A1(n12722), .A2(n15353), .ZN(n12267) );
  NAND2_X1 U15540 ( .A1(n20683), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15167) );
  OAI21_X1 U15541 ( .B1(n15362), .B2(n12267), .A(n15167), .ZN(n12268) );
  NOR2_X1 U15542 ( .A1(n12283), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12273) );
  AND2_X4 U15543 ( .A1(n13148), .A2(n12273), .ZN(n12480) );
  NAND2_X1 U15544 ( .A1(n12480), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12279) );
  NAND2_X1 U15545 ( .A1(n12283), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12277) );
  INV_X1 U15546 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12274) );
  NOR2_X1 U15547 ( .A1(n19806), .A2(n12274), .ZN(n12275) );
  NOR2_X1 U15548 ( .A1(n12275), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12276) );
  MUX2_X1 U15549 ( .A(n19806), .B(n20248), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12284) );
  NAND2_X1 U15550 ( .A1(n12282), .A2(n9597), .ZN(n12299) );
  OAI211_X1 U15551 ( .C1(n12285), .C2(n12448), .A(n12284), .B(n12299), .ZN(
        n13930) );
  NAND2_X1 U15552 ( .A1(n13929), .A2(n13930), .ZN(n12296) );
  AOI22_X1 U15553 ( .A1(n9594), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n9598), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12288) );
  XNOR2_X1 U15554 ( .A(n12296), .B(n12294), .ZN(n13926) );
  NAND2_X1 U15555 ( .A1(n12289), .A2(n19806), .ZN(n12290) );
  MUX2_X1 U15556 ( .A(n12290), .B(n20176), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12293) );
  NAND2_X1 U15557 ( .A1(n12431), .A2(n12291), .ZN(n12292) );
  AND2_X1 U15558 ( .A1(n12293), .A2(n12292), .ZN(n13925) );
  INV_X1 U15559 ( .A(n12294), .ZN(n12295) );
  NAND2_X1 U15560 ( .A1(n12296), .A2(n12295), .ZN(n12297) );
  NAND2_X1 U15561 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12298) );
  OAI211_X1 U15562 ( .C1(n12448), .C2(n12300), .A(n12299), .B(n12298), .ZN(
        n12303) );
  XNOR2_X1 U15563 ( .A(n12305), .B(n12303), .ZN(n13923) );
  NAND2_X1 U15564 ( .A1(n12480), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U15565 ( .A1(n9594), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n9598), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12301) );
  AND2_X1 U15566 ( .A1(n12302), .A2(n12301), .ZN(n13922) );
  INV_X1 U15567 ( .A(n12303), .ZN(n12304) );
  AOI22_X1 U15568 ( .A1(n12431), .A2(n11166), .B1(n9594), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n12308) );
  NAND2_X1 U15569 ( .A1(n12480), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12307) );
  AOI22_X1 U15570 ( .A1(n9598), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12306) );
  AND3_X1 U15571 ( .A1(n12308), .A2(n12307), .A3(n12306), .ZN(n14666) );
  INV_X1 U15572 ( .A(n14666), .ZN(n12309) );
  NAND2_X1 U15573 ( .A1(n9594), .A2(P2_EAX_REG_4__SCAN_IN), .ZN(n12311) );
  NAND2_X1 U15574 ( .A1(n9597), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12310) );
  OAI211_X1 U15575 ( .C1(n12448), .C2(n12312), .A(n12311), .B(n12310), .ZN(
        n12313) );
  INV_X1 U15576 ( .A(n12313), .ZN(n12315) );
  NAND2_X1 U15577 ( .A1(n12480), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12314) );
  AND2_X1 U15578 ( .A1(n12315), .A2(n12314), .ZN(n15882) );
  NAND2_X1 U15579 ( .A1(n13921), .A2(n12316), .ZN(n15881) );
  NAND2_X1 U15580 ( .A1(n9594), .A2(P2_EAX_REG_5__SCAN_IN), .ZN(n12318) );
  NAND2_X1 U15581 ( .A1(n9597), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12317) );
  OAI211_X1 U15582 ( .C1(n12448), .C2(n12319), .A(n12318), .B(n12317), .ZN(
        n12320) );
  INV_X1 U15583 ( .A(n12320), .ZN(n12322) );
  NAND2_X1 U15584 ( .A1(n12480), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12321) );
  AND2_X1 U15585 ( .A1(n12322), .A2(n12321), .ZN(n16146) );
  INV_X1 U15586 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20400) );
  AOI22_X1 U15587 ( .A1(n9594), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n9598), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12324) );
  OAI21_X1 U15588 ( .B1(n12479), .B2(n20400), .A(n12324), .ZN(n13146) );
  NAND2_X1 U15589 ( .A1(n12431), .A2(n11025), .ZN(n12325) );
  INV_X1 U15590 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20402) );
  AOI22_X1 U15591 ( .A1(n9594), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n9597), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12326) );
  OAI21_X1 U15592 ( .B1(n12479), .B2(n20402), .A(n12326), .ZN(n13158) );
  AOI22_X1 U15593 ( .A1(n14479), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10835), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12330) );
  AOI22_X1 U15594 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n9579), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U15595 ( .A1(n9585), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U15596 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10818), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12327) );
  NAND4_X1 U15597 ( .A1(n12330), .A2(n12329), .A3(n12328), .A4(n12327), .ZN(
        n12336) );
  AOI22_X1 U15598 ( .A1(n14435), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12334) );
  AOI22_X1 U15599 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9589), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12333) );
  AOI22_X1 U15600 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n9587), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12332) );
  AOI22_X1 U15601 ( .A1(n9591), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n9592), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12331) );
  NAND4_X1 U15602 ( .A1(n12334), .A2(n12333), .A3(n12332), .A4(n12331), .ZN(
        n12335) );
  INV_X1 U15603 ( .A(n13899), .ZN(n14238) );
  NAND2_X1 U15604 ( .A1(n9594), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n12338) );
  NAND2_X1 U15605 ( .A1(n9597), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12337) );
  OAI211_X1 U15606 ( .C1(n12448), .C2(n14238), .A(n12338), .B(n12337), .ZN(
        n12339) );
  INV_X1 U15607 ( .A(n12339), .ZN(n12341) );
  NAND2_X1 U15608 ( .A1(n12480), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U15609 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10699), .B1(
        n14435), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U15610 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9578), .B1(n9579), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U15611 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10806), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12345) );
  AOI22_X1 U15612 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10818), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12344) );
  NAND4_X1 U15613 ( .A1(n12347), .A2(n12346), .A3(n12345), .A4(n12344), .ZN(
        n12353) );
  AOI22_X1 U15614 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14479), .B1(
        n10835), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U15615 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n9591), .B1(n9590), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12350) );
  AOI22_X1 U15616 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n9588), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12349) );
  AOI22_X1 U15617 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10823), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12348) );
  NAND4_X1 U15618 ( .A1(n12351), .A2(n12350), .A3(n12349), .A4(n12348), .ZN(
        n12352) );
  INV_X1 U15619 ( .A(n14080), .ZN(n12356) );
  NAND2_X1 U15620 ( .A1(n9594), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n12355) );
  NAND2_X1 U15621 ( .A1(n9598), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12354) );
  OAI211_X1 U15622 ( .C1(n12448), .C2(n12356), .A(n12355), .B(n12354), .ZN(
        n12357) );
  INV_X1 U15623 ( .A(n12357), .ZN(n12359) );
  NAND2_X1 U15624 ( .A1(n12480), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12358) );
  INV_X1 U15625 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12372) );
  AOI22_X1 U15626 ( .A1(n9594), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n9598), .B2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U15627 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n10699), .B1(
        n14435), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U15628 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10818), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U15629 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10806), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15630 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12360) );
  NAND4_X1 U15631 ( .A1(n12363), .A2(n12362), .A3(n12361), .A4(n12360), .ZN(
        n12369) );
  AOI22_X1 U15632 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n14479), .B1(
        n10835), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12367) );
  AOI22_X1 U15633 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n9588), .B1(n9591), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12366) );
  AOI22_X1 U15634 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n14473), .B1(
        n9590), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12365) );
  AOI22_X1 U15635 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10823), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12364) );
  NAND4_X1 U15636 ( .A1(n12367), .A2(n12366), .A3(n12365), .A4(n12364), .ZN(
        n12368) );
  NAND2_X1 U15637 ( .A1(n12431), .A2(n13905), .ZN(n12370) );
  OAI211_X1 U15638 ( .C1(n12479), .C2(n12372), .A(n12371), .B(n12370), .ZN(
        n13287) );
  NAND2_X1 U15639 ( .A1(n13286), .A2(n13287), .ZN(n13285) );
  INV_X1 U15640 ( .A(n13285), .ZN(n12389) );
  AOI22_X1 U15641 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n10699), .B1(
        n14435), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15642 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n9578), .B1(n9579), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U15643 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10806), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12374) );
  AOI22_X1 U15644 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10818), .B1(
        n9585), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12373) );
  NAND4_X1 U15645 ( .A1(n12376), .A2(n12375), .A3(n12374), .A4(n12373), .ZN(
        n12382) );
  AOI22_X1 U15646 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n14479), .B1(
        n10835), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12380) );
  AOI22_X1 U15647 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n9591), .B1(n9589), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12379) );
  AOI22_X1 U15648 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n9588), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U15649 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n9587), .B1(n9592), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12377) );
  NAND4_X1 U15650 ( .A1(n12380), .A2(n12379), .A3(n12378), .A4(n12377), .ZN(
        n12381) );
  NAND2_X1 U15651 ( .A1(n9594), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n12384) );
  NAND2_X1 U15652 ( .A1(n9598), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12383) );
  OAI211_X1 U15653 ( .C1(n12448), .C2(n13964), .A(n12384), .B(n12383), .ZN(
        n12385) );
  INV_X1 U15654 ( .A(n12385), .ZN(n12387) );
  NAND2_X1 U15655 ( .A1(n12480), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U15656 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n14479), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12393) );
  AOI22_X1 U15657 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10818), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12392) );
  AOI22_X1 U15658 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n9584), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12391) );
  AOI22_X1 U15659 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12390) );
  NAND4_X1 U15660 ( .A1(n12393), .A2(n12392), .A3(n12391), .A4(n12390), .ZN(
        n12399) );
  AOI22_X1 U15661 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10835), .B1(
        n14435), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12397) );
  AOI22_X1 U15662 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n9591), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12396) );
  AOI22_X1 U15663 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n9588), .B1(n9590), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12395) );
  AOI22_X1 U15664 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10823), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12394) );
  NAND4_X1 U15665 ( .A1(n12397), .A2(n12396), .A3(n12395), .A4(n12394), .ZN(
        n12398) );
  INV_X1 U15666 ( .A(n14391), .ZN(n14207) );
  NAND2_X1 U15667 ( .A1(n9594), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n12401) );
  NAND2_X1 U15668 ( .A1(n9598), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12400) );
  OAI211_X1 U15669 ( .C1(n12448), .C2(n14207), .A(n12401), .B(n12400), .ZN(
        n12402) );
  INV_X1 U15670 ( .A(n12402), .ZN(n12404) );
  NAND2_X1 U15671 ( .A1(n12480), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U15672 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n10699), .B1(
        n14435), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15673 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n9578), .B1(n9579), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12407) );
  AOI22_X1 U15674 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n10806), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12406) );
  AOI22_X1 U15675 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10818), .B1(
        n9585), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12405) );
  NAND4_X1 U15676 ( .A1(n12408), .A2(n12407), .A3(n12406), .A4(n12405), .ZN(
        n12414) );
  AOI22_X1 U15677 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n14479), .B1(
        n10835), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12412) );
  AOI22_X1 U15678 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n9591), .B1(n9589), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12411) );
  AOI22_X1 U15679 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n9588), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U15680 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n9587), .B1(n9592), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12409) );
  NAND4_X1 U15681 ( .A1(n12412), .A2(n12411), .A3(n12410), .A4(n12409), .ZN(
        n12413) );
  INV_X1 U15682 ( .A(n16039), .ZN(n12417) );
  NAND2_X1 U15683 ( .A1(n9594), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n12416) );
  NAND2_X1 U15684 ( .A1(n9597), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12415) );
  OAI211_X1 U15685 ( .C1(n12448), .C2(n12417), .A(n12416), .B(n12415), .ZN(
        n12418) );
  INV_X1 U15686 ( .A(n12418), .ZN(n12420) );
  NAND2_X1 U15687 ( .A1(n12480), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12419) );
  INV_X1 U15688 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n12434) );
  AOI22_X1 U15689 ( .A1(n9594), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n9598), .B2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12433) );
  AOI22_X1 U15690 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n14479), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12424) );
  AOI22_X1 U15691 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n9578), .B1(n9579), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12423) );
  AOI22_X1 U15692 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10806), .B1(
        n9585), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12422) );
  AOI22_X1 U15693 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10818), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12421) );
  NAND4_X1 U15694 ( .A1(n12424), .A2(n12423), .A3(n12422), .A4(n12421), .ZN(
        n12430) );
  AOI22_X1 U15695 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10835), .B1(
        n14435), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12428) );
  AOI22_X1 U15696 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n9588), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12427) );
  AOI22_X1 U15697 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n9592), .B1(
        n9589), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U15698 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n9591), .B1(n9587), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12425) );
  NAND4_X1 U15699 ( .A1(n12428), .A2(n12427), .A3(n12426), .A4(n12425), .ZN(
        n12429) );
  NAND2_X1 U15700 ( .A1(n12431), .A2(n16033), .ZN(n12432) );
  OAI211_X1 U15701 ( .C1(n12479), .C2(n12434), .A(n12433), .B(n12432), .ZN(
        n13789) );
  AOI22_X1 U15702 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n10699), .B1(
        n14435), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15703 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n9578), .B1(n9579), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U15704 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10806), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U15705 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10818), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12435) );
  NAND4_X1 U15706 ( .A1(n12438), .A2(n12437), .A3(n12436), .A4(n12435), .ZN(
        n12444) );
  AOI22_X1 U15707 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n14479), .B1(
        n10835), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12442) );
  AOI22_X1 U15708 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n9591), .B1(n9590), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12441) );
  AOI22_X1 U15709 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n9588), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12440) );
  AOI22_X1 U15710 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n9587), .B1(n9592), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12439) );
  NAND4_X1 U15711 ( .A1(n12442), .A2(n12441), .A3(n12440), .A4(n12439), .ZN(
        n12443) );
  INV_X1 U15712 ( .A(n16027), .ZN(n12447) );
  NAND2_X1 U15713 ( .A1(n9594), .A2(P2_EAX_REG_15__SCAN_IN), .ZN(n12446) );
  NAND2_X1 U15714 ( .A1(n9598), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12445) );
  OAI211_X1 U15715 ( .C1(n12448), .C2(n12447), .A(n12446), .B(n12445), .ZN(
        n12449) );
  INV_X1 U15716 ( .A(n12449), .ZN(n12451) );
  NAND2_X1 U15717 ( .A1(n12480), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12450) );
  NAND2_X1 U15718 ( .A1(n12480), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U15719 ( .A1(n9594), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n9598), .B2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12454) );
  INV_X1 U15720 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20420) );
  AOI22_X1 U15721 ( .A1(n9594), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n9597), .B2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12456) );
  OAI21_X1 U15722 ( .B1(n12479), .B2(n20420), .A(n12456), .ZN(n12802) );
  NAND2_X1 U15723 ( .A1(n12799), .A2(n12802), .ZN(n12800) );
  INV_X1 U15724 ( .A(n12800), .ZN(n12460) );
  NAND2_X1 U15725 ( .A1(n12480), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U15726 ( .A1(n9594), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n9598), .B2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12457) );
  INV_X1 U15727 ( .A(n15749), .ZN(n12459) );
  NAND2_X1 U15728 ( .A1(n12480), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U15729 ( .A1(n9594), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n9598), .B2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12461) );
  NAND2_X1 U15730 ( .A1(n12480), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15731 ( .A1(n9594), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n9598), .B2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12463) );
  INV_X1 U15732 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20426) );
  AOI22_X1 U15733 ( .A1(n9594), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n9598), .B2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12465) );
  OAI21_X1 U15734 ( .B1(n12479), .B2(n20426), .A(n12465), .ZN(n12821) );
  NAND2_X1 U15735 ( .A1(n12480), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12467) );
  AOI22_X1 U15736 ( .A1(n9594), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n9598), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12466) );
  NAND2_X1 U15737 ( .A1(n12480), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U15738 ( .A1(n9594), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n9598), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12468) );
  AND2_X1 U15739 ( .A1(n12469), .A2(n12468), .ZN(n15679) );
  INV_X1 U15740 ( .A(n15679), .ZN(n12470) );
  INV_X1 U15741 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20431) );
  AOI22_X1 U15742 ( .A1(n9594), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n9597), .B2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12471) );
  OAI21_X1 U15743 ( .B1(n12479), .B2(n20431), .A(n12471), .ZN(n15667) );
  NAND2_X1 U15744 ( .A1(n12480), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12473) );
  AOI22_X1 U15745 ( .A1(n9594), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n9598), .B2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12472) );
  AND2_X1 U15746 ( .A1(n12473), .A2(n12472), .ZN(n15650) );
  NAND2_X1 U15747 ( .A1(n12480), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U15748 ( .A1(n9594), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n9598), .B2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12474) );
  INV_X1 U15749 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20438) );
  AOI22_X1 U15750 ( .A1(n9594), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n9598), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12476) );
  OAI21_X1 U15751 ( .B1(n12479), .B2(n20438), .A(n12476), .ZN(n15621) );
  INV_X1 U15752 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20439) );
  AOI22_X1 U15753 ( .A1(n9594), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n9598), .B2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12478) );
  OAI21_X1 U15754 ( .B1(n12479), .B2(n20439), .A(n12478), .ZN(n14355) );
  INV_X1 U15755 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14168) );
  OAI222_X1 U15756 ( .A1(n14168), .A2(n9639), .B1(n20441), .B2(n12479), .C1(
        n12287), .C2(n21478), .ZN(n15599) );
  NAND2_X2 U15757 ( .A1(n14353), .A2(n15599), .ZN(n15600) );
  AOI222_X1 U15758 ( .A1(n12480), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n9594), 
        .B2(P2_EAX_REG_30__SCAN_IN), .C1(n9598), .C2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12754) );
  AOI222_X1 U15759 ( .A1(n12480), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n9594), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n9598), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12481) );
  NAND2_X1 U15760 ( .A1(n12494), .A2(n15978), .ZN(n12483) );
  MUX2_X1 U15761 ( .A(n12483), .B(n12482), .S(n12484), .Z(n12491) );
  NAND2_X1 U15762 ( .A1(n14120), .A2(n12484), .ZN(n12488) );
  OAI211_X1 U15763 ( .C1(n15978), .C2(n12486), .A(n12558), .B(n12485), .ZN(
        n12487) );
  OAI211_X1 U15764 ( .C1(n12482), .C2(n12489), .A(n12488), .B(n12487), .ZN(
        n12490) );
  NAND2_X1 U15765 ( .A1(n12491), .A2(n12490), .ZN(n12493) );
  INV_X1 U15766 ( .A(n12495), .ZN(n12496) );
  NOR2_X1 U15767 ( .A1(n19777), .A2(n15978), .ZN(n12506) );
  OAI21_X1 U15768 ( .B1(n12506), .B2(n10323), .A(n12499), .ZN(n12500) );
  NAND2_X1 U15769 ( .A1(n12498), .A2(n12500), .ZN(n12505) );
  NAND2_X1 U15770 ( .A1(n12501), .A2(n19806), .ZN(n12503) );
  NOR2_X1 U15771 ( .A1(n12558), .A2(n15978), .ZN(n12502) );
  NAND2_X1 U15772 ( .A1(n12503), .A2(n12502), .ZN(n12557) );
  AND3_X1 U15773 ( .A1(n12505), .A2(n12504), .A3(n12557), .ZN(n12536) );
  AND2_X1 U15774 ( .A1(n12282), .A2(n12506), .ZN(n12507) );
  NAND2_X1 U15775 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20369) );
  AND2_X1 U15776 ( .A1(n15586), .A2(n20369), .ZN(n12948) );
  NAND2_X1 U15777 ( .A1(n12509), .A2(n12951), .ZN(n12950) );
  INV_X1 U15778 ( .A(n12950), .ZN(n12510) );
  NAND3_X1 U15779 ( .A1(n12513), .A2(n12559), .A3(n14120), .ZN(n12514) );
  NAND2_X1 U15780 ( .A1(n12692), .A2(n19648), .ZN(n12531) );
  AND2_X1 U15781 ( .A1(n10593), .A2(n19806), .ZN(n12515) );
  NOR4_X1 U15782 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12519) );
  NOR4_X1 U15783 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12518) );
  NOR4_X1 U15784 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12517) );
  NOR4_X1 U15785 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12516) );
  AND4_X1 U15786 ( .A1(n12519), .A2(n12518), .A3(n12517), .A4(n12516), .ZN(
        n12524) );
  NOR4_X1 U15787 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12522) );
  NOR4_X1 U15788 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12521) );
  NOR4_X1 U15789 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12520) );
  INV_X1 U15790 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20395) );
  AND4_X1 U15791 ( .A1(n12522), .A2(n12521), .A3(n12520), .A4(n20395), .ZN(
        n12523) );
  NAND2_X1 U15792 ( .A1(n12524), .A2(n12523), .ZN(n12525) );
  AOI22_X1 U15793 ( .A1(n16136), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19647), .ZN(n12526) );
  INV_X1 U15794 ( .A(n12526), .ZN(n12529) );
  INV_X1 U15795 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n17433) );
  NOR2_X1 U15796 ( .A1(n16140), .A2(n17433), .ZN(n12528) );
  NOR2_X1 U15797 ( .A1(n12529), .A2(n12528), .ZN(n12530) );
  NAND2_X1 U15798 ( .A1(n12531), .A2(n12530), .ZN(P2_U2888) );
  NOR2_X1 U15799 ( .A1(n20370), .A2(n20391), .ZN(n20380) );
  NOR2_X1 U15800 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20383) );
  NOR3_X1 U15801 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20380), .A3(n20383), 
        .ZN(n15582) );
  NAND2_X1 U15802 ( .A1(n20369), .A2(n15582), .ZN(n13820) );
  INV_X1 U15803 ( .A(n13820), .ZN(n12949) );
  NAND2_X1 U15804 ( .A1(n10584), .A2(n12949), .ZN(n12544) );
  AOI21_X1 U15805 ( .B1(n12532), .B2(n12558), .A(n19777), .ZN(n12542) );
  INV_X1 U15806 ( .A(n12533), .ZN(n12540) );
  NAND3_X1 U15807 ( .A1(n12534), .A2(n12951), .A3(n12949), .ZN(n12535) );
  AND3_X1 U15808 ( .A1(n12537), .A2(n12536), .A3(n12535), .ZN(n13821) );
  MUX2_X1 U15809 ( .A(n12534), .B(n10584), .S(n9595), .Z(n12538) );
  NAND3_X1 U15810 ( .A1(n12538), .A2(n12951), .A3(n20369), .ZN(n12539) );
  NAND3_X1 U15811 ( .A1(n12540), .A2(n13821), .A3(n12539), .ZN(n12541) );
  AOI21_X1 U15812 ( .B1(n14151), .B2(n12542), .A(n12541), .ZN(n12543) );
  OAI21_X1 U15813 ( .B1(n14151), .B2(n12544), .A(n12543), .ZN(n12545) );
  INV_X1 U15814 ( .A(n12587), .ZN(n12552) );
  NAND2_X1 U15815 ( .A1(n14108), .A2(n9596), .ZN(n12550) );
  NAND2_X1 U15816 ( .A1(n12550), .A2(n12549), .ZN(n12551) );
  NAND2_X1 U15817 ( .A1(n12553), .A2(n15586), .ZN(n12555) );
  NAND2_X1 U15818 ( .A1(n12555), .A2(n12554), .ZN(n12565) );
  NAND2_X1 U15819 ( .A1(n12556), .A2(n15978), .ZN(n14102) );
  NAND2_X1 U15820 ( .A1(n14102), .A2(n12557), .ZN(n12563) );
  OAI22_X1 U15821 ( .A1(n15586), .A2(n19777), .B1(n12559), .B2(n12558), .ZN(
        n12560) );
  INV_X1 U15822 ( .A(n12560), .ZN(n12561) );
  AOI21_X1 U15823 ( .B1(n12563), .B2(n10585), .A(n12562), .ZN(n12564) );
  NAND2_X1 U15824 ( .A1(n12565), .A2(n12564), .ZN(n14111) );
  NOR2_X1 U15825 ( .A1(n14111), .A2(n9566), .ZN(n12566) );
  OR2_X2 U15826 ( .A1(n19719), .A2(n12791), .ZN(n16733) );
  NAND2_X1 U15827 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19729) );
  NAND2_X1 U15828 ( .A1(n12791), .A2(n19729), .ZN(n12567) );
  INV_X1 U15829 ( .A(n19604), .ZN(n16416) );
  NAND2_X1 U15830 ( .A1(n12587), .A2(n16416), .ZN(n16729) );
  AND2_X1 U15831 ( .A1(n12567), .A2(n16729), .ZN(n19723) );
  NAND2_X1 U15832 ( .A1(n17413), .A2(n19723), .ZN(n16713) );
  NAND3_X1 U15833 ( .A1(n19719), .A2(n19722), .A3(n19729), .ZN(n19736) );
  NAND2_X1 U15834 ( .A1(n12791), .A2(n19722), .ZN(n19730) );
  NAND3_X1 U15835 ( .A1(n19723), .A2(n19736), .A3(n19730), .ZN(n16714) );
  NOR3_X1 U15836 ( .A1(n19717), .A2(n16715), .A3(n16717), .ZN(n16698) );
  NAND2_X1 U15837 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16698), .ZN(
        n12575) );
  NOR2_X1 U15838 ( .A1(n16714), .A2(n9664), .ZN(n16688) );
  NOR2_X1 U15839 ( .A1(n16687), .A2(n16677), .ZN(n16673) );
  INV_X1 U15840 ( .A(n16673), .ZN(n12568) );
  NAND2_X1 U15841 ( .A1(n16733), .A2(n12568), .ZN(n12569) );
  INV_X1 U15842 ( .A(n12576), .ZN(n12570) );
  NAND2_X1 U15843 ( .A1(n16733), .A2(n12570), .ZN(n12571) );
  AOI21_X1 U15844 ( .B1(n16733), .B2(n16492), .A(n16479), .ZN(n12572) );
  NAND2_X1 U15845 ( .A1(n16509), .A2(n12572), .ZN(n16482) );
  NAND2_X1 U15846 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12577) );
  OR2_X1 U15847 ( .A1(n16482), .A2(n12577), .ZN(n12573) );
  AND2_X1 U15848 ( .A1(n12573), .A2(n16713), .ZN(n16443) );
  AOI21_X1 U15849 ( .B1(n12759), .B2(n16713), .A(n16443), .ZN(n12758) );
  OAI21_X1 U15850 ( .B1(n17413), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12758), .ZN(n12580) );
  NOR2_X1 U15851 ( .A1(n19722), .A2(n19729), .ZN(n19718) );
  NAND2_X1 U15852 ( .A1(n19722), .A2(n19729), .ZN(n12574) );
  OAI211_X1 U15853 ( .C1(n19719), .C2(n19718), .A(n12574), .B(n16733), .ZN(
        n14669) );
  INV_X1 U15854 ( .A(n12577), .ZN(n14347) );
  NOR4_X1 U15855 ( .A1(n16446), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12766), .A4(n12759), .ZN(n12578) );
  AOI211_X1 U15856 ( .C1(n12580), .C2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n12579), .B(n12578), .ZN(n12581) );
  OAI21_X1 U15857 ( .B1(n15946), .B2(n19728), .A(n12581), .ZN(n12582) );
  INV_X1 U15858 ( .A(n12582), .ZN(n12589) );
  NAND2_X1 U15859 ( .A1(n12509), .A2(n15978), .ZN(n12585) );
  AND2_X1 U15860 ( .A1(n12585), .A2(n13807), .ZN(n12586) );
  NAND2_X1 U15861 ( .A1(n12692), .A2(n16731), .ZN(n12588) );
  INV_X1 U15862 ( .A(n12803), .ZN(n12591) );
  INV_X1 U15863 ( .A(n16524), .ZN(n16523) );
  AND2_X1 U15864 ( .A1(n12796), .A2(n12592), .ZN(n12593) );
  OR2_X1 U15865 ( .A1(n12593), .A2(n9714), .ZN(n16552) );
  INV_X1 U15866 ( .A(n12594), .ZN(n12650) );
  NAND2_X1 U15867 ( .A1(n12595), .A2(n12597), .ZN(n12596) );
  AND2_X1 U15868 ( .A1(n12650), .A2(n12596), .ZN(n15745) );
  INV_X1 U15869 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15751) );
  NOR2_X1 U15870 ( .A1(n19705), .A2(n15751), .ZN(n16547) );
  NOR2_X1 U15871 ( .A1(n16419), .A2(n12597), .ZN(n12598) );
  AOI211_X1 U15872 ( .C1(n15745), .C2(n16425), .A(n16547), .B(n12598), .ZN(
        n12599) );
  OAI21_X1 U15873 ( .B1(n16552), .B2(n16429), .A(n12599), .ZN(n12600) );
  AOI21_X1 U15874 ( .B1(n16554), .B2(n16415), .A(n12600), .ZN(n12616) );
  INV_X1 U15875 ( .A(n16307), .ZN(n12603) );
  INV_X1 U15876 ( .A(n16300), .ZN(n12604) );
  INV_X1 U15877 ( .A(n12605), .ZN(n16271) );
  INV_X1 U15878 ( .A(n12606), .ZN(n16558) );
  NAND2_X1 U15879 ( .A1(n12609), .A2(n12608), .ZN(n12808) );
  INV_X1 U15880 ( .A(n12609), .ZN(n12610) );
  INV_X1 U15881 ( .A(n12611), .ZN(n16244) );
  NOR2_X1 U15882 ( .A1(n16244), .A2(n12811), .ZN(n12613) );
  XNOR2_X1 U15883 ( .A(n12812), .B(n12613), .ZN(n16555) );
  NAND2_X1 U15884 ( .A1(n12616), .A2(n12615), .ZN(P2_U2996) );
  NAND2_X1 U15885 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12618) );
  NAND2_X2 U15886 ( .A1(n12619), .A2(n12618), .ZN(n9609) );
  MUX2_X1 U15887 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n14299) );
  INV_X1 U15888 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12620) );
  MUX2_X1 U15889 ( .A(n12620), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n14274) );
  NOR2_X1 U15890 ( .A1(n14299), .A2(n14274), .ZN(n15915) );
  OAI21_X1 U15891 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n9711), .ZN(n15916) );
  AND2_X1 U15892 ( .A1(n15915), .A2(n15916), .ZN(n15903) );
  INV_X1 U15893 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15898) );
  NAND2_X1 U15894 ( .A1(n9711), .A2(n15898), .ZN(n12622) );
  NAND2_X1 U15895 ( .A1(n12621), .A2(n12622), .ZN(n15904) );
  NAND2_X1 U15896 ( .A1(n15903), .A2(n15904), .ZN(n15891) );
  NAND2_X1 U15897 ( .A1(n12621), .A2(n16418), .ZN(n12623) );
  AND2_X1 U15898 ( .A1(n9718), .A2(n12623), .ZN(n16426) );
  NOR2_X1 U15899 ( .A1(n15891), .A2(n16426), .ZN(n19613) );
  INV_X1 U15900 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12624) );
  NAND2_X1 U15901 ( .A1(n9718), .A2(n12624), .ZN(n12625) );
  NAND2_X1 U15902 ( .A1(n12627), .A2(n12625), .ZN(n19615) );
  NAND2_X1 U15903 ( .A1(n19613), .A2(n19615), .ZN(n15868) );
  NAND2_X1 U15904 ( .A1(n12627), .A2(n10302), .ZN(n12628) );
  AND2_X1 U15905 ( .A1(n12626), .A2(n12628), .ZN(n16391) );
  OR2_X1 U15906 ( .A1(n15868), .A2(n16391), .ZN(n15855) );
  NAND2_X1 U15907 ( .A1(n12626), .A2(n15861), .ZN(n12629) );
  AND2_X1 U15908 ( .A1(n10303), .A2(n12629), .ZN(n16378) );
  OR2_X1 U15909 ( .A1(n15855), .A2(n16378), .ZN(n14250) );
  INV_X1 U15910 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16368) );
  NAND2_X1 U15911 ( .A1(n10303), .A2(n16368), .ZN(n12630) );
  AND2_X1 U15912 ( .A1(n9721), .A2(n12630), .ZN(n16372) );
  NOR2_X1 U15913 ( .A1(n14250), .A2(n16372), .ZN(n15842) );
  INV_X1 U15914 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15847) );
  NAND2_X1 U15915 ( .A1(n9721), .A2(n15847), .ZN(n12632) );
  NAND2_X1 U15916 ( .A1(n12631), .A2(n12632), .ZN(n16356) );
  AND2_X1 U15917 ( .A1(n15842), .A2(n16356), .ZN(n15828) );
  NAND2_X1 U15918 ( .A1(n12631), .A2(n15834), .ZN(n12633) );
  NAND2_X1 U15919 ( .A1(n12634), .A2(n12633), .ZN(n16344) );
  AND2_X1 U15920 ( .A1(n15828), .A2(n16344), .ZN(n14286) );
  NAND2_X1 U15921 ( .A1(n12634), .A2(n14292), .ZN(n12635) );
  NAND2_X1 U15922 ( .A1(n9710), .A2(n12635), .ZN(n16327) );
  NAND2_X1 U15923 ( .A1(n14286), .A2(n16327), .ZN(n14265) );
  AOI21_X1 U15924 ( .B1(n16311), .B2(n9710), .A(n12637), .ZN(n16314) );
  NOR2_X1 U15925 ( .A1(n14265), .A2(n16314), .ZN(n15821) );
  OAI21_X1 U15926 ( .B1(n12637), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n12636), .ZN(n16299) );
  NAND2_X1 U15927 ( .A1(n15821), .A2(n16299), .ZN(n15799) );
  INV_X1 U15928 ( .A(n12638), .ZN(n12639) );
  NAND2_X1 U15929 ( .A1(n12636), .A2(n16292), .ZN(n12640) );
  AND2_X1 U15930 ( .A1(n12639), .A2(n12640), .ZN(n16294) );
  INV_X1 U15931 ( .A(n12641), .ZN(n12645) );
  NAND2_X1 U15932 ( .A1(n12639), .A2(n15790), .ZN(n12642) );
  NAND2_X1 U15933 ( .A1(n12645), .A2(n12642), .ZN(n16281) );
  INV_X1 U15934 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12644) );
  NAND2_X1 U15935 ( .A1(n12645), .A2(n12644), .ZN(n12646) );
  AND2_X1 U15936 ( .A1(n10459), .A2(n12646), .ZN(n16266) );
  INV_X1 U15937 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12647) );
  NAND2_X1 U15938 ( .A1(n10459), .A2(n12647), .ZN(n12648) );
  NAND2_X1 U15939 ( .A1(n12595), .A2(n12648), .ZN(n16259) );
  INV_X1 U15940 ( .A(n12649), .ZN(n12652) );
  NAND2_X1 U15941 ( .A1(n12650), .A2(n15739), .ZN(n12651) );
  NAND2_X1 U15942 ( .A1(n12652), .A2(n12651), .ZN(n16252) );
  INV_X1 U15943 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15719) );
  NAND2_X1 U15944 ( .A1(n12652), .A2(n15719), .ZN(n12653) );
  AND2_X1 U15945 ( .A1(n9719), .A2(n12653), .ZN(n16237) );
  INV_X1 U15946 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12655) );
  NAND2_X1 U15947 ( .A1(n9719), .A2(n12655), .ZN(n12656) );
  NAND2_X1 U15948 ( .A1(n12654), .A2(n12656), .ZN(n15703) );
  NAND2_X1 U15949 ( .A1(n12654), .A2(n16222), .ZN(n12657) );
  AND2_X1 U15950 ( .A1(n9722), .A2(n12657), .ZN(n16225) );
  NAND2_X1 U15951 ( .A1(n9722), .A2(n10317), .ZN(n12659) );
  NAND2_X1 U15952 ( .A1(n15663), .A2(n9609), .ZN(n12662) );
  INV_X1 U15953 ( .A(n12660), .ZN(n12664) );
  NAND2_X1 U15954 ( .A1(n12658), .A2(n16206), .ZN(n12661) );
  NAND2_X1 U15955 ( .A1(n12664), .A2(n12661), .ZN(n15664) );
  NAND2_X1 U15956 ( .A1(n12664), .A2(n10282), .ZN(n12665) );
  NAND2_X1 U15957 ( .A1(n12663), .A2(n12665), .ZN(n16194) );
  NAND2_X1 U15958 ( .A1(n12663), .A2(n16180), .ZN(n12667) );
  NAND2_X1 U15959 ( .A1(n12666), .A2(n12667), .ZN(n15633) );
  NAND2_X1 U15960 ( .A1(n12668), .A2(n15633), .ZN(n15617) );
  INV_X1 U15961 ( .A(n12669), .ZN(n12671) );
  NAND2_X1 U15962 ( .A1(n12666), .A2(n16170), .ZN(n12670) );
  NAND2_X1 U15963 ( .A1(n12671), .A2(n12670), .ZN(n15618) );
  INV_X1 U15964 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15610) );
  NAND2_X1 U15965 ( .A1(n12671), .A2(n15610), .ZN(n12672) );
  NAND2_X1 U15966 ( .A1(n15594), .A2(n9609), .ZN(n12675) );
  NAND2_X1 U15967 ( .A1(n10467), .A2(n16162), .ZN(n12674) );
  NAND2_X1 U15968 ( .A1(n12673), .A2(n12674), .ZN(n15595) );
  NAND2_X1 U15969 ( .A1(n12675), .A2(n15595), .ZN(n15596) );
  INV_X1 U15970 ( .A(n15944), .ZN(n12679) );
  XNOR2_X1 U15971 ( .A(n12673), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14682) );
  INV_X1 U15972 ( .A(n14682), .ZN(n12678) );
  NAND2_X1 U15973 ( .A1(n12679), .A2(n12678), .ZN(n14693) );
  INV_X1 U15974 ( .A(n20369), .ZN(n20381) );
  NAND2_X1 U15975 ( .A1(n13703), .A2(n15978), .ZN(n13704) );
  NOR2_X1 U15976 ( .A1(n15946), .A2(n15937), .ZN(n12690) );
  AND2_X1 U15977 ( .A1(n20369), .A2(n20122), .ZN(n12681) );
  NOR2_X1 U15978 ( .A1(n12941), .A2(n12681), .ZN(n14253) );
  AND2_X1 U15979 ( .A1(n15978), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12682) );
  INV_X1 U15980 ( .A(n15791), .ZN(n15914) );
  INV_X1 U15981 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20302) );
  AND2_X1 U15982 ( .A1(n20302), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12946) );
  NOR2_X1 U15983 ( .A1(n20304), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12683) );
  NAND2_X1 U15984 ( .A1(n12946), .A2(n12683), .ZN(n17416) );
  AND3_X1 U15985 ( .A1(n15914), .A2(n17416), .A3(n19705), .ZN(n12684) );
  NAND2_X1 U15986 ( .A1(n20122), .A2(n12949), .ZN(n14135) );
  NAND2_X1 U15987 ( .A1(n13877), .A2(n14135), .ZN(n14255) );
  OAI22_X1 U15988 ( .A1(n20448), .A2(n15816), .B1(n14255), .B2(n14252), .ZN(
        n12686) );
  AOI21_X1 U15989 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n15930), .A(
        n12686), .ZN(n12687) );
  OAI21_X1 U15990 ( .B1(n12688), .B2(n15875), .A(n12687), .ZN(n12689) );
  NOR2_X1 U15991 ( .A1(n12690), .A2(n12689), .ZN(n12694) );
  INV_X1 U15992 ( .A(n14135), .ZN(n12691) );
  NOR2_X1 U15993 ( .A1(n15430), .A2(n15412), .ZN(n12701) );
  NAND2_X1 U15994 ( .A1(n15232), .A2(n15423), .ZN(n12696) );
  NAND2_X1 U15995 ( .A1(n12697), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12698) );
  NAND2_X1 U15996 ( .A1(n12769), .A2(n20650), .ZN(n12716) );
  AND3_X1 U15997 ( .A1(n10072), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n14061) );
  NOR2_X2 U15998 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21163) );
  INV_X1 U15999 ( .A(n12704), .ZN(n14872) );
  AND2_X1 U16000 ( .A1(n12704), .A2(n12703), .ZN(n14808) );
  AOI21_X1 U16001 ( .B1(n12705), .B2(n14836), .A(n14808), .ZN(n12706) );
  NAND2_X1 U16002 ( .A1(n21377), .A2(n21376), .ZN(n12707) );
  NAND2_X1 U16003 ( .A1(n12707), .A2(n10072), .ZN(n12708) );
  NAND2_X1 U16004 ( .A1(n10072), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15579) );
  NAND2_X1 U16005 ( .A1(n21191), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12709) );
  NAND2_X1 U16006 ( .A1(n15579), .A2(n12709), .ZN(n13465) );
  INV_X1 U16007 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n14826) );
  NOR2_X1 U16008 ( .A1(n20667), .A2(n14826), .ZN(n12772) );
  NOR2_X1 U16009 ( .A1(n15344), .A2(n12710), .ZN(n12711) );
  AOI211_X1 U16010 ( .C1(n14825), .C2(n15347), .A(n12772), .B(n12711), .ZN(
        n12712) );
  INV_X1 U16011 ( .A(n12712), .ZN(n12713) );
  NAND2_X1 U16012 ( .A1(n12716), .A2(n12715), .ZN(P1_U2978) );
  INV_X1 U16013 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15371) );
  NAND3_X1 U16014 ( .A1(n12717), .A2(n15394), .A3(n15371), .ZN(n12718) );
  INV_X1 U16015 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15355) );
  INV_X1 U16016 ( .A(n15353), .ZN(n12723) );
  NAND2_X1 U16017 ( .A1(n12723), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12739) );
  NOR2_X1 U16018 ( .A1(n15324), .A2(n12739), .ZN(n12724) );
  XNOR2_X1 U16019 ( .A(n12725), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14712) );
  OR2_X1 U16020 ( .A1(n13240), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12728) );
  INV_X1 U16021 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15025) );
  NAND2_X1 U16022 ( .A1(n12726), .A2(n15025), .ZN(n12727) );
  NAND2_X1 U16023 ( .A1(n12728), .A2(n12727), .ZN(n12730) );
  OAI22_X1 U16024 ( .A1(n12730), .A2(n12782), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n12729), .ZN(n14732) );
  NAND2_X1 U16025 ( .A1(n14731), .A2(n12782), .ZN(n12734) );
  INV_X1 U16026 ( .A(n12730), .ZN(n12731) );
  NAND2_X1 U16027 ( .A1(n12732), .A2(n12731), .ZN(n12733) );
  NAND2_X1 U16028 ( .A1(n12734), .A2(n12733), .ZN(n12737) );
  AND2_X1 U16029 ( .A1(n13625), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12735) );
  AOI21_X1 U16030 ( .B1(n13240), .B2(P1_EBX_REG_30__SCAN_IN), .A(n12735), .ZN(
        n12781) );
  INV_X1 U16031 ( .A(n12781), .ZN(n12736) );
  INV_X1 U16032 ( .A(n14379), .ZN(n12738) );
  OAI21_X1 U16033 ( .B1(n12740), .B2(n12739), .A(n15352), .ZN(n12741) );
  INV_X1 U16034 ( .A(n12786), .ZN(n12743) );
  NOR2_X1 U16035 ( .A1(n15362), .A2(n15353), .ZN(n15356) );
  AOI21_X1 U16036 ( .B1(n15356), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12742) );
  NAND2_X1 U16037 ( .A1(n20683), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14707) );
  OAI21_X1 U16038 ( .B1(n12743), .B2(n12742), .A(n14707), .ZN(n12744) );
  INV_X1 U16039 ( .A(n12744), .ZN(n12745) );
  OAI211_X1 U16040 ( .C1(n14712), .C2(n20666), .A(n12746), .B(n12745), .ZN(
        P1_U3001) );
  NOR2_X1 U16041 ( .A1(n12747), .A2(n16160), .ZN(n12752) );
  INV_X1 U16042 ( .A(n12748), .ZN(n12750) );
  NOR2_X1 U16043 ( .A1(n12750), .A2(n12749), .ZN(n12751) );
  XNOR2_X1 U16044 ( .A(n12752), .B(n12751), .ZN(n12832) );
  NAND2_X1 U16045 ( .A1(n12832), .A2(n19726), .ZN(n12768) );
  AOI21_X1 U16046 ( .B1(n12754), .B2(n15600), .A(n12753), .ZN(n14690) );
  INV_X1 U16047 ( .A(n12758), .ZN(n12761) );
  INV_X1 U16048 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20445) );
  NOR2_X1 U16049 ( .A1(n19705), .A2(n20445), .ZN(n12835) );
  NOR3_X1 U16050 ( .A1(n16446), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n12759), .ZN(n12760) );
  AOI211_X1 U16051 ( .C1(n12761), .C2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12835), .B(n12760), .ZN(n12762) );
  NAND3_X1 U16052 ( .A1(n12768), .A2(n10473), .A3(n12767), .ZN(P2_U3016) );
  NAND2_X1 U16053 ( .A1(n12769), .A2(n20699), .ZN(n12775) );
  OAI21_X1 U16054 ( .B1(n14839), .B2(n12770), .A(n14812), .ZN(n15033) );
  OR2_X1 U16055 ( .A1(n15033), .A2(n20668), .ZN(n12774) );
  NOR2_X1 U16056 ( .A1(n15403), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12771) );
  AOI211_X1 U16057 ( .C1(n15406), .C2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12772), .B(n12771), .ZN(n12773) );
  NAND2_X1 U16058 ( .A1(n12775), .A2(n10464), .ZN(P1_U3010) );
  INV_X1 U16059 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12776) );
  XNOR2_X1 U16060 ( .A(n12779), .B(n12778), .ZN(n12912) );
  AND2_X1 U16061 ( .A1(n13625), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12780) );
  AOI21_X1 U16062 ( .B1(n13240), .B2(P1_EBX_REG_31__SCAN_IN), .A(n12780), .ZN(
        n12783) );
  XOR2_X1 U16063 ( .A(n12783), .B(n12781), .Z(n12785) );
  NOR2_X1 U16064 ( .A1(n12783), .A2(n12782), .ZN(n12784) );
  MUX2_X1 U16065 ( .A(n12785), .B(n12784), .S(n14731), .Z(n15022) );
  INV_X1 U16066 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21358) );
  NOR2_X1 U16067 ( .A1(n20667), .A2(n21358), .ZN(n12907) );
  NAND4_X1 U16068 ( .A1(n15356), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n12778), .ZN(n12787) );
  OAI21_X1 U16069 ( .B1(n12912), .B2(n20666), .A(n12788), .ZN(P1_U3000) );
  INV_X1 U16070 ( .A(n19719), .ZN(n12789) );
  NAND2_X1 U16071 ( .A1(n16733), .A2(n12803), .ZN(n12790) );
  NAND2_X1 U16072 ( .A1(n16635), .A2(n12790), .ZN(n16572) );
  AOI21_X1 U16073 ( .B1(n12792), .B2(n12791), .A(n16572), .ZN(n12793) );
  INV_X1 U16074 ( .A(n12796), .ZN(n12797) );
  AOI21_X1 U16075 ( .B1(n12798), .B2(n12795), .A(n12797), .ZN(n16261) );
  OAI21_X1 U16076 ( .B1(n12799), .B2(n12802), .A(n12801), .ZN(n16127) );
  OR2_X1 U16077 ( .A1(n19705), .A2(n20420), .ZN(n16258) );
  OAI21_X1 U16078 ( .B1(n16127), .B2(n16722), .A(n16258), .ZN(n12805) );
  NOR2_X1 U16079 ( .A1(n12803), .A2(n16662), .ZN(n16545) );
  INV_X1 U16080 ( .A(n16545), .ZN(n16569) );
  OAI21_X1 U16081 ( .B1(n16286), .B2(n16710), .A(n16569), .ZN(n12804) );
  AOI21_X1 U16082 ( .B1(n12808), .B2(n12807), .A(n12806), .ZN(n16265) );
  XNOR2_X1 U16083 ( .A(n12815), .B(n10448), .ZN(n12841) );
  NAND2_X1 U16084 ( .A1(n12841), .A2(n19726), .ZN(n12831) );
  INV_X1 U16085 ( .A(n12816), .ZN(n12823) );
  NOR2_X1 U16086 ( .A1(n16353), .A2(n12823), .ZN(n16235) );
  OAI21_X1 U16087 ( .B1(n16235), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16227), .ZN(n12846) );
  NAND2_X1 U16088 ( .A1(n12817), .A2(n15714), .ZN(n15713) );
  INV_X1 U16089 ( .A(n15688), .ZN(n12818) );
  AOI21_X1 U16090 ( .B1(n12819), .B2(n15713), .A(n12818), .ZN(n15701) );
  OR2_X1 U16091 ( .A1(n15720), .A2(n12821), .ZN(n12822) );
  NAND2_X1 U16092 ( .A1(n12820), .A2(n12822), .ZN(n15706) );
  INV_X1 U16093 ( .A(n16509), .ZN(n12825) );
  NOR2_X1 U16094 ( .A1(n19705), .A2(n20426), .ZN(n12842) );
  NOR3_X1 U16095 ( .A1(n12823), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n16662), .ZN(n12824) );
  AOI211_X1 U16096 ( .C1(n12825), .C2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12842), .B(n12824), .ZN(n12826) );
  OAI21_X1 U16097 ( .B1(n15706), .B2(n16722), .A(n12826), .ZN(n12827) );
  AOI21_X1 U16098 ( .B1(n15701), .B2(n19712), .A(n12827), .ZN(n12828) );
  NAND2_X1 U16099 ( .A1(n12831), .A2(n12830), .ZN(P2_U3025) );
  NAND2_X1 U16100 ( .A1(n12832), .A2(n16394), .ZN(n12840) );
  INV_X1 U16101 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12833) );
  NOR2_X1 U16102 ( .A1(n16419), .A2(n12833), .ZN(n12834) );
  AOI211_X1 U16103 ( .C1(n14682), .C2(n16425), .A(n12835), .B(n12834), .ZN(
        n12836) );
  OAI21_X1 U16104 ( .B1(n14687), .B2(n16429), .A(n12836), .ZN(n12837) );
  INV_X1 U16105 ( .A(n12837), .ZN(n12838) );
  NAND3_X1 U16106 ( .A1(n12840), .A2(n12839), .A3(n12838), .ZN(P2_U2984) );
  NAND2_X1 U16107 ( .A1(n12841), .A2(n16394), .ZN(n12849) );
  AOI21_X1 U16108 ( .B1(n16354), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n12842), .ZN(n12843) );
  OAI21_X1 U16109 ( .B1(n15703), .B2(n16406), .A(n12843), .ZN(n12844) );
  AOI21_X1 U16110 ( .B1(n15701), .B2(n16409), .A(n12844), .ZN(n12845) );
  NAND2_X1 U16111 ( .A1(n12849), .A2(n12848), .ZN(P2_U2993) );
  NAND2_X1 U16112 ( .A1(n12850), .A2(n14734), .ZN(n12851) );
  NAND2_X1 U16113 ( .A1(n12872), .A2(n12851), .ZN(n15159) );
  AOI22_X1 U16114 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12885), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12856) );
  AOI22_X1 U16115 ( .A1(n11410), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12855) );
  AOI22_X1 U16116 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12854) );
  AOI22_X1 U16117 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12853) );
  NAND4_X1 U16118 ( .A1(n12856), .A2(n12855), .A3(n12854), .A4(n12853), .ZN(
        n12863) );
  AOI22_X1 U16119 ( .A1(n11411), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12861) );
  AOI22_X1 U16120 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12860) );
  AOI22_X1 U16121 ( .A1(n12887), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12859) );
  AOI22_X1 U16122 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12857), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12858) );
  NAND4_X1 U16123 ( .A1(n12861), .A2(n12860), .A3(n12859), .A4(n12858), .ZN(
        n12862) );
  NOR2_X1 U16124 ( .A1(n12863), .A2(n12862), .ZN(n12875) );
  NAND2_X1 U16125 ( .A1(n12865), .A2(n12864), .ZN(n12874) );
  XNOR2_X1 U16126 ( .A(n12875), .B(n12874), .ZN(n12869) );
  NAND2_X1 U16127 ( .A1(n21239), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12867) );
  NAND2_X1 U16128 ( .A1(n12904), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12866) );
  OAI211_X1 U16129 ( .C1(n12869), .C2(n12868), .A(n12867), .B(n12866), .ZN(
        n12870) );
  MUX2_X1 U16130 ( .A(n15159), .B(n12870), .S(n12902), .Z(n14730) );
  INV_X1 U16131 ( .A(n12872), .ZN(n12873) );
  XNOR2_X1 U16132 ( .A(n12873), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14708) );
  INV_X1 U16133 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n15067) );
  NOR2_X1 U16134 ( .A1(n12875), .A2(n12874), .ZN(n12895) );
  AOI22_X1 U16135 ( .A1(n11411), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11431), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12884) );
  AOI22_X1 U16136 ( .A1(n12877), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12876), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12883) );
  AOI22_X1 U16137 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12878), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12882) );
  AOI22_X1 U16138 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12880), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12881) );
  NAND4_X1 U16139 ( .A1(n12884), .A2(n12883), .A3(n12882), .A4(n12881), .ZN(
        n12893) );
  AOI22_X1 U16140 ( .A1(n11423), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12891) );
  AOI22_X1 U16141 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U16142 ( .A1(n12885), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12852), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12889) );
  AOI22_X1 U16143 ( .A1(n12887), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12886), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12888) );
  NAND4_X1 U16144 ( .A1(n12891), .A2(n12890), .A3(n12889), .A4(n12888), .ZN(
        n12892) );
  NOR2_X1 U16145 ( .A1(n12893), .A2(n12892), .ZN(n12894) );
  XNOR2_X1 U16146 ( .A(n12895), .B(n12894), .ZN(n12897) );
  NAND2_X1 U16147 ( .A1(n12897), .A2(n12896), .ZN(n12899) );
  OAI21_X1 U16148 ( .B1(n21191), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n21239), .ZN(n12898) );
  OAI211_X1 U16149 ( .C1(n12900), .C2(n15067), .A(n12899), .B(n12898), .ZN(
        n12901) );
  OAI21_X1 U16150 ( .B1(n14708), .B2(n12902), .A(n12901), .ZN(n14369) );
  AOI22_X1 U16151 ( .A1(n12904), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12903), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12905) );
  INV_X1 U16152 ( .A(n20712), .ZN(n20649) );
  AOI21_X1 U16153 ( .B1(n20641), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n12907), .ZN(n12908) );
  OAI21_X1 U16154 ( .B1(n20654), .B2(n12909), .A(n12908), .ZN(n12910) );
  AOI21_X1 U16155 ( .B1(n14721), .B2(n20649), .A(n12910), .ZN(n12911) );
  OAI21_X1 U16156 ( .B1(n12912), .B2(n15339), .A(n12911), .ZN(P1_U2968) );
  NAND2_X1 U16157 ( .A1(n15177), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15200) );
  INV_X1 U16158 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15385) );
  NAND2_X1 U16159 ( .A1(n15196), .A2(n20699), .ZN(n12922) );
  OAI21_X1 U16160 ( .B1(n14787), .B2(n12915), .A(n12914), .ZN(n15029) );
  INV_X1 U16161 ( .A(n12916), .ZN(n15370) );
  AND2_X1 U16162 ( .A1(n20683), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15195) );
  INV_X1 U16163 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12917) );
  AND3_X1 U16164 ( .A1(n12917), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12918) );
  AND2_X1 U16165 ( .A1(n15391), .A2(n12918), .ZN(n15369) );
  AOI211_X1 U16166 ( .C1(n15370), .C2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15195), .B(n15369), .ZN(n12919) );
  NAND2_X1 U16167 ( .A1(n12922), .A2(n12921), .ZN(P1_U3006) );
  NOR2_X1 U16168 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12924) );
  NOR4_X1 U16169 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12923) );
  NAND4_X1 U16170 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12924), .A4(n12923), .ZN(n12937) );
  NOR4_X1 U16171 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(
        P1_ADDRESS_REG_16__SCAN_IN), .A3(P1_ADDRESS_REG_15__SCAN_IN), .A4(
        P1_ADDRESS_REG_14__SCAN_IN), .ZN(n12928) );
  NOR4_X1 U16172 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(
        P1_ADDRESS_REG_20__SCAN_IN), .A3(P1_ADDRESS_REG_19__SCAN_IN), .A4(
        P1_ADDRESS_REG_18__SCAN_IN), .ZN(n12927) );
  NOR4_X1 U16173 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(
        P1_ADDRESS_REG_8__SCAN_IN), .A3(P1_ADDRESS_REG_7__SCAN_IN), .A4(
        P1_ADDRESS_REG_5__SCAN_IN), .ZN(n12926) );
  NOR4_X1 U16174 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(
        P1_ADDRESS_REG_12__SCAN_IN), .A3(P1_ADDRESS_REG_11__SCAN_IN), .A4(
        P1_ADDRESS_REG_10__SCAN_IN), .ZN(n12925) );
  AND4_X1 U16175 ( .A1(n12928), .A2(n12927), .A3(n12926), .A4(n12925), .ZN(
        n12933) );
  NOR4_X1 U16176 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_6__SCAN_IN), .A4(
        P1_ADDRESS_REG_2__SCAN_IN), .ZN(n12931) );
  NOR4_X1 U16177 ( .A1(P1_ADDRESS_REG_25__SCAN_IN), .A2(
        P1_ADDRESS_REG_24__SCAN_IN), .A3(P1_ADDRESS_REG_23__SCAN_IN), .A4(
        P1_ADDRESS_REG_22__SCAN_IN), .ZN(n12930) );
  NOR4_X1 U16178 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(
        P1_ADDRESS_REG_28__SCAN_IN), .A3(P1_ADDRESS_REG_27__SCAN_IN), .A4(
        P1_ADDRESS_REG_26__SCAN_IN), .ZN(n12929) );
  INV_X1 U16179 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n21319) );
  AND4_X1 U16180 ( .A1(n12931), .A2(n12930), .A3(n12929), .A4(n21319), .ZN(
        n12932) );
  NAND2_X1 U16181 ( .A1(n12933), .A2(n12932), .ZN(n12934) );
  INV_X1 U16182 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21374) );
  NOR3_X1 U16183 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21374), .ZN(n12936) );
  NOR4_X1 U16184 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12935) );
  NAND4_X1 U16185 ( .A1(n20709), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12936), .A4(
        n12935), .ZN(U214) );
  NOR2_X1 U16186 ( .A1(n16770), .A2(n12937), .ZN(n17432) );
  NAND2_X1 U16187 ( .A1(n17432), .A2(U214), .ZN(U212) );
  AND2_X1 U16188 ( .A1(n12946), .A2(n20381), .ZN(n17418) );
  NAND2_X1 U16189 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n14155) );
  NAND2_X1 U16190 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16742), .ZN(n14140) );
  INV_X1 U16191 ( .A(n14140), .ZN(n17419) );
  AOI221_X1 U16192 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .C1(P2_STATE2_REG_0__SCAN_IN), .C2(
        P2_STATE2_REG_1__SCAN_IN), .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n12938)
         );
  NOR3_X1 U16193 ( .A1(n17418), .A2(n17419), .A3(n12938), .ZN(P2_U3178) );
  INV_X1 U16194 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21304) );
  INV_X1 U16195 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21310) );
  NOR2_X1 U16196 ( .A1(n21312), .A2(n21310), .ZN(n21306) );
  INV_X1 U16197 ( .A(HOLD), .ZN(n21300) );
  NOR2_X1 U16198 ( .A1(n21304), .A2(n21300), .ZN(n21302) );
  OAI22_X1 U16199 ( .A1(n21306), .A2(n21302), .B1(n21315), .B2(n21300), .ZN(
        n12939) );
  OAI211_X1 U16200 ( .C1(n21304), .C2(n21308), .A(n12939), .B(n14051), .ZN(
        P1_U3195) );
  NOR2_X1 U16201 ( .A1(n12498), .A2(n17428), .ZN(n14149) );
  NAND2_X1 U16202 ( .A1(n14149), .A2(n12951), .ZN(n15927) );
  INV_X1 U16203 ( .A(n15927), .ZN(n15940) );
  INV_X1 U16204 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12942) );
  AND2_X1 U16205 ( .A1(n20463), .A2(n16757), .ZN(n12943) );
  INV_X1 U16206 ( .A(n12943), .ZN(n12940) );
  OAI211_X1 U16207 ( .C1(n15940), .C2(n12942), .A(n12941), .B(n12940), .ZN(
        P2_U2814) );
  INV_X1 U16208 ( .A(n15586), .ZN(n12945) );
  OAI21_X1 U16209 ( .B1(n12943), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n15590), 
        .ZN(n12944) );
  OAI21_X1 U16210 ( .B1(n12945), .B2(n15590), .A(n12944), .ZN(P2_U3612) );
  AOI22_X1 U16211 ( .A1(n15590), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n20462), 
        .B2(n12946), .ZN(n12947) );
  INV_X1 U16212 ( .A(n12947), .ZN(P2_U2816) );
  NOR3_X1 U16213 ( .A1(n12950), .A2(n12949), .A3(n12948), .ZN(n14125) );
  NOR2_X1 U16214 ( .A1(n14125), .A2(n17428), .ZN(n19581) );
  INV_X1 U16215 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n12959) );
  INV_X1 U16216 ( .A(n13807), .ZN(n12953) );
  INV_X1 U16217 ( .A(n12951), .ZN(n12952) );
  AOI22_X1 U16218 ( .A1(n13806), .A2(n12953), .B1(n12952), .B2(n12509), .ZN(
        n12954) );
  OAI21_X1 U16219 ( .B1(n13806), .B2(n13808), .A(n12954), .ZN(n14124) );
  AOI21_X1 U16220 ( .B1(n12955), .B2(n9595), .A(n17415), .ZN(n12956) );
  NOR2_X1 U16221 ( .A1(n12956), .A2(n14119), .ZN(n12957) );
  OAI21_X1 U16222 ( .B1(n14124), .B2(n12957), .A(n19581), .ZN(n12958) );
  OAI21_X1 U16223 ( .B1(n19581), .B2(n12959), .A(n12958), .ZN(P2_U3609) );
  NAND2_X1 U16224 ( .A1(n21239), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14060) );
  INV_X1 U16225 ( .A(n15565), .ZN(n15575) );
  NAND2_X1 U16226 ( .A1(n14213), .A2(n15002), .ZN(n12962) );
  NAND2_X1 U16227 ( .A1(n12960), .A2(n11979), .ZN(n12961) );
  NAND2_X1 U16228 ( .A1(n12962), .A2(n12961), .ZN(n12968) );
  OAI21_X1 U16229 ( .B1(n12968), .B2(n14227), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n12963) );
  OAI21_X1 U16230 ( .B1(n14060), .B2(n15575), .A(n12963), .ZN(P1_U2803) );
  AND2_X1 U16231 ( .A1(n21163), .A2(n14650), .ZN(n14718) );
  AOI211_X1 U16232 ( .C1(P1_MEMORYFETCH_REG_SCAN_IN), .C2(n12965), .A(n14718), 
        .B(n12980), .ZN(n12966) );
  INV_X1 U16233 ( .A(n12966), .ZN(P1_U2801) );
  NAND3_X1 U16234 ( .A1(n15002), .A2(n14051), .A3(n13625), .ZN(n12967) );
  AND2_X1 U16235 ( .A1(n12967), .A2(n21308), .ZN(n21383) );
  OR2_X1 U16236 ( .A1(n12968), .A2(n21383), .ZN(n14044) );
  NAND2_X1 U16237 ( .A1(n14044), .A2(n13609), .ZN(n20489) );
  INV_X1 U16238 ( .A(n20489), .ZN(n12978) );
  INV_X1 U16239 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n12977) );
  AND3_X1 U16240 ( .A1(n13981), .A2(n9764), .A3(n12969), .ZN(n12970) );
  MUX2_X1 U16241 ( .A(n13982), .B(n12970), .S(n14213), .Z(n12974) );
  NAND2_X1 U16242 ( .A1(n12972), .A2(n12971), .ZN(n12973) );
  NAND2_X1 U16243 ( .A1(n12974), .A2(n12973), .ZN(n12975) );
  OR2_X1 U16244 ( .A1(n14043), .A2(n20489), .ZN(n12976) );
  OAI21_X1 U16245 ( .B1(n12978), .B2(n12977), .A(n12976), .ZN(P1_U3484) );
  NAND2_X1 U16246 ( .A1(n12980), .A2(n20733), .ZN(n20639) );
  INV_X1 U16247 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20602) );
  INV_X1 U16248 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n12982) );
  INV_X1 U16249 ( .A(DATAI_15_), .ZN(n12981) );
  INV_X1 U16250 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13971) );
  MUX2_X1 U16251 ( .A(n12981), .B(n13971), .S(n20709), .Z(n15140) );
  OAI222_X1 U16252 ( .A1(n20639), .A2(n20602), .B1(n12982), .B2(n13550), .C1(
        n20633), .C2(n15140), .ZN(P1_U2967) );
  NOR2_X1 U16253 ( .A1(n17217), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12983) );
  AND2_X2 U16254 ( .A1(n13426), .A2(n12983), .ZN(n13507) );
  INV_X4 U16255 ( .A(n18006), .ZN(n18108) );
  AND2_X2 U16256 ( .A1(n13426), .A2(n12984), .ZN(n18002) );
  INV_X2 U16257 ( .A(n18002), .ZN(n17276) );
  AOI22_X1 U16258 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18107), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12990) );
  INV_X1 U16259 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12985) );
  OR2_X1 U16260 ( .A1(n14333), .A2(n12985), .ZN(n12989) );
  INV_X2 U16261 ( .A(n13034), .ZN(n18106) );
  NAND2_X1 U16262 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12988) );
  NAND2_X1 U16263 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12987) );
  NAND4_X1 U16264 ( .A1(n12990), .A2(n12989), .A3(n12988), .A4(n12987), .ZN(
        n12995) );
  NAND2_X1 U16265 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12993) );
  NAND2_X2 U16266 ( .A1(n12991), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n18077) );
  NAND2_X1 U16267 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12992) );
  OAI211_X1 U16268 ( .C1(n9640), .C2(n18127), .A(n12993), .B(n12992), .ZN(
        n12994) );
  NOR2_X1 U16269 ( .A1(n12995), .A2(n12994), .ZN(n13006) );
  AOI22_X1 U16270 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13004) );
  AOI22_X1 U16271 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17312), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13003) );
  NOR2_X1 U16272 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12998) );
  INV_X2 U16273 ( .A(n13095), .ZN(n18101) );
  AOI22_X1 U16274 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13002) );
  INV_X2 U16275 ( .A(n18085), .ZN(n17300) );
  AOI22_X1 U16276 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13001) );
  AND2_X2 U16277 ( .A1(n13006), .A2(n13005), .ZN(n16838) );
  INV_X1 U16278 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13009) );
  NAND2_X1 U16279 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13008) );
  NAND2_X1 U16280 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n13007) );
  OAI211_X1 U16281 ( .C1(n13009), .C2(n14333), .A(n13008), .B(n13007), .ZN(
        n13010) );
  INV_X1 U16282 ( .A(n13010), .ZN(n13014) );
  AOI22_X1 U16283 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13061), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13013) );
  INV_X2 U16284 ( .A(n17276), .ZN(n17953) );
  AOI22_X1 U16285 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13012) );
  NAND2_X1 U16286 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n13011) );
  NAND4_X1 U16287 ( .A1(n13014), .A2(n13013), .A3(n13012), .A4(n13011), .ZN(
        n13020) );
  INV_X1 U16288 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17320) );
  AOI22_X1 U16289 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17312), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13018) );
  INV_X2 U16290 ( .A(n10444), .ZN(n18100) );
  AOI22_X1 U16291 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13017) );
  AOI22_X1 U16292 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13016) );
  AOI22_X1 U16293 ( .A1(n13361), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13015) );
  NAND4_X1 U16294 ( .A1(n13018), .A2(n13017), .A3(n13016), .A4(n13015), .ZN(
        n13019) );
  OR2_X2 U16295 ( .A1(n13020), .A2(n13019), .ZN(n18996) );
  INV_X2 U16296 ( .A(n14333), .ZN(n13207) );
  AOI22_X1 U16297 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13061), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13027) );
  NAND2_X1 U16298 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n13023) );
  NAND2_X1 U16299 ( .A1(n17953), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n13022) );
  NAND2_X1 U16300 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n13021) );
  AOI22_X1 U16301 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13025) );
  NAND2_X1 U16302 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n13024) );
  NAND4_X1 U16303 ( .A1(n13027), .A2(n13026), .A3(n13025), .A4(n13024), .ZN(
        n13033) );
  AOI22_X1 U16304 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13031) );
  AOI22_X1 U16305 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17312), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13030) );
  AOI22_X1 U16306 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13029) );
  INV_X2 U16307 ( .A(n10444), .ZN(n17266) );
  AOI22_X1 U16308 ( .A1(n17266), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13028) );
  NAND4_X1 U16309 ( .A1(n13031), .A2(n13030), .A3(n13029), .A4(n13028), .ZN(
        n13032) );
  INV_X1 U16310 ( .A(n13061), .ZN(n13034) );
  AOI22_X1 U16311 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17322), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13041) );
  NAND2_X1 U16312 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n13037) );
  NAND2_X1 U16313 ( .A1(n17953), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n13036) );
  NAND2_X1 U16314 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n13035) );
  AOI22_X1 U16315 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13039) );
  NAND2_X1 U16316 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n13038) );
  NAND4_X1 U16317 ( .A1(n13041), .A2(n13040), .A3(n13039), .A4(n13038), .ZN(
        n13047) );
  AOI22_X1 U16318 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13045) );
  AOI22_X1 U16319 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17312), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13044) );
  AOI22_X1 U16320 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13043) );
  AOI22_X1 U16321 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17266), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13042) );
  NAND4_X1 U16322 ( .A1(n13045), .A2(n13044), .A3(n13043), .A4(n13042), .ZN(
        n13046) );
  OR2_X2 U16323 ( .A1(n13047), .A2(n13046), .ZN(n19010) );
  NAND2_X1 U16324 ( .A1(n18992), .A2(n19010), .ZN(n13369) );
  AOI22_X1 U16325 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13052) );
  AOI22_X1 U16326 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13051) );
  INV_X1 U16327 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18075) );
  NAND2_X1 U16328 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n13048) );
  NAND2_X1 U16329 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13049) );
  AOI22_X1 U16330 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13057) );
  INV_X4 U16331 ( .A(n10446), .ZN(n18099) );
  INV_X2 U16332 ( .A(n13229), .ZN(n17299) );
  AOI22_X1 U16333 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13056) );
  AOI22_X1 U16334 ( .A1(n13053), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U16335 ( .A1(n17266), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13054) );
  NAND2_X1 U16336 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n13060) );
  NAND2_X1 U16337 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13059) );
  NAND2_X1 U16338 ( .A1(n14312), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n13058) );
  AOI22_X1 U16339 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13061), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13064) );
  AOI22_X1 U16340 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18107), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13063) );
  NAND2_X1 U16341 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n13062) );
  NAND4_X1 U16342 ( .A1(n13065), .A2(n13064), .A3(n13063), .A4(n13062), .ZN(
        n13071) );
  AOI22_X1 U16343 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13069) );
  AOI22_X1 U16344 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17312), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13068) );
  AOI22_X1 U16345 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13067) );
  AOI22_X1 U16346 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13066) );
  NAND4_X1 U16347 ( .A1(n13069), .A2(n13068), .A3(n13067), .A4(n13066), .ZN(
        n13070) );
  MUX2_X1 U16348 ( .A(n13074), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n13182) );
  NAND2_X1 U16349 ( .A1(n19407), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13082) );
  NAND2_X1 U16350 ( .A1(n13182), .A2(n13181), .ZN(n13076) );
  NAND2_X1 U16351 ( .A1(n13074), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13075) );
  NAND2_X1 U16352 ( .A1(n13076), .A2(n13075), .ZN(n13085) );
  MUX2_X1 U16353 ( .A(n13077), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13084) );
  NAND2_X1 U16354 ( .A1(n13085), .A2(n13084), .ZN(n13079) );
  NAND2_X1 U16355 ( .A1(n13077), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13078) );
  NAND2_X1 U16356 ( .A1(n13079), .A2(n13078), .ZN(n13080) );
  OAI22_X1 U16357 ( .A1(n13080), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n19395), .ZN(n13087) );
  NOR2_X1 U16358 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19395), .ZN(
        n13081) );
  NAND2_X1 U16359 ( .A1(n13080), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13086) );
  AOI22_X1 U16360 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13087), .B1(
        n13081), .B2(n13086), .ZN(n13093) );
  OAI21_X1 U16361 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19407), .A(
        n13082), .ZN(n13083) );
  INV_X1 U16362 ( .A(n13083), .ZN(n13386) );
  XNOR2_X1 U16363 ( .A(n13085), .B(n13084), .ZN(n13092) );
  INV_X1 U16364 ( .A(n13093), .ZN(n13091) );
  NAND2_X1 U16365 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13086), .ZN(
        n13090) );
  INV_X1 U16366 ( .A(n13087), .ZN(n13089) );
  NAND2_X1 U16367 ( .A1(n13186), .A2(n13392), .ZN(n13370) );
  NOR2_X1 U16368 ( .A1(n16838), .A2(n19001), .ZN(n13196) );
  INV_X1 U16369 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13661) );
  AOI22_X1 U16370 ( .A1(n17299), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18100), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13099) );
  AOI22_X1 U16371 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13098) );
  AOI22_X1 U16372 ( .A1(n9568), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13053), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13097) );
  AOI22_X1 U16373 ( .A1(n14312), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13096) );
  AOI22_X1 U16374 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13103) );
  INV_X1 U16375 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17275) );
  OR2_X1 U16376 ( .A1(n14333), .A2(n17275), .ZN(n13102) );
  NAND2_X1 U16377 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13101) );
  NAND2_X1 U16378 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13100) );
  NAND2_X1 U16379 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13106) );
  NAND2_X1 U16380 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13105) );
  NAND2_X1 U16381 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13104) );
  AOI22_X1 U16382 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17322), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13115) );
  AOI22_X1 U16383 ( .A1(n18008), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13114) );
  INV_X1 U16384 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17291) );
  NAND2_X1 U16385 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13110) );
  NAND2_X1 U16386 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13109) );
  OAI211_X1 U16387 ( .C1(n14333), .C2(n17291), .A(n13110), .B(n13109), .ZN(
        n13111) );
  INV_X1 U16388 ( .A(n13111), .ZN(n13113) );
  NAND2_X1 U16389 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13112) );
  NAND4_X1 U16390 ( .A1(n13115), .A2(n13114), .A3(n13113), .A4(n13112), .ZN(
        n13121) );
  AOI22_X1 U16391 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18100), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U16392 ( .A1(n17299), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13118) );
  AOI22_X1 U16393 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13117) );
  AOI22_X1 U16394 ( .A1(n13361), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13053), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13116) );
  NAND4_X1 U16395 ( .A1(n13119), .A2(n13118), .A3(n13117), .A4(n13116), .ZN(
        n13120) );
  NAND2_X1 U16396 ( .A1(n18985), .A2(n19561), .ZN(n13122) );
  NOR2_X1 U16397 ( .A1(n19554), .A2(n13122), .ZN(n13123) );
  INV_X1 U16398 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13227) );
  INV_X1 U16399 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17916) );
  NAND2_X1 U16400 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n18144) );
  OAI21_X1 U16401 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n18144), .ZN(n17920) );
  OAI222_X1 U16402 ( .A1(n18148), .A2(n13227), .B1(n18154), .B2(n17916), .C1(
        n17233), .C2(n17920), .ZN(P3_U2702) );
  AOI22_X1 U16403 ( .A1(n13207), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13125) );
  AOI22_X1 U16404 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18107), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13124) );
  OAI211_X1 U16405 ( .C1(n18112), .C2(n17320), .A(n13125), .B(n13124), .ZN(
        n13133) );
  INV_X1 U16406 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18135) );
  AOI22_X1 U16407 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13126) );
  OAI21_X1 U16408 ( .B1(n17239), .B2(n18135), .A(n13126), .ZN(n13132) );
  AOI22_X1 U16409 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13130) );
  AOI22_X1 U16410 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13129) );
  AOI22_X1 U16411 ( .A1(n13053), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13128) );
  AOI22_X1 U16412 ( .A1(n17266), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13127) );
  NAND4_X1 U16413 ( .A1(n13130), .A2(n13129), .A3(n13128), .A4(n13127), .ZN(
        n13131) );
  NOR3_X1 U16414 ( .A1(n13133), .A2(n13132), .A3(n13131), .ZN(n16857) );
  NAND4_X1 U16415 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_9__SCAN_IN), .A4(P3_EBX_REG_8__SCAN_IN), .ZN(n13135) );
  INV_X1 U16416 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n18143) );
  NOR2_X1 U16417 ( .A1(n18143), .A2(n18144), .ZN(n18134) );
  NAND3_X1 U16418 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n18134), .ZN(n13134) );
  NAND4_X1 U16419 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(n18137), .ZN(n18122) );
  NOR2_X1 U16420 ( .A1(n13135), .A2(n18122), .ZN(n13537) );
  INV_X1 U16421 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17779) );
  NOR2_X1 U16422 ( .A1(n18151), .A2(n9653), .ZN(n13312) );
  OAI21_X1 U16423 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n13537), .A(n13312), .ZN(
        n13136) );
  OAI21_X1 U16424 ( .B1(n16857), .B2(n18148), .A(n13136), .ZN(P3_U2691) );
  XNOR2_X1 U16425 ( .A(n13137), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16728) );
  NOR2_X1 U16426 ( .A1(n16416), .A2(n10612), .ZN(n16730) );
  INV_X1 U16427 ( .A(n13138), .ZN(n13140) );
  NAND2_X1 U16428 ( .A1(n13140), .A2(n13139), .ZN(n13141) );
  XNOR2_X1 U16429 ( .A(n13141), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16727) );
  AND2_X1 U16430 ( .A1(n16394), .A2(n16727), .ZN(n13142) );
  AOI211_X1 U16431 ( .C1(n16728), .C2(n16415), .A(n16730), .B(n13142), .ZN(
        n13144) );
  MUX2_X1 U16432 ( .A(n16406), .B(n16419), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13143) );
  OAI211_X1 U16433 ( .C1(n13720), .C2(n16429), .A(n13144), .B(n13143), .ZN(
        P2_U3013) );
  INV_X1 U16434 ( .A(n13146), .ZN(n13147) );
  XNOR2_X1 U16435 ( .A(n13145), .B(n13147), .ZN(n16701) );
  INV_X1 U16436 ( .A(n16701), .ZN(n13155) );
  INV_X1 U16437 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19682) );
  INV_X1 U16438 ( .A(n16137), .ZN(n13151) );
  INV_X1 U16439 ( .A(n13149), .ZN(n13150) );
  INV_X1 U16440 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n13257) );
  OR2_X1 U16441 ( .A1(n16770), .A2(n13257), .ZN(n13153) );
  NAND2_X1 U16442 ( .A1(n16770), .A2(BUF2_REG_6__SCAN_IN), .ZN(n13152) );
  NAND2_X1 U16443 ( .A1(n13153), .A2(n13152), .ZN(n19797) );
  INV_X1 U16444 ( .A(n19797), .ZN(n13154) );
  OAI222_X1 U16445 ( .A1(n13155), .A2(n16156), .B1(n19682), .B2(n16151), .C1(
        n19655), .C2(n13154), .ZN(P2_U2913) );
  OR2_X1 U16446 ( .A1(n13159), .A2(n13158), .ZN(n13160) );
  NAND2_X1 U16447 ( .A1(n13157), .A2(n13160), .ZN(n16686) );
  INV_X1 U16448 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19680) );
  INV_X1 U16449 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13161) );
  OR2_X1 U16450 ( .A1(n16772), .A2(n13161), .ZN(n13163) );
  NAND2_X1 U16451 ( .A1(n16770), .A2(BUF2_REG_7__SCAN_IN), .ZN(n13162) );
  NAND2_X1 U16452 ( .A1(n13163), .A2(n13162), .ZN(n19810) );
  INV_X1 U16453 ( .A(n19810), .ZN(n13164) );
  OAI222_X1 U16454 ( .A1(n16686), .A2(n16156), .B1(n19680), .B2(n16151), .C1(
        n19655), .C2(n13164), .ZN(P2_U2912) );
  INV_X1 U16455 ( .A(n13165), .ZN(n13166) );
  AOI21_X1 U16456 ( .B1(n13167), .B2(n13157), .A(n13166), .ZN(n16675) );
  INV_X1 U16457 ( .A(n16675), .ZN(n13172) );
  INV_X1 U16458 ( .A(n19655), .ZN(n13793) );
  INV_X1 U16459 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n13168) );
  OR2_X1 U16460 ( .A1(n16770), .A2(n13168), .ZN(n13170) );
  NAND2_X1 U16461 ( .A1(n16772), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13169) );
  NAND2_X1 U16462 ( .A1(n13170), .A2(n13169), .ZN(n16083) );
  AOI22_X1 U16463 ( .A1(n13793), .A2(n16083), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n19647), .ZN(n13171) );
  OAI21_X1 U16464 ( .B1(n13172), .B2(n16156), .A(n13171), .ZN(P2_U2911) );
  NAND2_X1 U16465 ( .A1(n10593), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13173) );
  AOI21_X1 U16466 ( .B1(n15978), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13175) );
  AND2_X1 U16467 ( .A1(n13629), .A2(n13175), .ZN(n13176) );
  NOR2_X1 U16468 ( .A1(n13806), .A2(n13807), .ZN(n13823) );
  INV_X2 U16469 ( .A(n15999), .ZN(n16043) );
  NOR2_X1 U16470 ( .A1(n15938), .A2(n16043), .ZN(n13178) );
  AOI21_X1 U16471 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n16043), .A(n13178), .ZN(
        n13179) );
  OAI21_X1 U16472 ( .B1(n16799), .B2(n16029), .A(n13179), .ZN(P2_U2887) );
  NAND3_X1 U16473 ( .A1(n13180), .A2(n19554), .A3(n18298), .ZN(n13203) );
  XNOR2_X1 U16474 ( .A(n13182), .B(n13181), .ZN(n13183) );
  NAND2_X1 U16475 ( .A1(n13184), .A2(n13183), .ZN(n13387) );
  NAND2_X1 U16476 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19386) );
  NAND2_X1 U16477 ( .A1(n19401), .A2(n19386), .ZN(n13435) );
  INV_X1 U16478 ( .A(n13435), .ZN(n13202) );
  INV_X1 U16479 ( .A(n19001), .ZN(n13185) );
  NAND2_X1 U16480 ( .A1(n18295), .A2(n18985), .ZN(n13200) );
  INV_X1 U16481 ( .A(n16838), .ZN(n19005) );
  NAND2_X1 U16482 ( .A1(n19005), .A2(n19001), .ZN(n13188) );
  INV_X1 U16483 ( .A(n13188), .ZN(n13385) );
  NAND4_X1 U16484 ( .A1(n13385), .A2(n13186), .A3(n13189), .A4(n13375), .ZN(
        n13197) );
  NAND2_X1 U16485 ( .A1(n13188), .A2(n19010), .ZN(n13187) );
  NAND2_X1 U16486 ( .A1(n13187), .A2(n18996), .ZN(n13192) );
  OAI21_X1 U16487 ( .B1(n13380), .B2(n18989), .A(n13188), .ZN(n13191) );
  AND2_X1 U16488 ( .A1(n16838), .A2(n19001), .ZN(n13372) );
  NAND2_X1 U16489 ( .A1(n13372), .A2(n13189), .ZN(n13190) );
  NAND3_X1 U16490 ( .A1(n13192), .A2(n13191), .A3(n13190), .ZN(n13193) );
  INV_X1 U16491 ( .A(n13395), .ZN(n13195) );
  NAND2_X1 U16492 ( .A1(n13380), .A2(n17523), .ZN(n13433) );
  NAND2_X1 U16493 ( .A1(n13382), .A2(n13384), .ZN(n16807) );
  NAND2_X1 U16494 ( .A1(n13200), .A2(n16807), .ZN(n13201) );
  NAND2_X1 U16495 ( .A1(n13202), .A2(n13201), .ZN(n13438) );
  INV_X1 U16496 ( .A(n13219), .ZN(n13218) );
  NAND2_X1 U16497 ( .A1(n13218), .A2(n19010), .ZN(n18251) );
  INV_X1 U16498 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n13222) );
  INV_X1 U16499 ( .A(n13372), .ZN(n17215) );
  NOR2_X2 U16500 ( .A1(n13219), .A2(n17215), .ZN(n18249) );
  AOI22_X1 U16501 ( .A1(n18008), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17322), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13211) );
  NAND2_X1 U16502 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n13206) );
  NAND2_X1 U16503 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13205) );
  NAND2_X1 U16504 ( .A1(n13507), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13204) );
  AND3_X1 U16505 ( .A1(n13206), .A2(n13205), .A3(n13204), .ZN(n13210) );
  AOI22_X1 U16506 ( .A1(n18061), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13209) );
  NAND2_X1 U16507 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n13208) );
  NAND4_X1 U16508 ( .A1(n13211), .A2(n13210), .A3(n13209), .A4(n13208), .ZN(
        n13217) );
  AOI22_X1 U16509 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13215) );
  AOI22_X1 U16510 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13214) );
  AOI22_X1 U16511 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13213) );
  AOI22_X1 U16512 ( .A1(n17299), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18101), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13212) );
  NAND4_X1 U16513 ( .A1(n13215), .A2(n13214), .A3(n13213), .A4(n13212), .ZN(
        n13216) );
  NAND2_X1 U16514 ( .A1(n13218), .A2(n18157), .ZN(n18203) );
  AOI21_X1 U16515 ( .B1(n18203), .B2(n21512), .A(n13540), .ZN(n13220) );
  AOI21_X1 U16516 ( .B1(n18249), .B2(n13495), .A(n13220), .ZN(n13221) );
  OAI21_X1 U16517 ( .B1(n18255), .B2(n13222), .A(n13221), .ZN(P3_U2735) );
  INV_X1 U16518 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13225) );
  AOI22_X1 U16519 ( .A1(n13207), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13224) );
  AOI22_X1 U16520 ( .A1(n13507), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13223) );
  OAI211_X1 U16521 ( .C1(n18112), .C2(n13225), .A(n13224), .B(n13223), .ZN(
        n13236) );
  AOI22_X1 U16522 ( .A1(n18008), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13226) );
  OAI21_X1 U16523 ( .B1(n17239), .B2(n13227), .A(n13226), .ZN(n13235) );
  AOI22_X1 U16524 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13233) );
  AOI22_X1 U16525 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13232) );
  AOI22_X1 U16526 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13231) );
  AOI22_X1 U16527 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13230) );
  NAND4_X1 U16528 ( .A1(n13233), .A2(n13232), .A3(n13231), .A4(n13230), .ZN(
        n13234) );
  NOR3_X1 U16529 ( .A1(n13236), .A2(n13235), .A3(n13234), .ZN(n13546) );
  INV_X1 U16530 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n18119) );
  NOR2_X1 U16531 ( .A1(n18119), .A2(n18118), .ZN(n13238) );
  INV_X1 U16532 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17816) );
  NOR3_X1 U16533 ( .A1(n17816), .A2(n18119), .A3(n18118), .ZN(n18094) );
  NOR2_X1 U16534 ( .A1(n18094), .A2(n18151), .ZN(n13237) );
  OAI21_X1 U16535 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n13238), .A(n13237), .ZN(
        n13239) );
  OAI21_X1 U16536 ( .B1(n13546), .B2(n18148), .A(n13239), .ZN(P3_U2694) );
  NOR2_X1 U16537 ( .A1(n13240), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13241) );
  OR2_X1 U16538 ( .A1(n13242), .A2(n13241), .ZN(n15012) );
  NAND2_X1 U16539 ( .A1(n14213), .A2(n13297), .ZN(n13245) );
  NAND4_X1 U16540 ( .A1(n13243), .A2(n13980), .A3(n20763), .A4(n11385), .ZN(
        n13604) );
  NAND2_X1 U16541 ( .A1(n13245), .A2(n13244), .ZN(n13246) );
  INV_X1 U16542 ( .A(n13247), .ZN(n13250) );
  OAI21_X1 U16543 ( .B1(n13250), .B2(n13249), .A(n13248), .ZN(n15020) );
  INV_X2 U16544 ( .A(n20596), .ZN(n15055) );
  OAI222_X1 U16545 ( .A1(n15012), .A2(n20594), .B1(n21464), .B2(n20599), .C1(
        n15020), .C2(n15055), .ZN(P1_U2872) );
  AOI22_X1 U16546 ( .A1(n13601), .A2(P1_EAX_REG_24__SCAN_IN), .B1(n13268), 
        .B2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13253) );
  INV_X1 U16547 ( .A(DATAI_8_), .ZN(n13252) );
  NAND2_X1 U16548 ( .A1(n20709), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13251) );
  OAI21_X1 U16549 ( .B1(n20709), .B2(n13252), .A(n13251), .ZN(n15152) );
  NAND2_X1 U16550 ( .A1(n13587), .A2(n15152), .ZN(n13577) );
  NAND2_X1 U16551 ( .A1(n13253), .A2(n13577), .ZN(P1_U2945) );
  AOI22_X1 U16552 ( .A1(n13601), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n13268), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13256) );
  INV_X1 U16553 ( .A(DATAI_4_), .ZN(n13255) );
  NAND2_X1 U16554 ( .A1(n20709), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13254) );
  OAI21_X1 U16555 ( .B1(n20709), .B2(n13255), .A(n13254), .ZN(n15113) );
  NAND2_X1 U16556 ( .A1(n13587), .A2(n15113), .ZN(n13599) );
  NAND2_X1 U16557 ( .A1(n13256), .A2(n13599), .ZN(P1_U2941) );
  AOI22_X1 U16558 ( .A1(n13601), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n13268), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13260) );
  INV_X1 U16559 ( .A(DATAI_6_), .ZN(n13258) );
  MUX2_X1 U16560 ( .A(n13258), .B(n13257), .S(n20709), .Z(n20759) );
  INV_X1 U16561 ( .A(n20759), .ZN(n13259) );
  NAND2_X1 U16562 ( .A1(n13587), .A2(n13259), .ZN(n13591) );
  NAND2_X1 U16563 ( .A1(n13260), .A2(n13591), .ZN(P1_U2943) );
  AOI22_X1 U16564 ( .A1(n13601), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n13268), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13263) );
  INV_X1 U16565 ( .A(DATAI_9_), .ZN(n13261) );
  INV_X1 U16566 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13490) );
  MUX2_X1 U16567 ( .A(n13261), .B(n13490), .S(n20709), .Z(n15150) );
  INV_X1 U16568 ( .A(n15150), .ZN(n13262) );
  NAND2_X1 U16569 ( .A1(n13587), .A2(n13262), .ZN(n13595) );
  NAND2_X1 U16570 ( .A1(n13263), .A2(n13595), .ZN(P1_U2946) );
  AOI22_X1 U16571 ( .A1(n13601), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n13268), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13267) );
  NAND2_X1 U16572 ( .A1(n20711), .A2(DATAI_7_), .ZN(n13265) );
  NAND2_X1 U16573 ( .A1(n20709), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13264) );
  AND2_X1 U16574 ( .A1(n13265), .A2(n13264), .ZN(n20767) );
  INV_X1 U16575 ( .A(n20767), .ZN(n13266) );
  NAND2_X1 U16576 ( .A1(n13587), .A2(n13266), .ZN(n13589) );
  NAND2_X1 U16577 ( .A1(n13267), .A2(n13589), .ZN(P1_U2944) );
  AOI22_X1 U16578 ( .A1(n13601), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n13268), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13272) );
  NAND2_X1 U16579 ( .A1(n20711), .A2(DATAI_5_), .ZN(n13270) );
  NAND2_X1 U16580 ( .A1(n20709), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13269) );
  AND2_X1 U16581 ( .A1(n13270), .A2(n13269), .ZN(n20754) );
  INV_X1 U16582 ( .A(n20754), .ZN(n13271) );
  NAND2_X1 U16583 ( .A1(n13587), .A2(n13271), .ZN(n13593) );
  NAND2_X1 U16584 ( .A1(n13272), .A2(n13593), .ZN(P1_U2942) );
  INV_X1 U16585 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13275) );
  AOI22_X1 U16586 ( .A1(n13207), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13274) );
  AOI22_X1 U16587 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18107), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13273) );
  OAI211_X1 U16588 ( .C1(n18112), .C2(n13275), .A(n13274), .B(n13273), .ZN(
        n13283) );
  INV_X1 U16589 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18133) );
  AOI22_X1 U16590 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13276) );
  OAI21_X1 U16591 ( .B1(n17239), .B2(n18133), .A(n13276), .ZN(n13282) );
  AOI22_X1 U16592 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13280) );
  AOI22_X1 U16593 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13279) );
  AOI22_X1 U16594 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13278) );
  AOI22_X1 U16595 ( .A1(n17266), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13277) );
  NAND4_X1 U16596 ( .A1(n13280), .A2(n13279), .A3(n13278), .A4(n13277), .ZN(
        n13281) );
  NOR3_X1 U16597 ( .A1(n13283), .A2(n13282), .A3(n13281), .ZN(n16855) );
  INV_X1 U16598 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17767) );
  AOI22_X1 U16599 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n13312), .B1(n13657), 
        .B2(n17767), .ZN(n13284) );
  OAI21_X1 U16600 ( .B1(n16855), .B2(n18148), .A(n13284), .ZN(P3_U2690) );
  OR2_X1 U16601 ( .A1(n13286), .A2(n13287), .ZN(n13288) );
  NAND2_X1 U16602 ( .A1(n13285), .A2(n13288), .ZN(n16647) );
  INV_X1 U16603 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n17461) );
  OR2_X1 U16604 ( .A1(n16770), .A2(n17461), .ZN(n13290) );
  NAND2_X1 U16605 ( .A1(n16772), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13289) );
  NAND2_X1 U16606 ( .A1(n13290), .A2(n13289), .ZN(n16069) );
  AOI22_X1 U16607 ( .A1(n13793), .A2(n16069), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n19647), .ZN(n13291) );
  OAI21_X1 U16608 ( .B1(n16647), .B2(n16156), .A(n13291), .ZN(P2_U2909) );
  INV_X1 U16609 ( .A(n14649), .ZN(n13674) );
  NOR2_X1 U16610 ( .A1(n13293), .A2(n13292), .ZN(n13296) );
  AOI21_X1 U16611 ( .B1(n14058), .B2(n13294), .A(n13293), .ZN(n13608) );
  AOI22_X1 U16612 ( .A1(n13674), .A2(n13296), .B1(n13608), .B2(n13295), .ZN(
        n13298) );
  MUX2_X1 U16613 ( .A(n13298), .B(n13297), .S(n14213), .Z(n13304) );
  INV_X1 U16614 ( .A(n13299), .ZN(n13302) );
  INV_X1 U16615 ( .A(n13300), .ZN(n14035) );
  NAND2_X1 U16616 ( .A1(n14035), .A2(n13301), .ZN(n13606) );
  OAI211_X1 U16617 ( .C1(n11381), .C2(n15004), .A(n13302), .B(n13606), .ZN(
        n13303) );
  INV_X1 U16618 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n14031) );
  NAND2_X1 U16619 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n14220) );
  INV_X1 U16620 ( .A(n14220), .ZN(n15537) );
  NAND2_X1 U16621 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15537), .ZN(n15540) );
  NOR2_X1 U16622 ( .A1(n14031), .A2(n15540), .ZN(n13305) );
  AOI21_X1 U16623 ( .B1(n14037), .B2(n13609), .A(n13305), .ZN(n13309) );
  NAND2_X1 U16624 ( .A1(n10072), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13306) );
  INV_X1 U16625 ( .A(n15577), .ZN(n13311) );
  INV_X1 U16626 ( .A(n20872), .ZN(n21126) );
  OR2_X1 U16627 ( .A1(n13307), .A2(n21126), .ZN(n13308) );
  XNOR2_X1 U16628 ( .A(n13308), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14036) );
  INV_X1 U16629 ( .A(n14036), .ZN(n20552) );
  OR4_X1 U16630 ( .A1(n20552), .A2(n13309), .A3(n15575), .A4(n13300), .ZN(
        n13310) );
  OAI21_X1 U16631 ( .B1(n14039), .B2(n13311), .A(n13310), .ZN(P1_U3468) );
  NAND2_X1 U16632 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .ZN(n14323) );
  AOI21_X1 U16633 ( .B1(n18150), .B2(n14323), .A(n13312), .ZN(n13327) );
  AOI21_X1 U16634 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n13657), .A(
        P3_EBX_REG_14__SCAN_IN), .ZN(n13326) );
  AOI22_X1 U16635 ( .A1(n13207), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13319) );
  NAND2_X1 U16636 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n13315) );
  NAND2_X1 U16637 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n13314) );
  NAND2_X1 U16638 ( .A1(n13507), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n13313) );
  AND3_X1 U16639 ( .A1(n13315), .A2(n13314), .A3(n13313), .ZN(n13318) );
  INV_X1 U16640 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16882) );
  AOI22_X1 U16641 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13317) );
  NAND2_X1 U16642 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n13316) );
  NAND4_X1 U16643 ( .A1(n13319), .A2(n13318), .A3(n13317), .A4(n13316), .ZN(
        n13325) );
  AOI22_X1 U16644 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13323) );
  AOI22_X1 U16645 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13322) );
  AOI22_X1 U16646 ( .A1(n13053), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13321) );
  AOI22_X1 U16647 ( .A1(n17266), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13320) );
  NAND4_X1 U16648 ( .A1(n13323), .A2(n13322), .A3(n13321), .A4(n13320), .ZN(
        n13324) );
  NOR2_X1 U16649 ( .A1(n13325), .A2(n13324), .ZN(n18234) );
  OAI22_X1 U16650 ( .A1(n13327), .A2(n13326), .B1(n18234), .B2(n18148), .ZN(
        P3_U2689) );
  AOI22_X1 U16651 ( .A1(n18061), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17322), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13334) );
  NAND2_X1 U16652 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n13330) );
  NAND2_X1 U16653 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n13329) );
  NAND2_X1 U16654 ( .A1(n13507), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n13328) );
  AND3_X1 U16655 ( .A1(n13330), .A2(n13329), .A3(n13328), .ZN(n13333) );
  AOI22_X1 U16656 ( .A1(n18008), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13332) );
  NAND2_X1 U16657 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n13331) );
  AOI22_X1 U16658 ( .A1(n13228), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13338) );
  AOI22_X1 U16659 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17312), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13337) );
  AOI22_X1 U16660 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13336) );
  AOI22_X1 U16661 ( .A1(n17266), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13335) );
  INV_X1 U16662 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n21444) );
  NAND2_X1 U16663 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n13540), .ZN(n13503) );
  INV_X1 U16664 ( .A(n13503), .ZN(n13339) );
  AOI22_X1 U16665 ( .A1(n18251), .A2(P3_EAX_REG_2__SCAN_IN), .B1(n18157), .B2(
        n13339), .ZN(n13340) );
  OAI222_X1 U16666 ( .A1(n18197), .A2(n16958), .B1(n18255), .B2(n21444), .C1(
        n13340), .C2(n13353), .ZN(P3_U2733) );
  INV_X1 U16667 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18993) );
  AOI22_X1 U16668 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17322), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13346) );
  NAND2_X1 U16669 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13343) );
  NAND2_X1 U16670 ( .A1(n13507), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n13342) );
  NAND2_X1 U16671 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n13341) );
  AOI22_X1 U16672 ( .A1(n18061), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18100), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13345) );
  NAND2_X1 U16673 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n13344) );
  NAND4_X1 U16674 ( .A1(n13346), .A2(n10454), .A3(n13345), .A4(n13344), .ZN(
        n13352) );
  AOI22_X1 U16675 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13350) );
  AOI22_X1 U16676 ( .A1(n13053), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13349) );
  AOI22_X1 U16677 ( .A1(n17299), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13348) );
  AOI22_X1 U16678 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13347) );
  NAND4_X1 U16679 ( .A1(n13350), .A2(n13349), .A3(n13348), .A4(n13347), .ZN(
        n13351) );
  INV_X1 U16680 ( .A(n16960), .ZN(n16966) );
  NAND2_X1 U16681 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n13353), .ZN(n13522) );
  INV_X1 U16682 ( .A(n13522), .ZN(n13521) );
  AOI21_X1 U16683 ( .B1(n18251), .B2(P3_EAX_REG_3__SCAN_IN), .A(n13353), .ZN(
        n13354) );
  OAI222_X1 U16684 ( .A1(n18255), .A2(n18993), .B1(n18197), .B2(n16966), .C1(
        n13521), .C2(n13354), .ZN(P3_U2732) );
  AOI22_X1 U16685 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17322), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13360) );
  NAND2_X1 U16686 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13357) );
  NAND2_X1 U16687 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13356) );
  NAND2_X1 U16688 ( .A1(n13507), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13355) );
  AOI22_X1 U16689 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17266), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13359) );
  NAND2_X1 U16690 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13358) );
  NAND4_X1 U16691 ( .A1(n13360), .A2(n9682), .A3(n13359), .A4(n13358), .ZN(
        n13367) );
  AOI22_X1 U16692 ( .A1(n13361), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17312), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13365) );
  AOI22_X1 U16693 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13364) );
  AOI22_X1 U16694 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13363) );
  AOI22_X1 U16695 ( .A1(n14312), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13053), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13362) );
  NAND4_X1 U16696 ( .A1(n13365), .A2(n13364), .A3(n13363), .A4(n13362), .ZN(
        n13366) );
  XNOR2_X1 U16697 ( .A(n16904), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n16902) );
  AND2_X1 U16698 ( .A1(n13495), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18677) );
  NAND2_X1 U16699 ( .A1(n18678), .A2(n18677), .ZN(n18676) );
  INV_X1 U16700 ( .A(n13404), .ZN(n13506) );
  NAND2_X1 U16701 ( .A1(n13506), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13368) );
  NAND2_X1 U16702 ( .A1(n18676), .A2(n13368), .ZN(n16903) );
  XNOR2_X1 U16703 ( .A(n16902), .B(n16903), .ZN(n18665) );
  NAND2_X1 U16704 ( .A1(n13369), .A2(n18985), .ZN(n13417) );
  NAND2_X1 U16705 ( .A1(n13417), .A2(n13370), .ZN(n13371) );
  NAND2_X1 U16706 ( .A1(n13384), .A2(n13371), .ZN(n13379) );
  NOR2_X1 U16707 ( .A1(n19554), .A2(n18985), .ZN(n19388) );
  OAI21_X1 U16708 ( .B1(n13372), .B2(n18157), .A(n19388), .ZN(n13394) );
  NAND2_X1 U16709 ( .A1(n18992), .A2(n13373), .ZN(n13374) );
  OAI21_X1 U16710 ( .B1(n13375), .B2(n18992), .A(n13374), .ZN(n13376) );
  INV_X1 U16711 ( .A(n13376), .ZN(n13377) );
  NOR2_X1 U16712 ( .A1(n13380), .A2(n19388), .ZN(n19571) );
  INV_X1 U16713 ( .A(n13382), .ZN(n13383) );
  OR2_X2 U16714 ( .A1(n19406), .A2(n18958), .ZN(n18875) );
  INV_X2 U16715 ( .A(n18875), .ZN(n18839) );
  XNOR2_X1 U16716 ( .A(n18298), .B(n18989), .ZN(n13397) );
  NAND2_X1 U16717 ( .A1(n13744), .A2(n13385), .ZN(n13391) );
  OR2_X1 U16718 ( .A1(n13387), .A2(n13386), .ZN(n13388) );
  NAND2_X1 U16719 ( .A1(n13389), .A2(n13388), .ZN(n19400) );
  NAND3_X1 U16720 ( .A1(n19400), .A2(n18985), .A3(n19005), .ZN(n13390) );
  NAND2_X1 U16721 ( .A1(n13391), .A2(n13390), .ZN(n13393) );
  NAND2_X1 U16722 ( .A1(n13393), .A2(n13392), .ZN(n13402) );
  OAI211_X1 U16723 ( .C1(n17523), .C2(n13396), .A(n13395), .B(n13394), .ZN(
        n13436) );
  AOI21_X1 U16724 ( .B1(n13744), .B2(n18996), .A(n13436), .ZN(n13401) );
  INV_X1 U16725 ( .A(n19401), .ZN(n13398) );
  NOR2_X2 U16726 ( .A1(n19452), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n19524) );
  NOR2_X1 U16727 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19450) );
  OAI21_X1 U16728 ( .B1(n19553), .B2(n13397), .A(n19386), .ZN(n17522) );
  OR3_X1 U16729 ( .A1(n13399), .A2(n13398), .A3(n17522), .ZN(n13400) );
  NAND3_X1 U16730 ( .A1(n13402), .A2(n13401), .A3(n13400), .ZN(n13403) );
  INV_X1 U16731 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13410) );
  NAND2_X1 U16732 ( .A1(n13404), .A2(n13495), .ZN(n16959) );
  NOR2_X1 U16733 ( .A1(n13405), .A2(n13410), .ZN(n16970) );
  OAI21_X1 U16734 ( .B1(n13495), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13406) );
  NAND2_X1 U16735 ( .A1(n13406), .A2(n13506), .ZN(n13407) );
  OAI211_X1 U16736 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n13407), .B(n16959), .ZN(n16969) );
  XNOR2_X1 U16737 ( .A(n16968), .B(n16969), .ZN(n18670) );
  INV_X1 U16738 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17216) );
  NAND2_X1 U16739 ( .A1(n18861), .A2(n17216), .ZN(n18758) );
  INV_X1 U16740 ( .A(n18958), .ZN(n18784) );
  NAND2_X1 U16741 ( .A1(n18784), .A2(n18868), .ZN(n18759) );
  AOI211_X1 U16742 ( .C1(n18758), .C2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n18766), .B(n13410), .ZN(n13409) );
  INV_X1 U16743 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18956) );
  OAI21_X1 U16744 ( .B1(n18956), .B2(n17216), .A(n13410), .ZN(n18895) );
  NOR2_X1 U16745 ( .A1(n13410), .A2(n18956), .ZN(n18782) );
  NAND2_X1 U16746 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18782), .ZN(
        n18786) );
  INV_X1 U16747 ( .A(n19406), .ZN(n18896) );
  AOI21_X1 U16748 ( .B1(n18895), .B2(n18786), .A(n18896), .ZN(n13408) );
  AOI211_X1 U16749 ( .C1(n18670), .C2(n19404), .A(n13409), .B(n13408), .ZN(
        n13412) );
  OAI21_X1 U16750 ( .B1(n18868), .B2(n17216), .A(n18784), .ZN(n17163) );
  NAND3_X1 U16751 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17163), .A3(
        n13410), .ZN(n13411) );
  AOI21_X1 U16752 ( .B1(n13412), .B2(n13411), .A(n18899), .ZN(n13413) );
  INV_X1 U16753 ( .A(n13413), .ZN(n13416) );
  NOR2_X1 U16754 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n17930) );
  NOR2_X1 U16755 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n13414) );
  INV_X2 U16756 ( .A(n13496), .ZN(n18840) );
  INV_X1 U16757 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19469) );
  NOR2_X1 U16758 ( .A1(n18840), .A2(n19469), .ZN(n18669) );
  AOI21_X1 U16759 ( .B1(n18955), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18669), .ZN(n13415) );
  OAI211_X1 U16760 ( .C1(n18665), .C2(n18906), .A(n13416), .B(n13415), .ZN(
        P3_U2860) );
  INV_X1 U16761 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16954) );
  OAI22_X1 U16762 ( .A1(n16954), .A2(n18956), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17225) );
  INV_X1 U16763 ( .A(n17225), .ZN(n13432) );
  NOR2_X1 U16764 ( .A1(n19444), .A2(n17216), .ZN(n17226) );
  NOR2_X1 U16765 ( .A1(n16808), .A2(n13417), .ZN(n13423) );
  NAND2_X1 U16766 ( .A1(n13419), .A2(n13418), .ZN(n13420) );
  NAND2_X1 U16767 ( .A1(n13421), .A2(n13420), .ZN(n13422) );
  OR2_X1 U16768 ( .A1(n13423), .A2(n13422), .ZN(n13448) );
  NOR2_X1 U16769 ( .A1(n17220), .A2(n19391), .ZN(n13424) );
  NAND2_X1 U16770 ( .A1(n13448), .A2(n13424), .ZN(n13430) );
  INV_X1 U16771 ( .A(n17220), .ZN(n13425) );
  NAND2_X1 U16772 ( .A1(n13425), .A2(n19391), .ZN(n13449) );
  NAND2_X1 U16773 ( .A1(n13451), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13453) );
  NAND2_X1 U16774 ( .A1(n13449), .A2(n13453), .ZN(n17898) );
  AOI21_X1 U16775 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18861), .A(
        n18958), .ZN(n13446) );
  NOR2_X1 U16776 ( .A1(n13426), .A2(n13446), .ZN(n13428) );
  AOI22_X1 U16777 ( .A1(n19406), .A2(n17898), .B1(n13428), .B2(n13427), .ZN(
        n13429) );
  AND2_X1 U16778 ( .A1(n13430), .A2(n13429), .ZN(n19390) );
  INV_X1 U16779 ( .A(n17930), .ZN(n19570) );
  NAND2_X1 U16780 ( .A1(n17886), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n14332) );
  OAI22_X1 U16781 ( .A1(n19390), .A2(n19570), .B1(n14332), .B2(n17898), .ZN(
        n13431) );
  AOI21_X1 U16782 ( .B1(n13432), .B2(n17226), .A(n13431), .ZN(n13445) );
  INV_X1 U16783 ( .A(n19561), .ZN(n19430) );
  INV_X1 U16784 ( .A(n13433), .ZN(n13434) );
  OAI221_X1 U16785 ( .B1(n13434), .B2(n19388), .C1(n13434), .C2(n9649), .A(
        n19553), .ZN(n18256) );
  OR2_X1 U16786 ( .A1(n13435), .A2(n18256), .ZN(n13442) );
  INV_X1 U16787 ( .A(n13436), .ZN(n13437) );
  NAND2_X1 U16788 ( .A1(n13438), .A2(n13437), .ZN(n13439) );
  NOR2_X1 U16789 ( .A1(n13440), .A2(n13439), .ZN(n13441) );
  INV_X1 U16790 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19558) );
  NAND2_X1 U16791 ( .A1(n19558), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18976) );
  INV_X1 U16792 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n17525) );
  NAND3_X1 U16793 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_1__SCAN_IN), .ZN(n19538)
         );
  OR2_X1 U16794 ( .A1(n17525), .A2(n19538), .ZN(n13443) );
  OAI211_X1 U16795 ( .C1(n19430), .C2(n19426), .A(n18976), .B(n13443), .ZN(
        n17229) );
  INV_X1 U16796 ( .A(n17229), .ZN(n14330) );
  NAND2_X1 U16797 ( .A1(n14330), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13444) );
  OAI21_X1 U16798 ( .B1(n13445), .B2(n14330), .A(n13444), .ZN(P3_U3288) );
  INV_X1 U16799 ( .A(n13446), .ZN(n17222) );
  AOI22_X1 U16800 ( .A1(n19406), .A2(n13449), .B1(n13451), .B2(n17222), .ZN(
        n13447) );
  NOR2_X1 U16801 ( .A1(n13447), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n19398) );
  NAND2_X1 U16802 ( .A1(n13448), .A2(n13453), .ZN(n13450) );
  OAI211_X1 U16803 ( .C1(n13451), .C2(n18784), .A(n13450), .B(n13449), .ZN(
        n19396) );
  AOI22_X1 U16804 ( .A1(n17229), .A2(n19398), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19396), .ZN(n13457) );
  NAND2_X1 U16805 ( .A1(n13453), .A2(n13452), .ZN(n13454) );
  NAND2_X1 U16806 ( .A1(n10445), .A2(n13454), .ZN(n16828) );
  NOR3_X1 U16807 ( .A1(n14330), .A2(n16828), .A3(n14332), .ZN(n13455) );
  AOI21_X1 U16808 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n14330), .A(
        n13455), .ZN(n13456) );
  OAI21_X1 U16809 ( .B1(n13457), .B2(n19570), .A(n13456), .ZN(P3_U3285) );
  NAND3_X1 U16810 ( .A1(n13460), .A2(n13459), .A3(n13458), .ZN(n13461) );
  AOI21_X1 U16811 ( .B1(n20713), .B2(n13462), .A(n13461), .ZN(n13464) );
  NOR2_X1 U16812 ( .A1(n13464), .A2(n13463), .ZN(n13655) );
  OAI21_X1 U16813 ( .B1(n20641), .B2(n13465), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13466) );
  NAND2_X1 U16814 ( .A1(n20683), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13646) );
  NAND2_X1 U16815 ( .A1(n13466), .A2(n13646), .ZN(n13467) );
  AOI21_X1 U16816 ( .B1(n13655), .B2(n20650), .A(n13467), .ZN(n13468) );
  OAI21_X1 U16817 ( .B1(n20712), .B2(n15020), .A(n13468), .ZN(P1_U2999) );
  INV_X1 U16818 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n21491) );
  INV_X1 U16819 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17736) );
  NOR2_X1 U16820 ( .A1(n17736), .A2(n14323), .ZN(n13658) );
  NAND4_X1 U16821 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(P3_EBX_REG_16__SCAN_IN), 
        .A3(n9653), .A4(n13658), .ZN(n18056) );
  OAI21_X1 U16822 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n13469), .A(n18021), .ZN(
        n13487) );
  INV_X1 U16823 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13471) );
  INV_X1 U16824 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13470) );
  OAI22_X1 U16825 ( .A1(n18077), .A2(n13471), .B1(n9640), .B2(n13470), .ZN(
        n13476) );
  INV_X1 U16826 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13474) );
  AOI22_X1 U16827 ( .A1(n18061), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13473) );
  AOI22_X1 U16828 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18107), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13472) );
  OAI211_X1 U16829 ( .C1(n18112), .C2(n13474), .A(n13473), .B(n13472), .ZN(
        n13475) );
  AOI211_X1 U16830 ( .C1(n17293), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n13476), .B(n13475), .ZN(n13485) );
  INV_X1 U16831 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13477) );
  NOR2_X1 U16832 ( .A1(n13478), .A2(n13477), .ZN(n13481) );
  INV_X1 U16833 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17311) );
  INV_X1 U16834 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13479) );
  OAI22_X1 U16835 ( .A1(n17311), .A2(n10445), .B1(n13095), .B2(n13479), .ZN(
        n13480) );
  AOI211_X1 U16836 ( .C1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .C2(n18098), .A(
        n13481), .B(n13480), .ZN(n13484) );
  AOI22_X1 U16837 ( .A1(n17266), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13483) );
  AOI22_X1 U16838 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13482) );
  NAND4_X1 U16839 ( .A1(n13485), .A2(n13484), .A3(n13483), .A4(n13482), .ZN(
        n16839) );
  NAND2_X1 U16840 ( .A1(n18151), .A2(n16839), .ZN(n13486) );
  OAI21_X1 U16841 ( .B1(n13487), .B2(n18151), .A(n13486), .ZN(P3_U2684) );
  AND2_X1 U16842 ( .A1(n13165), .A2(n13488), .ZN(n13489) );
  NOR2_X1 U16843 ( .A1(n13286), .A2(n13489), .ZN(n16659) );
  INV_X1 U16844 ( .A(n16659), .ZN(n13494) );
  INV_X1 U16845 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19676) );
  OR2_X1 U16846 ( .A1(n16770), .A2(n13490), .ZN(n13492) );
  NAND2_X1 U16847 ( .A1(n16772), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13491) );
  NAND2_X1 U16848 ( .A1(n13492), .A2(n13491), .ZN(n16076) );
  INV_X1 U16849 ( .A(n16076), .ZN(n13493) );
  OAI222_X1 U16850 ( .A1(n13494), .A2(n16156), .B1(n16151), .B2(n19676), .C1(
        n19655), .C2(n13493), .ZN(P2_U2910) );
  NOR2_X1 U16851 ( .A1(n13495), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18674) );
  NOR2_X1 U16852 ( .A1(n18674), .A2(n18677), .ZN(n13753) );
  AOI21_X1 U16853 ( .B1(n18784), .B2(n18944), .A(n17216), .ZN(n13500) );
  INV_X1 U16854 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n13497) );
  NOR2_X1 U16855 ( .A1(n18840), .A2(n13497), .ZN(n13749) );
  INV_X1 U16856 ( .A(n13753), .ZN(n13498) );
  NOR2_X1 U16857 ( .A1(n18906), .A2(n13498), .ZN(n13499) );
  AOI211_X1 U16858 ( .C1(n13500), .C2(n18840), .A(n13749), .B(n13499), .ZN(
        n13502) );
  NAND2_X1 U16859 ( .A1(n18896), .A2(n18868), .ZN(n18816) );
  INV_X1 U16860 ( .A(n18816), .ZN(n18747) );
  NOR3_X1 U16861 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18747), .A3(
        n18899), .ZN(n18954) );
  INV_X1 U16862 ( .A(n18954), .ZN(n13501) );
  OAI211_X1 U16863 ( .C1(n13753), .C2(n18923), .A(n13502), .B(n13501), .ZN(
        P3_U2862) );
  INV_X1 U16864 ( .A(n18255), .ZN(n18236) );
  NAND2_X1 U16865 ( .A1(n18236), .A2(BUF2_REG_1__SCAN_IN), .ZN(n13505) );
  OAI211_X1 U16866 ( .C1(n13540), .C2(P3_EAX_REG_1__SCAN_IN), .A(n18251), .B(
        n13503), .ZN(n13504) );
  OAI211_X1 U16867 ( .C1(n13506), .C2(n18197), .A(n13505), .B(n13504), .ZN(
        P3_U2734) );
  AOI22_X1 U16868 ( .A1(n18061), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13514) );
  NAND2_X1 U16869 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n13510) );
  NAND2_X1 U16870 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n13509) );
  NAND2_X1 U16871 ( .A1(n13507), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n13508) );
  AND3_X1 U16872 ( .A1(n13510), .A2(n13509), .A3(n13508), .ZN(n13513) );
  AOI22_X1 U16873 ( .A1(n18008), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13512) );
  NAND2_X1 U16874 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n13511) );
  NAND4_X1 U16875 ( .A1(n13514), .A2(n13513), .A3(n13512), .A4(n13511), .ZN(
        n13520) );
  AOI22_X1 U16876 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13518) );
  AOI22_X1 U16877 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17312), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13517) );
  AOI22_X1 U16878 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13516) );
  AOI22_X1 U16879 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13515) );
  NAND4_X1 U16880 ( .A1(n13518), .A2(n13517), .A3(n13516), .A4(n13515), .ZN(
        n13519) );
  INV_X1 U16881 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18997) );
  AOI21_X1 U16882 ( .B1(n18251), .B2(P3_EAX_REG_4__SCAN_IN), .A(n13521), .ZN(
        n13523) );
  INV_X1 U16883 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18332) );
  NOR2_X1 U16884 ( .A1(n18332), .A2(n13522), .ZN(n13697) );
  OAI222_X1 U16885 ( .A1(n18197), .A2(n16964), .B1(n18255), .B2(n18997), .C1(
        n13523), .C2(n13697), .ZN(P3_U2731) );
  AOI22_X1 U16886 ( .A1(n13507), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18107), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13525) );
  NAND2_X1 U16887 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n13524) );
  AND2_X1 U16888 ( .A1(n13525), .A2(n13524), .ZN(n13529) );
  AOI22_X1 U16889 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13528) );
  AOI22_X1 U16890 ( .A1(n13207), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13527) );
  NAND2_X1 U16891 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13526) );
  NAND4_X1 U16892 ( .A1(n13529), .A2(n13528), .A3(n13527), .A4(n13526), .ZN(
        n13535) );
  AOI22_X1 U16893 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13533) );
  AOI22_X1 U16894 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13532) );
  AOI22_X1 U16895 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13531) );
  AOI22_X1 U16896 ( .A1(n17266), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13530) );
  NAND4_X1 U16897 ( .A1(n13533), .A2(n13532), .A3(n13531), .A4(n13530), .ZN(
        n13534) );
  OR2_X1 U16898 ( .A1(n13535), .A2(n13534), .ZN(n16860) );
  AOI21_X1 U16899 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n18094), .A(
        P3_EBX_REG_11__SCAN_IN), .ZN(n13536) );
  NOR3_X1 U16900 ( .A1(n13537), .A2(n13536), .A3(n18151), .ZN(n13538) );
  AOI21_X1 U16901 ( .B1(n18151), .B2(n16860), .A(n13538), .ZN(n13539) );
  INV_X1 U16902 ( .A(n13539), .ZN(P3_U2692) );
  INV_X1 U16903 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17485) );
  NAND3_X1 U16904 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .ZN(n13542) );
  NAND4_X1 U16905 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .A4(P3_EAX_REG_3__SCAN_IN), .ZN(n13541) );
  INV_X1 U16906 ( .A(n16833), .ZN(n18250) );
  NOR2_X1 U16907 ( .A1(n18250), .A2(n19010), .ZN(n18247) );
  AOI22_X1 U16908 ( .A1(n18247), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n18251), .ZN(n13545) );
  NAND3_X1 U16909 ( .A1(n18247), .A2(P3_EAX_REG_8__SCAN_IN), .A3(
        P3_EAX_REG_9__SCAN_IN), .ZN(n18242) );
  INV_X1 U16910 ( .A(n18242), .ZN(n13544) );
  OAI222_X1 U16911 ( .A1(n18255), .A2(n17485), .B1(n18197), .B2(n13546), .C1(
        n13545), .C2(n13544), .ZN(P3_U2726) );
  NAND2_X1 U16912 ( .A1(n20711), .A2(DATAI_3_), .ZN(n13548) );
  NAND2_X1 U16913 ( .A1(n20709), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13547) );
  INV_X1 U16914 ( .A(n20744), .ZN(n13549) );
  NAND2_X1 U16915 ( .A1(n13587), .A2(n13549), .ZN(n13568) );
  NAND2_X1 U16916 ( .A1(n20637), .A2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13551) );
  OAI211_X1 U16917 ( .C1(n20639), .C2(n15117), .A(n13568), .B(n13551), .ZN(
        P1_U2940) );
  NAND2_X1 U16918 ( .A1(n20711), .A2(DATAI_1_), .ZN(n13553) );
  NAND2_X1 U16919 ( .A1(n20709), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13552) );
  AND2_X1 U16920 ( .A1(n13553), .A2(n13552), .ZN(n20735) );
  INV_X1 U16921 ( .A(n20735), .ZN(n13554) );
  NAND2_X1 U16922 ( .A1(n13587), .A2(n13554), .ZN(n13560) );
  NAND2_X1 U16923 ( .A1(n20637), .A2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13555) );
  OAI211_X1 U16924 ( .C1(n20639), .C2(n15126), .A(n13560), .B(n13555), .ZN(
        P1_U2938) );
  INV_X1 U16925 ( .A(DATAI_2_), .ZN(n13557) );
  NAND2_X1 U16926 ( .A1(n20709), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13556) );
  OAI21_X1 U16927 ( .B1(n20709), .B2(n13557), .A(n13556), .ZN(n15122) );
  NAND2_X1 U16928 ( .A1(n13587), .A2(n15122), .ZN(n13575) );
  NAND2_X1 U16929 ( .A1(n20637), .A2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13558) );
  OAI211_X1 U16930 ( .C1(n20639), .C2(n13559), .A(n13575), .B(n13558), .ZN(
        P1_U2939) );
  AOI22_X1 U16931 ( .A1(n13601), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20637), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13561) );
  NAND2_X1 U16932 ( .A1(n13561), .A2(n13560), .ZN(P1_U2953) );
  AOI22_X1 U16933 ( .A1(n13601), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20637), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n13564) );
  INV_X1 U16934 ( .A(DATAI_11_), .ZN(n13562) );
  INV_X1 U16935 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13620) );
  MUX2_X1 U16936 ( .A(n13562), .B(n13620), .S(n20709), .Z(n15147) );
  INV_X1 U16937 ( .A(n15147), .ZN(n13563) );
  NAND2_X1 U16938 ( .A1(n13587), .A2(n13563), .ZN(n13602) );
  NAND2_X1 U16939 ( .A1(n13564), .A2(n13602), .ZN(P1_U2963) );
  AOI22_X1 U16940 ( .A1(n13601), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20637), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n13567) );
  INV_X1 U16941 ( .A(DATAI_14_), .ZN(n13565) );
  INV_X1 U16942 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n13790) );
  MUX2_X1 U16943 ( .A(n13565), .B(n13790), .S(n20709), .Z(n15141) );
  INV_X1 U16944 ( .A(n15141), .ZN(n13566) );
  NAND2_X1 U16945 ( .A1(n13587), .A2(n13566), .ZN(n13583) );
  NAND2_X1 U16946 ( .A1(n13567), .A2(n13583), .ZN(P1_U2966) );
  AOI22_X1 U16947 ( .A1(n13601), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20637), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13569) );
  NAND2_X1 U16948 ( .A1(n13569), .A2(n13568), .ZN(P1_U2955) );
  AOI22_X1 U16949 ( .A1(n13601), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20637), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13572) );
  INV_X1 U16950 ( .A(DATAI_12_), .ZN(n13570) );
  INV_X1 U16951 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n17458) );
  MUX2_X1 U16952 ( .A(n13570), .B(n17458), .S(n20709), .Z(n15146) );
  INV_X1 U16953 ( .A(n15146), .ZN(n13571) );
  NAND2_X1 U16954 ( .A1(n13587), .A2(n13571), .ZN(n13573) );
  NAND2_X1 U16955 ( .A1(n13572), .A2(n13573), .ZN(P1_U2949) );
  AOI22_X1 U16956 ( .A1(n13601), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20637), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n13574) );
  NAND2_X1 U16957 ( .A1(n13574), .A2(n13573), .ZN(P1_U2964) );
  AOI22_X1 U16958 ( .A1(n13601), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20637), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13576) );
  NAND2_X1 U16959 ( .A1(n13576), .A2(n13575), .ZN(P1_U2954) );
  AOI22_X1 U16960 ( .A1(n13601), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20637), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n13578) );
  NAND2_X1 U16961 ( .A1(n13578), .A2(n13577), .ZN(P1_U2960) );
  AOI22_X1 U16962 ( .A1(n13601), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20637), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13582) );
  INV_X1 U16963 ( .A(DATAI_0_), .ZN(n13580) );
  NAND2_X1 U16964 ( .A1(n20709), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13579) );
  OAI21_X1 U16965 ( .B1(n20709), .B2(n13580), .A(n13579), .ZN(n15132) );
  INV_X1 U16966 ( .A(n15132), .ZN(n20725) );
  NOR2_X1 U16967 ( .A1(n20633), .A2(n20725), .ZN(n20628) );
  INV_X1 U16968 ( .A(n20628), .ZN(n13581) );
  NAND2_X1 U16969 ( .A1(n13582), .A2(n13581), .ZN(P1_U2952) );
  AOI22_X1 U16970 ( .A1(n13601), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20637), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13584) );
  NAND2_X1 U16971 ( .A1(n13584), .A2(n13583), .ZN(P1_U2951) );
  AOI22_X1 U16972 ( .A1(n13601), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20637), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n13588) );
  INV_X1 U16973 ( .A(DATAI_10_), .ZN(n13585) );
  MUX2_X1 U16974 ( .A(n13585), .B(n17461), .S(n20709), .Z(n15149) );
  INV_X1 U16975 ( .A(n15149), .ZN(n13586) );
  NAND2_X1 U16976 ( .A1(n13587), .A2(n13586), .ZN(n13597) );
  NAND2_X1 U16977 ( .A1(n13588), .A2(n13597), .ZN(P1_U2962) );
  AOI22_X1 U16978 ( .A1(n13601), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20637), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13590) );
  NAND2_X1 U16979 ( .A1(n13590), .A2(n13589), .ZN(P1_U2959) );
  AOI22_X1 U16980 ( .A1(n13601), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20637), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13592) );
  NAND2_X1 U16981 ( .A1(n13592), .A2(n13591), .ZN(P1_U2958) );
  AOI22_X1 U16982 ( .A1(n13601), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20637), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13594) );
  NAND2_X1 U16983 ( .A1(n13594), .A2(n13593), .ZN(P1_U2957) );
  AOI22_X1 U16984 ( .A1(n13601), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20637), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n13596) );
  NAND2_X1 U16985 ( .A1(n13596), .A2(n13595), .ZN(P1_U2961) );
  AOI22_X1 U16986 ( .A1(n13601), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20637), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13598) );
  NAND2_X1 U16987 ( .A1(n13598), .A2(n13597), .ZN(P1_U2947) );
  AOI22_X1 U16988 ( .A1(n13601), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20637), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13600) );
  NAND2_X1 U16989 ( .A1(n13600), .A2(n13599), .ZN(P1_U2956) );
  AOI22_X1 U16990 ( .A1(n13601), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20637), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13603) );
  NAND2_X1 U16991 ( .A1(n13603), .A2(n13602), .ZN(P1_U2948) );
  OR2_X1 U16992 ( .A1(n13604), .A2(n15002), .ZN(n13605) );
  OR2_X1 U16993 ( .A1(n13611), .A2(n20763), .ZN(n13612) );
  INV_X1 U16994 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20627) );
  INV_X1 U16995 ( .A(n13612), .ZN(n13613) );
  OAI222_X1 U16996 ( .A1(n15020), .A2(n15158), .B1(n15157), .B2(n20627), .C1(
        n15156), .C2(n20725), .ZN(P1_U2904) );
  OAI21_X1 U16997 ( .B1(n13616), .B2(n13615), .A(n13614), .ZN(n15011) );
  OAI222_X1 U16998 ( .A1(n15011), .A2(n15158), .B1(n15157), .B2(n11580), .C1(
        n15156), .C2(n20735), .ZN(P1_U2903) );
  NAND2_X1 U16999 ( .A1(n13285), .A2(n13618), .ZN(n13619) );
  NAND2_X1 U17000 ( .A1(n13617), .A2(n13619), .ZN(n16634) );
  INV_X1 U17001 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19672) );
  OR2_X1 U17002 ( .A1(n16770), .A2(n13620), .ZN(n13622) );
  NAND2_X1 U17003 ( .A1(n16770), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13621) );
  NAND2_X1 U17004 ( .A1(n13622), .A2(n13621), .ZN(n16062) );
  INV_X1 U17005 ( .A(n16062), .ZN(n13623) );
  OAI222_X1 U17006 ( .A1(n16634), .A2(n16156), .B1(n16151), .B2(n19672), .C1(
        n19655), .C2(n13623), .ZN(P2_U2908) );
  XNOR2_X1 U17007 ( .A(n13624), .B(n13625), .ZN(n20692) );
  INV_X1 U17008 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13626) );
  OAI222_X1 U17009 ( .A1(n20692), .A2(n20594), .B1(n13626), .B2(n20599), .C1(
        n15011), .C2(n15055), .ZN(P1_U2871) );
  NAND2_X1 U17010 ( .A1(n19873), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19743) );
  INV_X1 U17011 ( .A(n19873), .ZN(n13633) );
  NAND2_X1 U17012 ( .A1(n13633), .A2(n20480), .ZN(n13627) );
  NAND2_X1 U17013 ( .A1(n19743), .A2(n13627), .ZN(n19917) );
  NOR2_X1 U17014 ( .A1(n19917), .A2(n20252), .ZN(n20180) );
  AOI21_X1 U17015 ( .B1(n13757), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n20180), .ZN(n13628) );
  OAI21_X2 U17016 ( .B1(n19727), .B2(n13632), .A(n13628), .ZN(n13764) );
  INV_X1 U17017 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13630) );
  INV_X1 U17018 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13631) );
  INV_X1 U17019 ( .A(n13632), .ZN(n13755) );
  NAND2_X1 U17020 ( .A1(n13757), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13635) );
  NAND2_X1 U17021 ( .A1(n20176), .A2(n20248), .ZN(n13634) );
  AND2_X1 U17022 ( .A1(n13634), .A2(n13633), .ZN(n19847) );
  NAND2_X1 U17023 ( .A1(n19847), .A2(n20463), .ZN(n20120) );
  NAND2_X1 U17024 ( .A1(n13635), .A2(n20120), .ZN(n13636) );
  INV_X1 U17025 ( .A(n16758), .ZN(n13638) );
  NAND2_X1 U17026 ( .A1(n13638), .A2(n13637), .ZN(n13639) );
  MUX2_X1 U17027 ( .A(n19727), .B(n13644), .S(n16043), .Z(n13645) );
  OAI21_X1 U17028 ( .B1(n20472), .B2(n16029), .A(n13645), .ZN(P2_U2885) );
  OAI21_X1 U17029 ( .B1(n20668), .B2(n15012), .A(n13646), .ZN(n13654) );
  NOR2_X1 U17030 ( .A1(n20676), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13647) );
  NOR2_X1 U17031 ( .A1(n20677), .A2(n13647), .ZN(n20697) );
  INV_X1 U17032 ( .A(n13648), .ZN(n13649) );
  NOR3_X1 U17033 ( .A1(n13650), .A2(n13649), .A3(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13651) );
  AOI21_X1 U17034 ( .B1(n20697), .B2(n13652), .A(n13651), .ZN(n13653) );
  AOI211_X1 U17035 ( .C1(n13655), .C2(n20699), .A(n13654), .B(n13653), .ZN(
        n13656) );
  INV_X1 U17036 ( .A(n13656), .ZN(P1_U3031) );
  NAND2_X1 U17037 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n14326), .ZN(n13729) );
  INV_X1 U17038 ( .A(n13729), .ZN(n13728) );
  AOI21_X1 U17039 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n18148), .A(n14326), .ZN(
        n13673) );
  NAND2_X1 U17040 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13660) );
  NAND2_X1 U17041 ( .A1(n13507), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n13659) );
  OAI211_X1 U17042 ( .C1(n17276), .C2(n13661), .A(n13660), .B(n13659), .ZN(
        n13662) );
  INV_X1 U17043 ( .A(n13662), .ZN(n13666) );
  AOI22_X1 U17044 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13665) );
  AOI22_X1 U17045 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13664) );
  NAND2_X1 U17046 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13663) );
  NAND4_X1 U17047 ( .A1(n13666), .A2(n13665), .A3(n13664), .A4(n13663), .ZN(
        n13672) );
  AOI22_X1 U17048 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13670) );
  AOI22_X1 U17049 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13669) );
  AOI22_X1 U17050 ( .A1(n13053), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13668) );
  AOI22_X1 U17051 ( .A1(n17266), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13667) );
  NAND4_X1 U17052 ( .A1(n13670), .A2(n13669), .A3(n13668), .A4(n13667), .ZN(
        n13671) );
  NOR2_X1 U17053 ( .A1(n13672), .A2(n13671), .ZN(n16848) );
  OAI22_X1 U17054 ( .A1(n13728), .A2(n13673), .B1(n16848), .B2(n18148), .ZN(
        P3_U2687) );
  INV_X1 U17055 ( .A(n14051), .ZN(n13676) );
  NAND2_X1 U17056 ( .A1(n20600), .A2(n11993), .ZN(n13958) );
  INV_X1 U17057 ( .A(n20612), .ZN(n21378) );
  NOR2_X4 U17058 ( .A1(n20600), .A2(n20624), .ZN(n20615) );
  AOI22_X1 U17059 ( .A1(n20624), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13678) );
  OAI21_X1 U17060 ( .B1(n15086), .B2(n13958), .A(n13678), .ZN(P1_U2910) );
  INV_X1 U17061 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13680) );
  AOI22_X1 U17062 ( .A1(n20624), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13679) );
  OAI21_X1 U17063 ( .B1(n13680), .B2(n13958), .A(n13679), .ZN(P1_U2912) );
  INV_X1 U17064 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n20635) );
  AOI22_X1 U17065 ( .A1(n20624), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13681) );
  OAI21_X1 U17066 ( .B1(n20635), .B2(n13958), .A(n13681), .ZN(P1_U2907) );
  AOI22_X1 U17067 ( .A1(n20624), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13682) );
  OAI21_X1 U17068 ( .B1(n15077), .B2(n13958), .A(n13682), .ZN(P1_U2908) );
  AOI22_X1 U17069 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13686) );
  NAND2_X1 U17070 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n13685) );
  NAND2_X1 U17071 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n13684) );
  NAND2_X1 U17072 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n13683) );
  NAND4_X1 U17073 ( .A1(n13686), .A2(n13685), .A3(n13684), .A4(n13683), .ZN(
        n13691) );
  INV_X1 U17074 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13689) );
  NAND2_X1 U17075 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n13688) );
  NAND2_X1 U17076 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n13687) );
  OAI211_X1 U17077 ( .C1(n14333), .C2(n13689), .A(n13688), .B(n13687), .ZN(
        n13690) );
  NOR2_X1 U17078 ( .A1(n13691), .A2(n13690), .ZN(n13696) );
  AOI22_X1 U17079 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13695) );
  AOI22_X1 U17080 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13694) );
  AOI22_X1 U17081 ( .A1(n13053), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13693) );
  AOI22_X1 U17082 ( .A1(n14312), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13692) );
  INV_X1 U17083 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n19002) );
  AOI21_X1 U17084 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n18251), .A(n13697), .ZN(
        n13698) );
  NAND2_X1 U17085 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n13697), .ZN(n16878) );
  INV_X1 U17086 ( .A(n16878), .ZN(n16894) );
  OAI222_X1 U17087 ( .A1(n18197), .A2(n16962), .B1(n18255), .B2(n19002), .C1(
        n13698), .C2(n16894), .ZN(P3_U2730) );
  INV_X1 U17088 ( .A(n13617), .ZN(n13699) );
  OAI21_X1 U17089 ( .B1(n13699), .B2(n9762), .A(n13885), .ZN(n16623) );
  OR2_X1 U17090 ( .A1(n16770), .A2(n17458), .ZN(n13701) );
  NAND2_X1 U17091 ( .A1(n16770), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13700) );
  NAND2_X1 U17092 ( .A1(n13701), .A2(n13700), .ZN(n16054) );
  AOI22_X1 U17093 ( .A1(n13793), .A2(n16054), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n19647), .ZN(n13702) );
  OAI21_X1 U17094 ( .B1(n16623), .B2(n16156), .A(n13702), .ZN(P2_U2907) );
  AOI22_X1 U17095 ( .A1(n13795), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n13877), .ZN(n13705) );
  NAND2_X1 U17096 ( .A1(n19698), .A2(n19797), .ZN(n13845) );
  NAND2_X1 U17097 ( .A1(n13705), .A2(n13845), .ZN(P2_U2958) );
  AOI22_X1 U17098 ( .A1(n13795), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(n13877), .ZN(n13709) );
  INV_X1 U17099 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n13706) );
  OR2_X1 U17100 ( .A1(n16772), .A2(n13706), .ZN(n13708) );
  NAND2_X1 U17101 ( .A1(n16772), .A2(BUF2_REG_5__SCAN_IN), .ZN(n13707) );
  NAND2_X1 U17102 ( .A1(n13708), .A2(n13707), .ZN(n19787) );
  NAND2_X1 U17103 ( .A1(n19698), .A2(n19787), .ZN(n13875) );
  NAND2_X1 U17104 ( .A1(n13709), .A2(n13875), .ZN(P2_U2957) );
  AOI22_X1 U17105 ( .A1(n13795), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n19700), .ZN(n13713) );
  INV_X1 U17106 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n13710) );
  OR2_X1 U17107 ( .A1(n16772), .A2(n13710), .ZN(n13712) );
  NAND2_X1 U17108 ( .A1(n16772), .A2(BUF2_REG_1__SCAN_IN), .ZN(n13711) );
  AND2_X1 U17109 ( .A1(n13712), .A2(n13711), .ZN(n19646) );
  INV_X1 U17110 ( .A(n19646), .ZN(n16784) );
  NAND2_X1 U17111 ( .A1(n19698), .A2(n16784), .ZN(n13882) );
  NAND2_X1 U17112 ( .A1(n13713), .A2(n13882), .ZN(P2_U2953) );
  AOI22_X1 U17113 ( .A1(n13795), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_23__SCAN_IN), .B2(n13877), .ZN(n13714) );
  NAND2_X1 U17114 ( .A1(n19698), .A2(n19810), .ZN(n13878) );
  NAND2_X1 U17115 ( .A1(n13714), .A2(n13878), .ZN(P2_U2959) );
  AOI22_X1 U17116 ( .A1(n13795), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n13877), .ZN(n13715) );
  NAND2_X1 U17117 ( .A1(n19698), .A2(n16076), .ZN(n13867) );
  NAND2_X1 U17118 ( .A1(n13715), .A2(n13867), .ZN(P2_U2961) );
  MUX2_X1 U17119 ( .A(n13720), .B(n14281), .S(n16043), .Z(n13721) );
  OAI21_X1 U17120 ( .B1(n19739), .B2(n16029), .A(n13721), .ZN(P2_U2886) );
  OR2_X1 U17121 ( .A1(n13722), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13724) );
  AND2_X1 U17122 ( .A1(n13724), .A2(n13723), .ZN(n20700) );
  MUX2_X1 U17123 ( .A(n20654), .B(n15344), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13725) );
  NAND2_X1 U17124 ( .A1(n20683), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20693) );
  NAND2_X1 U17125 ( .A1(n13725), .A2(n20693), .ZN(n13726) );
  AOI21_X1 U17126 ( .B1(n20700), .B2(n20650), .A(n13726), .ZN(n13727) );
  OAI21_X1 U17127 ( .B1(n15011), .B2(n20712), .A(n13727), .ZN(P1_U2998) );
  AOI21_X1 U17128 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n18148), .A(n13728), .ZN(
        n13743) );
  INV_X1 U17129 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17717) );
  NOR2_X1 U17130 ( .A1(n17717), .A2(n13729), .ZN(n18072) );
  INV_X1 U17131 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17298) );
  NAND2_X1 U17132 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13731) );
  NAND2_X1 U17133 ( .A1(n13507), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13730) );
  OAI211_X1 U17134 ( .C1(n17276), .C2(n17298), .A(n13731), .B(n13730), .ZN(
        n13732) );
  INV_X1 U17135 ( .A(n13732), .ZN(n13736) );
  AOI22_X1 U17136 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13735) );
  AOI22_X1 U17137 ( .A1(n13207), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13734) );
  NAND2_X1 U17138 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13733) );
  NAND4_X1 U17139 ( .A1(n13736), .A2(n13735), .A3(n13734), .A4(n13733), .ZN(
        n13742) );
  AOI22_X1 U17140 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13740) );
  AOI22_X1 U17141 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13739) );
  AOI22_X1 U17142 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13738) );
  AOI22_X1 U17143 ( .A1(n17266), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13737) );
  NAND4_X1 U17144 ( .A1(n13740), .A2(n13739), .A3(n13738), .A4(n13737), .ZN(
        n13741) );
  NOR2_X1 U17145 ( .A1(n13742), .A2(n13741), .ZN(n16847) );
  OAI22_X1 U17146 ( .A1(n13743), .A2(n18072), .B1(n16847), .B2(n18148), .ZN(
        P3_U2686) );
  NAND2_X1 U17147 ( .A1(n19404), .A2(n13744), .ZN(n13747) );
  INV_X1 U17148 ( .A(n19400), .ZN(n13745) );
  OR2_X4 U17149 ( .A1(n19421), .A2(n19430), .ZN(n17524) );
  NAND2_X1 U17150 ( .A1(n19558), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18439) );
  NAND2_X1 U17151 ( .A1(n19555), .A2(n19539), .ZN(n17519) );
  NAND2_X1 U17152 ( .A1(n19570), .A2(n17519), .ZN(n18965) );
  NAND2_X1 U17153 ( .A1(n18965), .A2(n19558), .ZN(n13748) );
  NAND3_X1 U17154 ( .A1(n19444), .A2(n18439), .A3(n18672), .ZN(n13750) );
  AOI21_X1 U17155 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13750), .A(
        n13749), .ZN(n13752) );
  NOR2_X4 U17156 ( .A1(n17524), .A2(n18298), .ZN(n18680) );
  NAND2_X1 U17157 ( .A1(n18680), .A2(n13753), .ZN(n13751) );
  OAI211_X1 U17158 ( .C1(n18612), .C2(n13753), .A(n13752), .B(n13751), .ZN(
        P3_U2830) );
  AND3_X1 U17159 ( .A1(n20471), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20009) );
  NAND2_X1 U17160 ( .A1(n20009), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20044) );
  NAND2_X1 U17161 ( .A1(n19743), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13756) );
  NAND2_X1 U17162 ( .A1(n20044), .A2(n13756), .ZN(n20178) );
  AOI22_X1 U17163 ( .A1(n13757), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20463), .B2(n20178), .ZN(n13758) );
  OR2_X1 U17164 ( .A1(n13760), .A2(n13759), .ZN(n13761) );
  INV_X1 U17165 ( .A(n13762), .ZN(n13763) );
  NAND2_X1 U17166 ( .A1(n13764), .A2(n13763), .ZN(n13765) );
  NAND2_X1 U17167 ( .A1(n13778), .A2(n13779), .ZN(n13769) );
  NAND2_X1 U17168 ( .A1(n10593), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13766) );
  AND2_X1 U17169 ( .A1(n13767), .A2(n13766), .ZN(n13768) );
  AND2_X1 U17170 ( .A1(n14571), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13770) );
  NAND2_X1 U17171 ( .A1(n13902), .A2(n13770), .ZN(n13910) );
  OR2_X1 U17172 ( .A1(n13902), .A2(n13770), .ZN(n13771) );
  NAND2_X1 U17173 ( .A1(n13910), .A2(n13771), .ZN(n19627) );
  AND2_X1 U17174 ( .A1(n11061), .A2(n13772), .ZN(n13775) );
  OAI21_X1 U17175 ( .B1(n13775), .B2(n13774), .A(n13773), .ZN(n16430) );
  MUX2_X1 U17176 ( .A(n13776), .B(n16430), .S(n15999), .Z(n13777) );
  OAI21_X1 U17177 ( .B1(n19627), .B2(n16029), .A(n13777), .ZN(P2_U2883) );
  INV_X1 U17178 ( .A(n20465), .ZN(n15911) );
  NOR2_X1 U17179 ( .A1(n13780), .A2(n16043), .ZN(n13781) );
  AOI21_X1 U17180 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n16043), .A(n13781), .ZN(
        n13782) );
  OAI21_X1 U17181 ( .B1(n15911), .B2(n16029), .A(n13782), .ZN(P2_U2884) );
  XOR2_X1 U17182 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13910), .Z(n13786)
         );
  NOR2_X1 U17183 ( .A1(n13773), .A2(n13783), .ZN(n13914) );
  AOI21_X1 U17184 ( .B1(n13783), .B2(n13773), .A(n13914), .ZN(n19622) );
  NOR2_X1 U17185 ( .A1(n15999), .A2(n11071), .ZN(n13784) );
  AOI21_X1 U17186 ( .B1(n19622), .B2(n15999), .A(n13784), .ZN(n13785) );
  OAI21_X1 U17187 ( .B1(n13786), .B2(n16029), .A(n13785), .ZN(P2_U2882) );
  OAI21_X1 U17188 ( .B1(n13887), .B2(n13789), .A(n13788), .ZN(n16585) );
  OR2_X1 U17189 ( .A1(n16772), .A2(n13790), .ZN(n13792) );
  NAND2_X1 U17190 ( .A1(n16772), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13791) );
  NAND2_X1 U17191 ( .A1(n13792), .A2(n13791), .ZN(n19697) );
  AOI22_X1 U17192 ( .A1(n13793), .A2(n19697), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19647), .ZN(n13794) );
  OAI21_X1 U17193 ( .B1(n16585), .B2(n16156), .A(n13794), .ZN(P2_U2905) );
  INV_X1 U17194 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14182) );
  NAND2_X1 U17195 ( .A1(n19701), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13796) );
  NAND2_X1 U17196 ( .A1(n19698), .A2(n16069), .ZN(n13798) );
  OAI211_X1 U17197 ( .C1(n14182), .C2(n13805), .A(n13796), .B(n13798), .ZN(
        P2_U2962) );
  INV_X1 U17198 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14172) );
  NAND2_X1 U17199 ( .A1(n19701), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13797) );
  NAND2_X1 U17200 ( .A1(n19698), .A2(n16083), .ZN(n13803) );
  OAI211_X1 U17201 ( .C1(n14172), .C2(n13805), .A(n13797), .B(n13803), .ZN(
        P2_U2960) );
  INV_X1 U17202 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19674) );
  NAND2_X1 U17203 ( .A1(n19701), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13799) );
  OAI211_X1 U17204 ( .C1(n19674), .C2(n13805), .A(n13799), .B(n13798), .ZN(
        P2_U2977) );
  INV_X1 U17205 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19670) );
  NAND2_X1 U17206 ( .A1(n19701), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13800) );
  NAND2_X1 U17207 ( .A1(n19698), .A2(n16054), .ZN(n13801) );
  OAI211_X1 U17208 ( .C1(n19670), .C2(n13805), .A(n13800), .B(n13801), .ZN(
        P2_U2979) );
  INV_X1 U17209 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14166) );
  NAND2_X1 U17210 ( .A1(n19701), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13802) );
  OAI211_X1 U17211 ( .C1(n14166), .C2(n13805), .A(n13802), .B(n13801), .ZN(
        P2_U2964) );
  INV_X1 U17212 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19678) );
  NAND2_X1 U17213 ( .A1(n19701), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13804) );
  OAI211_X1 U17214 ( .C1(n19678), .C2(n13805), .A(n13804), .B(n13803), .ZN(
        P2_U2975) );
  INV_X1 U17215 ( .A(n16765), .ZN(n17422) );
  INV_X1 U17216 ( .A(n14111), .ZN(n14095) );
  INV_X1 U17217 ( .A(n9589), .ZN(n13819) );
  NAND2_X1 U17218 ( .A1(n13808), .A2(n13807), .ZN(n14093) );
  INV_X1 U17219 ( .A(n14103), .ZN(n13811) );
  NAND2_X1 U17220 ( .A1(n13811), .A2(n13810), .ZN(n14087) );
  AOI22_X1 U17221 ( .A1(n14093), .A2(n14087), .B1(n11046), .B2(n14108), .ZN(
        n13817) );
  NOR2_X1 U17222 ( .A1(n13812), .A2(n9566), .ZN(n14090) );
  AOI21_X1 U17223 ( .B1(n14090), .B2(n14087), .A(n14604), .ZN(n13815) );
  INV_X1 U17224 ( .A(n11046), .ZN(n13813) );
  NAND2_X1 U17225 ( .A1(n14108), .A2(n13813), .ZN(n14089) );
  INV_X1 U17226 ( .A(n14089), .ZN(n13814) );
  NOR2_X1 U17227 ( .A1(n13815), .A2(n13814), .ZN(n13816) );
  MUX2_X1 U17228 ( .A(n13817), .B(n13816), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13818) );
  OAI211_X1 U17229 ( .C1(n13780), .C2(n14095), .A(n13819), .B(n13818), .ZN(
        n14098) );
  AOI22_X1 U17230 ( .A1(n20465), .A2(n17422), .B1(n20462), .B2(n14098), .ZN(
        n13831) );
  OR2_X1 U17231 ( .A1(n12498), .A2(n13820), .ZN(n13826) );
  INV_X1 U17232 ( .A(n13821), .ZN(n13822) );
  NOR2_X1 U17233 ( .A1(n13823), .A2(n13822), .ZN(n13824) );
  OAI211_X1 U17234 ( .C1(n14151), .C2(n13826), .A(n13825), .B(n13824), .ZN(
        n14130) );
  NAND2_X1 U17235 ( .A1(n14130), .A2(n14187), .ZN(n13828) );
  AOI22_X1 U17236 ( .A1(n17419), .A2(P2_FLUSH_REG_SCAN_IN), .B1(
        P2_STATE2_REG_3__SCAN_IN), .B2(n15584), .ZN(n13827) );
  INV_X1 U17237 ( .A(n17344), .ZN(n13830) );
  NAND2_X1 U17238 ( .A1(n13830), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13829) );
  OAI21_X1 U17239 ( .B1(n13831), .B2(n13830), .A(n13829), .ZN(P2_U3596) );
  NAND2_X1 U17240 ( .A1(n13833), .A2(n13614), .ZN(n13834) );
  AND2_X1 U17241 ( .A1(n13832), .A2(n13834), .ZN(n20586) );
  INV_X1 U17242 ( .A(n20586), .ZN(n13892) );
  INV_X1 U17243 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n21525) );
  INV_X1 U17244 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13835) );
  OAI22_X1 U17245 ( .A1(n15344), .A2(n21525), .B1(n20667), .B2(n13835), .ZN(
        n13836) );
  AOI21_X1 U17246 ( .B1(n15347), .B2(n20576), .A(n13836), .ZN(n13840) );
  OR2_X1 U17247 ( .A1(n13838), .A2(n13837), .ZN(n20681) );
  NAND3_X1 U17248 ( .A1(n20681), .A2(n20680), .A3(n20650), .ZN(n13839) );
  OAI211_X1 U17249 ( .C1(n13892), .C2(n20712), .A(n13840), .B(n13839), .ZN(
        P1_U2997) );
  AOI22_X1 U17250 ( .A1(n19701), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n13877), .ZN(n13844) );
  INV_X1 U17251 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n13841) );
  OR2_X1 U17252 ( .A1(n16772), .A2(n13841), .ZN(n13843) );
  NAND2_X1 U17253 ( .A1(n16772), .A2(BUF2_REG_0__SCAN_IN), .ZN(n13842) );
  AND2_X1 U17254 ( .A1(n13843), .A2(n13842), .ZN(n19656) );
  INV_X1 U17255 ( .A(n19656), .ZN(n16769) );
  NAND2_X1 U17256 ( .A1(n19698), .A2(n16769), .ZN(n13880) );
  NAND2_X1 U17257 ( .A1(n13844), .A2(n13880), .ZN(P2_U2967) );
  AOI22_X1 U17258 ( .A1(n19701), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_6__SCAN_IN), .B2(n13877), .ZN(n13846) );
  NAND2_X1 U17259 ( .A1(n13846), .A2(n13845), .ZN(P2_U2973) );
  AOI22_X1 U17260 ( .A1(n19701), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n13877), .ZN(n13847) );
  NAND2_X1 U17261 ( .A1(n19698), .A2(n16062), .ZN(n13859) );
  NAND2_X1 U17262 ( .A1(n13847), .A2(n13859), .ZN(P2_U2978) );
  AOI22_X1 U17263 ( .A1(n19701), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n13877), .ZN(n13850) );
  OR2_X1 U17264 ( .A1(n16770), .A2(n17468), .ZN(n13849) );
  NAND2_X1 U17265 ( .A1(n16772), .A2(BUF2_REG_4__SCAN_IN), .ZN(n13848) );
  AND2_X1 U17266 ( .A1(n13849), .A2(n13848), .ZN(n19632) );
  INV_X1 U17267 ( .A(n19632), .ZN(n19779) );
  NAND2_X1 U17268 ( .A1(n19698), .A2(n19779), .ZN(n13869) );
  NAND2_X1 U17269 ( .A1(n13850), .A2(n13869), .ZN(P2_U2956) );
  AOI22_X1 U17270 ( .A1(n19701), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n13877), .ZN(n13854) );
  INV_X1 U17271 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13851) );
  OR2_X1 U17272 ( .A1(n16770), .A2(n13851), .ZN(n13853) );
  NAND2_X1 U17273 ( .A1(n16770), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13852) );
  NAND2_X1 U17274 ( .A1(n13853), .A2(n13852), .ZN(n16047) );
  NAND2_X1 U17275 ( .A1(n19698), .A2(n16047), .ZN(n13873) );
  NAND2_X1 U17276 ( .A1(n13854), .A2(n13873), .ZN(P2_U2965) );
  AOI22_X1 U17277 ( .A1(n19701), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n19700), .ZN(n13858) );
  INV_X1 U17278 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n13855) );
  OR2_X1 U17279 ( .A1(n16772), .A2(n13855), .ZN(n13857) );
  NAND2_X1 U17280 ( .A1(n16772), .A2(BUF2_REG_2__SCAN_IN), .ZN(n13856) );
  NAND2_X1 U17281 ( .A1(n13857), .A2(n13856), .ZN(n19762) );
  NAND2_X1 U17282 ( .A1(n19698), .A2(n19762), .ZN(n13871) );
  NAND2_X1 U17283 ( .A1(n13858), .A2(n13871), .ZN(P2_U2969) );
  AOI22_X1 U17284 ( .A1(n19701), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n13877), .ZN(n13860) );
  NAND2_X1 U17285 ( .A1(n13860), .A2(n13859), .ZN(P2_U2963) );
  AOI22_X1 U17286 ( .A1(n19701), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n19700), .ZN(n13864) );
  INV_X1 U17287 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n13861) );
  OR2_X1 U17288 ( .A1(n16772), .A2(n13861), .ZN(n13863) );
  NAND2_X1 U17289 ( .A1(n16772), .A2(BUF2_REG_3__SCAN_IN), .ZN(n13862) );
  AND2_X1 U17290 ( .A1(n13863), .A2(n13862), .ZN(n19639) );
  INV_X1 U17291 ( .A(n19639), .ZN(n19770) );
  NAND2_X1 U17292 ( .A1(n19698), .A2(n19770), .ZN(n13865) );
  NAND2_X1 U17293 ( .A1(n13864), .A2(n13865), .ZN(P2_U2970) );
  AOI22_X1 U17294 ( .A1(n19701), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n19700), .ZN(n13866) );
  NAND2_X1 U17295 ( .A1(n13866), .A2(n13865), .ZN(P2_U2955) );
  AOI22_X1 U17296 ( .A1(n19701), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n13877), .ZN(n13868) );
  NAND2_X1 U17297 ( .A1(n13868), .A2(n13867), .ZN(P2_U2976) );
  AOI22_X1 U17298 ( .A1(n19701), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n19700), .ZN(n13870) );
  NAND2_X1 U17299 ( .A1(n13870), .A2(n13869), .ZN(P2_U2971) );
  AOI22_X1 U17300 ( .A1(n19701), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n19700), .ZN(n13872) );
  NAND2_X1 U17301 ( .A1(n13872), .A2(n13871), .ZN(P2_U2954) );
  AOI22_X1 U17302 ( .A1(n19701), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n13877), .ZN(n13874) );
  NAND2_X1 U17303 ( .A1(n13874), .A2(n13873), .ZN(P2_U2980) );
  AOI22_X1 U17304 ( .A1(n19701), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n19700), .ZN(n13876) );
  NAND2_X1 U17305 ( .A1(n13876), .A2(n13875), .ZN(P2_U2972) );
  AOI22_X1 U17306 ( .A1(n19701), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_7__SCAN_IN), .B2(n13877), .ZN(n13879) );
  NAND2_X1 U17307 ( .A1(n13879), .A2(n13878), .ZN(P2_U2974) );
  AOI22_X1 U17308 ( .A1(n19701), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n19700), .ZN(n13881) );
  NAND2_X1 U17309 ( .A1(n13881), .A2(n13880), .ZN(P2_U2952) );
  AOI22_X1 U17310 ( .A1(n19701), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_1__SCAN_IN), .B2(n19700), .ZN(n13883) );
  NAND2_X1 U17311 ( .A1(n13883), .A2(n13882), .ZN(P2_U2968) );
  INV_X1 U17312 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n21432) );
  INV_X1 U17313 ( .A(n15122), .ZN(n20739) );
  OAI222_X1 U17314 ( .A1(n13892), .A2(n15158), .B1(n15157), .B2(n21432), .C1(
        n15156), .C2(n20739), .ZN(P1_U2902) );
  AND2_X1 U17315 ( .A1(n13885), .A2(n13884), .ZN(n13886) );
  NOR2_X1 U17316 ( .A1(n13887), .A2(n13886), .ZN(n16598) );
  INV_X1 U17317 ( .A(n16598), .ZN(n13889) );
  INV_X1 U17318 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19668) );
  INV_X1 U17319 ( .A(n16047), .ZN(n13888) );
  OAI222_X1 U17320 ( .A1(n13889), .A2(n16156), .B1(n16151), .B2(n19668), .C1(
        n19655), .C2(n13888), .ZN(P2_U2906) );
  XNOR2_X1 U17321 ( .A(n13891), .B(n13890), .ZN(n20682) );
  INV_X1 U17322 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13893) );
  OAI222_X1 U17323 ( .A1(n20682), .A2(n20594), .B1(n20599), .B2(n13893), .C1(
        n13892), .C2(n15055), .ZN(P1_U2870) );
  AND2_X1 U17324 ( .A1(n14084), .A2(n13894), .ZN(n13896) );
  OR2_X1 U17325 ( .A1(n13896), .A2(n13895), .ZN(n16342) );
  NAND2_X1 U17326 ( .A1(n16652), .A2(n15999), .ZN(n13907) );
  NAND2_X1 U17327 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13909) );
  NAND2_X1 U17328 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13897) );
  NOR2_X1 U17329 ( .A1(n13909), .A2(n13897), .ZN(n13898) );
  NAND3_X1 U17330 ( .A1(n13899), .A2(n14080), .A3(n13898), .ZN(n13900) );
  NOR2_X1 U17331 ( .A1(n14549), .A2(n13900), .ZN(n13901) );
  INV_X1 U17332 ( .A(n13903), .ZN(n13904) );
  OAI211_X1 U17333 ( .C1(n13904), .C2(n13905), .A(n16037), .B(n13965), .ZN(
        n13906) );
  OAI211_X1 U17334 ( .C1(n15999), .C2(n11085), .A(n13907), .B(n13906), .ZN(
        P2_U2877) );
  NOR2_X1 U17335 ( .A1(n13910), .A2(n13908), .ZN(n13912) );
  NOR2_X1 U17336 ( .A1(n13910), .A2(n13909), .ZN(n14079) );
  INV_X1 U17337 ( .A(n14079), .ZN(n13911) );
  OAI211_X1 U17338 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13912), .A(
        n13911), .B(n16037), .ZN(n13920) );
  INV_X1 U17339 ( .A(n13914), .ZN(n13916) );
  NAND2_X1 U17340 ( .A1(n13916), .A2(n13915), .ZN(n13917) );
  NAND2_X1 U17341 ( .A1(n13913), .A2(n13917), .ZN(n16704) );
  MUX2_X1 U17342 ( .A(n16704), .B(n13918), .S(n16043), .Z(n13919) );
  NAND2_X1 U17343 ( .A1(n13920), .A2(n13919), .ZN(P2_U2881) );
  INV_X1 U17344 ( .A(n19762), .ZN(n13939) );
  OR2_X1 U17345 ( .A1(n13923), .A2(n13922), .ZN(n13924) );
  NAND2_X1 U17346 ( .A1(n14665), .A2(n13924), .ZN(n20477) );
  XNOR2_X1 U17347 ( .A(n20472), .B(n20477), .ZN(n13935) );
  OR2_X1 U17348 ( .A1(n13926), .A2(n13925), .ZN(n13927) );
  NAND2_X1 U17349 ( .A1(n13928), .A2(n13927), .ZN(n19640) );
  NOR2_X1 U17350 ( .A1(n20461), .A2(n19640), .ZN(n13932) );
  AOI21_X1 U17351 ( .B1(n20461), .B2(n19640), .A(n13932), .ZN(n19642) );
  INV_X1 U17352 ( .A(n13930), .ZN(n13931) );
  XNOR2_X1 U17353 ( .A(n13929), .B(n13931), .ZN(n19651) );
  NAND2_X1 U17354 ( .A1(n19652), .A2(n19651), .ZN(n19650) );
  NAND2_X1 U17355 ( .A1(n19642), .A2(n19650), .ZN(n19641) );
  INV_X1 U17356 ( .A(n13932), .ZN(n13933) );
  NAND2_X1 U17357 ( .A1(n19641), .A2(n13933), .ZN(n13934) );
  NAND2_X1 U17358 ( .A1(n13934), .A2(n13935), .ZN(n16147) );
  OAI21_X1 U17359 ( .B1(n13935), .B2(n13934), .A(n16147), .ZN(n13936) );
  NAND2_X1 U17360 ( .A1(n13936), .A2(n19649), .ZN(n13938) );
  AOI22_X1 U17361 ( .A1(n19648), .A2(n20477), .B1(n19647), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13937) );
  OAI211_X1 U17362 ( .C1(n13939), .C2(n19655), .A(n13938), .B(n13937), .ZN(
        P2_U2917) );
  XNOR2_X1 U17363 ( .A(n14079), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13945) );
  AND2_X1 U17364 ( .A1(n13913), .A2(n13941), .ZN(n13942) );
  NOR2_X1 U17365 ( .A1(n13940), .A2(n13942), .ZN(n16691) );
  NOR2_X1 U17366 ( .A1(n15999), .A2(n11076), .ZN(n13943) );
  AOI21_X1 U17367 ( .B1(n16691), .B2(n15999), .A(n13943), .ZN(n13944) );
  OAI21_X1 U17368 ( .B1(n13945), .B2(n16029), .A(n13944), .ZN(P2_U2880) );
  AOI22_X1 U17369 ( .A1(n20624), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13946) );
  OAI21_X1 U17370 ( .B1(n15091), .B2(n13958), .A(n13946), .ZN(P1_U2911) );
  AOI22_X1 U17371 ( .A1(n20624), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13947) );
  OAI21_X1 U17372 ( .B1(n15099), .B2(n13958), .A(n13947), .ZN(P1_U2913) );
  INV_X1 U17373 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13949) );
  AOI22_X1 U17374 ( .A1(n20624), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13948) );
  OAI21_X1 U17375 ( .B1(n13949), .B2(n13958), .A(n13948), .ZN(P1_U2916) );
  AOI22_X1 U17376 ( .A1(n20624), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13950) );
  OAI21_X1 U17377 ( .B1(n15082), .B2(n13958), .A(n13950), .ZN(P1_U2909) );
  AOI22_X1 U17378 ( .A1(n20624), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13951) );
  OAI21_X1 U17379 ( .B1(n15067), .B2(n13958), .A(n13951), .ZN(P1_U2906) );
  AOI22_X1 U17380 ( .A1(n20624), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13952) );
  OAI21_X1 U17381 ( .B1(n15108), .B2(n13958), .A(n13952), .ZN(P1_U2915) );
  INV_X1 U17382 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n20630) );
  AOI22_X1 U17383 ( .A1(n20624), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13953) );
  OAI21_X1 U17384 ( .B1(n20630), .B2(n13958), .A(n13953), .ZN(P1_U2920) );
  AOI22_X1 U17385 ( .A1(n20624), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13954) );
  OAI21_X1 U17386 ( .B1(n15104), .B2(n13958), .A(n13954), .ZN(P1_U2914) );
  AOI22_X1 U17387 ( .A1(n20612), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13955) );
  OAI21_X1 U17388 ( .B1(n15126), .B2(n13958), .A(n13955), .ZN(P1_U2919) );
  AOI22_X1 U17389 ( .A1(n20612), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13956) );
  OAI21_X1 U17390 ( .B1(n15117), .B2(n13958), .A(n13956), .ZN(P1_U2917) );
  AOI22_X1 U17391 ( .A1(n20612), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13957) );
  OAI21_X1 U17392 ( .B1(n13559), .B2(n13958), .A(n13957), .ZN(P1_U2918) );
  XNOR2_X1 U17393 ( .A(n13959), .B(n13960), .ZN(n14231) );
  INV_X1 U17394 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20621) );
  OAI222_X1 U17395 ( .A1(n14231), .A2(n15158), .B1(n15157), .B2(n20621), .C1(
        n15156), .C2(n20744), .ZN(P1_U2901) );
  INV_X1 U17396 ( .A(n13961), .ZN(n13963) );
  INV_X1 U17397 ( .A(n13895), .ZN(n13962) );
  NOR2_X1 U17398 ( .A1(n13962), .A2(n13963), .ZN(n14206) );
  AOI21_X1 U17399 ( .B1(n13963), .B2(n13962), .A(n14206), .ZN(n16641) );
  NAND2_X1 U17400 ( .A1(n16641), .A2(n15999), .ZN(n13969) );
  INV_X1 U17401 ( .A(n13965), .ZN(n13967) );
  OAI211_X1 U17402 ( .C1(n13967), .C2(n13966), .A(n16037), .B(n14393), .ZN(
        n13968) );
  OAI211_X1 U17403 ( .C1(n15999), .C2(n13970), .A(n13969), .B(n13968), .ZN(
        P2_U2876) );
  OR2_X1 U17404 ( .A1(n16770), .A2(n13971), .ZN(n13973) );
  NAND2_X1 U17405 ( .A1(n16772), .A2(BUF2_REG_15__SCAN_IN), .ZN(n13972) );
  NAND2_X1 U17406 ( .A1(n13973), .A2(n13972), .ZN(n14069) );
  AOI222_X1 U17407 ( .A1(n14069), .A2(n19698), .B1(P2_LWORD_REG_15__SCAN_IN), 
        .B2(n19701), .C1(P2_EAX_REG_15__SCAN_IN), .C2(n19700), .ZN(n13974) );
  INV_X1 U17408 ( .A(n13974), .ZN(P2_U2982) );
  NAND4_X1 U17409 ( .A1(n13300), .A2(n13975), .A3(n12207), .A4(n12243), .ZN(
        n13976) );
  OR2_X1 U17410 ( .A1(n13977), .A2(n13976), .ZN(n14011) );
  INV_X1 U17411 ( .A(n14011), .ZN(n13993) );
  OR2_X1 U17412 ( .A1(n21127), .A2(n13993), .ZN(n13988) );
  XNOR2_X1 U17413 ( .A(n13978), .B(n13979), .ZN(n13983) );
  NAND3_X1 U17414 ( .A1(n13993), .A2(n13980), .A3(n13983), .ZN(n13986) );
  XNOR2_X1 U17415 ( .A(n11465), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13984) );
  NAND2_X1 U17416 ( .A1(n13982), .A2(n13981), .ZN(n14017) );
  INV_X1 U17417 ( .A(n13983), .ZN(n15571) );
  AOI22_X1 U17418 ( .A1(n14649), .A2(n13984), .B1(n14017), .B2(n15571), .ZN(
        n13985) );
  AND2_X1 U17419 ( .A1(n13986), .A2(n13985), .ZN(n13987) );
  NAND2_X1 U17420 ( .A1(n13988), .A2(n13987), .ZN(n15566) );
  MUX2_X1 U17421 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15566), .S(
        n14037), .Z(n14030) );
  NAND2_X1 U17422 ( .A1(n11586), .A2(n14011), .ZN(n13990) );
  NAND2_X1 U17423 ( .A1(n13995), .A2(n10177), .ZN(n13989) );
  NAND2_X1 U17424 ( .A1(n13990), .A2(n13989), .ZN(n14652) );
  NAND2_X1 U17425 ( .A1(n14649), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13991) );
  NAND2_X1 U17426 ( .A1(n13991), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13992) );
  OR2_X1 U17427 ( .A1(n14652), .A2(n13992), .ZN(n13999) );
  INV_X1 U17428 ( .A(n13999), .ZN(n14001) );
  OR2_X1 U17429 ( .A1(n21188), .A2(n13993), .ZN(n13997) );
  NOR2_X1 U17430 ( .A1(n13994), .A2(n13978), .ZN(n15559) );
  AOI22_X1 U17431 ( .A1(n14649), .A2(n11465), .B1(n15559), .B2(n13995), .ZN(
        n13996) );
  NAND2_X1 U17432 ( .A1(n13997), .A2(n13996), .ZN(n15560) );
  OAI211_X1 U17433 ( .C1(n13999), .C2(n13998), .A(n14037), .B(n15560), .ZN(
        n14000) );
  OAI21_X1 U17434 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n14001), .A(
        n14000), .ZN(n14002) );
  AOI21_X1 U17435 ( .B1(n14030), .B2(n21123), .A(n14002), .ZN(n14003) );
  INV_X1 U17436 ( .A(n14003), .ZN(n14006) );
  INV_X1 U17437 ( .A(n14030), .ZN(n14004) );
  NAND2_X1 U17438 ( .A1(n14004), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14005) );
  NAND2_X1 U17439 ( .A1(n14006), .A2(n14005), .ZN(n14028) );
  INV_X1 U17440 ( .A(n14007), .ZN(n14008) );
  OAI21_X1 U17441 ( .B1(n13978), .B2(n14025), .A(n14008), .ZN(n14009) );
  NOR2_X1 U17442 ( .A1(n14009), .A2(n11808), .ZN(n15574) );
  NOR2_X1 U17443 ( .A1(n14010), .A2(n15574), .ZN(n14012) );
  MUX2_X1 U17444 ( .A(n14012), .B(n20720), .S(n14011), .Z(n14024) );
  INV_X1 U17445 ( .A(n14013), .ZN(n14032) );
  INV_X1 U17446 ( .A(n14014), .ZN(n14015) );
  MUX2_X1 U17447 ( .A(n14015), .B(n14025), .S(n13978), .Z(n14016) );
  NAND3_X1 U17448 ( .A1(n14017), .A2(n14032), .A3(n14016), .ZN(n14022) );
  NAND2_X1 U17449 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14018) );
  INV_X1 U17450 ( .A(n14018), .ZN(n14019) );
  MUX2_X1 U17451 ( .A(n14019), .B(n14018), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14020) );
  NAND2_X1 U17452 ( .A1(n14649), .A2(n14020), .ZN(n14021) );
  NAND2_X1 U17453 ( .A1(n14022), .A2(n14021), .ZN(n14023) );
  NOR2_X1 U17454 ( .A1(n14024), .A2(n14023), .ZN(n15576) );
  MUX2_X1 U17455 ( .A(n14025), .B(n15576), .S(n14037), .Z(n14034) );
  NAND2_X1 U17456 ( .A1(n14028), .A2(n14034), .ZN(n14026) );
  NAND2_X1 U17457 ( .A1(n14026), .A2(n21186), .ZN(n14027) );
  OAI21_X1 U17458 ( .B1(n14028), .B2(n14034), .A(n14027), .ZN(n14029) );
  NAND2_X1 U17459 ( .A1(n14029), .A2(n20708), .ZN(n14049) );
  NAND2_X1 U17460 ( .A1(n14030), .A2(n14650), .ZN(n14033) );
  NAND2_X1 U17461 ( .A1(n14031), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14040) );
  OAI22_X1 U17462 ( .A1(n14034), .A2(n14033), .B1(n14032), .B2(n14040), .ZN(
        n14218) );
  NAND2_X1 U17463 ( .A1(n14036), .A2(n14035), .ZN(n14038) );
  MUX2_X1 U17464 ( .A(n14039), .B(n14038), .S(n14037), .Z(n14041) );
  OAI22_X1 U17465 ( .A1(n14041), .A2(P1_STATE2_REG_1__SCAN_IN), .B1(n14040), 
        .B2(n14039), .ZN(n14216) );
  NOR2_X1 U17466 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n14045) );
  OAI211_X1 U17467 ( .C1(n14045), .C2(n14044), .A(n14043), .B(n14042), .ZN(
        n14046) );
  OR2_X1 U17468 ( .A1(n14216), .A2(n14046), .ZN(n14047) );
  NOR2_X1 U17469 ( .A1(n14218), .A2(n14047), .ZN(n14048) );
  NAND2_X1 U17470 ( .A1(n14049), .A2(n14048), .ZN(n14212) );
  OAI21_X1 U17471 ( .B1(n14212), .B2(n10072), .A(n14650), .ZN(n14059) );
  OR2_X1 U17472 ( .A1(n14051), .A2(n14050), .ZN(n14052) );
  NOR2_X1 U17473 ( .A1(n14053), .A2(n14052), .ZN(n14057) );
  INV_X1 U17474 ( .A(n15579), .ZN(n14055) );
  AOI21_X1 U17475 ( .B1(n21379), .B2(n14055), .A(n14054), .ZN(n14056) );
  AOI21_X1 U17476 ( .B1(n14058), .B2(n14057), .A(n14056), .ZN(n14063) );
  NAND2_X1 U17477 ( .A1(n14214), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14142) );
  NOR3_X1 U17478 ( .A1(n21379), .A2(n14060), .A3(n14650), .ZN(n14062) );
  NOR2_X1 U17479 ( .A1(n14062), .A2(n14061), .ZN(n15581) );
  AOI21_X1 U17480 ( .B1(n15581), .B2(n14220), .A(n14063), .ZN(n14065) );
  INV_X1 U17481 ( .A(n21384), .ZN(n14215) );
  AOI21_X1 U17482 ( .B1(n21000), .B2(n21308), .A(n14215), .ZN(n14064) );
  AOI211_X1 U17483 ( .C1(n14142), .C2(n14650), .A(n14065), .B(n14064), .ZN(
        P1_U3162) );
  INV_X1 U17484 ( .A(n14066), .ZN(n14067) );
  AOI21_X1 U17485 ( .B1(n14068), .B2(n13788), .A(n14067), .ZN(n16573) );
  INV_X1 U17486 ( .A(n16573), .ZN(n14071) );
  INV_X1 U17487 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19664) );
  INV_X1 U17488 ( .A(n14069), .ZN(n14070) );
  OAI222_X1 U17489 ( .A1(n14071), .A2(n16156), .B1(n16151), .B2(n19664), .C1(
        n14070), .C2(n19655), .ZN(P2_U2904) );
  INV_X1 U17490 ( .A(n14231), .ZN(n20571) );
  NOR2_X1 U17491 ( .A1(n14073), .A2(n14074), .ZN(n14075) );
  OR2_X1 U17492 ( .A1(n14072), .A2(n14075), .ZN(n20669) );
  OAI22_X1 U17493 ( .A1(n20594), .A2(n20669), .B1(n14076), .B2(n20599), .ZN(
        n14077) );
  AOI21_X1 U17494 ( .B1(n20571), .B2(n20596), .A(n14077), .ZN(n14078) );
  INV_X1 U17495 ( .A(n14078), .ZN(P1_U2869) );
  NAND2_X1 U17496 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14237) );
  NOR2_X1 U17497 ( .A1(n14237), .A2(n14238), .ZN(n14236) );
  OAI211_X1 U17498 ( .C1(n14236), .C2(n14080), .A(n16037), .B(n13903), .ZN(
        n14086) );
  NAND2_X1 U17499 ( .A1(n14081), .A2(n14082), .ZN(n14083) );
  NAND2_X1 U17500 ( .A1(n14084), .A2(n14083), .ZN(n16658) );
  INV_X1 U17501 ( .A(n16658), .ZN(n16358) );
  NAND2_X1 U17502 ( .A1(n16358), .A2(n15999), .ZN(n14085) );
  OAI211_X1 U17503 ( .C1(n15999), .C2(n10247), .A(n14086), .B(n14085), .ZN(
        P2_U2878) );
  NAND2_X1 U17504 ( .A1(n20471), .A2(n20480), .ZN(n19848) );
  NAND2_X1 U17505 ( .A1(n9582), .A2(n14087), .ZN(n14092) );
  AOI21_X1 U17506 ( .B1(n14093), .B2(n14092), .A(n14091), .ZN(n14094) );
  OAI21_X1 U17507 ( .B1(n19727), .B2(n14095), .A(n14094), .ZN(n16762) );
  INV_X1 U17508 ( .A(n14130), .ZN(n14097) );
  OAI22_X1 U17509 ( .A1(n14130), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16762), .B2(n14097), .ZN(n14128) );
  NAND2_X1 U17510 ( .A1(n14097), .A2(n10551), .ZN(n14096) );
  OAI21_X1 U17511 ( .B1(n14098), .B2(n14097), .A(n14096), .ZN(n14129) );
  OAI22_X1 U17512 ( .A1(n19848), .A2(n14128), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n14129), .ZN(n14099) );
  INV_X1 U17513 ( .A(n14099), .ZN(n14118) );
  INV_X1 U17514 ( .A(n19848), .ZN(n19876) );
  OAI22_X1 U17515 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n14129), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n14128), .ZN(n14116) );
  INV_X1 U17516 ( .A(n14108), .ZN(n14100) );
  NOR2_X1 U17517 ( .A1(n14100), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14106) );
  INV_X1 U17518 ( .A(n12584), .ZN(n14101) );
  AND2_X1 U17519 ( .A1(n14102), .A2(n14101), .ZN(n14107) );
  NOR3_X1 U17520 ( .A1(n14107), .A2(n14104), .A3(n14103), .ZN(n14105) );
  AOI211_X1 U17521 ( .C1(n16732), .C2(n14111), .A(n14106), .B(n14105), .ZN(
        n14303) );
  INV_X1 U17522 ( .A(n14303), .ZN(n14113) );
  INV_X1 U17523 ( .A(n15938), .ZN(n17406) );
  INV_X1 U17524 ( .A(n14107), .ZN(n14109) );
  MUX2_X1 U17525 ( .A(n14109), .B(n14108), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n14110) );
  AOI21_X1 U17526 ( .B1(n17406), .B2(n14111), .A(n14110), .ZN(n16755) );
  INV_X1 U17527 ( .A(n16755), .ZN(n14112) );
  OAI22_X1 U17528 ( .A1(n14113), .A2(n20176), .B1(n20248), .B2(n14112), .ZN(
        n14114) );
  OAI21_X1 U17529 ( .B1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n14303), .A(
        n14114), .ZN(n14115) );
  OAI211_X1 U17530 ( .C1(n19876), .C2(n14116), .A(n14130), .B(n14115), .ZN(
        n14117) );
  AOI21_X1 U17531 ( .B1(n14118), .B2(n14117), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n14134) );
  INV_X1 U17532 ( .A(n14119), .ZN(n14123) );
  NOR3_X1 U17533 ( .A1(n14122), .A2(n14121), .A3(n10574), .ZN(n17341) );
  NOR3_X1 U17534 ( .A1(n14124), .A2(n14123), .A3(n17341), .ZN(n14127) );
  OAI21_X1 U17535 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n14125), .ZN(n14126) );
  OAI211_X1 U17536 ( .C1(n14129), .C2(n14128), .A(n14127), .B(n14126), .ZN(
        n14132) );
  NOR2_X1 U17537 ( .A1(n14130), .A2(n17343), .ZN(n14131) );
  OR2_X1 U17538 ( .A1(n14132), .A2(n14131), .ZN(n14133) );
  OAI21_X1 U17539 ( .B1(n17414), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n14139) );
  NOR2_X1 U17540 ( .A1(n15978), .A2(n14135), .ZN(n14137) );
  OR2_X1 U17541 ( .A1(n14136), .A2(n20302), .ZN(n15588) );
  AOI21_X1 U17542 ( .B1(n12680), .B2(n14137), .A(n15588), .ZN(n14138) );
  OAI21_X1 U17543 ( .B1(n17425), .B2(n15584), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n14141) );
  NAND2_X1 U17544 ( .A1(n14141), .A2(n14140), .ZN(P2_U3593) );
  INV_X1 U17545 ( .A(n14142), .ZN(n14143) );
  OAI21_X1 U17546 ( .B1(n14143), .B2(n21000), .A(n15540), .ZN(P1_U3466) );
  NAND2_X1 U17547 ( .A1(n14146), .A2(n14145), .ZN(n14147) );
  AND2_X1 U17548 ( .A1(n14144), .A2(n14147), .ZN(n20648) );
  INV_X1 U17549 ( .A(n20648), .ZN(n14148) );
  INV_X1 U17550 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20619) );
  INV_X1 U17551 ( .A(n15113), .ZN(n20749) );
  OAI222_X1 U17552 ( .A1(n15158), .A2(n14148), .B1(n15157), .B2(n20619), .C1(
        n15156), .C2(n20749), .ZN(P1_U2900) );
  INV_X1 U17553 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n14158) );
  INV_X1 U17554 ( .A(n14149), .ZN(n14150) );
  INV_X1 U17555 ( .A(n19696), .ZN(n14154) );
  OR2_X1 U17556 ( .A1(n14155), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14156) );
  INV_X2 U17557 ( .A(n14156), .ZN(n19694) );
  AOI22_X1 U17558 ( .A1(n19694), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n14157) );
  OAI21_X1 U17559 ( .B1(n14158), .B2(n19658), .A(n14157), .ZN(P2_U2933) );
  INV_X1 U17560 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n14160) );
  AOI22_X1 U17561 ( .A1(n19694), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n14159) );
  OAI21_X1 U17562 ( .B1(n14160), .B2(n19658), .A(n14159), .ZN(P2_U2935) );
  INV_X1 U17563 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n14162) );
  AOI22_X1 U17564 ( .A1(n19694), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14161) );
  OAI21_X1 U17565 ( .B1(n14162), .B2(n19658), .A(n14161), .ZN(P2_U2931) );
  INV_X1 U17566 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14164) );
  AOI22_X1 U17567 ( .A1(n19694), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14163) );
  OAI21_X1 U17568 ( .B1(n14164), .B2(n19658), .A(n14163), .ZN(P2_U2928) );
  AOI22_X1 U17569 ( .A1(n19694), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14165) );
  OAI21_X1 U17570 ( .B1(n14166), .B2(n19658), .A(n14165), .ZN(P2_U2923) );
  AOI22_X1 U17571 ( .A1(n19694), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14167) );
  OAI21_X1 U17572 ( .B1(n14168), .B2(n19658), .A(n14167), .ZN(P2_U2922) );
  INV_X1 U17573 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14170) );
  AOI22_X1 U17574 ( .A1(n19694), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n14169) );
  OAI21_X1 U17575 ( .B1(n14170), .B2(n19658), .A(n14169), .ZN(P2_U2934) );
  AOI22_X1 U17576 ( .A1(n19694), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14171) );
  OAI21_X1 U17577 ( .B1(n14172), .B2(n19658), .A(n14171), .ZN(P2_U2927) );
  INV_X1 U17578 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14174) );
  AOI22_X1 U17579 ( .A1(n19694), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14173) );
  OAI21_X1 U17580 ( .B1(n14174), .B2(n19658), .A(n14173), .ZN(P2_U2932) );
  INV_X1 U17581 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14176) );
  AOI22_X1 U17582 ( .A1(n19694), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14175) );
  OAI21_X1 U17583 ( .B1(n14176), .B2(n19658), .A(n14175), .ZN(P2_U2924) );
  INV_X1 U17584 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14178) );
  AOI22_X1 U17585 ( .A1(n19694), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14177) );
  OAI21_X1 U17586 ( .B1(n14178), .B2(n19658), .A(n14177), .ZN(P2_U2930) );
  INV_X1 U17587 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14180) );
  AOI22_X1 U17588 ( .A1(n19694), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n14179) );
  OAI21_X1 U17589 ( .B1(n14180), .B2(n19658), .A(n14179), .ZN(P2_U2929) );
  AOI22_X1 U17590 ( .A1(n19694), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14181) );
  OAI21_X1 U17591 ( .B1(n14182), .B2(n19658), .A(n14181), .ZN(P2_U2925) );
  INV_X1 U17592 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14184) );
  AOI22_X1 U17593 ( .A1(n19694), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14183) );
  OAI21_X1 U17594 ( .B1(n14184), .B2(n19658), .A(n14183), .ZN(P2_U2926) );
  AOI21_X1 U17595 ( .B1(n17425), .B2(n20381), .A(n17418), .ZN(n14189) );
  INV_X1 U17596 ( .A(n15791), .ZN(n19616) );
  INV_X1 U17597 ( .A(n20462), .ZN(n16756) );
  NOR3_X1 U17598 ( .A1(n20381), .A2(n16756), .A3(n15584), .ZN(n14186) );
  INV_X1 U17599 ( .A(n17425), .ZN(n14185) );
  OAI21_X1 U17600 ( .B1(n14187), .B2(n14186), .A(n14185), .ZN(n14188) );
  OAI211_X1 U17601 ( .C1(n14189), .C2(n16757), .A(n19616), .B(n14188), .ZN(
        P2_U3177) );
  OAI21_X1 U17602 ( .B1(n14192), .B2(n14191), .A(n14190), .ZN(n17372) );
  NAND2_X1 U17603 ( .A1(n14194), .A2(n14195), .ZN(n14196) );
  NAND2_X1 U17604 ( .A1(n14193), .A2(n14196), .ZN(n20542) );
  INV_X1 U17605 ( .A(n20542), .ZN(n14203) );
  AND2_X1 U17606 ( .A1(n20683), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n17371) );
  INV_X1 U17607 ( .A(n20677), .ZN(n15516) );
  INV_X1 U17608 ( .A(n15467), .ZN(n14197) );
  OR2_X1 U17609 ( .A1(n20676), .A2(n14197), .ZN(n14198) );
  NAND2_X1 U17610 ( .A1(n15516), .A2(n14198), .ZN(n15492) );
  AOI21_X1 U17611 ( .B1(n20679), .B2(n14199), .A(n15492), .ZN(n17377) );
  NAND2_X1 U17612 ( .A1(n20675), .A2(n14200), .ZN(n17379) );
  NAND2_X1 U17613 ( .A1(n17379), .A2(n20676), .ZN(n15468) );
  NAND2_X1 U17614 ( .A1(n15514), .A2(n15468), .ZN(n20674) );
  NAND2_X1 U17615 ( .A1(n20658), .A2(n14201), .ZN(n17378) );
  OAI22_X1 U17616 ( .A1(n17377), .A2(n14201), .B1(n20674), .B2(n17378), .ZN(
        n14202) );
  AOI211_X1 U17617 ( .C1(n20696), .C2(n14203), .A(n17371), .B(n14202), .ZN(
        n14204) );
  OAI21_X1 U17618 ( .B1(n20666), .B2(n17372), .A(n14204), .ZN(P1_U3026) );
  OAI21_X1 U17619 ( .B1(n14206), .B2(n14205), .A(n15812), .ZN(n16617) );
  INV_X1 U17620 ( .A(n14393), .ZN(n14209) );
  NOR2_X1 U17621 ( .A1(n14393), .A2(n14207), .ZN(n16040) );
  INV_X1 U17622 ( .A(n16040), .ZN(n14208) );
  OAI211_X1 U17623 ( .C1(n14209), .C2(n14391), .A(n14208), .B(n16037), .ZN(
        n14211) );
  NAND2_X1 U17624 ( .A1(n16043), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14210) );
  OAI211_X1 U17625 ( .C1(n16617), .C2(n16043), .A(n14211), .B(n14210), .ZN(
        P2_U2875) );
  INV_X1 U17626 ( .A(n14212), .ZN(n14228) );
  OAI21_X1 U17627 ( .B1(n14215), .B2(n15573), .A(n14214), .ZN(n14225) );
  INV_X1 U17628 ( .A(n13994), .ZN(n14217) );
  AOI21_X1 U17629 ( .B1(n14218), .B2(n14217), .A(n14216), .ZN(n14219) );
  INV_X1 U17630 ( .A(n14219), .ZN(n15536) );
  NOR2_X1 U17631 ( .A1(n15536), .A2(n14220), .ZN(n15533) );
  NOR2_X1 U17632 ( .A1(n21308), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14221) );
  NOR4_X1 U17633 ( .A1(n15533), .A2(n14223), .A3(n14222), .A4(n14221), .ZN(
        n14224) );
  MUX2_X1 U17634 ( .A(n14225), .B(n14224), .S(P1_STATE2_REG_0__SCAN_IN), .Z(
        n14226) );
  OAI21_X1 U17635 ( .B1(n14228), .B2(n14227), .A(n14226), .ZN(P1_U3161) );
  XNOR2_X1 U17636 ( .A(n20642), .B(n20673), .ZN(n14229) );
  NAND2_X1 U17637 ( .A1(n14229), .A2(n12143), .ZN(n20644) );
  OAI21_X1 U17638 ( .B1(n14229), .B2(n12143), .A(n20644), .ZN(n20665) );
  INV_X1 U17639 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n14230) );
  OAI22_X1 U17640 ( .A1(n15344), .A2(n20566), .B1(n20667), .B2(n14230), .ZN(
        n14233) );
  NOR2_X1 U17641 ( .A1(n14231), .A2(n20712), .ZN(n14232) );
  AOI211_X1 U17642 ( .C1(n15347), .C2(n20561), .A(n14233), .B(n14232), .ZN(
        n14234) );
  OAI21_X1 U17643 ( .B1(n15339), .B2(n20665), .A(n14234), .ZN(P1_U2996) );
  OAI21_X1 U17644 ( .B1(n13940), .B2(n14235), .A(n14081), .ZN(n16369) );
  NOR2_X1 U17645 ( .A1(n16369), .A2(n16043), .ZN(n14240) );
  AOI211_X1 U17646 ( .C1(n14238), .C2(n14237), .A(n16029), .B(n14236), .ZN(
        n14239) );
  AOI211_X1 U17647 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n16043), .A(n14240), .B(
        n14239), .ZN(n14241) );
  INV_X1 U17648 ( .A(n14241), .ZN(P2_U2879) );
  OAI21_X1 U17649 ( .B1(n14242), .B2(n14244), .A(n14243), .ZN(n17362) );
  INV_X1 U17650 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14249) );
  NOR2_X1 U17651 ( .A1(n14246), .A2(n14247), .ZN(n14248) );
  OR2_X1 U17652 ( .A1(n14245), .A2(n14248), .ZN(n20526) );
  OAI222_X1 U17653 ( .A1(n17362), .A2(n15055), .B1(n14249), .B2(n20599), .C1(
        n20594), .C2(n20526), .ZN(P1_U2865) );
  OAI222_X1 U17654 ( .A1(n15158), .A2(n17362), .B1(n15157), .B2(n11619), .C1(
        n15156), .C2(n20767), .ZN(P1_U2897) );
  NAND2_X1 U17655 ( .A1(n9609), .A2(n14250), .ZN(n14251) );
  XOR2_X1 U17656 ( .A(n14251), .B(n16372), .Z(n14264) );
  INV_X1 U17657 ( .A(n15937), .ZN(n19621) );
  INV_X1 U17658 ( .A(n16369), .ZN(n16679) );
  NAND2_X1 U17659 ( .A1(n16675), .A2(n15933), .ZN(n14260) );
  NAND2_X1 U17660 ( .A1(n14253), .A2(n14252), .ZN(n14254) );
  INV_X1 U17661 ( .A(n15934), .ZN(n19607) );
  INV_X2 U17662 ( .A(n15816), .ZN(n19605) );
  AOI21_X1 U17663 ( .B1(n19605), .B2(P2_REIP_REG_8__SCAN_IN), .A(n19604), .ZN(
        n14256) );
  OAI21_X1 U17664 ( .B1(n19607), .B2(n14257), .A(n14256), .ZN(n14258) );
  AOI21_X1 U17665 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n15930), .A(
        n14258), .ZN(n14259) );
  OAI211_X1 U17666 ( .C1(n15875), .C2(n14261), .A(n14260), .B(n14259), .ZN(
        n14262) );
  AOI21_X1 U17667 ( .B1(n19621), .B2(n16679), .A(n14262), .ZN(n14263) );
  OAI21_X1 U17668 ( .B1(n14264), .B2(n19616), .A(n14263), .ZN(P2_U2847) );
  NAND2_X1 U17669 ( .A1(n9609), .A2(n14265), .ZN(n14288) );
  XNOR2_X1 U17670 ( .A(n14288), .B(n16314), .ZN(n14272) );
  INV_X1 U17671 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20411) );
  NAND2_X1 U17672 ( .A1(n15934), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14266) );
  OAI211_X1 U17673 ( .C1(n20411), .C2(n15816), .A(n14266), .B(n16416), .ZN(
        n14269) );
  NOR2_X1 U17674 ( .A1(n14267), .A2(n15875), .ZN(n14268) );
  AOI211_X1 U17675 ( .C1(n15930), .C2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n14269), .B(n14268), .ZN(n14270) );
  OAI21_X1 U17676 ( .B1(n16623), .B2(n19611), .A(n14270), .ZN(n14271) );
  AOI21_X1 U17677 ( .B1(n14272), .B2(n15791), .A(n14271), .ZN(n14273) );
  OAI21_X1 U17678 ( .B1(n15937), .B2(n16617), .A(n14273), .ZN(P2_U2843) );
  AND2_X1 U17679 ( .A1(n14274), .A2(n14299), .ZN(n14275) );
  NOR2_X1 U17680 ( .A1(n15915), .A2(n14275), .ZN(n14276) );
  NAND2_X1 U17681 ( .A1(n9609), .A2(n14276), .ZN(n14301) );
  MUX2_X1 U17682 ( .A(n15912), .B(n19625), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n14285) );
  AOI22_X1 U17683 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19605), .B1(n19609), 
        .B2(n14278), .ZN(n14280) );
  NAND2_X1 U17684 ( .A1(n15933), .A2(n19640), .ZN(n14279) );
  OAI211_X1 U17685 ( .C1(n19607), .C2(n14281), .A(n14280), .B(n14279), .ZN(
        n14283) );
  NOR2_X1 U17686 ( .A1(n19739), .A2(n15927), .ZN(n14282) );
  AOI211_X1 U17687 ( .C1(n19621), .C2(n16732), .A(n14283), .B(n14282), .ZN(
        n14284) );
  OAI211_X1 U17688 ( .C1(n14301), .C2(n19616), .A(n14285), .B(n14284), .ZN(
        P2_U2854) );
  INV_X1 U17689 ( .A(n16641), .ZN(n14298) );
  OAI21_X1 U17690 ( .B1(n14286), .B2(n16327), .A(n15791), .ZN(n14287) );
  OAI22_X1 U17691 ( .A1(n15912), .A2(n16327), .B1(n14288), .B2(n14287), .ZN(
        n14296) );
  NOR2_X1 U17692 ( .A1(n16634), .A2(n19611), .ZN(n14295) );
  NOR2_X1 U17693 ( .A1(n14289), .A2(n15875), .ZN(n14294) );
  AOI21_X1 U17694 ( .B1(n19605), .B2(P2_REIP_REG_11__SCAN_IN), .A(n19604), 
        .ZN(n14291) );
  NAND2_X1 U17695 ( .A1(n15934), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n14290) );
  OAI211_X1 U17696 ( .C1(n19625), .C2(n14292), .A(n14291), .B(n14290), .ZN(
        n14293) );
  NOR4_X1 U17697 ( .A1(n14296), .A2(n14295), .A3(n14294), .A4(n14293), .ZN(
        n14297) );
  OAI21_X1 U17698 ( .B1(n15937), .B2(n14298), .A(n14297), .ZN(P2_U2844) );
  INV_X1 U17699 ( .A(n14299), .ZN(n15943) );
  MUX2_X1 U17700 ( .A(n14300), .B(n15943), .S(n9609), .Z(n16754) );
  OAI21_X1 U17701 ( .B1(n9609), .B2(n14302), .A(n14301), .ZN(n16760) );
  NOR3_X1 U17702 ( .A1(n16754), .A2(n16760), .A3(n16757), .ZN(n14305) );
  OAI22_X1 U17703 ( .A1(n19739), .A2(n16765), .B1(n14303), .B2(n16756), .ZN(
        n14304) );
  OAI21_X1 U17704 ( .B1(n14305), .B2(n14304), .A(n17344), .ZN(n14306) );
  OAI21_X1 U17705 ( .B1(n17344), .B2(n14307), .A(n14306), .ZN(P2_U3600) );
  INV_X1 U17706 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14310) );
  NAND2_X1 U17707 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n14309) );
  NAND2_X1 U17708 ( .A1(n13507), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n14308) );
  OAI211_X1 U17709 ( .C1(n17276), .C2(n14310), .A(n14309), .B(n14308), .ZN(
        n14311) );
  INV_X1 U17710 ( .A(n14311), .ZN(n14316) );
  AOI22_X1 U17711 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14315) );
  AOI22_X1 U17712 ( .A1(n13207), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14314) );
  NAND2_X1 U17713 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14313) );
  NAND4_X1 U17714 ( .A1(n14316), .A2(n14315), .A3(n14314), .A4(n14313), .ZN(
        n14322) );
  AOI22_X1 U17715 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14320) );
  AOI22_X1 U17716 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14319) );
  AOI22_X1 U17717 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14318) );
  AOI22_X1 U17718 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14317) );
  NAND4_X1 U17719 ( .A1(n14320), .A2(n14319), .A3(n14318), .A4(n14317), .ZN(
        n14321) );
  OR2_X1 U17720 ( .A1(n14322), .A2(n14321), .ZN(n18230) );
  INV_X1 U17721 ( .A(n14323), .ZN(n14324) );
  AOI21_X1 U17722 ( .B1(n9653), .B2(n14324), .A(P3_EBX_REG_15__SCAN_IN), .ZN(
        n14325) );
  NOR2_X1 U17723 ( .A1(n14326), .A2(n14325), .ZN(n14327) );
  MUX2_X1 U17724 ( .A(n18230), .B(n14327), .S(n18148), .Z(P3_U2688) );
  INV_X1 U17725 ( .A(n14328), .ZN(n14334) );
  AOI21_X1 U17726 ( .B1(n14334), .B2(n17886), .A(n16807), .ZN(n14329) );
  INV_X1 U17727 ( .A(n14329), .ZN(n19420) );
  NOR2_X1 U17728 ( .A1(n19570), .A2(n19420), .ZN(n14331) );
  MUX2_X1 U17729 ( .A(n14331), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n14330), .Z(P3_U3284) );
  NAND3_X1 U17730 ( .A1(n14334), .A2(n14333), .A3(n17886), .ZN(n18963) );
  INV_X1 U17731 ( .A(n19538), .ZN(n14335) );
  OAI21_X1 U17732 ( .B1(n18963), .B2(P3_FLUSH_REG_SCAN_IN), .A(n14335), .ZN(
        n14336) );
  AND2_X1 U17733 ( .A1(n19011), .A2(n14336), .ZN(n18967) );
  INV_X1 U17734 ( .A(n18965), .ZN(n19560) );
  NOR2_X1 U17735 ( .A1(n19444), .A2(n17521), .ZN(n18579) );
  NOR2_X1 U17736 ( .A1(n19560), .A2(n18579), .ZN(n18969) );
  AOI21_X1 U17737 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18969), .ZN(n18970) );
  NOR2_X1 U17738 ( .A1(n18967), .A2(n18970), .ZN(n14338) );
  NAND3_X1 U17739 ( .A1(n19555), .A2(n19539), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n19085) );
  INV_X1 U17740 ( .A(n19085), .ZN(n19309) );
  NAND2_X1 U17741 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19407), .ZN(n19019) );
  INV_X1 U17742 ( .A(n18967), .ZN(n18975) );
  NAND2_X1 U17743 ( .A1(n19019), .A2(n18975), .ZN(n18968) );
  OR2_X1 U17744 ( .A1(n19309), .A2(n18968), .ZN(n14337) );
  MUX2_X1 U17745 ( .A(n14338), .B(n14337), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  OAI222_X1 U17746 ( .A1(n15055), .A2(n15081), .B1(n14340), .B2(n20599), .C1(
        n14339), .C2(n20594), .ZN(P1_U2844) );
  XNOR2_X1 U17747 ( .A(n10870), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17410) );
  INV_X1 U17748 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19595) );
  NOR2_X1 U17749 ( .A1(n16416), .A2(n19595), .ZN(n17405) );
  OAI21_X1 U17750 ( .B1(n15932), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14341), .ZN(n17408) );
  OAI21_X1 U17751 ( .B1(n16354), .B2(n14342), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14343) );
  OAI21_X1 U17752 ( .B1(n16422), .B2(n17408), .A(n14343), .ZN(n14344) );
  AOI211_X1 U17753 ( .C1(n17410), .C2(n16415), .A(n17405), .B(n14344), .ZN(
        n14345) );
  OAI21_X1 U17754 ( .B1(n15938), .B2(n16429), .A(n14345), .ZN(P2_U3014) );
  XOR2_X1 U17755 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14351), .Z(
        n14352) );
  NOR2_X1 U17756 ( .A1(n14354), .A2(n14355), .ZN(n14356) );
  INV_X1 U17757 ( .A(n16443), .ZN(n14357) );
  INV_X1 U17758 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21531) );
  OAI21_X1 U17759 ( .B1(n16446), .B2(n16173), .A(n21531), .ZN(n14358) );
  NOR2_X1 U17760 ( .A1(n19705), .A2(n20439), .ZN(n14364) );
  AOI21_X1 U17761 ( .B1(n16435), .B2(n14358), .A(n14364), .ZN(n14359) );
  OAI21_X1 U17762 ( .B1(n16057), .B2(n16722), .A(n14359), .ZN(n14363) );
  NAND2_X1 U17763 ( .A1(n15616), .A2(n14360), .ZN(n14361) );
  NAND2_X1 U17764 ( .A1(n9607), .A2(n14361), .ZN(n15955) );
  NOR2_X1 U17765 ( .A1(n15955), .A2(n19728), .ZN(n14362) );
  AOI21_X1 U17766 ( .B1(n16354), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14364), .ZN(n14366) );
  NAND2_X1 U17767 ( .A1(n9761), .A2(n16425), .ZN(n14365) );
  OAI211_X1 U17768 ( .C1(n15955), .C2(n16429), .A(n14366), .B(n14365), .ZN(
        n14367) );
  NAND2_X1 U17769 ( .A1(n14710), .A2(n20536), .ZN(n14378) );
  OAI22_X1 U17770 ( .A1(n20560), .A2(n14708), .B1(n14370), .B2(n20565), .ZN(
        n14376) );
  INV_X1 U17771 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14374) );
  INV_X1 U17772 ( .A(n14371), .ZN(n14735) );
  INV_X1 U17773 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21354) );
  NOR3_X1 U17774 ( .A1(n14950), .A2(n14735), .A3(n21354), .ZN(n14722) );
  INV_X1 U17775 ( .A(n14722), .ZN(n14373) );
  NAND2_X1 U17776 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14372) );
  AOI21_X1 U17777 ( .B1(n20517), .B2(n14372), .A(n14733), .ZN(n14725) );
  AOI21_X1 U17778 ( .B1(n14374), .B2(n14373), .A(n14725), .ZN(n14375) );
  AOI211_X1 U17779 ( .C1(n20574), .C2(P1_EBX_REG_30__SCAN_IN), .A(n14376), .B(
        n14375), .ZN(n14377) );
  OAI211_X1 U17780 ( .C1(n20589), .C2(n14379), .A(n14378), .B(n14377), .ZN(
        P1_U2810) );
  INV_X1 U17781 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14380) );
  OAI222_X1 U17782 ( .A1(n15055), .A2(n15071), .B1(n14380), .B2(n20599), .C1(
        n14379), .C2(n20594), .ZN(P1_U2842) );
  AOI22_X1 U17783 ( .A1(n14435), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14384) );
  AOI22_X1 U17784 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14383) );
  AOI22_X1 U17785 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14382) );
  AOI22_X1 U17786 ( .A1(n10818), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14381) );
  NAND4_X1 U17787 ( .A1(n14384), .A2(n14383), .A3(n14382), .A4(n14381), .ZN(
        n14390) );
  AOI22_X1 U17788 ( .A1(n14479), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10835), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14388) );
  AOI22_X1 U17789 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9591), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14387) );
  AOI22_X1 U17790 ( .A1(n9588), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14386) );
  AOI22_X1 U17791 ( .A1(n9587), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n9592), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14385) );
  NAND4_X1 U17792 ( .A1(n14388), .A2(n14387), .A3(n14386), .A4(n14385), .ZN(
        n14389) );
  OR2_X1 U17793 ( .A1(n14390), .A2(n14389), .ZN(n16022) );
  AND2_X1 U17794 ( .A1(n16027), .A2(n16022), .ZN(n14392) );
  AOI22_X1 U17795 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n14435), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14397) );
  AOI22_X1 U17796 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9578), .B1(n9579), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14396) );
  AOI22_X1 U17797 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10806), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14395) );
  AOI22_X1 U17798 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10818), .B1(
        n9585), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14394) );
  NAND4_X1 U17799 ( .A1(n14397), .A2(n14396), .A3(n14395), .A4(n14394), .ZN(
        n14403) );
  AOI22_X1 U17800 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10835), .B1(
        n14479), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14401) );
  AOI22_X1 U17801 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n9591), .B1(n9589), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14400) );
  AOI22_X1 U17802 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9588), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14399) );
  AOI22_X1 U17803 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10823), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14398) );
  NAND4_X1 U17804 ( .A1(n14401), .A2(n14400), .A3(n14399), .A4(n14398), .ZN(
        n14402) );
  OR2_X1 U17805 ( .A1(n14403), .A2(n14402), .ZN(n16017) );
  INV_X1 U17806 ( .A(n16013), .ZN(n14414) );
  AOI22_X1 U17807 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n14435), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14407) );
  AOI22_X1 U17808 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n9578), .B1(n9579), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14406) );
  AOI22_X1 U17809 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10806), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14405) );
  AOI22_X1 U17810 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10818), .B1(
        n9585), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14404) );
  NAND4_X1 U17811 ( .A1(n14407), .A2(n14406), .A3(n14405), .A4(n14404), .ZN(
        n14413) );
  AOI22_X1 U17812 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10835), .B1(
        n14479), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14411) );
  AOI22_X1 U17813 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n9591), .B1(n9589), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14410) );
  AOI22_X1 U17814 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n9588), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14409) );
  AOI22_X1 U17815 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10823), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14408) );
  NAND4_X1 U17816 ( .A1(n14411), .A2(n14410), .A3(n14409), .A4(n14408), .ZN(
        n14412) );
  AOI22_X1 U17817 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n14435), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14418) );
  AOI22_X1 U17818 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n9578), .B1(n9579), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14417) );
  AOI22_X1 U17819 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10806), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14416) );
  AOI22_X1 U17820 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10818), .B1(
        n9585), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14415) );
  NAND4_X1 U17821 ( .A1(n14418), .A2(n14417), .A3(n14416), .A4(n14415), .ZN(
        n14424) );
  AOI22_X1 U17822 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10835), .B1(
        n14479), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14422) );
  AOI22_X1 U17823 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n9591), .B1(n9589), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14421) );
  AOI22_X1 U17824 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n9588), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14420) );
  AOI22_X1 U17825 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10823), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14419) );
  NAND4_X1 U17826 ( .A1(n14422), .A2(n14421), .A3(n14420), .A4(n14419), .ZN(
        n14423) );
  NOR2_X1 U17827 ( .A1(n14424), .A2(n14423), .ZN(n16009) );
  AOI22_X1 U17828 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n14435), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14428) );
  AOI22_X1 U17829 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n9578), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14427) );
  AOI22_X1 U17830 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10806), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14426) );
  AOI22_X1 U17831 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10818), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14425) );
  NAND4_X1 U17832 ( .A1(n14428), .A2(n14427), .A3(n14426), .A4(n14425), .ZN(
        n14434) );
  AOI22_X1 U17833 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10835), .B1(
        n14479), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14432) );
  AOI22_X1 U17834 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n9591), .B1(n9589), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14431) );
  AOI22_X1 U17835 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n9588), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14430) );
  AOI22_X1 U17836 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10823), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14429) );
  NAND4_X1 U17837 ( .A1(n14432), .A2(n14431), .A3(n14430), .A4(n14429), .ZN(
        n14433) );
  OR2_X1 U17838 ( .A1(n14434), .A2(n14433), .ZN(n16004) );
  AOI22_X1 U17839 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n14435), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14439) );
  AOI22_X1 U17840 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n9578), .B1(n9579), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14438) );
  AOI22_X1 U17841 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n10806), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14437) );
  AOI22_X1 U17842 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n10818), .B1(
        n9585), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14436) );
  NAND4_X1 U17843 ( .A1(n14439), .A2(n14438), .A3(n14437), .A4(n14436), .ZN(
        n14445) );
  AOI22_X1 U17844 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10835), .B1(
        n14479), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14443) );
  AOI22_X1 U17845 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n9591), .B1(n9590), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14442) );
  AOI22_X1 U17846 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n9588), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14441) );
  AOI22_X1 U17847 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n9587), .B1(n9592), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14440) );
  NAND4_X1 U17848 ( .A1(n14443), .A2(n14442), .A3(n14441), .A4(n14440), .ZN(
        n14444) );
  OR2_X1 U17849 ( .A1(n14445), .A2(n14444), .ZN(n15998) );
  AOI22_X1 U17850 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n14435), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14449) );
  AOI22_X1 U17851 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n9578), .B1(
        n10805), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14448) );
  AOI22_X1 U17852 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10806), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14447) );
  AOI22_X1 U17853 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10818), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14446) );
  NAND4_X1 U17854 ( .A1(n14449), .A2(n14448), .A3(n14447), .A4(n14446), .ZN(
        n14455) );
  AOI22_X1 U17855 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10835), .B1(
        n14479), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14453) );
  AOI22_X1 U17856 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n9591), .B1(n9590), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14452) );
  AOI22_X1 U17857 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n9588), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14451) );
  AOI22_X1 U17858 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10823), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14450) );
  NAND4_X1 U17859 ( .A1(n14453), .A2(n14452), .A3(n14451), .A4(n14450), .ZN(
        n14454) );
  OR2_X1 U17860 ( .A1(n14455), .A2(n14454), .ZN(n15993) );
  NAND2_X1 U17861 ( .A1(n14624), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n14459) );
  NAND2_X1 U17862 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14458) );
  NAND2_X1 U17863 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n14457) );
  NAND2_X1 U17864 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14456) );
  AND4_X1 U17865 ( .A1(n14459), .A2(n14458), .A3(n14457), .A4(n14456), .ZN(
        n14462) );
  AOI22_X1 U17866 ( .A1(n14629), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14628), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14460) );
  XNOR2_X1 U17867 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14621) );
  NAND4_X1 U17868 ( .A1(n14462), .A2(n14461), .A3(n14460), .A4(n14621), .ZN(
        n14471) );
  NAND2_X1 U17869 ( .A1(n14624), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n14466) );
  NAND2_X1 U17870 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n14465) );
  NAND2_X1 U17871 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n14464) );
  NAND2_X1 U17872 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n14463) );
  AND4_X1 U17873 ( .A1(n14466), .A2(n14465), .A3(n14464), .A4(n14463), .ZN(
        n14469) );
  INV_X1 U17874 ( .A(n14621), .ZN(n14631) );
  AOI22_X1 U17875 ( .A1(n14629), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9570), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14467) );
  NAND4_X1 U17876 ( .A1(n14469), .A2(n14631), .A3(n14468), .A4(n14467), .ZN(
        n14470) );
  AND2_X1 U17877 ( .A1(n14471), .A2(n14470), .ZN(n14508) );
  INV_X1 U17878 ( .A(n14508), .ZN(n14511) );
  AOI22_X1 U17879 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10835), .B1(
        n14435), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14478) );
  AOI22_X1 U17880 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n9588), .B1(n9592), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14477) );
  AOI22_X1 U17881 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n9590), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14476) );
  AOI22_X1 U17882 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n9587), .B1(n9591), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14475) );
  NAND4_X1 U17883 ( .A1(n14478), .A2(n14477), .A3(n14476), .A4(n14475), .ZN(
        n14487) );
  AOI22_X1 U17884 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14479), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14485) );
  AOI22_X1 U17885 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10806), .B1(
        n9577), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14484) );
  AOI22_X1 U17886 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(n9584), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14483) );
  AOI22_X1 U17887 ( .A1(n10805), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10818), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14482) );
  NAND4_X1 U17888 ( .A1(n14485), .A2(n14484), .A3(n14483), .A4(n14482), .ZN(
        n14486) );
  OR2_X1 U17889 ( .A1(n14487), .A2(n14486), .ZN(n14506) );
  NAND2_X1 U17890 ( .A1(n14560), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n14491) );
  NAND2_X1 U17891 ( .A1(n10019), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14490) );
  NAND2_X1 U17892 ( .A1(n14628), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n14488) );
  AND4_X1 U17893 ( .A1(n14491), .A2(n14490), .A3(n14489), .A4(n14488), .ZN(
        n14494) );
  AOI22_X1 U17894 ( .A1(n14624), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14604), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14493) );
  AOI22_X1 U17895 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14492) );
  NAND4_X1 U17896 ( .A1(n14494), .A2(n14493), .A3(n14492), .A4(n14621), .ZN(
        n14503) );
  NAND2_X1 U17897 ( .A1(n14560), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n14498) );
  NAND2_X1 U17898 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n14497) );
  NAND2_X1 U17899 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n14496) );
  NAND2_X1 U17900 ( .A1(n9581), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14495) );
  AND4_X1 U17901 ( .A1(n14498), .A2(n14497), .A3(n14496), .A4(n14495), .ZN(
        n14501) );
  AOI22_X1 U17902 ( .A1(n14624), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9569), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14499) );
  NAND4_X1 U17903 ( .A1(n14501), .A2(n14631), .A3(n14500), .A4(n14499), .ZN(
        n14502) );
  NAND2_X1 U17904 ( .A1(n14503), .A2(n14502), .ZN(n15977) );
  INV_X1 U17905 ( .A(n15977), .ZN(n14504) );
  NAND2_X1 U17906 ( .A1(n14506), .A2(n14504), .ZN(n14512) );
  XOR2_X1 U17907 ( .A(n14511), .B(n14512), .Z(n14505) );
  NAND2_X1 U17908 ( .A1(n14505), .A2(n14571), .ZN(n15980) );
  NOR2_X1 U17909 ( .A1(n9596), .A2(n15977), .ZN(n14507) );
  OAI22_X1 U17910 ( .A1(n14507), .A2(n14506), .B1(n14512), .B2(n9595), .ZN(
        n15979) );
  NOR2_X1 U17911 ( .A1(n15980), .A2(n15979), .ZN(n14510) );
  NAND2_X1 U17912 ( .A1(n9595), .A2(n14508), .ZN(n15981) );
  NOR3_X1 U17913 ( .A1(n15979), .A2(n15977), .A3(n15981), .ZN(n14509) );
  NOR2_X1 U17914 ( .A1(n14512), .A2(n14511), .ZN(n14529) );
  NAND2_X1 U17915 ( .A1(n14624), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n14516) );
  NAND2_X1 U17916 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14515) );
  NAND2_X1 U17917 ( .A1(n9581), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n14514) );
  NAND2_X1 U17918 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n14513) );
  AND4_X1 U17919 ( .A1(n14516), .A2(n14515), .A3(n14514), .A4(n14513), .ZN(
        n14519) );
  AOI22_X1 U17920 ( .A1(n14629), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14628), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14517) );
  NAND4_X1 U17921 ( .A1(n14519), .A2(n14518), .A3(n14517), .A4(n14621), .ZN(
        n14528) );
  NAND2_X1 U17922 ( .A1(n14624), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n14523) );
  NAND2_X1 U17923 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n14522) );
  NAND2_X1 U17924 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14521) );
  NAND2_X1 U17925 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n14520) );
  AND4_X1 U17926 ( .A1(n14523), .A2(n14522), .A3(n14521), .A4(n14520), .ZN(
        n14526) );
  AOI22_X1 U17927 ( .A1(n14629), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14628), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14524) );
  NAND4_X1 U17928 ( .A1(n14526), .A2(n14631), .A3(n14525), .A4(n14524), .ZN(
        n14527) );
  AND2_X1 U17929 ( .A1(n14528), .A2(n14527), .ZN(n14530) );
  NAND2_X1 U17930 ( .A1(n14529), .A2(n14530), .ZN(n14552) );
  OAI211_X1 U17931 ( .C1(n14529), .C2(n14530), .A(n14552), .B(n14571), .ZN(
        n14547) );
  NAND2_X1 U17932 ( .A1(n9596), .A2(n14530), .ZN(n15972) );
  NAND2_X1 U17933 ( .A1(n14624), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n14534) );
  NAND2_X1 U17934 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14533) );
  NAND2_X1 U17935 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n14532) );
  NAND2_X1 U17936 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n14531) );
  AND4_X1 U17937 ( .A1(n14534), .A2(n14533), .A3(n14532), .A4(n14531), .ZN(
        n14537) );
  AOI22_X1 U17938 ( .A1(n14629), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9569), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14535) );
  NAND4_X1 U17939 ( .A1(n14537), .A2(n14536), .A3(n14535), .A4(n14621), .ZN(
        n14546) );
  NAND2_X1 U17940 ( .A1(n14624), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n14541) );
  NAND2_X1 U17941 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n14540) );
  NAND2_X1 U17942 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14539) );
  NAND2_X1 U17943 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n14538) );
  AND4_X1 U17944 ( .A1(n14541), .A2(n14540), .A3(n14539), .A4(n14538), .ZN(
        n14544) );
  AOI22_X1 U17945 ( .A1(n14629), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9570), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14542) );
  NAND4_X1 U17946 ( .A1(n14544), .A2(n14631), .A3(n14543), .A4(n14542), .ZN(
        n14545) );
  NAND2_X1 U17947 ( .A1(n14546), .A2(n14545), .ZN(n15964) );
  NOR2_X2 U17948 ( .A1(n14548), .A2(n14547), .ZN(n15963) );
  XNOR2_X1 U17949 ( .A(n14552), .B(n15964), .ZN(n14550) );
  NOR2_X1 U17950 ( .A1(n14550), .A2(n14549), .ZN(n15966) );
  NAND2_X1 U17951 ( .A1(n15963), .A2(n15966), .ZN(n14551) );
  OAI21_X2 U17952 ( .B1(n15973), .B2(n10471), .A(n14551), .ZN(n14576) );
  INV_X1 U17953 ( .A(n14570), .ZN(n14573) );
  NAND2_X1 U17954 ( .A1(n14560), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n14556) );
  NAND2_X1 U17955 ( .A1(n10019), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14555) );
  NAND2_X1 U17956 ( .A1(n9570), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n14553) );
  AND4_X1 U17957 ( .A1(n14556), .A2(n14555), .A3(n14554), .A4(n14553), .ZN(
        n14559) );
  AOI22_X1 U17958 ( .A1(n14624), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9580), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14558) );
  INV_X1 U17959 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n20029) );
  AOI22_X1 U17960 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14557) );
  NAND4_X1 U17961 ( .A1(n14559), .A2(n14558), .A3(n14557), .A4(n14621), .ZN(
        n14569) );
  NAND2_X1 U17962 ( .A1(n14560), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n14564) );
  NAND2_X1 U17963 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n14563) );
  NAND2_X1 U17964 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n14562) );
  NAND2_X1 U17965 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14561) );
  AND4_X1 U17966 ( .A1(n14564), .A2(n14563), .A3(n14562), .A4(n14561), .ZN(
        n14567) );
  AOI22_X1 U17967 ( .A1(n14596), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9570), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14566) );
  NAND4_X1 U17968 ( .A1(n14567), .A2(n14631), .A3(n14566), .A4(n14565), .ZN(
        n14568) );
  NAND2_X1 U17969 ( .A1(n14569), .A2(n14568), .ZN(n14578) );
  INV_X1 U17970 ( .A(n14578), .ZN(n14572) );
  OAI211_X1 U17971 ( .C1(n14573), .C2(n14572), .A(n14571), .B(n14611), .ZN(
        n14575) );
  AND2_X2 U17972 ( .A1(n14576), .A2(n14574), .ZN(n15952) );
  NOR2_X1 U17973 ( .A1(n14576), .A2(n14574), .ZN(n14577) );
  NOR2_X2 U17974 ( .A1(n15952), .A2(n14577), .ZN(n15960) );
  NOR2_X1 U17975 ( .A1(n15978), .A2(n14578), .ZN(n15959) );
  INV_X1 U17976 ( .A(n15952), .ZN(n14595) );
  NAND2_X1 U17977 ( .A1(n14624), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n14582) );
  NAND2_X1 U17978 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14581) );
  NAND2_X1 U17979 ( .A1(n14604), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n14580) );
  NAND2_X1 U17980 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14579) );
  AND4_X1 U17981 ( .A1(n14582), .A2(n14581), .A3(n14580), .A4(n14579), .ZN(
        n14585) );
  AOI22_X1 U17982 ( .A1(n14629), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9570), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14583) );
  NAND4_X1 U17983 ( .A1(n14585), .A2(n14584), .A3(n14583), .A4(n14621), .ZN(
        n14594) );
  NAND2_X1 U17984 ( .A1(n14624), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n14589) );
  NAND2_X1 U17985 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n14588) );
  NAND2_X1 U17986 ( .A1(n9581), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n14587) );
  NAND2_X1 U17987 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n14586) );
  AND4_X1 U17988 ( .A1(n14589), .A2(n14588), .A3(n14587), .A4(n14586), .ZN(
        n14592) );
  AOI22_X1 U17989 ( .A1(n14629), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14628), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14590) );
  NAND4_X1 U17990 ( .A1(n14592), .A2(n14631), .A3(n14591), .A4(n14590), .ZN(
        n14593) );
  NAND2_X1 U17991 ( .A1(n14594), .A2(n14593), .ZN(n15953) );
  AOI22_X1 U17992 ( .A1(n14624), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14628), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14598) );
  AND2_X1 U17993 ( .A1(n14598), .A2(n14597), .ZN(n14601) );
  AOI22_X1 U17994 ( .A1(n14629), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14600) );
  AOI22_X1 U17995 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14604), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14599) );
  NAND4_X1 U17996 ( .A1(n14601), .A2(n14631), .A3(n14600), .A4(n14599), .ZN(
        n14610) );
  AOI22_X1 U17997 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9569), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14602) );
  AND2_X1 U17998 ( .A1(n14603), .A2(n14602), .ZN(n14608) );
  AOI22_X1 U17999 ( .A1(n14605), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14604), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14607) );
  AOI22_X1 U18000 ( .A1(n14618), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14606) );
  NAND4_X1 U18001 ( .A1(n14608), .A2(n14607), .A3(n14606), .A4(n14621), .ZN(
        n14609) );
  NAND2_X1 U18002 ( .A1(n14610), .A2(n14609), .ZN(n14615) );
  INV_X1 U18003 ( .A(n14611), .ZN(n15951) );
  INV_X1 U18004 ( .A(n15953), .ZN(n14612) );
  AND2_X1 U18005 ( .A1(n15978), .A2(n14612), .ZN(n14613) );
  NAND2_X1 U18006 ( .A1(n15951), .A2(n14613), .ZN(n14614) );
  NOR2_X1 U18007 ( .A1(n14614), .A2(n14615), .ZN(n14616) );
  AOI21_X1 U18008 ( .B1(n14615), .B2(n14614), .A(n14616), .ZN(n15947) );
  INV_X1 U18009 ( .A(n14616), .ZN(n14617) );
  AOI22_X1 U18010 ( .A1(n14624), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14620) );
  AOI22_X1 U18011 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14619) );
  NAND2_X1 U18012 ( .A1(n14620), .A2(n14619), .ZN(n14637) );
  AOI22_X1 U18013 ( .A1(n14629), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9569), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14623) );
  NAND3_X1 U18014 ( .A1(n14623), .A2(n14622), .A3(n14621), .ZN(n14636) );
  AOI22_X1 U18015 ( .A1(n14624), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14618), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14627) );
  AOI22_X1 U18016 ( .A1(n9580), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14626) );
  NAND2_X1 U18017 ( .A1(n14627), .A2(n14626), .ZN(n14635) );
  AOI22_X1 U18018 ( .A1(n14629), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9570), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14633) );
  NAND3_X1 U18019 ( .A1(n14633), .A2(n14632), .A3(n14631), .ZN(n14634) );
  OAI22_X1 U18020 ( .A1(n14637), .A2(n14636), .B1(n14635), .B2(n14634), .ZN(
        n14638) );
  INV_X1 U18021 ( .A(n14638), .ZN(n14639) );
  XNOR2_X1 U18022 ( .A(n14640), .B(n14639), .ZN(n14648) );
  INV_X1 U18023 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14643) );
  NAND2_X1 U18024 ( .A1(n16136), .A2(BUF2_REG_30__SCAN_IN), .ZN(n14642) );
  AOI22_X1 U18025 ( .A1(n16137), .A2(n19697), .B1(n19647), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14641) );
  OAI211_X1 U18026 ( .C1(n16140), .C2(n14643), .A(n14642), .B(n14641), .ZN(
        n14644) );
  AOI21_X1 U18027 ( .B1(n14690), .B2(n19648), .A(n14644), .ZN(n14645) );
  OAI21_X1 U18028 ( .B1(n14648), .B2(n16144), .A(n14645), .ZN(P2_U2889) );
  NOR2_X1 U18029 ( .A1(n14687), .A2(n16043), .ZN(n14646) );
  AOI21_X1 U18030 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n16043), .A(n14646), .ZN(
        n14647) );
  OAI21_X1 U18031 ( .B1(n14648), .B2(n16029), .A(n14647), .ZN(P2_U2857) );
  AOI21_X1 U18032 ( .B1(n14649), .B2(n15565), .A(n15577), .ZN(n14654) );
  OAI22_X1 U18033 ( .A1(n15573), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n14650), .ZN(n14651) );
  AOI21_X1 U18034 ( .B1(n14652), .B2(n15565), .A(n14651), .ZN(n14653) );
  OAI22_X1 U18035 ( .A1(n14654), .A2(n10177), .B1(n15577), .B2(n14653), .ZN(
        P1_U3474) );
  OR2_X1 U18036 ( .A1(n14656), .A2(n14655), .ZN(n14676) );
  NAND3_X1 U18037 ( .A1(n14676), .A2(n14675), .A3(n19721), .ZN(n14674) );
  NAND2_X1 U18038 ( .A1(n14659), .A2(n14658), .ZN(n14661) );
  XOR2_X1 U18039 ( .A(n14661), .B(n14660), .Z(n14679) );
  INV_X1 U18040 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20396) );
  INV_X1 U18041 ( .A(n14662), .ZN(n14663) );
  NAND2_X1 U18042 ( .A1(n14665), .A2(n14663), .ZN(n15883) );
  NAND2_X1 U18043 ( .A1(n14665), .A2(n14664), .ZN(n14667) );
  NAND2_X1 U18044 ( .A1(n14667), .A2(n14666), .ZN(n14668) );
  NAND2_X1 U18045 ( .A1(n15883), .A2(n14668), .ZN(n16148) );
  INV_X1 U18046 ( .A(n16148), .ZN(n20469) );
  NAND2_X1 U18047 ( .A1(n16731), .A2(n20469), .ZN(n14671) );
  INV_X1 U18048 ( .A(n14669), .ZN(n16716) );
  AOI22_X1 U18049 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16714), .B1(
        n16716), .B2(n16715), .ZN(n14670) );
  OAI211_X1 U18050 ( .C1(n20396), .C2(n16416), .A(n14671), .B(n14670), .ZN(
        n14672) );
  AOI21_X1 U18051 ( .B1(n14679), .B2(n19726), .A(n14672), .ZN(n14673) );
  OAI211_X1 U18052 ( .C1(n19728), .C2(n13780), .A(n14674), .B(n14673), .ZN(
        P2_U3043) );
  NAND3_X1 U18053 ( .A1(n14676), .A2(n14675), .A3(n16415), .ZN(n14681) );
  AOI22_X1 U18054 ( .A1(n16354), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_REIP_REG_3__SCAN_IN), .B2(n19604), .ZN(n14677) );
  OAI21_X1 U18055 ( .B1(n16406), .B2(n15904), .A(n14677), .ZN(n14678) );
  AOI21_X1 U18056 ( .B1(n14679), .B2(n16394), .A(n14678), .ZN(n14680) );
  OAI211_X1 U18057 ( .C1(n16429), .C2(n13780), .A(n14681), .B(n14680), .ZN(
        P2_U3011) );
  INV_X1 U18058 ( .A(n15596), .ZN(n14694) );
  OAI21_X1 U18059 ( .B1(n15596), .B2(n19616), .A(n15912), .ZN(n14683) );
  NAND2_X1 U18060 ( .A1(n14683), .A2(n14682), .ZN(n14692) );
  AOI22_X1 U18061 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n19605), .B1(n15934), 
        .B2(P2_EBX_REG_30__SCAN_IN), .ZN(n14685) );
  NAND2_X1 U18062 ( .A1(n15930), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14684) );
  OAI211_X1 U18063 ( .C1(n14686), .C2(n15875), .A(n14685), .B(n14684), .ZN(
        n14689) );
  NOR2_X1 U18064 ( .A1(n14687), .A2(n15937), .ZN(n14688) );
  AOI211_X1 U18065 ( .C1(n14690), .C2(n15933), .A(n14689), .B(n14688), .ZN(
        n14691) );
  OAI211_X1 U18066 ( .C1(n14694), .C2(n14693), .A(n14692), .B(n14691), .ZN(
        P2_U2825) );
  INV_X1 U18067 ( .A(n14695), .ZN(n14696) );
  XNOR2_X1 U18068 ( .A(n14697), .B(n14696), .ZN(n19725) );
  OAI21_X1 U18069 ( .B1(n14700), .B2(n14699), .A(n14698), .ZN(n14701) );
  INV_X1 U18070 ( .A(n14701), .ZN(n19720) );
  INV_X1 U18071 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15920) );
  NAND2_X1 U18072 ( .A1(n19604), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n19735) );
  OAI21_X1 U18073 ( .B1(n16419), .B2(n15920), .A(n19735), .ZN(n14702) );
  AOI21_X1 U18074 ( .B1(n19720), .B2(n16415), .A(n14702), .ZN(n14703) );
  OAI21_X1 U18075 ( .B1(n16406), .B2(n15916), .A(n14703), .ZN(n14704) );
  AOI21_X1 U18076 ( .B1(n16394), .B2(n19725), .A(n14704), .ZN(n14705) );
  OAI21_X1 U18077 ( .B1(n19727), .B2(n16429), .A(n14705), .ZN(P2_U3012) );
  NAND2_X1 U18078 ( .A1(n20641), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14706) );
  OAI211_X1 U18079 ( .C1(n20654), .C2(n14708), .A(n14707), .B(n14706), .ZN(
        n14709) );
  AOI21_X1 U18080 ( .B1(n14710), .B2(n20649), .A(n14709), .ZN(n14711) );
  OAI21_X1 U18081 ( .B1(n14712), .B2(n15339), .A(n14711), .ZN(P1_U2969) );
  OR2_X1 U18082 ( .A1(n15142), .A2(n14713), .ZN(n14715) );
  NAND2_X1 U18083 ( .A1(n14721), .A2(n14714), .ZN(n14717) );
  AOI22_X1 U18084 ( .A1(n15137), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15142), .ZN(n14716) );
  OAI211_X1 U18085 ( .C1(n15135), .C2(n17433), .A(n14717), .B(n14716), .ZN(
        P1_U2873) );
  NAND2_X1 U18086 ( .A1(n15002), .A2(n12013), .ZN(n14720) );
  OR2_X1 U18087 ( .A1(n14718), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n14719) );
  MUX2_X1 U18088 ( .A(n14720), .B(n14719), .S(n21382), .Z(P1_U3487) );
  INV_X1 U18089 ( .A(n14721), .ZN(n14728) );
  AOI22_X1 U18090 ( .A1(n20541), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20579), .ZN(n14724) );
  NAND3_X1 U18091 ( .A1(n14722), .A2(P1_REIP_REG_30__SCAN_IN), .A3(n21358), 
        .ZN(n14723) );
  OAI211_X1 U18092 ( .C1(n14725), .C2(n21358), .A(n14724), .B(n14723), .ZN(
        n14726) );
  AOI21_X1 U18093 ( .B1(n15022), .B2(n20532), .A(n14726), .ZN(n14727) );
  OAI21_X1 U18094 ( .B1(n14728), .B2(n17350), .A(n14727), .ZN(P1_U2809) );
  OAI21_X1 U18095 ( .B1(n12732), .B2(n14732), .A(n14731), .ZN(n15359) );
  INV_X1 U18096 ( .A(n15359), .ZN(n14741) );
  INV_X1 U18097 ( .A(n14733), .ZN(n14739) );
  OAI22_X1 U18098 ( .A1(n20560), .A2(n15159), .B1(n14734), .B2(n20565), .ZN(
        n14737) );
  NOR3_X1 U18099 ( .A1(n14950), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n14735), 
        .ZN(n14736) );
  AOI211_X1 U18100 ( .C1(P1_EBX_REG_29__SCAN_IN), .C2(n20541), .A(n14737), .B(
        n14736), .ZN(n14738) );
  OAI21_X1 U18101 ( .B1(n14739), .B2(n21354), .A(n14738), .ZN(n14740) );
  AOI21_X1 U18102 ( .B1(n14741), .B2(n20532), .A(n14740), .ZN(n14742) );
  OAI21_X1 U18103 ( .B1(n15165), .B2(n17350), .A(n14742), .ZN(P1_U2811) );
  AOI21_X1 U18104 ( .B1(n14746), .B2(n14761), .A(n14745), .ZN(n15360) );
  INV_X1 U18105 ( .A(n14747), .ZN(n14750) );
  INV_X1 U18106 ( .A(n20562), .ZN(n14748) );
  AOI21_X1 U18107 ( .B1(n20555), .B2(n14750), .A(n14748), .ZN(n14766) );
  INV_X1 U18108 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n14754) );
  OAI22_X1 U18109 ( .A1(n20560), .A2(n15174), .B1(n14749), .B2(n20565), .ZN(
        n14752) );
  NOR3_X1 U18110 ( .A1(n14950), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14750), 
        .ZN(n14751) );
  AOI211_X1 U18111 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n20541), .A(n14752), .B(
        n14751), .ZN(n14753) );
  OAI21_X1 U18112 ( .B1(n14766), .B2(n14754), .A(n14753), .ZN(n14755) );
  AOI21_X1 U18113 ( .B1(n15360), .B2(n20532), .A(n14755), .ZN(n14756) );
  OAI21_X1 U18114 ( .B1(n15181), .B2(n17350), .A(n14756), .ZN(P1_U2813) );
  AOI21_X1 U18115 ( .B1(n14758), .B2(n14757), .A(n14743), .ZN(n15191) );
  INV_X1 U18116 ( .A(n15191), .ZN(n15090) );
  NAND2_X1 U18117 ( .A1(n12914), .A2(n14759), .ZN(n14760) );
  NAND2_X1 U18118 ( .A1(n14761), .A2(n14760), .ZN(n15027) );
  INV_X1 U18119 ( .A(n15027), .ZN(n15377) );
  AOI21_X1 U18120 ( .B1(n20555), .B2(n14762), .A(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14765) );
  AOI22_X1 U18121 ( .A1(n20575), .A2(n15187), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20579), .ZN(n14764) );
  NAND2_X1 U18122 ( .A1(n20541), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14763) );
  OAI211_X1 U18123 ( .C1(n14766), .C2(n14765), .A(n14764), .B(n14763), .ZN(
        n14767) );
  AOI21_X1 U18124 ( .B1(n15377), .B2(n20532), .A(n14767), .ZN(n14768) );
  OAI21_X1 U18125 ( .B1(n15090), .B2(n17350), .A(n14768), .ZN(P1_U2814) );
  OAI21_X1 U18126 ( .B1(n14769), .B2(n14770), .A(n14757), .ZN(n15199) );
  INV_X1 U18127 ( .A(n14771), .ZN(n14782) );
  AOI21_X1 U18128 ( .B1(n20562), .B2(n14782), .A(n14856), .ZN(n14798) );
  INV_X1 U18129 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n21524) );
  INV_X1 U18130 ( .A(n15193), .ZN(n14772) );
  AOI22_X1 U18131 ( .A1(n20575), .A2(n14772), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20579), .ZN(n14776) );
  NAND2_X1 U18132 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14773) );
  OAI211_X1 U18133 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14774), .A(n20555), 
        .B(n14773), .ZN(n14775) );
  OAI211_X1 U18134 ( .C1(n20553), .C2(n21524), .A(n14776), .B(n14775), .ZN(
        n14778) );
  NOR2_X1 U18135 ( .A1(n15029), .A2(n20589), .ZN(n14777) );
  AOI211_X1 U18136 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14798), .A(n14778), 
        .B(n14777), .ZN(n14779) );
  OAI21_X1 U18137 ( .B1(n15199), .B2(n17350), .A(n14779), .ZN(P1_U2815) );
  INV_X1 U18138 ( .A(n14780), .ZN(n14793) );
  AOI21_X1 U18139 ( .B1(n14781), .B2(n14793), .A(n14769), .ZN(n15207) );
  INV_X1 U18140 ( .A(n15207), .ZN(n15098) );
  INV_X1 U18141 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14785) );
  AOI22_X1 U18142 ( .A1(n20575), .A2(n15203), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20579), .ZN(n14784) );
  NAND3_X1 U18143 ( .A1(n20555), .A2(n21344), .A3(n14782), .ZN(n14783) );
  OAI211_X1 U18144 ( .C1(n20553), .C2(n14785), .A(n14784), .B(n14783), .ZN(
        n14786) );
  AOI21_X1 U18145 ( .B1(n14798), .B2(P1_REIP_REG_24__SCAN_IN), .A(n14786), 
        .ZN(n14790) );
  AOI21_X1 U18146 ( .B1(n14788), .B2(n14795), .A(n14787), .ZN(n15388) );
  NAND2_X1 U18147 ( .A1(n15388), .A2(n20532), .ZN(n14789) );
  OAI211_X1 U18148 ( .C1(n15098), .C2(n17350), .A(n14790), .B(n14789), .ZN(
        P1_U2816) );
  AOI21_X1 U18149 ( .B1(n14794), .B2(n14792), .A(n14780), .ZN(n15214) );
  INV_X1 U18150 ( .A(n15214), .ZN(n15103) );
  INV_X1 U18151 ( .A(n14795), .ZN(n14796) );
  AOI21_X1 U18152 ( .B1(n14797), .B2(n14809), .A(n14796), .ZN(n15397) );
  INV_X1 U18153 ( .A(n14798), .ZN(n14804) );
  AOI21_X1 U18154 ( .B1(n20555), .B2(n14799), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14803) );
  OAI22_X1 U18155 ( .A1(n20560), .A2(n15212), .B1(n14800), .B2(n20565), .ZN(
        n14801) );
  AOI21_X1 U18156 ( .B1(n20574), .B2(P1_EBX_REG_23__SCAN_IN), .A(n14801), .ZN(
        n14802) );
  OAI21_X1 U18157 ( .B1(n14804), .B2(n14803), .A(n14802), .ZN(n14805) );
  AOI21_X1 U18158 ( .B1(n15397), .B2(n20532), .A(n14805), .ZN(n14806) );
  OAI21_X1 U18159 ( .B1(n15103), .B2(n17350), .A(n14806), .ZN(P1_U2817) );
  OAI21_X1 U18160 ( .B1(n14808), .B2(n14807), .A(n14792), .ZN(n15223) );
  INV_X1 U18161 ( .A(n14809), .ZN(n14810) );
  AOI21_X1 U18162 ( .B1(n14812), .B2(n14811), .A(n14810), .ZN(n15400) );
  NAND2_X1 U18163 ( .A1(n20562), .A2(n14813), .ZN(n20518) );
  NAND2_X1 U18164 ( .A1(n14858), .A2(n14814), .ZN(n14815) );
  OR2_X1 U18165 ( .A1(n20518), .A2(n14815), .ZN(n14816) );
  NAND2_X1 U18166 ( .A1(n20517), .A2(n14816), .ZN(n14846) );
  OAI22_X1 U18167 ( .A1(n20560), .A2(n15216), .B1(n14817), .B2(n20565), .ZN(
        n14821) );
  NOR2_X1 U18168 ( .A1(n14826), .A2(n21340), .ZN(n14818) );
  AOI211_X1 U18169 ( .C1(n14819), .C2(n21340), .A(n14818), .B(n14950), .ZN(
        n14820) );
  AOI211_X1 U18170 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n20541), .A(n14821), .B(
        n14820), .ZN(n14822) );
  OAI21_X1 U18171 ( .B1(n21340), .B2(n14846), .A(n14822), .ZN(n14823) );
  AOI21_X1 U18172 ( .B1(n15400), .B2(n20532), .A(n14823), .ZN(n14824) );
  OAI21_X1 U18173 ( .B1(n15223), .B2(n17350), .A(n14824), .ZN(P1_U2818) );
  INV_X1 U18174 ( .A(n15033), .ZN(n14832) );
  NOR2_X1 U18175 ( .A1(n14846), .A2(n14826), .ZN(n14831) );
  INV_X1 U18176 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15034) );
  AOI22_X1 U18177 ( .A1(n20575), .A2(n14825), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20579), .ZN(n14829) );
  NAND3_X1 U18178 ( .A1(n20555), .A2(n14827), .A3(n14826), .ZN(n14828) );
  OAI211_X1 U18179 ( .C1(n20553), .C2(n15034), .A(n14829), .B(n14828), .ZN(
        n14830) );
  AOI211_X1 U18180 ( .C1(n14832), .C2(n20532), .A(n14831), .B(n14830), .ZN(
        n14833) );
  OAI21_X1 U18181 ( .B1(n15112), .B2(n17350), .A(n14833), .ZN(P1_U2819) );
  NAND2_X1 U18182 ( .A1(n14850), .A2(n14834), .ZN(n14835) );
  NAND2_X1 U18183 ( .A1(n14836), .A2(n14835), .ZN(n15225) );
  NOR2_X1 U18184 ( .A1(n14854), .A2(n14837), .ZN(n14838) );
  OR2_X1 U18185 ( .A1(n14839), .A2(n14838), .ZN(n15035) );
  INV_X1 U18186 ( .A(n15035), .ZN(n15417) );
  INV_X1 U18187 ( .A(n14947), .ZN(n14841) );
  INV_X1 U18188 ( .A(n20505), .ZN(n14972) );
  NOR2_X1 U18189 ( .A1(n14972), .A2(n14842), .ZN(n14903) );
  NAND3_X1 U18190 ( .A1(n14903), .A2(P1_REIP_REG_14__SCAN_IN), .A3(
        P1_REIP_REG_15__SCAN_IN), .ZN(n14908) );
  INV_X1 U18191 ( .A(n14857), .ZN(n14843) );
  NOR2_X1 U18192 ( .A1(n14908), .A2(n14843), .ZN(n14876) );
  AOI21_X1 U18193 ( .B1(n14876), .B2(n14862), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n14847) );
  OAI22_X1 U18194 ( .A1(n20560), .A2(n15227), .B1(n21510), .B2(n20565), .ZN(
        n14844) );
  AOI21_X1 U18195 ( .B1(n20574), .B2(P1_EBX_REG_20__SCAN_IN), .A(n14844), .ZN(
        n14845) );
  OAI21_X1 U18196 ( .B1(n14847), .B2(n14846), .A(n14845), .ZN(n14848) );
  AOI21_X1 U18197 ( .B1(n15417), .B2(n20532), .A(n14848), .ZN(n14849) );
  OAI21_X1 U18198 ( .B1(n15225), .B2(n17350), .A(n14849), .ZN(P1_U2820) );
  INV_X1 U18199 ( .A(n14850), .ZN(n14851) );
  AOI21_X1 U18200 ( .B1(n14852), .B2(n14872), .A(n14851), .ZN(n15237) );
  INV_X1 U18201 ( .A(n15237), .ZN(n15121) );
  INV_X1 U18202 ( .A(n14853), .ZN(n14874) );
  AOI21_X1 U18203 ( .B1(n14855), .B2(n14874), .A(n14854), .ZN(n15426) );
  AOI21_X1 U18204 ( .B1(n14857), .B2(P1_REIP_REG_15__SCAN_IN), .A(n14856), 
        .ZN(n14861) );
  NAND2_X1 U18205 ( .A1(n20517), .A2(n20518), .ZN(n20545) );
  INV_X1 U18206 ( .A(n14858), .ZN(n14859) );
  NAND2_X1 U18207 ( .A1(n20517), .A2(n14859), .ZN(n14860) );
  NAND2_X1 U18208 ( .A1(n20545), .A2(n14860), .ZN(n14929) );
  NOR2_X1 U18209 ( .A1(n14861), .A2(n14929), .ZN(n14895) );
  INV_X1 U18210 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14868) );
  INV_X1 U18211 ( .A(n14862), .ZN(n14863) );
  OAI211_X1 U18212 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(P1_REIP_REG_18__SCAN_IN), .A(n14876), .B(n14863), .ZN(n14867) );
  NAND2_X1 U18213 ( .A1(n20575), .A2(n15233), .ZN(n14864) );
  OAI211_X1 U18214 ( .C1(n20565), .C2(n15235), .A(n14864), .B(n20667), .ZN(
        n14865) );
  AOI21_X1 U18215 ( .B1(n20541), .B2(P1_EBX_REG_19__SCAN_IN), .A(n14865), .ZN(
        n14866) );
  OAI211_X1 U18216 ( .C1(n14895), .C2(n14868), .A(n14867), .B(n14866), .ZN(
        n14869) );
  AOI21_X1 U18217 ( .B1(n15426), .B2(n20532), .A(n14869), .ZN(n14870) );
  OAI21_X1 U18218 ( .B1(n15121), .B2(n17350), .A(n14870), .ZN(P1_U2821) );
  OAI21_X1 U18219 ( .B1(n14871), .B2(n14873), .A(n14872), .ZN(n15245) );
  AOI21_X1 U18220 ( .B1(n14875), .B2(n14890), .A(n14853), .ZN(n15429) );
  INV_X1 U18221 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n14881) );
  NAND2_X1 U18222 ( .A1(n14876), .A2(n14881), .ZN(n14880) );
  AOI21_X1 U18223 ( .B1(n20579), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20683), .ZN(n14877) );
  OAI21_X1 U18224 ( .B1(n20560), .B2(n15239), .A(n14877), .ZN(n14878) );
  AOI21_X1 U18225 ( .B1(n20574), .B2(P1_EBX_REG_18__SCAN_IN), .A(n14878), .ZN(
        n14879) );
  OAI211_X1 U18226 ( .C1(n14895), .C2(n14881), .A(n14880), .B(n14879), .ZN(
        n14882) );
  AOI21_X1 U18227 ( .B1(n15429), .B2(n20532), .A(n14882), .ZN(n14883) );
  OAI21_X1 U18228 ( .B1(n15245), .B2(n17350), .A(n14883), .ZN(P1_U2822) );
  INV_X1 U18229 ( .A(n14871), .ZN(n14885) );
  OAI21_X1 U18230 ( .B1(n14884), .B2(n14886), .A(n14885), .ZN(n15252) );
  OR2_X1 U18231 ( .A1(n14887), .A2(n14888), .ZN(n14889) );
  AND2_X1 U18232 ( .A1(n14890), .A2(n14889), .ZN(n15445) );
  INV_X1 U18233 ( .A(n14908), .ZN(n14891) );
  AOI21_X1 U18234 ( .B1(n14891), .B2(P1_REIP_REG_16__SCAN_IN), .A(
        P1_REIP_REG_17__SCAN_IN), .ZN(n14896) );
  NAND2_X1 U18235 ( .A1(n20575), .A2(n15255), .ZN(n14892) );
  OAI211_X1 U18236 ( .C1(n20565), .C2(n15251), .A(n14892), .B(n20667), .ZN(
        n14893) );
  AOI21_X1 U18237 ( .B1(n20541), .B2(P1_EBX_REG_17__SCAN_IN), .A(n14893), .ZN(
        n14894) );
  OAI21_X1 U18238 ( .B1(n14896), .B2(n14895), .A(n14894), .ZN(n14897) );
  AOI21_X1 U18239 ( .B1(n20532), .B2(n15445), .A(n14897), .ZN(n14898) );
  OAI21_X1 U18240 ( .B1(n15252), .B2(n17350), .A(n14898), .ZN(P1_U2823) );
  AOI21_X1 U18241 ( .B1(n14900), .B2(n14915), .A(n14884), .ZN(n15269) );
  INV_X1 U18242 ( .A(n15269), .ZN(n15139) );
  NOR2_X1 U18243 ( .A1(n9742), .A2(n14901), .ZN(n14902) );
  OR2_X1 U18244 ( .A1(n14887), .A2(n14902), .ZN(n15040) );
  INV_X1 U18245 ( .A(n15040), .ZN(n15455) );
  INV_X1 U18246 ( .A(n14903), .ZN(n14931) );
  NOR3_X1 U18247 ( .A1(n14931), .A2(P1_REIP_REG_15__SCAN_IN), .A3(n21330), 
        .ZN(n14921) );
  OAI21_X1 U18248 ( .B1(n14921), .B2(n14929), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n14907) );
  NAND2_X1 U18249 ( .A1(n20575), .A2(n15265), .ZN(n14904) );
  OAI211_X1 U18250 ( .C1(n20565), .C2(n15267), .A(n14904), .B(n20667), .ZN(
        n14905) );
  AOI21_X1 U18251 ( .B1(n20541), .B2(P1_EBX_REG_16__SCAN_IN), .A(n14905), .ZN(
        n14906) );
  OAI211_X1 U18252 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(n14908), .A(n14907), 
        .B(n14906), .ZN(n14909) );
  AOI21_X1 U18253 ( .B1(n20532), .B2(n15455), .A(n14909), .ZN(n14910) );
  OAI21_X1 U18254 ( .B1(n15139), .B2(n17350), .A(n14910), .ZN(P1_U2824) );
  INV_X1 U18255 ( .A(n14941), .ZN(n14912) );
  INV_X1 U18256 ( .A(n14977), .ZN(n14943) );
  OR2_X1 U18257 ( .A1(n14911), .A2(n14943), .ZN(n14914) );
  AND2_X1 U18258 ( .A1(n14945), .A2(n14928), .ZN(n14926) );
  OAI21_X1 U18259 ( .B1(n14926), .B2(n14916), .A(n14915), .ZN(n15279) );
  NAND2_X1 U18260 ( .A1(n20541), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n14920) );
  INV_X1 U18261 ( .A(n15272), .ZN(n14917) );
  NAND2_X1 U18262 ( .A1(n20575), .A2(n14917), .ZN(n14919) );
  NAND2_X1 U18263 ( .A1(n20579), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14918) );
  NAND4_X1 U18264 ( .A1(n14920), .A2(n20667), .A3(n14919), .A4(n14918), .ZN(
        n14922) );
  AOI211_X1 U18265 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n14929), .A(n14922), 
        .B(n14921), .ZN(n14925) );
  AOI21_X1 U18266 ( .B1(n14923), .B2(n14933), .A(n9742), .ZN(n15458) );
  NAND2_X1 U18267 ( .A1(n15458), .A2(n20532), .ZN(n14924) );
  OAI211_X1 U18268 ( .C1(n15279), .C2(n17350), .A(n14925), .B(n14924), .ZN(
        P1_U2825) );
  INV_X1 U18269 ( .A(n14926), .ZN(n14927) );
  INV_X1 U18270 ( .A(n15280), .ZN(n14939) );
  INV_X1 U18271 ( .A(n14929), .ZN(n14930) );
  AOI21_X1 U18272 ( .B1(n14931), .B2(n21330), .A(n14930), .ZN(n14938) );
  INV_X1 U18273 ( .A(n14933), .ZN(n14934) );
  AOI21_X1 U18274 ( .B1(n14935), .B2(n14932), .A(n14934), .ZN(n15472) );
  AOI22_X1 U18275 ( .A1(P1_EBX_REG_14__SCAN_IN), .A2(n20574), .B1(n20532), 
        .B2(n15472), .ZN(n14936) );
  OAI211_X1 U18276 ( .C1(n20565), .C2(n11712), .A(n14936), .B(n20667), .ZN(
        n14937) );
  AOI211_X1 U18277 ( .C1(n20575), .C2(n14939), .A(n14938), .B(n14937), .ZN(
        n14940) );
  OAI21_X1 U18278 ( .B1(n15290), .B2(n17350), .A(n14940), .ZN(P1_U2826) );
  INV_X1 U18279 ( .A(n14911), .ZN(n15049) );
  OAI21_X1 U18280 ( .B1(n15049), .B2(n14941), .A(n14942), .ZN(n14978) );
  OAI21_X1 U18281 ( .B1(n14978), .B2(n14943), .A(n14942), .ZN(n14963) );
  NAND2_X1 U18282 ( .A1(n14963), .A2(n14962), .ZN(n14961) );
  INV_X1 U18283 ( .A(n14944), .ZN(n14946) );
  AOI21_X1 U18284 ( .B1(n14961), .B2(n14946), .A(n14945), .ZN(n15302) );
  INV_X1 U18285 ( .A(n15302), .ZN(n15145) );
  NOR2_X1 U18286 ( .A1(n21328), .A2(n14988), .ZN(n14951) );
  NAND2_X1 U18287 ( .A1(n20517), .A2(n14947), .ZN(n14948) );
  NAND2_X1 U18288 ( .A1(n20517), .A2(n14980), .ZN(n14949) );
  OAI21_X1 U18289 ( .B1(n14951), .B2(n14950), .A(n17357), .ZN(n14973) );
  OAI21_X1 U18290 ( .B1(n14968), .B2(n14952), .A(n14932), .ZN(n15477) );
  AOI21_X1 U18291 ( .B1(n20579), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n20683), .ZN(n14953) );
  OAI21_X1 U18292 ( .B1(n20560), .B2(n15300), .A(n14953), .ZN(n14954) );
  AOI21_X1 U18293 ( .B1(n20574), .B2(P1_EBX_REG_13__SCAN_IN), .A(n14954), .ZN(
        n14958) );
  INV_X1 U18294 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n14955) );
  NAND3_X1 U18295 ( .A1(n20505), .A2(n14956), .A3(n14955), .ZN(n14957) );
  OAI211_X1 U18296 ( .C1(n15477), .C2(n20589), .A(n14958), .B(n14957), .ZN(
        n14959) );
  AOI21_X1 U18297 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n14973), .A(n14959), 
        .ZN(n14960) );
  OAI21_X1 U18298 ( .B1(n15145), .B2(n17350), .A(n14960), .ZN(P1_U2827) );
  OAI21_X1 U18299 ( .B1(n14963), .B2(n14962), .A(n14961), .ZN(n15311) );
  AOI21_X1 U18300 ( .B1(n20579), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n20683), .ZN(n14964) );
  OAI21_X1 U18301 ( .B1(n20560), .B2(n15304), .A(n14964), .ZN(n14971) );
  INV_X1 U18302 ( .A(n14965), .ZN(n14967) );
  AOI21_X1 U18303 ( .B1(n14967), .B2(n14979), .A(n14966), .ZN(n14969) );
  OR2_X1 U18304 ( .A1(n14969), .A2(n14968), .ZN(n15494) );
  NOR2_X1 U18305 ( .A1(n15494), .A2(n20589), .ZN(n14970) );
  AOI211_X1 U18306 ( .C1(P1_EBX_REG_12__SCAN_IN), .C2(n20541), .A(n14971), .B(
        n14970), .ZN(n14976) );
  NOR3_X1 U18307 ( .A1(n14972), .A2(n14988), .A3(n14980), .ZN(n14974) );
  OAI21_X1 U18308 ( .B1(n14974), .B2(P1_REIP_REG_12__SCAN_IN), .A(n14973), 
        .ZN(n14975) );
  OAI211_X1 U18309 ( .C1(n15311), .C2(n17350), .A(n14976), .B(n14975), .ZN(
        P1_U2828) );
  XNOR2_X1 U18310 ( .A(n14978), .B(n14977), .ZN(n15320) );
  XNOR2_X1 U18311 ( .A(n14965), .B(n14979), .ZN(n15505) );
  NOR2_X1 U18312 ( .A1(n14980), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n14986) );
  NAND2_X1 U18313 ( .A1(n20541), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n14984) );
  INV_X1 U18314 ( .A(n15318), .ZN(n14981) );
  NAND2_X1 U18315 ( .A1(n20575), .A2(n14981), .ZN(n14983) );
  NAND2_X1 U18316 ( .A1(n20579), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14982) );
  NAND4_X1 U18317 ( .A1(n14984), .A2(n20667), .A3(n14983), .A4(n14982), .ZN(
        n14985) );
  AOI21_X1 U18318 ( .B1(n20505), .B2(n14986), .A(n14985), .ZN(n14987) );
  OAI21_X1 U18319 ( .B1(n17357), .B2(n14988), .A(n14987), .ZN(n14989) );
  AOI21_X1 U18320 ( .B1(n20532), .B2(n15505), .A(n14989), .ZN(n14990) );
  OAI21_X1 U18321 ( .B1(n15148), .B2(n17350), .A(n14990), .ZN(P1_U2829) );
  OAI21_X1 U18322 ( .B1(n10434), .B2(n9756), .A(n14991), .ZN(n15350) );
  INV_X1 U18323 ( .A(n20511), .ZN(n15000) );
  OAI21_X1 U18324 ( .B1(n14245), .B2(n14993), .A(n15059), .ZN(n14994) );
  INV_X1 U18325 ( .A(n14994), .ZN(n17382) );
  AOI22_X1 U18326 ( .A1(n15346), .A2(n20575), .B1(n20532), .B2(n17382), .ZN(
        n14995) );
  OAI211_X1 U18327 ( .C1(n20565), .C2(n15343), .A(n14995), .B(n20667), .ZN(
        n14999) );
  NAND4_X1 U18328 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .A4(n20540), .ZN(n14997) );
  OAI22_X1 U18329 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14997), .B1(n14996), 
        .B2(n20553), .ZN(n14998) );
  AOI211_X1 U18330 ( .C1(P1_REIP_REG_8__SCAN_IN), .C2(n15000), .A(n14999), .B(
        n14998), .ZN(n15001) );
  OAI21_X1 U18331 ( .B1(n15350), .B2(n17350), .A(n15001), .ZN(P1_U2832) );
  OR2_X1 U18332 ( .A1(n21382), .A2(n15002), .ZN(n15003) );
  NAND2_X1 U18333 ( .A1(n17350), .A2(n15003), .ZN(n20585) );
  INV_X1 U18334 ( .A(n20585), .ZN(n15021) );
  OR2_X1 U18335 ( .A1(n21382), .A2(n15004), .ZN(n20578) );
  INV_X1 U18336 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n15005) );
  OAI22_X1 U18337 ( .A1(n20578), .A2(n21188), .B1(n20562), .B2(n15005), .ZN(
        n15007) );
  NAND2_X1 U18338 ( .A1(n20555), .A2(n15005), .ZN(n20563) );
  OAI21_X1 U18339 ( .B1(n20589), .B2(n20692), .A(n20563), .ZN(n15006) );
  AOI211_X1 U18340 ( .C1(n20574), .C2(P1_EBX_REG_1__SCAN_IN), .A(n15007), .B(
        n15006), .ZN(n15010) );
  MUX2_X1 U18341 ( .A(n20565), .B(n20560), .S(n15008), .Z(n15009) );
  OAI211_X1 U18342 ( .C1(n15011), .C2(n15021), .A(n15010), .B(n15009), .ZN(
        P1_U2839) );
  INV_X1 U18343 ( .A(n15012), .ZN(n15013) );
  AND2_X1 U18344 ( .A1(n20532), .A2(n15013), .ZN(n15018) );
  INV_X1 U18345 ( .A(n11586), .ZN(n15016) );
  NAND2_X1 U18346 ( .A1(n20541), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n15015) );
  OAI21_X1 U18347 ( .B1(n20575), .B2(n20579), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15014) );
  OAI211_X1 U18348 ( .C1(n20578), .C2(n15016), .A(n15015), .B(n15014), .ZN(
        n15017) );
  AOI211_X1 U18349 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(n20517), .A(n15018), .B(
        n15017), .ZN(n15019) );
  OAI21_X1 U18350 ( .B1(n15021), .B2(n15020), .A(n15019), .ZN(P1_U2840) );
  INV_X1 U18351 ( .A(n15022), .ZN(n15024) );
  INV_X1 U18352 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15023) );
  OAI22_X1 U18353 ( .A1(n15024), .A2(n20594), .B1(n20599), .B2(n15023), .ZN(
        P1_U2841) );
  OAI222_X1 U18354 ( .A1(n15165), .A2(n15055), .B1(n15025), .B2(n20599), .C1(
        n15359), .C2(n20594), .ZN(P1_U2843) );
  AOI22_X1 U18355 ( .A1(n15360), .A2(n20590), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n15062), .ZN(n15026) );
  OAI21_X1 U18356 ( .B1(n15181), .B2(n15055), .A(n15026), .ZN(P1_U2845) );
  INV_X1 U18357 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15028) );
  OAI222_X1 U18358 ( .A1(n15090), .A2(n15055), .B1(n15028), .B2(n20599), .C1(
        n15027), .C2(n20594), .ZN(P1_U2846) );
  OAI222_X1 U18359 ( .A1(n15055), .A2(n15199), .B1(n21524), .B2(n20599), .C1(
        n15029), .C2(n20594), .ZN(P1_U2847) );
  AOI22_X1 U18360 ( .A1(n15388), .A2(n20590), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n15062), .ZN(n15030) );
  OAI21_X1 U18361 ( .B1(n15098), .B2(n15055), .A(n15030), .ZN(P1_U2848) );
  AOI22_X1 U18362 ( .A1(n15397), .A2(n20590), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n15062), .ZN(n15031) );
  OAI21_X1 U18363 ( .B1(n15103), .B2(n15055), .A(n15031), .ZN(P1_U2849) );
  AOI22_X1 U18364 ( .A1(n15400), .A2(n20590), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n15062), .ZN(n15032) );
  OAI21_X1 U18365 ( .B1(n15223), .B2(n15055), .A(n15032), .ZN(P1_U2850) );
  OAI222_X1 U18366 ( .A1(n15055), .A2(n15112), .B1(n15034), .B2(n20599), .C1(
        n15033), .C2(n20594), .ZN(P1_U2851) );
  OAI222_X1 U18367 ( .A1(n15225), .A2(n15055), .B1(n15036), .B2(n20599), .C1(
        n15035), .C2(n20594), .ZN(P1_U2852) );
  AOI22_X1 U18368 ( .A1(n15426), .A2(n20590), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n15062), .ZN(n15037) );
  OAI21_X1 U18369 ( .B1(n15121), .B2(n15055), .A(n15037), .ZN(P1_U2853) );
  AOI22_X1 U18370 ( .A1(n15429), .A2(n20590), .B1(P1_EBX_REG_18__SCAN_IN), 
        .B2(n15062), .ZN(n15038) );
  OAI21_X1 U18371 ( .B1(n15245), .B2(n15055), .A(n15038), .ZN(P1_U2854) );
  AOI22_X1 U18372 ( .A1(n15445), .A2(n20590), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n15062), .ZN(n15039) );
  OAI21_X1 U18373 ( .B1(n15252), .B2(n15055), .A(n15039), .ZN(P1_U2855) );
  OAI222_X1 U18374 ( .A1(n15139), .A2(n15055), .B1(n15041), .B2(n20599), .C1(
        n15040), .C2(n20594), .ZN(P1_U2856) );
  AOI22_X1 U18375 ( .A1(n15458), .A2(n20590), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n15062), .ZN(n15042) );
  OAI21_X1 U18376 ( .B1(n15279), .B2(n15055), .A(n15042), .ZN(P1_U2857) );
  AOI22_X1 U18377 ( .A1(n15472), .A2(n20590), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n15062), .ZN(n15043) );
  OAI21_X1 U18378 ( .B1(n15290), .B2(n15055), .A(n15043), .ZN(P1_U2858) );
  INV_X1 U18379 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15044) );
  OAI222_X1 U18380 ( .A1(n15145), .A2(n15055), .B1(n15044), .B2(n20599), .C1(
        n15477), .C2(n20594), .ZN(P1_U2859) );
  OAI222_X1 U18381 ( .A1(n15311), .A2(n15055), .B1(n15045), .B2(n20599), .C1(
        n15494), .C2(n20594), .ZN(P1_U2860) );
  AOI22_X1 U18382 ( .A1(n15505), .A2(n20590), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n15062), .ZN(n15046) );
  OAI21_X1 U18383 ( .B1(n15148), .B2(n15055), .A(n15046), .ZN(P1_U2861) );
  INV_X1 U18384 ( .A(n15048), .ZN(n15050) );
  AOI21_X1 U18385 ( .B1(n10433), .B2(n15050), .A(n15049), .ZN(n15328) );
  INV_X1 U18386 ( .A(n15328), .ZN(n17351) );
  NAND2_X1 U18387 ( .A1(n15051), .A2(n15052), .ZN(n15053) );
  AND2_X1 U18388 ( .A1(n14965), .A2(n15053), .ZN(n17346) );
  AOI22_X1 U18389 ( .A1(n17346), .A2(n20590), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n15062), .ZN(n15054) );
  OAI21_X1 U18390 ( .B1(n17351), .B2(n15055), .A(n15054), .ZN(P1_U2862) );
  AND2_X1 U18391 ( .A1(n14991), .A2(n15056), .ZN(n15057) );
  NOR2_X1 U18392 ( .A1(n15048), .A2(n15057), .ZN(n20513) );
  INV_X1 U18393 ( .A(n20513), .ZN(n15151) );
  INV_X1 U18394 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n15061) );
  NAND2_X1 U18395 ( .A1(n15059), .A2(n15058), .ZN(n15060) );
  NAND2_X1 U18396 ( .A1(n15051), .A2(n15060), .ZN(n20507) );
  OAI222_X1 U18397 ( .A1(n15151), .A2(n15055), .B1(n15061), .B2(n20599), .C1(
        n20594), .C2(n20507), .ZN(P1_U2863) );
  AOI22_X1 U18398 ( .A1(n17382), .A2(n20590), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n15062), .ZN(n15063) );
  OAI21_X1 U18399 ( .B1(n15350), .B2(n15055), .A(n15063), .ZN(P1_U2864) );
  NAND2_X1 U18400 ( .A1(n14144), .A2(n15064), .ZN(n15065) );
  NAND2_X1 U18401 ( .A1(n10450), .A2(n15065), .ZN(n17373) );
  INV_X1 U18402 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n15066) );
  OAI222_X1 U18403 ( .A1(n17373), .A2(n15055), .B1(n15066), .B2(n20599), .C1(
        n20594), .C2(n20542), .ZN(P1_U2867) );
  OAI22_X1 U18404 ( .A1(n15127), .A2(n15141), .B1(n15157), .B2(n15067), .ZN(
        n15068) );
  AOI21_X1 U18405 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n15129), .A(n15068), .ZN(
        n15070) );
  NAND2_X1 U18406 ( .A1(n15137), .A2(DATAI_30_), .ZN(n15069) );
  OAI211_X1 U18407 ( .C1(n15071), .C2(n15158), .A(n15070), .B(n15069), .ZN(
        P1_U2874) );
  INV_X1 U18408 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16049) );
  INV_X1 U18409 ( .A(n15127), .ZN(n15133) );
  INV_X1 U18410 ( .A(DATAI_13_), .ZN(n15073) );
  NAND2_X1 U18411 ( .A1(n20709), .A2(BUF1_REG_13__SCAN_IN), .ZN(n15072) );
  OAI21_X1 U18412 ( .B1(n20709), .B2(n15073), .A(n15072), .ZN(n20631) );
  AOI22_X1 U18413 ( .A1(n15133), .A2(n20631), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n15142), .ZN(n15074) );
  OAI21_X1 U18414 ( .B1(n16049), .B2(n15135), .A(n15074), .ZN(n15075) );
  AOI21_X1 U18415 ( .B1(n15137), .B2(DATAI_29_), .A(n15075), .ZN(n15076) );
  OAI21_X1 U18416 ( .B1(n15165), .B2(n15158), .A(n15076), .ZN(P1_U2875) );
  OAI22_X1 U18417 ( .A1(n15127), .A2(n15146), .B1(n15157), .B2(n15077), .ZN(
        n15078) );
  AOI21_X1 U18418 ( .B1(n15129), .B2(BUF1_REG_28__SCAN_IN), .A(n15078), .ZN(
        n15080) );
  NAND2_X1 U18419 ( .A1(n15137), .A2(DATAI_28_), .ZN(n15079) );
  OAI211_X1 U18420 ( .C1(n15081), .C2(n15158), .A(n15080), .B(n15079), .ZN(
        P1_U2876) );
  OAI22_X1 U18421 ( .A1(n15127), .A2(n15147), .B1(n15157), .B2(n15082), .ZN(
        n15083) );
  AOI21_X1 U18422 ( .B1(n15129), .B2(BUF1_REG_27__SCAN_IN), .A(n15083), .ZN(
        n15085) );
  NAND2_X1 U18423 ( .A1(n15137), .A2(DATAI_27_), .ZN(n15084) );
  OAI211_X1 U18424 ( .C1(n15181), .C2(n15158), .A(n15085), .B(n15084), .ZN(
        P1_U2877) );
  OAI22_X1 U18425 ( .A1(n15127), .A2(n15149), .B1(n15157), .B2(n15086), .ZN(
        n15088) );
  INV_X1 U18426 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n17440) );
  NOR2_X1 U18427 ( .A1(n15135), .A2(n17440), .ZN(n15087) );
  AOI211_X1 U18428 ( .C1(DATAI_26_), .C2(n15137), .A(n15088), .B(n15087), .ZN(
        n15089) );
  OAI21_X1 U18429 ( .B1(n15090), .B2(n15158), .A(n15089), .ZN(P1_U2878) );
  OAI22_X1 U18430 ( .A1(n15127), .A2(n15150), .B1(n15157), .B2(n15091), .ZN(
        n15092) );
  AOI21_X1 U18431 ( .B1(n15129), .B2(BUF1_REG_25__SCAN_IN), .A(n15092), .ZN(
        n15094) );
  NAND2_X1 U18432 ( .A1(n15137), .A2(DATAI_25_), .ZN(n15093) );
  OAI211_X1 U18433 ( .C1(n15199), .C2(n15158), .A(n15094), .B(n15093), .ZN(
        P1_U2879) );
  AOI22_X1 U18434 ( .A1(n15133), .A2(n15152), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n15142), .ZN(n15095) );
  OAI21_X1 U18435 ( .B1(n15135), .B2(n17443), .A(n15095), .ZN(n15096) );
  AOI21_X1 U18436 ( .B1(n15137), .B2(DATAI_24_), .A(n15096), .ZN(n15097) );
  OAI21_X1 U18437 ( .B1(n15098), .B2(n15158), .A(n15097), .ZN(P1_U2880) );
  OAI22_X1 U18438 ( .A1(n15127), .A2(n20767), .B1(n15157), .B2(n15099), .ZN(
        n15100) );
  AOI21_X1 U18439 ( .B1(n15129), .B2(BUF1_REG_23__SCAN_IN), .A(n15100), .ZN(
        n15102) );
  NAND2_X1 U18440 ( .A1(n15137), .A2(DATAI_23_), .ZN(n15101) );
  OAI211_X1 U18441 ( .C1(n15103), .C2(n15158), .A(n15102), .B(n15101), .ZN(
        P1_U2881) );
  OAI22_X1 U18442 ( .A1(n15127), .A2(n20759), .B1(n15157), .B2(n15104), .ZN(
        n15105) );
  AOI21_X1 U18443 ( .B1(n15129), .B2(BUF1_REG_22__SCAN_IN), .A(n15105), .ZN(
        n15107) );
  NAND2_X1 U18444 ( .A1(n15137), .A2(DATAI_22_), .ZN(n15106) );
  OAI211_X1 U18445 ( .C1(n15223), .C2(n15158), .A(n15107), .B(n15106), .ZN(
        P1_U2882) );
  OAI22_X1 U18446 ( .A1(n15127), .A2(n20754), .B1(n15157), .B2(n15108), .ZN(
        n15109) );
  AOI21_X1 U18447 ( .B1(n15129), .B2(BUF1_REG_21__SCAN_IN), .A(n15109), .ZN(
        n15111) );
  NAND2_X1 U18448 ( .A1(n15137), .A2(DATAI_21_), .ZN(n15110) );
  OAI211_X1 U18449 ( .C1(n15112), .C2(n15158), .A(n15111), .B(n15110), .ZN(
        P1_U2883) );
  INV_X1 U18450 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16110) );
  AOI22_X1 U18451 ( .A1(n15133), .A2(n15113), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n15142), .ZN(n15114) );
  OAI21_X1 U18452 ( .B1(n15135), .B2(n16110), .A(n15114), .ZN(n15115) );
  AOI21_X1 U18453 ( .B1(n15137), .B2(DATAI_20_), .A(n15115), .ZN(n15116) );
  OAI21_X1 U18454 ( .B1(n15225), .B2(n15158), .A(n15116), .ZN(P1_U2884) );
  OAI22_X1 U18455 ( .A1(n15127), .A2(n20744), .B1(n15157), .B2(n15117), .ZN(
        n15118) );
  AOI21_X1 U18456 ( .B1(n15129), .B2(BUF1_REG_19__SCAN_IN), .A(n15118), .ZN(
        n15120) );
  NAND2_X1 U18457 ( .A1(n15137), .A2(DATAI_19_), .ZN(n15119) );
  OAI211_X1 U18458 ( .C1(n15121), .C2(n15158), .A(n15120), .B(n15119), .ZN(
        P1_U2885) );
  INV_X1 U18459 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n17450) );
  AOI22_X1 U18460 ( .A1(n15133), .A2(n15122), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n15142), .ZN(n15123) );
  OAI21_X1 U18461 ( .B1(n15135), .B2(n17450), .A(n15123), .ZN(n15124) );
  AOI21_X1 U18462 ( .B1(n15137), .B2(DATAI_18_), .A(n15124), .ZN(n15125) );
  OAI21_X1 U18463 ( .B1(n15245), .B2(n15158), .A(n15125), .ZN(P1_U2886) );
  OAI22_X1 U18464 ( .A1(n15127), .A2(n20735), .B1(n15157), .B2(n15126), .ZN(
        n15128) );
  AOI21_X1 U18465 ( .B1(n15129), .B2(BUF1_REG_17__SCAN_IN), .A(n15128), .ZN(
        n15131) );
  NAND2_X1 U18466 ( .A1(n15137), .A2(DATAI_17_), .ZN(n15130) );
  OAI211_X1 U18467 ( .C1(n15252), .C2(n15158), .A(n15131), .B(n15130), .ZN(
        P1_U2887) );
  INV_X1 U18468 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16141) );
  AOI22_X1 U18469 ( .A1(n15133), .A2(n15132), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n15142), .ZN(n15134) );
  OAI21_X1 U18470 ( .B1(n15135), .B2(n16141), .A(n15134), .ZN(n15136) );
  AOI21_X1 U18471 ( .B1(n15137), .B2(DATAI_16_), .A(n15136), .ZN(n15138) );
  OAI21_X1 U18472 ( .B1(n15139), .B2(n15158), .A(n15138), .ZN(P1_U2888) );
  OAI222_X1 U18473 ( .A1(n15158), .A2(n15279), .B1(n15156), .B2(n15140), .C1(
        n20602), .C2(n15157), .ZN(P1_U2889) );
  INV_X1 U18474 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20604) );
  OAI222_X1 U18475 ( .A1(n15158), .A2(n15290), .B1(n15157), .B2(n20604), .C1(
        n15156), .C2(n15141), .ZN(P1_U2890) );
  AOI22_X1 U18476 ( .A1(n15143), .A2(n20631), .B1(n15142), .B2(
        P1_EAX_REG_13__SCAN_IN), .ZN(n15144) );
  OAI21_X1 U18477 ( .B1(n15145), .B2(n15158), .A(n15144), .ZN(P1_U2891) );
  INV_X1 U18478 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20607) );
  OAI222_X1 U18479 ( .A1(n15311), .A2(n15158), .B1(n20607), .B2(n15157), .C1(
        n15156), .C2(n15146), .ZN(P1_U2892) );
  OAI222_X1 U18480 ( .A1(n15158), .A2(n15148), .B1(n15157), .B2(n11687), .C1(
        n15156), .C2(n15147), .ZN(P1_U2893) );
  INV_X1 U18481 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20610) );
  OAI222_X1 U18482 ( .A1(n15158), .A2(n17351), .B1(n15157), .B2(n20610), .C1(
        n15156), .C2(n15149), .ZN(P1_U2894) );
  OAI222_X1 U18483 ( .A1(n15158), .A2(n15151), .B1(n15157), .B2(n11653), .C1(
        n15156), .C2(n15150), .ZN(P1_U2895) );
  INV_X1 U18484 ( .A(n15152), .ZN(n15153) );
  OAI222_X1 U18485 ( .A1(n15158), .A2(n15350), .B1(n15157), .B2(n11637), .C1(
        n15156), .C2(n15153), .ZN(P1_U2896) );
  XOR2_X1 U18486 ( .A(n15154), .B(n10450), .Z(n20591) );
  INV_X1 U18487 ( .A(n20591), .ZN(n15155) );
  OAI222_X1 U18488 ( .A1(n15156), .A2(n20759), .B1(n15158), .B2(n15155), .C1(
        n11568), .C2(n15157), .ZN(P1_U2898) );
  OAI222_X1 U18489 ( .A1(n15158), .A2(n17373), .B1(n15157), .B2(n11552), .C1(
        n15156), .C2(n20754), .ZN(P1_U2899) );
  NOR2_X1 U18490 ( .A1(n20667), .A2(n21354), .ZN(n15354) );
  NOR2_X1 U18491 ( .A1(n20654), .A2(n15159), .ZN(n15160) );
  AOI211_X1 U18492 ( .C1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n20641), .A(
        n15354), .B(n15160), .ZN(n15164) );
  XNOR2_X1 U18493 ( .A(n15332), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15161) );
  NAND2_X1 U18494 ( .A1(n15351), .A2(n20650), .ZN(n15163) );
  OAI211_X1 U18495 ( .C1(n15165), .C2(n20712), .A(n15164), .B(n15163), .ZN(
        P1_U2970) );
  NAND2_X1 U18496 ( .A1(n15347), .A2(n15166), .ZN(n15168) );
  OAI211_X1 U18497 ( .C1(n15169), .C2(n15344), .A(n15168), .B(n15167), .ZN(
        n15170) );
  AOI21_X1 U18498 ( .B1(n15171), .B2(n20649), .A(n15170), .ZN(n15172) );
  OAI21_X1 U18499 ( .B1(n15339), .B2(n15173), .A(n15172), .ZN(P1_U2971) );
  AND2_X1 U18500 ( .A1(n20683), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n15364) );
  NOR2_X1 U18501 ( .A1(n20654), .A2(n15174), .ZN(n15175) );
  AOI211_X1 U18502 ( .C1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n20641), .A(
        n15364), .B(n15175), .ZN(n15180) );
  NAND2_X1 U18503 ( .A1(n15177), .A2(n15176), .ZN(n15178) );
  OAI211_X1 U18504 ( .C1(n15181), .C2(n20712), .A(n15180), .B(n15179), .ZN(
        P1_U2972) );
  OAI21_X1 U18505 ( .B1(n15210), .B2(n15182), .A(n15324), .ZN(n15184) );
  OAI211_X1 U18506 ( .C1(n15185), .C2(n15210), .A(n15184), .B(n15183), .ZN(
        n15186) );
  XNOR2_X1 U18507 ( .A(n15186), .B(n15371), .ZN(n15379) );
  NAND2_X1 U18508 ( .A1(n15347), .A2(n15187), .ZN(n15188) );
  NAND2_X1 U18509 ( .A1(n20683), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15374) );
  OAI211_X1 U18510 ( .C1(n15189), .C2(n15344), .A(n15188), .B(n15374), .ZN(
        n15190) );
  AOI21_X1 U18511 ( .B1(n15191), .B2(n20649), .A(n15190), .ZN(n15192) );
  OAI21_X1 U18512 ( .B1(n15339), .B2(n15379), .A(n15192), .ZN(P1_U2973) );
  NOR2_X1 U18513 ( .A1(n20654), .A2(n15193), .ZN(n15194) );
  AOI211_X1 U18514 ( .C1(n20641), .C2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15195), .B(n15194), .ZN(n15198) );
  NAND2_X1 U18515 ( .A1(n15196), .A2(n20650), .ZN(n15197) );
  OAI211_X1 U18516 ( .C1(n15199), .C2(n20712), .A(n15198), .B(n15197), .ZN(
        P1_U2974) );
  NOR2_X1 U18517 ( .A1(n15210), .A2(n10416), .ZN(n15201) );
  MUX2_X1 U18518 ( .A(n15332), .B(n15201), .S(n15200), .Z(n15202) );
  XNOR2_X1 U18519 ( .A(n15202), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15390) );
  INV_X1 U18520 ( .A(n15203), .ZN(n15205) );
  NAND2_X1 U18521 ( .A1(n20683), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15384) );
  NAND2_X1 U18522 ( .A1(n20641), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15204) );
  OAI211_X1 U18523 ( .C1(n20654), .C2(n15205), .A(n15384), .B(n15204), .ZN(
        n15206) );
  AOI21_X1 U18524 ( .B1(n15207), .B2(n20649), .A(n15206), .ZN(n15208) );
  OAI21_X1 U18525 ( .B1(n15390), .B2(n15339), .A(n15208), .ZN(P1_U2975) );
  XNOR2_X1 U18526 ( .A(n15332), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15209) );
  XNOR2_X1 U18527 ( .A(n15210), .B(n15209), .ZN(n15399) );
  NAND2_X1 U18528 ( .A1(n20683), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15392) );
  NAND2_X1 U18529 ( .A1(n20641), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15211) );
  OAI211_X1 U18530 ( .C1(n20654), .C2(n15212), .A(n15392), .B(n15211), .ZN(
        n15213) );
  AOI21_X1 U18531 ( .B1(n15214), .B2(n20649), .A(n15213), .ZN(n15215) );
  OAI21_X1 U18532 ( .B1(n15399), .B2(n15339), .A(n15215), .ZN(P1_U2976) );
  AND2_X1 U18533 ( .A1(n20683), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15404) );
  NOR2_X1 U18534 ( .A1(n20654), .A2(n15216), .ZN(n15217) );
  AOI211_X1 U18535 ( .C1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n20641), .A(
        n15404), .B(n15217), .ZN(n15222) );
  NAND2_X1 U18536 ( .A1(n15219), .A2(n15218), .ZN(n15220) );
  XNOR2_X1 U18537 ( .A(n15220), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15401) );
  NAND2_X1 U18538 ( .A1(n15401), .A2(n20650), .ZN(n15221) );
  OAI211_X1 U18539 ( .C1(n15223), .C2(n20712), .A(n15222), .B(n15221), .ZN(
        P1_U2977) );
  XNOR2_X1 U18540 ( .A(n15224), .B(n15415), .ZN(n15419) );
  INV_X1 U18541 ( .A(n15225), .ZN(n15229) );
  NAND2_X1 U18542 ( .A1(n20683), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15413) );
  NAND2_X1 U18543 ( .A1(n20641), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15226) );
  OAI211_X1 U18544 ( .C1(n20654), .C2(n15227), .A(n15413), .B(n15226), .ZN(
        n15228) );
  AOI21_X1 U18545 ( .B1(n15229), .B2(n20649), .A(n15228), .ZN(n15230) );
  OAI21_X1 U18546 ( .B1(n15419), .B2(n15339), .A(n15230), .ZN(P1_U2979) );
  XNOR2_X1 U18547 ( .A(n15332), .B(n15423), .ZN(n15231) );
  XNOR2_X1 U18548 ( .A(n15232), .B(n15231), .ZN(n15428) );
  NAND2_X1 U18549 ( .A1(n15347), .A2(n15233), .ZN(n15234) );
  NAND2_X1 U18550 ( .A1(n20683), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15421) );
  OAI211_X1 U18551 ( .C1(n15344), .C2(n15235), .A(n15234), .B(n15421), .ZN(
        n15236) );
  AOI21_X1 U18552 ( .B1(n15237), .B2(n20649), .A(n15236), .ZN(n15238) );
  OAI21_X1 U18553 ( .B1(n15428), .B2(n15339), .A(n15238), .ZN(P1_U2980) );
  AND2_X1 U18554 ( .A1(n20683), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15435) );
  NOR2_X1 U18555 ( .A1(n20654), .A2(n15239), .ZN(n15240) );
  AOI211_X1 U18556 ( .C1(n20641), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15435), .B(n15240), .ZN(n15244) );
  OR2_X1 U18557 ( .A1(n15242), .A2(n15241), .ZN(n15431) );
  NAND3_X1 U18558 ( .A1(n15431), .A2(n15430), .A3(n20650), .ZN(n15243) );
  OAI211_X1 U18559 ( .C1(n15245), .C2(n20712), .A(n15244), .B(n15243), .ZN(
        P1_U2981) );
  NOR2_X1 U18560 ( .A1(n10416), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15249) );
  AOI21_X1 U18561 ( .B1(n15322), .B2(n15247), .A(n15246), .ZN(n15248) );
  MUX2_X1 U18562 ( .A(n15249), .B(n15332), .S(n15248), .Z(n15250) );
  XNOR2_X1 U18563 ( .A(n15250), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15447) );
  NAND2_X1 U18564 ( .A1(n20683), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15441) );
  OAI21_X1 U18565 ( .B1(n15344), .B2(n15251), .A(n15441), .ZN(n15254) );
  NOR2_X1 U18566 ( .A1(n15252), .A2(n20712), .ZN(n15253) );
  AOI211_X1 U18567 ( .C1(n15347), .C2(n15255), .A(n15254), .B(n15253), .ZN(
        n15256) );
  OAI21_X1 U18568 ( .B1(n15447), .B2(n15339), .A(n15256), .ZN(P1_U2982) );
  INV_X1 U18569 ( .A(n15322), .ZN(n15294) );
  INV_X1 U18570 ( .A(n15257), .ZN(n15259) );
  AOI211_X1 U18571 ( .C1(n15294), .C2(n15259), .A(n15258), .B(n15283), .ZN(
        n15276) );
  INV_X1 U18572 ( .A(n15262), .ZN(n15260) );
  NOR2_X1 U18573 ( .A1(n15261), .A2(n15260), .ZN(n15275) );
  NAND2_X1 U18574 ( .A1(n15276), .A2(n15275), .ZN(n15274) );
  NAND2_X1 U18575 ( .A1(n15274), .A2(n15262), .ZN(n15263) );
  XOR2_X1 U18576 ( .A(n15264), .B(n15263), .Z(n15457) );
  NAND2_X1 U18577 ( .A1(n15347), .A2(n15265), .ZN(n15266) );
  NAND2_X1 U18578 ( .A1(n20683), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15451) );
  OAI211_X1 U18579 ( .C1(n15344), .C2(n15267), .A(n15266), .B(n15451), .ZN(
        n15268) );
  AOI21_X1 U18580 ( .B1(n15269), .B2(n20649), .A(n15268), .ZN(n15270) );
  OAI21_X1 U18581 ( .B1(n15457), .B2(n15339), .A(n15270), .ZN(P1_U2983) );
  INV_X1 U18582 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n15271) );
  NOR2_X1 U18583 ( .A1(n20667), .A2(n15271), .ZN(n15461) );
  NOR2_X1 U18584 ( .A1(n20654), .A2(n15272), .ZN(n15273) );
  AOI211_X1 U18585 ( .C1(n20641), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15461), .B(n15273), .ZN(n15278) );
  OAI21_X1 U18586 ( .B1(n15276), .B2(n15275), .A(n15274), .ZN(n15459) );
  NAND2_X1 U18587 ( .A1(n15459), .A2(n20650), .ZN(n15277) );
  OAI211_X1 U18588 ( .C1(n15279), .C2(n20712), .A(n15278), .B(n15277), .ZN(
        P1_U2984) );
  NOR2_X1 U18589 ( .A1(n20667), .A2(n21330), .ZN(n15471) );
  NOR2_X1 U18590 ( .A1(n20654), .A2(n15280), .ZN(n15281) );
  AOI211_X1 U18591 ( .C1(n20641), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15471), .B(n15281), .ZN(n15289) );
  OAI21_X1 U18592 ( .B1(n15294), .B2(n15283), .A(n15282), .ZN(n15285) );
  NAND2_X1 U18593 ( .A1(n15285), .A2(n15284), .ZN(n15287) );
  XNOR2_X1 U18594 ( .A(n15332), .B(n21509), .ZN(n15286) );
  XNOR2_X1 U18595 ( .A(n15287), .B(n15286), .ZN(n15469) );
  NAND2_X1 U18596 ( .A1(n15469), .A2(n20650), .ZN(n15288) );
  OAI211_X1 U18597 ( .C1(n15290), .C2(n20712), .A(n15289), .B(n15288), .ZN(
        P1_U2985) );
  INV_X1 U18598 ( .A(n15291), .ZN(n15292) );
  AOI21_X1 U18599 ( .B1(n15294), .B2(n15293), .A(n15292), .ZN(n15308) );
  AND2_X1 U18600 ( .A1(n15295), .A2(n15296), .ZN(n15307) );
  NAND2_X1 U18601 ( .A1(n15308), .A2(n15307), .ZN(n15306) );
  NAND2_X1 U18602 ( .A1(n15306), .A2(n15296), .ZN(n15298) );
  XNOR2_X1 U18603 ( .A(n15298), .B(n15297), .ZN(n15485) );
  NAND2_X1 U18604 ( .A1(n20683), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15478) );
  NAND2_X1 U18605 ( .A1(n20641), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15299) );
  OAI211_X1 U18606 ( .C1(n20654), .C2(n15300), .A(n15478), .B(n15299), .ZN(
        n15301) );
  AOI21_X1 U18607 ( .B1(n15302), .B2(n20649), .A(n15301), .ZN(n15303) );
  OAI21_X1 U18608 ( .B1(n15339), .B2(n15485), .A(n15303), .ZN(P1_U2986) );
  NOR2_X1 U18609 ( .A1(n20667), .A2(n21328), .ZN(n15496) );
  NOR2_X1 U18610 ( .A1(n20654), .A2(n15304), .ZN(n15305) );
  AOI211_X1 U18611 ( .C1(n20641), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15496), .B(n15305), .ZN(n15310) );
  OAI21_X1 U18612 ( .B1(n15308), .B2(n15307), .A(n15306), .ZN(n15486) );
  NAND2_X1 U18613 ( .A1(n15486), .A2(n20650), .ZN(n15309) );
  OAI211_X1 U18614 ( .C1(n15311), .C2(n20712), .A(n15310), .B(n15309), .ZN(
        P1_U2987) );
  INV_X1 U18615 ( .A(n15342), .ZN(n15313) );
  NOR2_X1 U18616 ( .A1(n15324), .A2(n15312), .ZN(n15340) );
  AOI21_X1 U18617 ( .B1(n15313), .B2(n17388), .A(n15340), .ZN(n15314) );
  AOI21_X1 U18618 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n15342), .A(
        n15314), .ZN(n15334) );
  INV_X1 U18619 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15331) );
  NOR3_X1 U18620 ( .A1(n15323), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n10416), .ZN(n15326) );
  INV_X1 U18621 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21428) );
  NOR3_X1 U18622 ( .A1(n15322), .A2(n15324), .A3(n21428), .ZN(n15315) );
  NOR2_X1 U18623 ( .A1(n15326), .A2(n15315), .ZN(n15316) );
  XNOR2_X1 U18624 ( .A(n15316), .B(n21437), .ZN(n15512) );
  NAND2_X1 U18625 ( .A1(n20683), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n15507) );
  NAND2_X1 U18626 ( .A1(n20641), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15317) );
  OAI211_X1 U18627 ( .C1(n20654), .C2(n15318), .A(n15507), .B(n15317), .ZN(
        n15319) );
  AOI21_X1 U18628 ( .B1(n15320), .B2(n20649), .A(n15319), .ZN(n15321) );
  OAI21_X1 U18629 ( .B1(n15512), .B2(n15339), .A(n15321), .ZN(P1_U2988) );
  XNOR2_X1 U18630 ( .A(n15322), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15325) );
  INV_X1 U18631 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n17356) );
  NOR2_X1 U18632 ( .A1(n20667), .A2(n17356), .ZN(n15520) );
  NOR2_X1 U18633 ( .A1(n15344), .A2(n17348), .ZN(n15327) );
  AOI211_X1 U18634 ( .C1(n15347), .C2(n17354), .A(n15520), .B(n15327), .ZN(
        n15330) );
  NAND2_X1 U18635 ( .A1(n15328), .A2(n20649), .ZN(n15329) );
  OAI211_X1 U18636 ( .C1(n9642), .C2(n15339), .A(n15330), .B(n15329), .ZN(
        P1_U2989) );
  XNOR2_X1 U18637 ( .A(n15332), .B(n15331), .ZN(n15333) );
  XNOR2_X1 U18638 ( .A(n15334), .B(n15333), .ZN(n15532) );
  INV_X1 U18639 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20510) );
  NOR2_X1 U18640 ( .A1(n20667), .A2(n20510), .ZN(n15525) );
  AOI21_X1 U18641 ( .B1(n20641), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n15525), .ZN(n15335) );
  OAI21_X1 U18642 ( .B1(n15336), .B2(n20654), .A(n15335), .ZN(n15337) );
  AOI21_X1 U18643 ( .B1(n20513), .B2(n20649), .A(n15337), .ZN(n15338) );
  OAI21_X1 U18644 ( .B1(n15532), .B2(n15339), .A(n15338), .ZN(P1_U2990) );
  XNOR2_X1 U18645 ( .A(n15340), .B(n17388), .ZN(n15341) );
  XNOR2_X1 U18646 ( .A(n15342), .B(n15341), .ZN(n17385) );
  NAND2_X1 U18647 ( .A1(n17385), .A2(n20650), .ZN(n15349) );
  NAND2_X1 U18648 ( .A1(n20683), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n17380) );
  OAI21_X1 U18649 ( .B1(n15344), .B2(n15343), .A(n17380), .ZN(n15345) );
  AOI21_X1 U18650 ( .B1(n15347), .B2(n15346), .A(n15345), .ZN(n15348) );
  OAI211_X1 U18651 ( .C1(n20712), .C2(n15350), .A(n15349), .B(n15348), .ZN(
        P1_U2991) );
  NAND2_X1 U18652 ( .A1(n15351), .A2(n20699), .ZN(n15358) );
  OAI211_X1 U18653 ( .C1(n20668), .C2(n15359), .A(n15358), .B(n15357), .ZN(
        P1_U3002) );
  INV_X1 U18654 ( .A(n15360), .ZN(n15368) );
  NAND2_X1 U18655 ( .A1(n15361), .A2(n20699), .ZN(n15367) );
  NOR2_X1 U18656 ( .A1(n15362), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15363) );
  AOI211_X1 U18657 ( .C1(n15365), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15364), .B(n15363), .ZN(n15366) );
  OAI211_X1 U18658 ( .C1(n20668), .C2(n15368), .A(n15367), .B(n15366), .ZN(
        P1_U3004) );
  OAI21_X1 U18659 ( .B1(n15370), .B2(n15369), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15375) );
  NAND3_X1 U18660 ( .A1(n15391), .A2(n15372), .A3(n15371), .ZN(n15373) );
  NAND3_X1 U18661 ( .A1(n15375), .A2(n15374), .A3(n15373), .ZN(n15376) );
  AOI21_X1 U18662 ( .B1(n15377), .B2(n20696), .A(n15376), .ZN(n15378) );
  OAI21_X1 U18663 ( .B1(n15379), .B2(n20666), .A(n15378), .ZN(P1_U3005) );
  INV_X1 U18664 ( .A(n15380), .ZN(n15382) );
  AOI21_X1 U18665 ( .B1(n15382), .B2(n15394), .A(n15381), .ZN(n15386) );
  NAND3_X1 U18666 ( .A1(n15391), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n15385), .ZN(n15383) );
  OAI211_X1 U18667 ( .C1(n15386), .C2(n15385), .A(n15384), .B(n15383), .ZN(
        n15387) );
  AOI21_X1 U18668 ( .B1(n15388), .B2(n20696), .A(n15387), .ZN(n15389) );
  OAI21_X1 U18669 ( .B1(n15390), .B2(n20666), .A(n15389), .ZN(P1_U3007) );
  NAND2_X1 U18670 ( .A1(n15391), .A2(n15394), .ZN(n15393) );
  OAI211_X1 U18671 ( .C1(n15395), .C2(n15394), .A(n15393), .B(n15392), .ZN(
        n15396) );
  AOI21_X1 U18672 ( .B1(n15397), .B2(n20696), .A(n15396), .ZN(n15398) );
  OAI21_X1 U18673 ( .B1(n15399), .B2(n20666), .A(n15398), .ZN(P1_U3008) );
  INV_X1 U18674 ( .A(n15400), .ZN(n15409) );
  NAND2_X1 U18675 ( .A1(n15401), .A2(n20699), .ZN(n15408) );
  XNOR2_X1 U18676 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15402) );
  NOR2_X1 U18677 ( .A1(n15403), .A2(n15402), .ZN(n15405) );
  AOI211_X1 U18678 ( .C1(n15406), .C2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15405), .B(n15404), .ZN(n15407) );
  OAI211_X1 U18679 ( .C1(n20668), .C2(n15409), .A(n15408), .B(n15407), .ZN(
        P1_U3009) );
  INV_X1 U18680 ( .A(n15410), .ZN(n15420) );
  NAND3_X1 U18681 ( .A1(n15420), .A2(n15412), .A3(n15411), .ZN(n15414) );
  OAI211_X1 U18682 ( .C1(n15424), .C2(n15415), .A(n15414), .B(n15413), .ZN(
        n15416) );
  AOI21_X1 U18683 ( .B1(n15417), .B2(n20696), .A(n15416), .ZN(n15418) );
  OAI21_X1 U18684 ( .B1(n15419), .B2(n20666), .A(n15418), .ZN(P1_U3011) );
  NAND2_X1 U18685 ( .A1(n15420), .A2(n15423), .ZN(n15422) );
  OAI211_X1 U18686 ( .C1(n15424), .C2(n15423), .A(n15422), .B(n15421), .ZN(
        n15425) );
  AOI21_X1 U18687 ( .B1(n15426), .B2(n20696), .A(n15425), .ZN(n15427) );
  OAI21_X1 U18688 ( .B1(n15428), .B2(n20666), .A(n15427), .ZN(P1_U3012) );
  INV_X1 U18689 ( .A(n15429), .ZN(n15439) );
  NAND3_X1 U18690 ( .A1(n15431), .A2(n15430), .A3(n20699), .ZN(n15438) );
  INV_X1 U18691 ( .A(n15432), .ZN(n15433) );
  AOI21_X1 U18692 ( .B1(n15433), .B2(n20702), .A(n15481), .ZN(n15443) );
  INV_X1 U18693 ( .A(n15443), .ZN(n15436) );
  NOR3_X1 U18694 ( .A1(n15450), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15433), .ZN(n15434) );
  AOI211_X1 U18695 ( .C1(n15436), .C2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15435), .B(n15434), .ZN(n15437) );
  OAI211_X1 U18696 ( .C1(n20668), .C2(n15439), .A(n15438), .B(n15437), .ZN(
        P1_U3013) );
  NOR2_X1 U18697 ( .A1(n15450), .A2(n15440), .ZN(n15448) );
  AOI21_X1 U18698 ( .B1(n15448), .B2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15442) );
  OAI21_X1 U18699 ( .B1(n15443), .B2(n15442), .A(n15441), .ZN(n15444) );
  AOI21_X1 U18700 ( .B1(n15445), .B2(n20696), .A(n15444), .ZN(n15446) );
  OAI21_X1 U18701 ( .B1(n15447), .B2(n20666), .A(n15446), .ZN(P1_U3014) );
  INV_X1 U18702 ( .A(n15448), .ZN(n15453) );
  OAI21_X1 U18703 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15449), .A(
        n9921), .ZN(n15462) );
  NOR3_X1 U18704 ( .A1(n15450), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n21509), .ZN(n15460) );
  OAI21_X1 U18705 ( .B1(n15462), .B2(n15460), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15452) );
  OAI211_X1 U18706 ( .C1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15453), .A(
        n15452), .B(n15451), .ZN(n15454) );
  AOI21_X1 U18707 ( .B1(n20696), .B2(n15455), .A(n15454), .ZN(n15456) );
  OAI21_X1 U18708 ( .B1(n15457), .B2(n20666), .A(n15456), .ZN(P1_U3015) );
  INV_X1 U18709 ( .A(n15458), .ZN(n15465) );
  NAND2_X1 U18710 ( .A1(n15459), .A2(n20699), .ZN(n15464) );
  AOI211_X1 U18711 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15462), .A(
        n15461), .B(n15460), .ZN(n15463) );
  OAI211_X1 U18712 ( .C1(n20668), .C2(n15465), .A(n15464), .B(n15463), .ZN(
        P1_U3016) );
  INV_X1 U18713 ( .A(n15466), .ZN(n15487) );
  NOR2_X1 U18714 ( .A1(n15467), .A2(n15487), .ZN(n15518) );
  NAND2_X1 U18715 ( .A1(n15468), .A2(n15518), .ZN(n15528) );
  NOR2_X1 U18716 ( .A1(n15528), .A2(n15519), .ZN(n15510) );
  INV_X1 U18717 ( .A(n15510), .ZN(n15476) );
  NAND4_X1 U18718 ( .A1(n21509), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15475) );
  NAND2_X1 U18719 ( .A1(n15469), .A2(n20699), .ZN(n15474) );
  NOR2_X1 U18720 ( .A1(n9921), .A2(n21509), .ZN(n15470) );
  AOI211_X1 U18721 ( .C1(n15472), .C2(n20696), .A(n15471), .B(n15470), .ZN(
        n15473) );
  OAI211_X1 U18722 ( .C1(n15476), .C2(n15475), .A(n15474), .B(n15473), .ZN(
        P1_U3017) );
  INV_X1 U18723 ( .A(n15477), .ZN(n15480) );
  INV_X1 U18724 ( .A(n15478), .ZN(n15479) );
  AOI21_X1 U18725 ( .B1(n15480), .B2(n20696), .A(n15479), .ZN(n15484) );
  OAI21_X1 U18726 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15482), .A(
        n15481), .ZN(n15483) );
  OAI211_X1 U18727 ( .C1(n15485), .C2(n20666), .A(n15484), .B(n15483), .ZN(
        P1_U3018) );
  INV_X1 U18728 ( .A(n15486), .ZN(n15504) );
  INV_X1 U18729 ( .A(n20675), .ZN(n15493) );
  INV_X1 U18730 ( .A(n20679), .ZN(n15490) );
  NOR3_X1 U18731 ( .A1(n15488), .A2(n15519), .A3(n15487), .ZN(n15489) );
  OAI22_X1 U18732 ( .A1(n15490), .A2(n15489), .B1(n15500), .B2(n20676), .ZN(
        n15491) );
  NOR2_X1 U18733 ( .A1(n15492), .A2(n15491), .ZN(n15508) );
  OAI21_X1 U18734 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15493), .A(
        n15508), .ZN(n15497) );
  NOR2_X1 U18735 ( .A1(n15494), .A2(n20668), .ZN(n15495) );
  AOI211_X1 U18736 ( .C1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15497), .A(
        n15496), .B(n15495), .ZN(n15503) );
  INV_X1 U18737 ( .A(n20674), .ZN(n15498) );
  NAND3_X1 U18738 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20658), .A3(
        n15498), .ZN(n17403) );
  INV_X1 U18739 ( .A(n17403), .ZN(n15501) );
  NAND3_X1 U18740 ( .A1(n15501), .A2(n15500), .A3(n15499), .ZN(n15502) );
  OAI211_X1 U18741 ( .C1(n15504), .C2(n20666), .A(n15503), .B(n15502), .ZN(
        P1_U3019) );
  NAND2_X1 U18742 ( .A1(n15505), .A2(n20696), .ZN(n15506) );
  OAI211_X1 U18743 ( .C1(n15508), .C2(n21437), .A(n15507), .B(n15506), .ZN(
        n15509) );
  AOI21_X1 U18744 ( .B1(n15510), .B2(n21437), .A(n15509), .ZN(n15511) );
  OAI21_X1 U18745 ( .B1(n15512), .B2(n20666), .A(n15511), .ZN(P1_U3020) );
  NAND2_X1 U18746 ( .A1(n20679), .A2(n15513), .ZN(n15515) );
  OR2_X1 U18747 ( .A1(n20676), .A2(n15514), .ZN(n20685) );
  AOI21_X1 U18748 ( .B1(n20672), .B2(n15518), .A(n15517), .ZN(n15530) );
  OAI21_X1 U18749 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15519), .ZN(n15522) );
  AOI21_X1 U18750 ( .B1(n17346), .B2(n20696), .A(n15520), .ZN(n15521) );
  OAI21_X1 U18751 ( .B1(n15528), .B2(n15522), .A(n15521), .ZN(n15523) );
  AOI21_X1 U18752 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n15530), .A(
        n15523), .ZN(n15524) );
  OAI21_X1 U18753 ( .B1(n9642), .B2(n20666), .A(n15524), .ZN(P1_U3021) );
  INV_X1 U18754 ( .A(n20507), .ZN(n15526) );
  AOI21_X1 U18755 ( .B1(n15526), .B2(n20696), .A(n15525), .ZN(n15527) );
  OAI21_X1 U18756 ( .B1(n15528), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15527), .ZN(n15529) );
  AOI21_X1 U18757 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15530), .A(
        n15529), .ZN(n15531) );
  OAI21_X1 U18758 ( .B1(n15532), .B2(n20666), .A(n15531), .ZN(P1_U3022) );
  INV_X1 U18759 ( .A(n15533), .ZN(n15535) );
  NAND2_X1 U18760 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21000), .ZN(n15544) );
  NAND2_X1 U18761 ( .A1(n11586), .A2(n15544), .ZN(n15534) );
  OAI211_X1 U18762 ( .C1(n21155), .C2(n21376), .A(n15535), .B(n15534), .ZN(
        n15542) );
  NOR2_X1 U18763 ( .A1(n15536), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n15541) );
  OR2_X1 U18764 ( .A1(n21384), .A2(n15537), .ZN(n15538) );
  MUX2_X1 U18765 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15542), .S(
        n20707), .Z(P1_U3478) );
  NAND2_X1 U18766 ( .A1(n15543), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21243) );
  NAND2_X1 U18767 ( .A1(n21243), .A2(n21163), .ZN(n20835) );
  NOR2_X1 U18768 ( .A1(n15543), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15545) );
  INV_X1 U18769 ( .A(n15544), .ZN(n15556) );
  OAI22_X1 U18770 ( .A1(n20835), .A2(n15545), .B1(n21188), .B2(n15556), .ZN(
        n15546) );
  MUX2_X1 U18771 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15546), .S(
        n20707), .Z(P1_U3477) );
  XNOR2_X1 U18772 ( .A(n15547), .B(n21243), .ZN(n15548) );
  OAI22_X1 U18773 ( .A1(n15548), .A2(n21376), .B1(n21127), .B2(n15556), .ZN(
        n15549) );
  MUX2_X1 U18774 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15549), .S(
        n20707), .Z(P1_U3476) );
  INV_X1 U18775 ( .A(n21092), .ZN(n21097) );
  INV_X1 U18776 ( .A(n15543), .ZN(n15552) );
  NAND2_X1 U18777 ( .A1(n20714), .A2(n15552), .ZN(n21156) );
  NAND3_X1 U18778 ( .A1(n21097), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(n21156), 
        .ZN(n15555) );
  INV_X1 U18779 ( .A(n15550), .ZN(n15554) );
  NOR2_X1 U18780 ( .A1(n20902), .A2(n21243), .ZN(n20966) );
  AOI21_X1 U18781 ( .B1(n15555), .B2(n15554), .A(n20966), .ZN(n15557) );
  INV_X1 U18782 ( .A(n20720), .ZN(n20994) );
  OAI22_X1 U18783 ( .A1(n15557), .A2(n21376), .B1(n20994), .B2(n15556), .ZN(
        n15558) );
  MUX2_X1 U18784 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15558), .S(
        n20707), .Z(P1_U3475) );
  INV_X1 U18785 ( .A(n15559), .ZN(n15563) );
  NAND2_X1 U18786 ( .A1(n15560), .A2(n15565), .ZN(n15562) );
  OAI22_X1 U18787 ( .A1(n12778), .A2(n20703), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15567) );
  NAND3_X1 U18788 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n15567), .A3(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15561) );
  OAI211_X1 U18789 ( .C1(n15573), .C2(n15563), .A(n15562), .B(n15561), .ZN(
        n15564) );
  MUX2_X1 U18790 ( .A(n15564), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15577), .Z(P1_U3473) );
  NAND2_X1 U18791 ( .A1(n15566), .A2(n15565), .ZN(n15570) );
  INV_X1 U18792 ( .A(n15567), .ZN(n15568) );
  NAND3_X1 U18793 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n15568), .A3(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15569) );
  OAI211_X1 U18794 ( .C1(n15573), .C2(n15571), .A(n15570), .B(n15569), .ZN(
        n15572) );
  MUX2_X1 U18795 ( .A(n15572), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15577), .Z(P1_U3472) );
  OAI22_X1 U18796 ( .A1(n15576), .A2(n15575), .B1(n15574), .B2(n15573), .ZN(
        n15578) );
  MUX2_X1 U18797 ( .A(n15578), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15577), .Z(P1_U3469) );
  NAND3_X1 U18798 ( .A1(n15581), .A2(n15580), .A3(n15579), .ZN(P1_U3163) );
  NOR2_X1 U18799 ( .A1(n15978), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n15583) );
  INV_X1 U18800 ( .A(n15582), .ZN(n20376) );
  OAI21_X1 U18801 ( .B1(n15583), .B2(n20376), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n15587) );
  OAI21_X1 U18802 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n15584), .ZN(n17421) );
  OAI21_X1 U18803 ( .B1(n20381), .B2(n20302), .A(n17421), .ZN(n15585) );
  OAI21_X1 U18804 ( .B1(n15587), .B2(n15586), .A(n15585), .ZN(n15592) );
  AOI22_X1 U18805 ( .A1(n15588), .A2(n20304), .B1(n20369), .B2(n19694), .ZN(
        n15589) );
  NAND2_X1 U18806 ( .A1(n15590), .A2(n15589), .ZN(n15591) );
  MUX2_X1 U18807 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n15592), .S(n15591), 
        .Z(P2_U3610) );
  AOI21_X1 U18808 ( .B1(n15593), .B2(n9607), .A(n12755), .ZN(n16431) );
  INV_X1 U18809 ( .A(n16431), .ZN(n16166) );
  INV_X1 U18810 ( .A(n15595), .ZN(n16164) );
  AOI21_X1 U18811 ( .B1(n15594), .B2(n16164), .A(n19616), .ZN(n15597) );
  OAI21_X1 U18812 ( .B1(n15597), .B2(n15931), .A(n15596), .ZN(n15606) );
  AOI22_X1 U18813 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19605), .B1(n15934), 
        .B2(P2_EBX_REG_29__SCAN_IN), .ZN(n15598) );
  OAI21_X1 U18814 ( .B1(n16162), .B2(n19625), .A(n15598), .ZN(n15603) );
  NOR2_X1 U18815 ( .A1(n16438), .A2(n19611), .ZN(n15602) );
  OAI211_X1 U18816 ( .C1(n15937), .C2(n16166), .A(n15606), .B(n15605), .ZN(
        P2_U2826) );
  AOI21_X1 U18817 ( .B1(n15607), .B2(n9761), .A(n19616), .ZN(n15608) );
  OAI21_X1 U18818 ( .B1(n15608), .B2(n15931), .A(n15594), .ZN(n15613) );
  AOI22_X1 U18819 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n19605), .B1(n15934), 
        .B2(P2_EBX_REG_28__SCAN_IN), .ZN(n15609) );
  OAI21_X1 U18820 ( .B1(n15610), .B2(n19625), .A(n15609), .ZN(n15611) );
  OR2_X1 U18821 ( .A1(n15630), .A2(n15614), .ZN(n15615) );
  NAND2_X1 U18822 ( .A1(n15616), .A2(n15615), .ZN(n16447) );
  AOI21_X1 U18823 ( .B1(n15617), .B2(n10274), .A(n19616), .ZN(n15619) );
  OAI21_X1 U18824 ( .B1(n15619), .B2(n15931), .A(n15607), .ZN(n15628) );
  NOR2_X1 U18825 ( .A1(n15620), .A2(n15621), .ZN(n15622) );
  AOI22_X1 U18826 ( .A1(P2_REIP_REG_27__SCAN_IN), .A2(n19605), .B1(n15934), 
        .B2(P2_EBX_REG_27__SCAN_IN), .ZN(n15624) );
  NAND2_X1 U18827 ( .A1(n15930), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15623) );
  OAI211_X1 U18828 ( .C1(n15625), .C2(n15875), .A(n15624), .B(n15623), .ZN(
        n15626) );
  AOI21_X1 U18829 ( .B1(n10453), .B2(n15933), .A(n15626), .ZN(n15627) );
  OAI211_X1 U18830 ( .C1(n15937), .C2(n16447), .A(n15628), .B(n15627), .ZN(
        P2_U2828) );
  AND2_X1 U18831 ( .A1(n15645), .A2(n15629), .ZN(n15631) );
  OR2_X1 U18832 ( .A1(n15631), .A2(n15630), .ZN(n16459) );
  INV_X1 U18833 ( .A(n15633), .ZN(n16183) );
  AOI21_X1 U18834 ( .B1(n15632), .B2(n16183), .A(n19616), .ZN(n15634) );
  OAI21_X1 U18835 ( .B1(n15634), .B2(n15931), .A(n15617), .ZN(n15642) );
  AND2_X1 U18836 ( .A1(n9657), .A2(n15635), .ZN(n15636) );
  AOI22_X1 U18837 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n19605), .B1(n15934), 
        .B2(P2_EBX_REG_26__SCAN_IN), .ZN(n15638) );
  NAND2_X1 U18838 ( .A1(n15930), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15637) );
  OAI211_X1 U18839 ( .C1(n15639), .C2(n15875), .A(n15638), .B(n15637), .ZN(
        n15640) );
  AOI21_X1 U18840 ( .B1(n10457), .B2(n15933), .A(n15640), .ZN(n15641) );
  OAI211_X1 U18841 ( .C1(n15937), .C2(n16459), .A(n15642), .B(n15641), .ZN(
        P2_U2829) );
  INV_X1 U18842 ( .A(n15643), .ZN(n15646) );
  OAI21_X1 U18843 ( .B1(n15646), .B2(n10236), .A(n15645), .ZN(n16192) );
  AOI21_X1 U18844 ( .B1(n15647), .B2(n10279), .A(n19616), .ZN(n15648) );
  OAI21_X1 U18845 ( .B1(n15648), .B2(n15931), .A(n15632), .ZN(n15659) );
  NAND2_X1 U18846 ( .A1(n15649), .A2(n15650), .ZN(n15651) );
  AND2_X1 U18847 ( .A1(n9657), .A2(n15651), .ZN(n16466) );
  XNOR2_X1 U18848 ( .A(n15653), .B(n15652), .ZN(n15656) );
  AOI22_X1 U18849 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19605), .B1(n15934), 
        .B2(P2_EBX_REG_25__SCAN_IN), .ZN(n15655) );
  NAND2_X1 U18850 ( .A1(n15930), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15654) );
  OAI211_X1 U18851 ( .C1(n15656), .C2(n15875), .A(n15655), .B(n15654), .ZN(
        n15657) );
  AOI21_X1 U18852 ( .B1(n16466), .B2(n15933), .A(n15657), .ZN(n15658) );
  OAI211_X1 U18853 ( .C1(n16192), .C2(n15937), .A(n15659), .B(n15658), .ZN(
        P2_U2830) );
  INV_X1 U18854 ( .A(n15660), .ZN(n15662) );
  OAI21_X1 U18855 ( .B1(n15662), .B2(n10237), .A(n15643), .ZN(n16486) );
  AOI21_X1 U18856 ( .B1(n15663), .B2(n10277), .A(n19616), .ZN(n15665) );
  OAI21_X1 U18857 ( .B1(n15665), .B2(n15931), .A(n15647), .ZN(n15674) );
  OR2_X1 U18858 ( .A1(n15666), .A2(n15667), .ZN(n15668) );
  AND2_X1 U18859 ( .A1(n15649), .A2(n15668), .ZN(n16483) );
  AOI22_X1 U18860 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n19605), .B1(n15934), 
        .B2(P2_EBX_REG_24__SCAN_IN), .ZN(n15670) );
  NAND2_X1 U18861 ( .A1(n15930), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15669) );
  OAI211_X1 U18862 ( .C1(n15671), .C2(n15875), .A(n15670), .B(n15669), .ZN(
        n15672) );
  AOI21_X1 U18863 ( .B1(n16483), .B2(n15933), .A(n15672), .ZN(n15673) );
  OAI211_X1 U18864 ( .C1(n16486), .C2(n15937), .A(n15674), .B(n15673), .ZN(
        P2_U2831) );
  OAI21_X1 U18865 ( .B1(n15675), .B2(n15676), .A(n15660), .ZN(n16496) );
  AOI21_X1 U18866 ( .B1(n9709), .B2(n9765), .A(n19616), .ZN(n15677) );
  OAI21_X1 U18867 ( .B1(n15677), .B2(n15931), .A(n15663), .ZN(n15686) );
  AND2_X1 U18868 ( .A1(n15694), .A2(n15679), .ZN(n15680) );
  NOR2_X1 U18869 ( .A1(n15666), .A2(n15680), .ZN(n16499) );
  NAND2_X1 U18870 ( .A1(n15681), .A2(n19609), .ZN(n15683) );
  AOI22_X1 U18871 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19605), .B1(n15934), 
        .B2(P2_EBX_REG_23__SCAN_IN), .ZN(n15682) );
  OAI211_X1 U18872 ( .C1(n19625), .C2(n10317), .A(n15683), .B(n15682), .ZN(
        n15684) );
  AOI21_X1 U18873 ( .B1(n16499), .B2(n15933), .A(n15684), .ZN(n15685) );
  OAI211_X1 U18874 ( .C1(n16496), .C2(n15937), .A(n15686), .B(n15685), .ZN(
        P2_U2832) );
  AND2_X1 U18875 ( .A1(n15688), .A2(n15687), .ZN(n15689) );
  OR2_X1 U18876 ( .A1(n15689), .A2(n15675), .ZN(n16510) );
  AOI21_X1 U18877 ( .B1(n15690), .B2(n16225), .A(n19616), .ZN(n15691) );
  OAI21_X1 U18878 ( .B1(n15931), .B2(n15691), .A(n9709), .ZN(n15700) );
  NAND2_X1 U18879 ( .A1(n12820), .A2(n15692), .ZN(n15693) );
  AND2_X1 U18880 ( .A1(n15694), .A2(n15693), .ZN(n16513) );
  AOI22_X1 U18881 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19605), .B1(n15934), 
        .B2(P2_EBX_REG_22__SCAN_IN), .ZN(n15696) );
  NAND2_X1 U18882 ( .A1(n15930), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15695) );
  OAI211_X1 U18883 ( .C1(n15697), .C2(n15875), .A(n15696), .B(n15695), .ZN(
        n15698) );
  AOI21_X1 U18884 ( .B1(n16513), .B2(n15933), .A(n15698), .ZN(n15699) );
  OAI211_X1 U18885 ( .C1(n16510), .C2(n15937), .A(n15700), .B(n15699), .ZN(
        P2_U2833) );
  INV_X1 U18886 ( .A(n15701), .ZN(n16000) );
  INV_X1 U18887 ( .A(n15702), .ZN(n15716) );
  INV_X1 U18888 ( .A(n15703), .ZN(n15704) );
  AOI21_X1 U18889 ( .B1(n15716), .B2(n15704), .A(n19616), .ZN(n15705) );
  OAI21_X1 U18890 ( .B1(n15705), .B2(n15931), .A(n15690), .ZN(n15712) );
  INV_X1 U18891 ( .A(n15706), .ZN(n16105) );
  AOI22_X1 U18892 ( .A1(P2_REIP_REG_21__SCAN_IN), .A2(n19605), .B1(n15934), 
        .B2(P2_EBX_REG_21__SCAN_IN), .ZN(n15708) );
  NAND2_X1 U18893 ( .A1(n15930), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15707) );
  OAI211_X1 U18894 ( .C1(n15709), .C2(n15875), .A(n15708), .B(n15707), .ZN(
        n15710) );
  AOI21_X1 U18895 ( .B1(n16105), .B2(n15933), .A(n15710), .ZN(n15711) );
  OAI211_X1 U18896 ( .C1(n15937), .C2(n16000), .A(n15712), .B(n15711), .ZN(
        P2_U2834) );
  OAI21_X1 U18897 ( .B1(n12817), .B2(n15714), .A(n15713), .ZN(n16519) );
  AOI21_X1 U18898 ( .B1(n15715), .B2(n16237), .A(n19616), .ZN(n15717) );
  OAI21_X1 U18899 ( .B1(n15931), .B2(n15717), .A(n15716), .ZN(n15728) );
  AOI22_X1 U18900 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n19605), .B1(n15934), 
        .B2(P2_EBX_REG_20__SCAN_IN), .ZN(n15718) );
  OAI21_X1 U18901 ( .B1(n15719), .B2(n19625), .A(n15718), .ZN(n15725) );
  INV_X1 U18902 ( .A(n15720), .ZN(n15723) );
  NAND2_X1 U18903 ( .A1(n15732), .A2(n15721), .ZN(n15722) );
  NAND2_X1 U18904 ( .A1(n15723), .A2(n15722), .ZN(n16527) );
  NOR2_X1 U18905 ( .A1(n16527), .A2(n19611), .ZN(n15724) );
  AOI211_X1 U18906 ( .C1(n19609), .C2(n15726), .A(n15725), .B(n15724), .ZN(
        n15727) );
  OAI211_X1 U18907 ( .C1(n15937), .C2(n16519), .A(n15728), .B(n15727), .ZN(
        P2_U2835) );
  NOR2_X1 U18908 ( .A1(n9714), .A2(n15729), .ZN(n15730) );
  OR2_X1 U18909 ( .A1(n12817), .A2(n15730), .ZN(n16538) );
  INV_X1 U18910 ( .A(n15732), .ZN(n15733) );
  AOI21_X1 U18911 ( .B1(n15734), .B2(n15731), .A(n15733), .ZN(n16535) );
  NAND2_X1 U18912 ( .A1(n15735), .A2(n19609), .ZN(n15738) );
  INV_X1 U18913 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20423) );
  OAI21_X1 U18914 ( .B1(n15816), .B2(n20423), .A(n16416), .ZN(n15736) );
  AOI21_X1 U18915 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n15934), .A(n15736), .ZN(
        n15737) );
  OAI211_X1 U18916 ( .C1(n19625), .C2(n15739), .A(n15738), .B(n15737), .ZN(
        n15743) );
  OAI21_X1 U18917 ( .B1(n15740), .B2(n16252), .A(n15791), .ZN(n15741) );
  AOI21_X1 U18918 ( .B1(n15912), .B2(n15741), .A(n10309), .ZN(n15742) );
  AOI211_X1 U18919 ( .C1(n15933), .C2(n16535), .A(n15743), .B(n15742), .ZN(
        n15744) );
  OAI21_X1 U18920 ( .B1(n16538), .B2(n15937), .A(n15744), .ZN(P2_U2836) );
  AOI21_X1 U18921 ( .B1(n15759), .B2(n15745), .A(n19616), .ZN(n15747) );
  INV_X1 U18922 ( .A(n15740), .ZN(n15746) );
  OAI21_X1 U18923 ( .B1(n15931), .B2(n15747), .A(n15746), .ZN(n15757) );
  INV_X1 U18924 ( .A(n15731), .ZN(n15748) );
  AOI21_X1 U18925 ( .B1(n15749), .B2(n12801), .A(n15748), .ZN(n16549) );
  NAND2_X1 U18926 ( .A1(n15934), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15750) );
  OAI211_X1 U18927 ( .C1(n15751), .C2(n15816), .A(n15750), .B(n16416), .ZN(
        n15752) );
  AOI21_X1 U18928 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n15930), .A(
        n15752), .ZN(n15753) );
  OAI21_X1 U18929 ( .B1(n15754), .B2(n15875), .A(n15753), .ZN(n15755) );
  AOI21_X1 U18930 ( .B1(n16549), .B2(n15933), .A(n15755), .ZN(n15756) );
  OAI211_X1 U18931 ( .C1(n15937), .C2(n16552), .A(n15757), .B(n15756), .ZN(
        P2_U2837) );
  INV_X1 U18932 ( .A(n16261), .ZN(n16018) );
  INV_X1 U18933 ( .A(n15758), .ZN(n15775) );
  AOI21_X1 U18934 ( .B1(n15775), .B2(n10294), .A(n19616), .ZN(n15760) );
  OAI21_X1 U18935 ( .B1(n15760), .B2(n15931), .A(n15759), .ZN(n15768) );
  NAND2_X1 U18936 ( .A1(n15930), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15762) );
  AOI21_X1 U18937 ( .B1(n19605), .B2(P2_REIP_REG_17__SCAN_IN), .A(n19604), 
        .ZN(n15761) );
  OAI211_X1 U18938 ( .C1(n19607), .C2(n15763), .A(n15762), .B(n15761), .ZN(
        n15765) );
  NOR2_X1 U18939 ( .A1(n16127), .A2(n19611), .ZN(n15764) );
  AOI211_X1 U18940 ( .C1(n19609), .C2(n15766), .A(n15765), .B(n15764), .ZN(
        n15767) );
  OAI211_X1 U18941 ( .C1(n15937), .C2(n16018), .A(n15768), .B(n15767), .ZN(
        P2_U2838) );
  OR2_X1 U18942 ( .A1(n15769), .A2(n15770), .ZN(n15771) );
  NAND2_X1 U18943 ( .A1(n12795), .A2(n15771), .ZN(n16563) );
  AND2_X1 U18944 ( .A1(n14066), .A2(n15772), .ZN(n15773) );
  NOR2_X1 U18945 ( .A1(n12799), .A2(n15773), .ZN(n16560) );
  AOI21_X1 U18946 ( .B1(n15774), .B2(n16266), .A(n19616), .ZN(n15776) );
  OAI21_X1 U18947 ( .B1(n15931), .B2(n15776), .A(n15775), .ZN(n15780) );
  AOI21_X1 U18948 ( .B1(n19605), .B2(P2_REIP_REG_16__SCAN_IN), .A(n19604), 
        .ZN(n15777) );
  OAI21_X1 U18949 ( .B1(n19607), .B2(n10938), .A(n15777), .ZN(n15778) );
  AOI21_X1 U18950 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n15930), .A(
        n15778), .ZN(n15779) );
  OAI211_X1 U18951 ( .C1(n15875), .C2(n15781), .A(n15780), .B(n15779), .ZN(
        n15782) );
  AOI21_X1 U18952 ( .B1(n15933), .B2(n16560), .A(n15782), .ZN(n15783) );
  OAI21_X1 U18953 ( .B1(n15937), .B2(n16563), .A(n15783), .ZN(P2_U2839) );
  AND2_X1 U18954 ( .A1(n9720), .A2(n15784), .ZN(n15785) );
  OR2_X1 U18955 ( .A1(n15785), .A2(n15769), .ZN(n16576) );
  NAND2_X1 U18956 ( .A1(n15786), .A2(n19609), .ZN(n15789) );
  NOR2_X1 U18957 ( .A1(n19607), .A2(n11097), .ZN(n15787) );
  AOI211_X1 U18958 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n19605), .A(n19604), 
        .B(n15787), .ZN(n15788) );
  OAI211_X1 U18959 ( .C1(n19625), .C2(n15790), .A(n15789), .B(n15788), .ZN(
        n15795) );
  OAI21_X1 U18960 ( .B1(n15800), .B2(n16281), .A(n15791), .ZN(n15793) );
  INV_X1 U18961 ( .A(n15774), .ZN(n15792) );
  AOI21_X1 U18962 ( .B1(n15912), .B2(n15793), .A(n15792), .ZN(n15794) );
  AOI211_X1 U18963 ( .C1(n16573), .C2(n15933), .A(n15795), .B(n15794), .ZN(
        n15796) );
  OAI21_X1 U18964 ( .B1(n15937), .B2(n16576), .A(n15796), .ZN(P2_U2840) );
  OR2_X1 U18965 ( .A1(n15812), .A2(n15811), .ZN(n15814) );
  NAND2_X1 U18966 ( .A1(n15814), .A2(n15797), .ZN(n15798) );
  NAND2_X1 U18967 ( .A1(n9720), .A2(n15798), .ZN(n16581) );
  INV_X1 U18968 ( .A(n16585), .ZN(n15809) );
  AOI21_X1 U18969 ( .B1(n15799), .B2(n16294), .A(n19616), .ZN(n15801) );
  OAI21_X1 U18970 ( .B1(n15931), .B2(n15801), .A(n10298), .ZN(n15806) );
  AOI21_X1 U18971 ( .B1(n19605), .B2(P2_REIP_REG_14__SCAN_IN), .A(n19604), 
        .ZN(n15802) );
  OAI21_X1 U18972 ( .B1(n19607), .B2(n15803), .A(n15802), .ZN(n15804) );
  AOI21_X1 U18973 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n15930), .A(
        n15804), .ZN(n15805) );
  OAI211_X1 U18974 ( .C1(n15875), .C2(n15807), .A(n15806), .B(n15805), .ZN(
        n15808) );
  AOI21_X1 U18975 ( .B1(n15809), .B2(n15933), .A(n15808), .ZN(n15810) );
  OAI21_X1 U18976 ( .B1(n16581), .B2(n15937), .A(n15810), .ZN(P2_U2841) );
  NAND2_X1 U18977 ( .A1(n15812), .A2(n15811), .ZN(n15813) );
  NAND2_X1 U18978 ( .A1(n15815), .A2(n19609), .ZN(n15819) );
  INV_X1 U18979 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n20413) );
  OAI21_X1 U18980 ( .B1(n15816), .B2(n20413), .A(n16416), .ZN(n15817) );
  AOI21_X1 U18981 ( .B1(P2_EBX_REG_13__SCAN_IN), .B2(n15934), .A(n15817), .ZN(
        n15818) );
  OAI211_X1 U18982 ( .C1(n19625), .C2(n10321), .A(n15819), .B(n15818), .ZN(
        n15825) );
  INV_X1 U18983 ( .A(n15821), .ZN(n15820) );
  OAI21_X1 U18984 ( .B1(n19616), .B2(n15820), .A(n15912), .ZN(n15823) );
  NOR2_X1 U18985 ( .A1(n15944), .A2(n15821), .ZN(n15822) );
  MUX2_X1 U18986 ( .A(n15823), .B(n15822), .S(n16299), .Z(n15824) );
  AOI211_X1 U18987 ( .C1(n15933), .C2(n16598), .A(n15825), .B(n15824), .ZN(
        n15826) );
  OAI21_X1 U18988 ( .B1(n16044), .B2(n15937), .A(n15826), .ZN(P2_U2842) );
  INV_X1 U18989 ( .A(n15828), .ZN(n15827) );
  OAI21_X1 U18990 ( .B1(n15914), .B2(n15827), .A(n15912), .ZN(n15830) );
  NOR2_X1 U18991 ( .A1(n15944), .A2(n15828), .ZN(n15829) );
  MUX2_X1 U18992 ( .A(n15830), .B(n15829), .S(n16344), .Z(n15831) );
  INV_X1 U18993 ( .A(n15831), .ZN(n15840) );
  AOI21_X1 U18994 ( .B1(n19605), .B2(P2_REIP_REG_10__SCAN_IN), .A(n19604), 
        .ZN(n15833) );
  NAND2_X1 U18995 ( .A1(n15934), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n15832) );
  OAI211_X1 U18996 ( .C1(n19625), .C2(n15834), .A(n15833), .B(n15832), .ZN(
        n15835) );
  AOI21_X1 U18997 ( .B1(n15836), .B2(n19609), .A(n15835), .ZN(n15837) );
  OAI21_X1 U18998 ( .B1(n16647), .B2(n19611), .A(n15837), .ZN(n15838) );
  AOI21_X1 U18999 ( .B1(n16652), .B2(n19621), .A(n15838), .ZN(n15839) );
  NAND2_X1 U19000 ( .A1(n15840), .A2(n15839), .ZN(P2_U2845) );
  INV_X1 U19001 ( .A(n15842), .ZN(n15841) );
  OAI21_X1 U19002 ( .B1(n15914), .B2(n15841), .A(n15912), .ZN(n15844) );
  NOR2_X1 U19003 ( .A1(n15944), .A2(n15842), .ZN(n15843) );
  MUX2_X1 U19004 ( .A(n15844), .B(n15843), .S(n16356), .Z(n15853) );
  AOI21_X1 U19005 ( .B1(n19605), .B2(P2_REIP_REG_9__SCAN_IN), .A(n19604), .ZN(
        n15846) );
  NAND2_X1 U19006 ( .A1(n15934), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n15845) );
  OAI211_X1 U19007 ( .C1(n19625), .C2(n15847), .A(n15846), .B(n15845), .ZN(
        n15848) );
  AOI21_X1 U19008 ( .B1(n15849), .B2(n19609), .A(n15848), .ZN(n15851) );
  NAND2_X1 U19009 ( .A1(n16659), .A2(n15933), .ZN(n15850) );
  OAI211_X1 U19010 ( .C1(n16658), .C2(n15937), .A(n15851), .B(n15850), .ZN(
        n15852) );
  INV_X1 U19011 ( .A(n15855), .ZN(n15854) );
  NOR2_X1 U19012 ( .A1(n15944), .A2(n15854), .ZN(n15857) );
  OAI21_X1 U19013 ( .B1(n15914), .B2(n15855), .A(n15912), .ZN(n15856) );
  MUX2_X1 U19014 ( .A(n15857), .B(n15856), .S(n16378), .Z(n15867) );
  NAND2_X1 U19015 ( .A1(n16691), .A2(n19621), .ZN(n15865) );
  INV_X1 U19016 ( .A(n15858), .ZN(n15863) );
  AOI21_X1 U19017 ( .B1(n19605), .B2(P2_REIP_REG_7__SCAN_IN), .A(n19604), .ZN(
        n15860) );
  NAND2_X1 U19018 ( .A1(n15934), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n15859) );
  OAI211_X1 U19019 ( .C1(n19625), .C2(n15861), .A(n15860), .B(n15859), .ZN(
        n15862) );
  AOI21_X1 U19020 ( .B1(n15863), .B2(n19609), .A(n15862), .ZN(n15864) );
  OAI211_X1 U19021 ( .C1(n16686), .C2(n19611), .A(n15865), .B(n15864), .ZN(
        n15866) );
  INV_X1 U19022 ( .A(n15868), .ZN(n19617) );
  NOR2_X1 U19023 ( .A1(n15944), .A2(n19617), .ZN(n15870) );
  OAI21_X1 U19024 ( .B1(n15914), .B2(n15868), .A(n15912), .ZN(n15869) );
  MUX2_X1 U19025 ( .A(n15870), .B(n15869), .S(n16391), .Z(n15880) );
  AOI21_X1 U19026 ( .B1(n19605), .B2(P2_REIP_REG_6__SCAN_IN), .A(n19604), .ZN(
        n15872) );
  NAND2_X1 U19027 ( .A1(n15934), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n15871) );
  OAI211_X1 U19028 ( .C1(n19625), .C2(n10302), .A(n15872), .B(n15871), .ZN(
        n15873) );
  INV_X1 U19029 ( .A(n15873), .ZN(n15874) );
  OAI21_X1 U19030 ( .B1(n15876), .B2(n15875), .A(n15874), .ZN(n15877) );
  AOI21_X1 U19031 ( .B1(n16701), .B2(n15933), .A(n15877), .ZN(n15878) );
  OAI21_X1 U19032 ( .B1(n16704), .B2(n15937), .A(n15878), .ZN(n15879) );
  INV_X1 U19033 ( .A(n16430), .ZN(n19711) );
  NAND2_X1 U19034 ( .A1(n15883), .A2(n15882), .ZN(n15884) );
  NAND2_X1 U19035 ( .A1(n15881), .A2(n15884), .ZN(n19626) );
  AOI21_X1 U19036 ( .B1(n19605), .B2(P2_REIP_REG_4__SCAN_IN), .A(n19604), .ZN(
        n15886) );
  NAND2_X1 U19037 ( .A1(n15934), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n15885) );
  OAI211_X1 U19038 ( .C1(n19625), .C2(n16418), .A(n15886), .B(n15885), .ZN(
        n15887) );
  AOI21_X1 U19039 ( .B1(n15888), .B2(n19609), .A(n15887), .ZN(n15889) );
  OAI21_X1 U19040 ( .B1(n19626), .B2(n19611), .A(n15889), .ZN(n15895) );
  INV_X1 U19041 ( .A(n15891), .ZN(n15890) );
  NOR2_X1 U19042 ( .A1(n15944), .A2(n15890), .ZN(n15893) );
  OAI21_X1 U19043 ( .B1(n15914), .B2(n15891), .A(n15912), .ZN(n15892) );
  MUX2_X1 U19044 ( .A(n15893), .B(n15892), .S(n16426), .Z(n15894) );
  AOI211_X1 U19045 ( .C1(n19711), .C2(n19621), .A(n15895), .B(n15894), .ZN(
        n15896) );
  OAI21_X1 U19046 ( .B1(n19627), .B2(n15927), .A(n15896), .ZN(P2_U2851) );
  AOI22_X1 U19047 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19605), .B1(n15934), 
        .B2(P2_EBX_REG_3__SCAN_IN), .ZN(n15897) );
  OAI21_X1 U19048 ( .B1(n15898), .B2(n19625), .A(n15897), .ZN(n15899) );
  AOI21_X1 U19049 ( .B1(n15900), .B2(n19609), .A(n15899), .ZN(n15901) );
  OAI21_X1 U19050 ( .B1(n16148), .B2(n19611), .A(n15901), .ZN(n15908) );
  INV_X1 U19051 ( .A(n15903), .ZN(n15902) );
  OAI21_X1 U19052 ( .B1(n15914), .B2(n15902), .A(n15912), .ZN(n15906) );
  NOR2_X1 U19053 ( .A1(n15944), .A2(n15903), .ZN(n15905) );
  MUX2_X1 U19054 ( .A(n15906), .B(n15905), .S(n15904), .Z(n15907) );
  AOI211_X1 U19055 ( .C1(n19621), .C2(n15909), .A(n15908), .B(n15907), .ZN(
        n15910) );
  OAI21_X1 U19056 ( .B1(n15911), .B2(n15927), .A(n15910), .ZN(P2_U2852) );
  INV_X1 U19057 ( .A(n15915), .ZN(n15913) );
  OAI21_X1 U19058 ( .B1(n15914), .B2(n15913), .A(n15912), .ZN(n15918) );
  NOR2_X1 U19059 ( .A1(n15944), .A2(n15915), .ZN(n15917) );
  MUX2_X1 U19060 ( .A(n15918), .B(n15917), .S(n15916), .Z(n15929) );
  NAND2_X1 U19061 ( .A1(n20477), .A2(n15933), .ZN(n15924) );
  AOI22_X1 U19062 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n19605), .B1(n15934), 
        .B2(P2_EBX_REG_2__SCAN_IN), .ZN(n15923) );
  NAND2_X1 U19063 ( .A1(n19609), .A2(n15919), .ZN(n15922) );
  OR2_X1 U19064 ( .A1(n19625), .A2(n15920), .ZN(n15921) );
  NAND4_X1 U19065 ( .A1(n15924), .A2(n15923), .A3(n15922), .A4(n15921), .ZN(
        n15925) );
  AOI21_X1 U19066 ( .B1(n10666), .B2(n19621), .A(n15925), .ZN(n15926) );
  OAI21_X1 U19067 ( .B1(n20472), .B2(n15927), .A(n15926), .ZN(n15928) );
  OAI21_X1 U19068 ( .B1(n15931), .B2(n15930), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15942) );
  AOI22_X1 U19069 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(n19605), .B1(n19609), 
        .B2(n15932), .ZN(n15936) );
  AOI22_X1 U19070 ( .A1(n15934), .A2(P2_EBX_REG_0__SCAN_IN), .B1(n15933), .B2(
        n19651), .ZN(n15935) );
  OAI211_X1 U19071 ( .C1(n15938), .C2(n15937), .A(n15936), .B(n15935), .ZN(
        n15939) );
  AOI21_X1 U19072 ( .B1(n19652), .B2(n15940), .A(n15939), .ZN(n15941) );
  OAI211_X1 U19073 ( .C1(n15944), .C2(n15943), .A(n15942), .B(n15941), .ZN(
        P2_U2855) );
  NAND2_X1 U19074 ( .A1(n16043), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n15945) );
  OAI21_X1 U19075 ( .B1(n15946), .B2(n16043), .A(n15945), .ZN(P2_U2856) );
  OR2_X1 U19076 ( .A1(n15948), .A2(n15947), .ZN(n16046) );
  NAND3_X1 U19077 ( .A1(n16046), .A2(n16045), .A3(n16037), .ZN(n15950) );
  NAND2_X1 U19078 ( .A1(n16043), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15949) );
  OAI211_X1 U19079 ( .C1(n16166), .C2(n16043), .A(n15950), .B(n15949), .ZN(
        P2_U2858) );
  NOR2_X1 U19080 ( .A1(n15952), .A2(n15951), .ZN(n15954) );
  XNOR2_X1 U19081 ( .A(n15954), .B(n15953), .ZN(n16061) );
  NOR2_X1 U19082 ( .A1(n15955), .A2(n16043), .ZN(n15956) );
  AOI21_X1 U19083 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16043), .A(n15956), .ZN(
        n15957) );
  OAI21_X1 U19084 ( .B1(n16061), .B2(n16029), .A(n15957), .ZN(P2_U2859) );
  OAI21_X1 U19085 ( .B1(n15960), .B2(n15959), .A(n15958), .ZN(n16068) );
  NOR2_X1 U19086 ( .A1(n16447), .A2(n16043), .ZN(n15961) );
  AOI21_X1 U19087 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n16043), .A(n15961), .ZN(
        n15962) );
  OAI21_X1 U19088 ( .B1(n16068), .B2(n16029), .A(n15962), .ZN(P2_U2860) );
  NOR2_X1 U19089 ( .A1(n15973), .A2(n15972), .ZN(n15971) );
  NOR2_X1 U19090 ( .A1(n15971), .A2(n15963), .ZN(n15968) );
  NOR2_X1 U19091 ( .A1(n15978), .A2(n15964), .ZN(n15965) );
  XNOR2_X1 U19092 ( .A(n15966), .B(n15965), .ZN(n15967) );
  XNOR2_X1 U19093 ( .A(n15968), .B(n15967), .ZN(n16074) );
  NOR2_X1 U19094 ( .A1(n16459), .A2(n16043), .ZN(n15969) );
  AOI21_X1 U19095 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n16043), .A(n15969), .ZN(
        n15970) );
  OAI21_X1 U19096 ( .B1(n16074), .B2(n16029), .A(n15970), .ZN(P2_U2861) );
  AOI21_X1 U19097 ( .B1(n15973), .B2(n15972), .A(n15971), .ZN(n16075) );
  NAND2_X1 U19098 ( .A1(n16075), .A2(n16037), .ZN(n15975) );
  NAND2_X1 U19099 ( .A1(n16043), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15974) );
  OAI211_X1 U19100 ( .C1(n16192), .C2(n16043), .A(n15975), .B(n15974), .ZN(
        P2_U2862) );
  INV_X1 U19101 ( .A(n15976), .ZN(n15992) );
  XNOR2_X1 U19102 ( .A(n15976), .B(n15979), .ZN(n15988) );
  NOR2_X1 U19103 ( .A1(n15978), .A2(n15977), .ZN(n15987) );
  NAND2_X1 U19104 ( .A1(n15988), .A2(n15987), .ZN(n15986) );
  OAI21_X1 U19105 ( .B1(n15992), .B2(n15979), .A(n15986), .ZN(n15983) );
  XOR2_X1 U19106 ( .A(n15981), .B(n15980), .Z(n15982) );
  XNOR2_X1 U19107 ( .A(n15983), .B(n15982), .ZN(n16088) );
  NOR2_X1 U19108 ( .A1(n16486), .A2(n16043), .ZN(n15984) );
  AOI21_X1 U19109 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n16043), .A(n15984), .ZN(
        n15985) );
  OAI21_X1 U19110 ( .B1(n16088), .B2(n16029), .A(n15985), .ZN(P2_U2863) );
  OAI21_X1 U19111 ( .B1(n15988), .B2(n15987), .A(n15986), .ZN(n16094) );
  NOR2_X1 U19112 ( .A1(n16496), .A2(n16043), .ZN(n15989) );
  AOI21_X1 U19113 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n16043), .A(n15989), .ZN(
        n15990) );
  OAI21_X1 U19114 ( .B1(n16029), .B2(n16094), .A(n15990), .ZN(P2_U2864) );
  OAI21_X1 U19115 ( .B1(n15991), .B2(n15993), .A(n15992), .ZN(n16100) );
  NOR2_X1 U19116 ( .A1(n16510), .A2(n16043), .ZN(n15994) );
  AOI21_X1 U19117 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n16043), .A(n15994), .ZN(
        n15995) );
  OAI21_X1 U19118 ( .B1(n16029), .B2(n16100), .A(n15995), .ZN(P2_U2865) );
  INV_X1 U19119 ( .A(n15991), .ZN(n15997) );
  OAI21_X1 U19120 ( .B1(n15996), .B2(n15998), .A(n15997), .ZN(n16107) );
  MUX2_X1 U19121 ( .A(n16001), .B(n16000), .S(n15999), .Z(n16002) );
  OAI21_X1 U19122 ( .B1(n16029), .B2(n16107), .A(n16002), .ZN(P2_U2866) );
  NOR2_X1 U19123 ( .A1(n16003), .A2(n16004), .ZN(n16005) );
  OR2_X1 U19124 ( .A1(n15996), .A2(n16005), .ZN(n16114) );
  NOR2_X1 U19125 ( .A1(n16519), .A2(n16043), .ZN(n16006) );
  AOI21_X1 U19126 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n16043), .A(n16006), .ZN(
        n16007) );
  OAI21_X1 U19127 ( .B1(n16029), .B2(n16114), .A(n16007), .ZN(P2_U2867) );
  AND2_X1 U19128 ( .A1(n16008), .A2(n16009), .ZN(n16010) );
  NOR2_X1 U19129 ( .A1(n16003), .A2(n16010), .ZN(n16115) );
  NAND2_X1 U19130 ( .A1(n16115), .A2(n16037), .ZN(n16012) );
  NAND2_X1 U19131 ( .A1(n16043), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n16011) );
  OAI211_X1 U19132 ( .C1(n16538), .C2(n16043), .A(n16012), .B(n16011), .ZN(
        P2_U2868) );
  OAI21_X1 U19133 ( .B1(n14414), .B2(n16014), .A(n16008), .ZN(n16126) );
  NOR2_X1 U19134 ( .A1(n16552), .A2(n16043), .ZN(n16015) );
  AOI21_X1 U19135 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n16043), .A(n16015), .ZN(
        n16016) );
  OAI21_X1 U19136 ( .B1(n16029), .B2(n16126), .A(n16016), .ZN(P2_U2869) );
  OAI21_X1 U19137 ( .B1(n16023), .B2(n16017), .A(n16013), .ZN(n16134) );
  NOR2_X1 U19138 ( .A1(n16018), .A2(n16043), .ZN(n16019) );
  AOI21_X1 U19139 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n16043), .A(n16019), .ZN(
        n16020) );
  OAI21_X1 U19140 ( .B1(n16029), .B2(n16134), .A(n16020), .ZN(P2_U2870) );
  NAND2_X1 U19141 ( .A1(n16040), .A2(n16039), .ZN(n16038) );
  INV_X1 U19142 ( .A(n16033), .ZN(n16021) );
  AOI21_X1 U19143 ( .B1(n16031), .B2(n16027), .A(n16022), .ZN(n16024) );
  NOR2_X1 U19144 ( .A1(n16024), .A2(n16023), .ZN(n16135) );
  NAND2_X1 U19145 ( .A1(n16135), .A2(n16037), .ZN(n16026) );
  NAND2_X1 U19146 ( .A1(n16043), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n16025) );
  OAI211_X1 U19147 ( .C1(n16563), .C2(n16043), .A(n16026), .B(n16025), .ZN(
        P2_U2871) );
  XNOR2_X1 U19148 ( .A(n16031), .B(n16027), .ZN(n16030) );
  MUX2_X1 U19149 ( .A(n16576), .B(n11097), .S(n16043), .Z(n16028) );
  OAI21_X1 U19150 ( .B1(n16030), .B2(n16029), .A(n16028), .ZN(P2_U2872) );
  INV_X1 U19151 ( .A(n16038), .ZN(n16034) );
  INV_X1 U19152 ( .A(n16031), .ZN(n16032) );
  OAI211_X1 U19153 ( .C1(n16034), .C2(n16033), .A(n16032), .B(n16037), .ZN(
        n16036) );
  NAND2_X1 U19154 ( .A1(n16043), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n16035) );
  OAI211_X1 U19155 ( .C1(n16581), .C2(n16043), .A(n16036), .B(n16035), .ZN(
        P2_U2873) );
  OAI211_X1 U19156 ( .C1(n16040), .C2(n16039), .A(n16038), .B(n16037), .ZN(
        n16042) );
  NAND2_X1 U19157 ( .A1(n16043), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n16041) );
  OAI211_X1 U19158 ( .C1(n16044), .C2(n16043), .A(n16042), .B(n16041), .ZN(
        P2_U2874) );
  NAND3_X1 U19159 ( .A1(n16046), .A2(n16045), .A3(n19649), .ZN(n16053) );
  AOI22_X1 U19160 ( .A1(n16137), .A2(n16047), .B1(n19647), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n16048) );
  OAI21_X1 U19161 ( .B1(n16140), .B2(n16049), .A(n16048), .ZN(n16051) );
  NOR2_X1 U19162 ( .A1(n16438), .A2(n16056), .ZN(n16050) );
  AOI211_X1 U19163 ( .C1(n16136), .C2(BUF2_REG_29__SCAN_IN), .A(n16051), .B(
        n16050), .ZN(n16052) );
  NAND2_X1 U19164 ( .A1(n16053), .A2(n16052), .ZN(P2_U2890) );
  AOI22_X1 U19165 ( .A1(n16137), .A2(n16054), .B1(n19647), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n16055) );
  OAI21_X1 U19166 ( .B1(n16140), .B2(n17437), .A(n16055), .ZN(n16059) );
  NOR2_X1 U19167 ( .A1(n16057), .A2(n16056), .ZN(n16058) );
  AOI211_X1 U19168 ( .C1(n16136), .C2(BUF2_REG_28__SCAN_IN), .A(n16059), .B(
        n16058), .ZN(n16060) );
  OAI21_X1 U19169 ( .B1(n16061), .B2(n16144), .A(n16060), .ZN(P2_U2891) );
  INV_X1 U19170 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16065) );
  NAND2_X1 U19171 ( .A1(n16136), .A2(BUF2_REG_27__SCAN_IN), .ZN(n16064) );
  AOI22_X1 U19172 ( .A1(n16137), .A2(n16062), .B1(n19647), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n16063) );
  OAI211_X1 U19173 ( .C1(n16140), .C2(n16065), .A(n16064), .B(n16063), .ZN(
        n16066) );
  AOI21_X1 U19174 ( .B1(n10453), .B2(n19648), .A(n16066), .ZN(n16067) );
  OAI21_X1 U19175 ( .B1(n16068), .B2(n16144), .A(n16067), .ZN(P2_U2892) );
  NAND2_X1 U19176 ( .A1(n16136), .A2(BUF2_REG_26__SCAN_IN), .ZN(n16071) );
  AOI22_X1 U19177 ( .A1(n16137), .A2(n16069), .B1(n19647), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n16070) );
  OAI211_X1 U19178 ( .C1(n16140), .C2(n17440), .A(n16071), .B(n16070), .ZN(
        n16072) );
  AOI21_X1 U19179 ( .B1(n10457), .B2(n19648), .A(n16072), .ZN(n16073) );
  OAI21_X1 U19180 ( .B1(n16074), .B2(n16144), .A(n16073), .ZN(P2_U2893) );
  INV_X1 U19181 ( .A(n16075), .ZN(n16082) );
  INV_X1 U19182 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16079) );
  NAND2_X1 U19183 ( .A1(n16136), .A2(BUF2_REG_25__SCAN_IN), .ZN(n16078) );
  AOI22_X1 U19184 ( .A1(n16137), .A2(n16076), .B1(n19647), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n16077) );
  OAI211_X1 U19185 ( .C1(n16140), .C2(n16079), .A(n16078), .B(n16077), .ZN(
        n16080) );
  AOI21_X1 U19186 ( .B1(n16466), .B2(n19648), .A(n16080), .ZN(n16081) );
  OAI21_X1 U19187 ( .B1(n16082), .B2(n16144), .A(n16081), .ZN(P2_U2894) );
  NAND2_X1 U19188 ( .A1(n16136), .A2(BUF2_REG_24__SCAN_IN), .ZN(n16085) );
  AOI22_X1 U19189 ( .A1(n16137), .A2(n16083), .B1(n19647), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n16084) );
  OAI211_X1 U19190 ( .C1(n16140), .C2(n17443), .A(n16085), .B(n16084), .ZN(
        n16086) );
  AOI21_X1 U19191 ( .B1(n16483), .B2(n19648), .A(n16086), .ZN(n16087) );
  OAI21_X1 U19192 ( .B1(n16088), .B2(n16144), .A(n16087), .ZN(P2_U2895) );
  INV_X1 U19193 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16091) );
  NAND2_X1 U19194 ( .A1(n16136), .A2(BUF2_REG_23__SCAN_IN), .ZN(n16090) );
  AOI22_X1 U19195 ( .A1(n16137), .A2(n19810), .B1(n19647), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16089) );
  OAI211_X1 U19196 ( .C1(n16091), .C2(n16140), .A(n16090), .B(n16089), .ZN(
        n16092) );
  AOI21_X1 U19197 ( .B1(n16499), .B2(n19648), .A(n16092), .ZN(n16093) );
  OAI21_X1 U19198 ( .B1(n16144), .B2(n16094), .A(n16093), .ZN(P2_U2896) );
  INV_X1 U19199 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16097) );
  NAND2_X1 U19200 ( .A1(n16136), .A2(BUF2_REG_22__SCAN_IN), .ZN(n16096) );
  AOI22_X1 U19201 ( .A1(n16137), .A2(n19797), .B1(n19647), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16095) );
  OAI211_X1 U19202 ( .C1(n16097), .C2(n16140), .A(n16096), .B(n16095), .ZN(
        n16098) );
  AOI21_X1 U19203 ( .B1(n16513), .B2(n19648), .A(n16098), .ZN(n16099) );
  OAI21_X1 U19204 ( .B1(n16144), .B2(n16100), .A(n16099), .ZN(P2_U2897) );
  INV_X1 U19205 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16103) );
  NAND2_X1 U19206 ( .A1(n16136), .A2(BUF2_REG_21__SCAN_IN), .ZN(n16102) );
  AOI22_X1 U19207 ( .A1(n16137), .A2(n19787), .B1(n19647), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n16101) );
  OAI211_X1 U19208 ( .C1(n16103), .C2(n16140), .A(n16102), .B(n16101), .ZN(
        n16104) );
  AOI21_X1 U19209 ( .B1(n16105), .B2(n19648), .A(n16104), .ZN(n16106) );
  OAI21_X1 U19210 ( .B1(n16144), .B2(n16107), .A(n16106), .ZN(P2_U2898) );
  INV_X1 U19211 ( .A(n16527), .ZN(n16112) );
  NAND2_X1 U19212 ( .A1(n16136), .A2(BUF2_REG_20__SCAN_IN), .ZN(n16109) );
  AOI22_X1 U19213 ( .A1(n16137), .A2(n19779), .B1(n19647), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16108) );
  OAI211_X1 U19214 ( .C1(n16110), .C2(n16140), .A(n16109), .B(n16108), .ZN(
        n16111) );
  AOI21_X1 U19215 ( .B1(n16112), .B2(n19648), .A(n16111), .ZN(n16113) );
  OAI21_X1 U19216 ( .B1(n16144), .B2(n16114), .A(n16113), .ZN(P2_U2899) );
  INV_X1 U19217 ( .A(n16115), .ZN(n16121) );
  INV_X1 U19218 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16118) );
  NAND2_X1 U19219 ( .A1(n16136), .A2(BUF2_REG_19__SCAN_IN), .ZN(n16117) );
  AOI22_X1 U19220 ( .A1(n16137), .A2(n19770), .B1(n19647), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n16116) );
  OAI211_X1 U19221 ( .C1(n16118), .C2(n16140), .A(n16117), .B(n16116), .ZN(
        n16119) );
  AOI21_X1 U19222 ( .B1(n16535), .B2(n19648), .A(n16119), .ZN(n16120) );
  OAI21_X1 U19223 ( .B1(n16144), .B2(n16121), .A(n16120), .ZN(P2_U2900) );
  NAND2_X1 U19224 ( .A1(n16136), .A2(BUF2_REG_18__SCAN_IN), .ZN(n16123) );
  AOI22_X1 U19225 ( .A1(n16137), .A2(n19762), .B1(n19647), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16122) );
  OAI211_X1 U19226 ( .C1(n17450), .C2(n16140), .A(n16123), .B(n16122), .ZN(
        n16124) );
  AOI21_X1 U19227 ( .B1(n16549), .B2(n19648), .A(n16124), .ZN(n16125) );
  OAI21_X1 U19228 ( .B1(n16144), .B2(n16126), .A(n16125), .ZN(P2_U2901) );
  INV_X1 U19229 ( .A(n16127), .ZN(n16132) );
  INV_X1 U19230 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16130) );
  NAND2_X1 U19231 ( .A1(n16136), .A2(BUF2_REG_17__SCAN_IN), .ZN(n16129) );
  AOI22_X1 U19232 ( .A1(n16137), .A2(n16784), .B1(n19647), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n16128) );
  OAI211_X1 U19233 ( .C1(n16130), .C2(n16140), .A(n16129), .B(n16128), .ZN(
        n16131) );
  AOI21_X1 U19234 ( .B1(n16132), .B2(n19648), .A(n16131), .ZN(n16133) );
  OAI21_X1 U19235 ( .B1(n16144), .B2(n16134), .A(n16133), .ZN(P2_U2902) );
  INV_X1 U19236 ( .A(n16135), .ZN(n16145) );
  NAND2_X1 U19237 ( .A1(n16136), .A2(BUF2_REG_16__SCAN_IN), .ZN(n16139) );
  AOI22_X1 U19238 ( .A1(n16137), .A2(n16769), .B1(n19647), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n16138) );
  OAI211_X1 U19239 ( .C1(n16141), .C2(n16140), .A(n16139), .B(n16138), .ZN(
        n16142) );
  AOI21_X1 U19240 ( .B1(n16560), .B2(n19648), .A(n16142), .ZN(n16143) );
  OAI21_X1 U19241 ( .B1(n16145), .B2(n16144), .A(n16143), .ZN(P2_U2903) );
  XNOR2_X1 U19242 ( .A(n15881), .B(n16146), .ZN(n19612) );
  OAI21_X1 U19243 ( .B1(n9823), .B2(n20477), .A(n16147), .ZN(n19634) );
  XNOR2_X1 U19244 ( .A(n20465), .B(n16148), .ZN(n19635) );
  NAND2_X1 U19245 ( .A1(n19634), .A2(n19635), .ZN(n19633) );
  OAI21_X1 U19246 ( .B1(n20469), .B2(n20465), .A(n19633), .ZN(n16149) );
  NAND2_X1 U19247 ( .A1(n16149), .A2(n19626), .ZN(n19628) );
  INV_X1 U19248 ( .A(n19627), .ZN(n16150) );
  NAND3_X1 U19249 ( .A1(n19628), .A2(n16150), .A3(n19649), .ZN(n16155) );
  INV_X1 U19250 ( .A(n19787), .ZN(n16152) );
  INV_X1 U19251 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19684) );
  OAI22_X1 U19252 ( .A1(n19655), .A2(n16152), .B1(n16151), .B2(n19684), .ZN(
        n16153) );
  INV_X1 U19253 ( .A(n16153), .ZN(n16154) );
  OAI211_X1 U19254 ( .C1(n19612), .C2(n16156), .A(n16155), .B(n16154), .ZN(
        P2_U2914) );
  NOR2_X1 U19255 ( .A1(n16451), .A2(n21531), .ZN(n16158) );
  OAI21_X1 U19256 ( .B1(n16158), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16157), .ZN(n16442) );
  NOR2_X1 U19257 ( .A1(n16160), .A2(n16159), .ZN(n16161) );
  XNOR2_X1 U19258 ( .A(n9605), .B(n16161), .ZN(n16440) );
  NOR2_X1 U19259 ( .A1(n19705), .A2(n20441), .ZN(n16434) );
  NOR2_X1 U19260 ( .A1(n16419), .A2(n16162), .ZN(n16163) );
  AOI211_X1 U19261 ( .C1(n16164), .C2(n16425), .A(n16434), .B(n16163), .ZN(
        n16165) );
  OAI21_X1 U19262 ( .B1(n16166), .B2(n16429), .A(n16165), .ZN(n16167) );
  AOI21_X1 U19263 ( .B1(n16394), .B2(n16440), .A(n16167), .ZN(n16168) );
  OAI21_X1 U19264 ( .B1(n16396), .B2(n16442), .A(n16168), .ZN(P2_U2985) );
  XNOR2_X1 U19265 ( .A(n16169), .B(n16173), .ZN(n16454) );
  OR2_X1 U19266 ( .A1(n19705), .A2(n20438), .ZN(n16444) );
  OAI21_X1 U19267 ( .B1(n16419), .B2(n16170), .A(n16444), .ZN(n16172) );
  NOR2_X1 U19268 ( .A1(n16447), .A2(n16429), .ZN(n16171) );
  AOI211_X1 U19269 ( .C1(n16425), .C2(n10274), .A(n16172), .B(n16171), .ZN(
        n16176) );
  INV_X1 U19270 ( .A(n16185), .ZN(n16174) );
  NAND2_X1 U19271 ( .A1(n16174), .A2(n16173), .ZN(n16450) );
  NAND3_X1 U19272 ( .A1(n16451), .A2(n16415), .A3(n16450), .ZN(n16175) );
  OAI211_X1 U19273 ( .C1(n16454), .C2(n16422), .A(n16176), .B(n16175), .ZN(
        P2_U2987) );
  OAI21_X1 U19274 ( .B1(n16177), .B2(n16189), .A(n16190), .ZN(n16178) );
  XOR2_X1 U19275 ( .A(n16179), .B(n16178), .Z(n16465) );
  NAND2_X1 U19276 ( .A1(n19604), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n16455) );
  OAI21_X1 U19277 ( .B1(n16419), .B2(n16180), .A(n16455), .ZN(n16182) );
  NOR2_X1 U19278 ( .A1(n16459), .A2(n16429), .ZN(n16181) );
  AOI211_X1 U19279 ( .C1(n16425), .C2(n16183), .A(n16182), .B(n16181), .ZN(
        n16188) );
  AOI21_X1 U19280 ( .B1(n16186), .B2(n16184), .A(n16185), .ZN(n16462) );
  NAND2_X1 U19281 ( .A1(n16462), .A2(n16415), .ZN(n16187) );
  OAI211_X1 U19282 ( .C1(n16465), .C2(n16422), .A(n16188), .B(n16187), .ZN(
        P2_U2988) );
  NAND2_X1 U19283 ( .A1(n10245), .A2(n16190), .ZN(n16191) );
  XNOR2_X1 U19284 ( .A(n16177), .B(n16191), .ZN(n16478) );
  INV_X1 U19285 ( .A(n16192), .ZN(n16474) );
  INV_X1 U19286 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20433) );
  NOR2_X1 U19287 ( .A1(n19705), .A2(n20433), .ZN(n16467) );
  AOI21_X1 U19288 ( .B1(n16354), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16467), .ZN(n16193) );
  OAI21_X1 U19289 ( .B1(n16194), .B2(n16406), .A(n16193), .ZN(n16195) );
  AOI21_X1 U19290 ( .B1(n16474), .B2(n16409), .A(n16195), .ZN(n16197) );
  INV_X1 U19291 ( .A(n14346), .ZN(n16198) );
  NAND2_X1 U19292 ( .A1(n16198), .A2(n16468), .ZN(n16475) );
  NAND3_X1 U19293 ( .A1(n16475), .A2(n16415), .A3(n16184), .ZN(n16196) );
  OAI211_X1 U19294 ( .C1(n16422), .C2(n16478), .A(n16197), .B(n16196), .ZN(
        P2_U2989) );
  NAND2_X1 U19295 ( .A1(n16199), .A2(n16219), .ZN(n16215) );
  XNOR2_X1 U19296 ( .A(n16200), .B(n16495), .ZN(n16214) );
  NAND2_X1 U19297 ( .A1(n16215), .A2(n16214), .ZN(n16500) );
  OAI21_X1 U19298 ( .B1(n16201), .B2(n16495), .A(n16500), .ZN(n16205) );
  NAND2_X1 U19299 ( .A1(n16203), .A2(n16202), .ZN(n16204) );
  XNOR2_X1 U19300 ( .A(n16205), .B(n16204), .ZN(n16488) );
  NOR2_X1 U19301 ( .A1(n19705), .A2(n20431), .ZN(n16480) );
  NOR2_X1 U19302 ( .A1(n16419), .A2(n16206), .ZN(n16207) );
  AOI211_X1 U19303 ( .C1(n10277), .C2(n16425), .A(n16480), .B(n16207), .ZN(
        n16208) );
  OAI21_X1 U19304 ( .B1(n16486), .B2(n16429), .A(n16208), .ZN(n16209) );
  AOI21_X1 U19305 ( .B1(n16394), .B2(n16488), .A(n16209), .ZN(n16210) );
  OAI21_X1 U19306 ( .B1(n16396), .B2(n16490), .A(n16210), .ZN(P2_U2990) );
  OAI21_X1 U19307 ( .B1(n16226), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16211), .ZN(n16504) );
  INV_X1 U19308 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20429) );
  OR2_X1 U19309 ( .A1(n19705), .A2(n20429), .ZN(n16493) );
  OAI21_X1 U19310 ( .B1(n16419), .B2(n10317), .A(n16493), .ZN(n16213) );
  NOR2_X1 U19311 ( .A1(n16496), .A2(n16429), .ZN(n16212) );
  AOI211_X1 U19312 ( .C1(n9765), .C2(n16425), .A(n16213), .B(n16212), .ZN(
        n16217) );
  OR2_X1 U19313 ( .A1(n16215), .A2(n16214), .ZN(n16501) );
  NAND3_X1 U19314 ( .A1(n16501), .A2(n16394), .A3(n16500), .ZN(n16216) );
  OAI211_X1 U19315 ( .C1(n16504), .C2(n16396), .A(n16217), .B(n16216), .ZN(
        P2_U2991) );
  NAND2_X1 U19316 ( .A1(n16219), .A2(n16218), .ZN(n16220) );
  XOR2_X1 U19317 ( .A(n16220), .B(n9669), .Z(n16518) );
  INV_X1 U19318 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n16221) );
  OR2_X1 U19319 ( .A1(n19705), .A2(n16221), .ZN(n16506) );
  OAI21_X1 U19320 ( .B1(n16419), .B2(n16222), .A(n16506), .ZN(n16224) );
  NOR2_X1 U19321 ( .A1(n16510), .A2(n16429), .ZN(n16223) );
  AOI211_X1 U19322 ( .C1(n16225), .C2(n16425), .A(n16224), .B(n16223), .ZN(
        n16229) );
  NAND2_X1 U19323 ( .A1(n16227), .A2(n16508), .ZN(n16514) );
  NAND3_X1 U19324 ( .A1(n16515), .A2(n16415), .A3(n16514), .ZN(n16228) );
  OAI211_X1 U19325 ( .C1(n16518), .C2(n16422), .A(n16229), .B(n16228), .ZN(
        P2_U2992) );
  NOR2_X1 U19326 ( .A1(n16232), .A2(n16231), .ZN(n16233) );
  XNOR2_X1 U19327 ( .A(n16234), .B(n16233), .ZN(n16532) );
  AOI21_X1 U19328 ( .B1(n21522), .B2(n16248), .A(n16235), .ZN(n16530) );
  INV_X1 U19329 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n16236) );
  NOR2_X1 U19330 ( .A1(n19705), .A2(n16236), .ZN(n16520) );
  AOI21_X1 U19331 ( .B1(n16354), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16520), .ZN(n16239) );
  NAND2_X1 U19332 ( .A1(n16237), .A2(n16425), .ZN(n16238) );
  OAI211_X1 U19333 ( .C1(n16519), .C2(n16429), .A(n16239), .B(n16238), .ZN(
        n16240) );
  AOI21_X1 U19334 ( .B1(n16530), .B2(n16415), .A(n16240), .ZN(n16241) );
  OAI21_X1 U19335 ( .B1(n16532), .B2(n16422), .A(n16241), .ZN(P2_U2994) );
  NAND2_X1 U19336 ( .A1(n16243), .A2(n16242), .ZN(n16247) );
  NOR2_X1 U19337 ( .A1(n16245), .A2(n16244), .ZN(n16246) );
  XOR2_X1 U19338 ( .A(n16247), .B(n16246), .Z(n16542) );
  INV_X1 U19339 ( .A(n16248), .ZN(n16249) );
  AOI21_X1 U19340 ( .B1(n16251), .B2(n16250), .A(n16249), .ZN(n16540) );
  NOR2_X1 U19341 ( .A1(n19705), .A2(n20423), .ZN(n16533) );
  NOR2_X1 U19342 ( .A1(n16252), .A2(n16406), .ZN(n16253) );
  AOI211_X1 U19343 ( .C1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n16354), .A(
        n16533), .B(n16253), .ZN(n16254) );
  OAI21_X1 U19344 ( .B1(n16538), .B2(n16429), .A(n16254), .ZN(n16255) );
  AOI21_X1 U19345 ( .B1(n16540), .B2(n16415), .A(n16255), .ZN(n16256) );
  OAI21_X1 U19346 ( .B1(n16542), .B2(n16422), .A(n16256), .ZN(P2_U2995) );
  NAND2_X1 U19347 ( .A1(n16354), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16257) );
  OAI211_X1 U19348 ( .C1(n16406), .C2(n16259), .A(n16258), .B(n16257), .ZN(
        n16260) );
  AOI21_X1 U19349 ( .B1(n16261), .B2(n16409), .A(n16260), .ZN(n16264) );
  OAI211_X1 U19350 ( .C1(n9567), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16262), .B(n16415), .ZN(n16263) );
  OAI211_X1 U19351 ( .C1(n16265), .C2(n16422), .A(n16264), .B(n16263), .ZN(
        P2_U2997) );
  INV_X1 U19352 ( .A(n16563), .ZN(n16269) );
  INV_X1 U19353 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20418) );
  NOR2_X1 U19354 ( .A1(n19705), .A2(n20418), .ZN(n16559) );
  AOI21_X1 U19355 ( .B1(n16354), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16559), .ZN(n16267) );
  OAI21_X1 U19356 ( .B1(n16406), .B2(n10299), .A(n16267), .ZN(n16268) );
  AOI21_X1 U19357 ( .B1(n16269), .B2(n16409), .A(n16268), .ZN(n16273) );
  NAND2_X1 U19358 ( .A1(n16270), .A2(n16271), .ZN(n16557) );
  NAND3_X1 U19359 ( .A1(n16558), .A2(n16557), .A3(n16394), .ZN(n16272) );
  OAI211_X1 U19360 ( .C1(n16274), .C2(n16396), .A(n16273), .B(n16272), .ZN(
        P2_U2998) );
  NAND2_X1 U19361 ( .A1(n16276), .A2(n16288), .ZN(n16280) );
  NAND2_X1 U19362 ( .A1(n16278), .A2(n16277), .ZN(n16279) );
  XNOR2_X1 U19363 ( .A(n16280), .B(n16279), .ZN(n16578) );
  INV_X1 U19364 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20416) );
  NOR2_X1 U19365 ( .A1(n19705), .A2(n20416), .ZN(n16571) );
  NOR2_X1 U19366 ( .A1(n16406), .A2(n16281), .ZN(n16282) );
  AOI211_X1 U19367 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16354), .A(
        n16571), .B(n16282), .ZN(n16283) );
  OAI21_X1 U19368 ( .B1(n16576), .B2(n16429), .A(n16283), .ZN(n16284) );
  AOI21_X1 U19369 ( .B1(n16578), .B2(n16394), .A(n16284), .ZN(n16285) );
  OAI21_X1 U19370 ( .B1(n16580), .B2(n16396), .A(n16285), .ZN(P2_U2999) );
  NAND2_X1 U19371 ( .A1(n16287), .A2(n16286), .ZN(n16597) );
  NAND2_X1 U19372 ( .A1(n16289), .A2(n16288), .ZN(n16290) );
  XNOR2_X1 U19373 ( .A(n16291), .B(n16290), .ZN(n16594) );
  NAND2_X1 U19374 ( .A1(n19604), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n16584) );
  OAI21_X1 U19375 ( .B1(n16419), .B2(n16292), .A(n16584), .ZN(n16293) );
  AOI21_X1 U19376 ( .B1(n16425), .B2(n16294), .A(n16293), .ZN(n16295) );
  OAI21_X1 U19377 ( .B1(n16581), .B2(n16429), .A(n16295), .ZN(n16296) );
  AOI21_X1 U19378 ( .B1(n16594), .B2(n16394), .A(n16296), .ZN(n16297) );
  OAI21_X1 U19379 ( .B1(n16597), .B2(n16396), .A(n16297), .ZN(P2_U3000) );
  XNOR2_X1 U19380 ( .A(n16615), .B(n16602), .ZN(n16614) );
  NOR2_X1 U19381 ( .A1(n19705), .A2(n20413), .ZN(n16599) );
  AOI21_X1 U19382 ( .B1(n16354), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16599), .ZN(n16298) );
  OAI21_X1 U19383 ( .B1(n16406), .B2(n16299), .A(n16298), .ZN(n16304) );
  NAND2_X1 U19384 ( .A1(n16301), .A2(n16300), .ZN(n16302) );
  NOR2_X1 U19385 ( .A1(n16611), .A2(n16422), .ZN(n16303) );
  AOI211_X1 U19386 ( .C1(n16409), .C2(n16608), .A(n16304), .B(n16303), .ZN(
        n16305) );
  OAI21_X1 U19387 ( .B1(n16614), .B2(n16396), .A(n16305), .ZN(P2_U3001) );
  AND2_X1 U19388 ( .A1(n16307), .A2(n16306), .ZN(n16308) );
  XNOR2_X1 U19389 ( .A(n16309), .B(n16308), .ZN(n16628) );
  INV_X1 U19390 ( .A(n16325), .ZN(n16310) );
  NAND2_X1 U19391 ( .A1(n16310), .A2(n16604), .ZN(n16616) );
  NAND3_X1 U19392 ( .A1(n16616), .A2(n16415), .A3(n16615), .ZN(n16316) );
  NAND2_X1 U19393 ( .A1(n19604), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n16618) );
  OAI21_X1 U19394 ( .B1(n16419), .B2(n16311), .A(n16618), .ZN(n16313) );
  NOR2_X1 U19395 ( .A1(n16617), .A2(n16429), .ZN(n16312) );
  AOI211_X1 U19396 ( .C1(n16314), .C2(n16425), .A(n16313), .B(n16312), .ZN(
        n16315) );
  OAI211_X1 U19397 ( .C1(n16628), .C2(n16422), .A(n16316), .B(n16315), .ZN(
        P2_U3002) );
  NAND2_X1 U19398 ( .A1(n16318), .A2(n16317), .ZN(n16324) );
  NAND2_X1 U19399 ( .A1(n16320), .A2(n16319), .ZN(n16322) );
  NAND2_X1 U19400 ( .A1(n16322), .A2(n16321), .ZN(n16323) );
  XOR2_X1 U19401 ( .A(n16324), .B(n16323), .Z(n16644) );
  NAND2_X1 U19402 ( .A1(n16629), .A2(n16415), .ZN(n16330) );
  INV_X1 U19403 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n20409) );
  NOR2_X1 U19404 ( .A1(n16416), .A2(n20409), .ZN(n16630) );
  AOI21_X1 U19405 ( .B1(n16354), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16630), .ZN(n16326) );
  OAI21_X1 U19406 ( .B1(n16406), .B2(n16327), .A(n16326), .ZN(n16328) );
  AOI21_X1 U19407 ( .B1(n16641), .B2(n16409), .A(n16328), .ZN(n16329) );
  OAI211_X1 U19408 ( .C1(n16644), .C2(n16422), .A(n16330), .B(n16329), .ZN(
        P2_U3003) );
  OAI21_X1 U19409 ( .B1(n16352), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16331), .ZN(n16656) );
  NAND2_X1 U19410 ( .A1(n16333), .A2(n16332), .ZN(n16382) );
  INV_X1 U19411 ( .A(n16334), .ZN(n16336) );
  OAI21_X1 U19412 ( .B1(n16382), .B2(n16336), .A(n16335), .ZN(n16351) );
  INV_X1 U19413 ( .A(n16349), .ZN(n16337) );
  OAI21_X1 U19414 ( .B1(n16351), .B2(n16337), .A(n16348), .ZN(n16341) );
  NAND2_X1 U19415 ( .A1(n16339), .A2(n16338), .ZN(n16340) );
  XNOR2_X1 U19416 ( .A(n16341), .B(n16340), .ZN(n16653) );
  NOR2_X1 U19417 ( .A1(n16342), .A2(n16429), .ZN(n16346) );
  NAND2_X1 U19418 ( .A1(n19604), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n16646) );
  NAND2_X1 U19419 ( .A1(n16354), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16343) );
  OAI211_X1 U19420 ( .C1(n16406), .C2(n16344), .A(n16646), .B(n16343), .ZN(
        n16345) );
  AOI211_X1 U19421 ( .C1(n16653), .C2(n16394), .A(n16346), .B(n16345), .ZN(
        n16347) );
  OAI21_X1 U19422 ( .B1(n16656), .B2(n16396), .A(n16347), .ZN(P2_U3004) );
  NAND2_X1 U19423 ( .A1(n16349), .A2(n16348), .ZN(n16350) );
  XNOR2_X1 U19424 ( .A(n16351), .B(n16350), .ZN(n16668) );
  AOI21_X1 U19425 ( .B1(n16353), .B2(n16636), .A(n16352), .ZN(n16657) );
  NAND2_X1 U19426 ( .A1(n16657), .A2(n16415), .ZN(n16360) );
  NAND2_X1 U19427 ( .A1(n19604), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n16660) );
  NAND2_X1 U19428 ( .A1(n16354), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16355) );
  OAI211_X1 U19429 ( .C1(n16406), .C2(n16356), .A(n16660), .B(n16355), .ZN(
        n16357) );
  AOI21_X1 U19430 ( .B1(n16358), .B2(n16409), .A(n16357), .ZN(n16359) );
  OAI211_X1 U19431 ( .C1(n16422), .C2(n16668), .A(n16360), .B(n16359), .ZN(
        P2_U3005) );
  INV_X1 U19432 ( .A(n16381), .ZN(n16361) );
  AOI21_X1 U19433 ( .B1(n16382), .B2(n16380), .A(n16361), .ZN(n16365) );
  NAND2_X1 U19434 ( .A1(n16363), .A2(n16362), .ZN(n16364) );
  XNOR2_X1 U19435 ( .A(n16365), .B(n16364), .ZN(n16682) );
  NAND3_X1 U19436 ( .A1(n16670), .A2(n16669), .A3(n16415), .ZN(n16374) );
  NAND2_X1 U19437 ( .A1(n19604), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n16671) );
  OAI21_X1 U19438 ( .B1(n16419), .B2(n16368), .A(n16671), .ZN(n16371) );
  NOR2_X1 U19439 ( .A1(n16369), .A2(n16429), .ZN(n16370) );
  AOI211_X1 U19440 ( .C1(n16372), .C2(n16425), .A(n16371), .B(n16370), .ZN(
        n16373) );
  OAI211_X1 U19441 ( .C1(n16682), .C2(n16422), .A(n16374), .B(n16373), .ZN(
        P2_U3006) );
  XNOR2_X1 U19442 ( .A(n16376), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16377) );
  XNOR2_X1 U19443 ( .A(n16375), .B(n16377), .ZN(n16695) );
  NAND2_X1 U19444 ( .A1(n16425), .A2(n16378), .ZN(n16379) );
  NAND2_X1 U19445 ( .A1(n19604), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n16685) );
  OAI211_X1 U19446 ( .C1(n15861), .C2(n16419), .A(n16379), .B(n16685), .ZN(
        n16385) );
  NAND2_X1 U19447 ( .A1(n16381), .A2(n16380), .ZN(n16383) );
  XOR2_X1 U19448 ( .A(n16383), .B(n16382), .Z(n16692) );
  NOR2_X1 U19449 ( .A1(n16692), .A2(n16422), .ZN(n16384) );
  AOI211_X1 U19450 ( .C1(n16409), .C2(n16691), .A(n16385), .B(n16384), .ZN(
        n16386) );
  OAI21_X1 U19451 ( .B1(n16695), .B2(n16396), .A(n16386), .ZN(P2_U3007) );
  XNOR2_X1 U19452 ( .A(n16387), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16711) );
  XOR2_X1 U19453 ( .A(n16389), .B(n16388), .Z(n16707) );
  NAND2_X1 U19454 ( .A1(n19604), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n16699) );
  OAI21_X1 U19455 ( .B1(n16419), .B2(n10302), .A(n16699), .ZN(n16390) );
  AOI21_X1 U19456 ( .B1(n16425), .B2(n16391), .A(n16390), .ZN(n16392) );
  OAI21_X1 U19457 ( .B1(n16704), .B2(n16429), .A(n16392), .ZN(n16393) );
  AOI21_X1 U19458 ( .B1(n16707), .B2(n16394), .A(n16393), .ZN(n16395) );
  OAI21_X1 U19459 ( .B1(n16711), .B2(n16396), .A(n16395), .ZN(P2_U3008) );
  OAI21_X1 U19460 ( .B1(n16397), .B2(n11025), .A(n19603), .ZN(n16400) );
  XNOR2_X1 U19461 ( .A(n16398), .B(n16717), .ZN(n16399) );
  XNOR2_X1 U19462 ( .A(n16400), .B(n16399), .ZN(n16726) );
  NOR2_X1 U19463 ( .A1(n16404), .A2(n16403), .ZN(n16405) );
  XNOR2_X1 U19464 ( .A(n16401), .B(n16405), .ZN(n16712) );
  NAND2_X1 U19465 ( .A1(n16712), .A2(n16415), .ZN(n16411) );
  NOR2_X1 U19466 ( .A1(n16406), .A2(n19615), .ZN(n16408) );
  NAND2_X1 U19467 ( .A1(n19604), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n16720) );
  OAI21_X1 U19468 ( .B1(n16419), .B2(n12624), .A(n16720), .ZN(n16407) );
  AOI211_X1 U19469 ( .C1(n19622), .C2(n16409), .A(n16408), .B(n16407), .ZN(
        n16410) );
  OAI211_X1 U19470 ( .C1(n16422), .C2(n16726), .A(n16411), .B(n16410), .ZN(
        P2_U3009) );
  XNOR2_X1 U19471 ( .A(n16412), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n16413) );
  XNOR2_X1 U19472 ( .A(n16414), .B(n16413), .ZN(n19713) );
  NAND2_X1 U19473 ( .A1(n19713), .A2(n16415), .ZN(n16428) );
  INV_X1 U19474 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n16417) );
  OAI22_X1 U19475 ( .A1(n16419), .A2(n16418), .B1(n16417), .B2(n16416), .ZN(
        n16424) );
  XNOR2_X1 U19476 ( .A(n16421), .B(n16420), .ZN(n19707) );
  NOR2_X1 U19477 ( .A1(n19707), .A2(n16422), .ZN(n16423) );
  AOI211_X1 U19478 ( .C1(n16426), .C2(n16425), .A(n16424), .B(n16423), .ZN(
        n16427) );
  OAI211_X1 U19479 ( .C1(n16430), .C2(n16429), .A(n16428), .B(n16427), .ZN(
        P2_U3010) );
  NAND2_X1 U19480 ( .A1(n16431), .A2(n19712), .ZN(n16437) );
  NOR3_X1 U19481 ( .A1(n16446), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n9941), .ZN(n16433) );
  AOI211_X1 U19482 ( .C1(n16435), .C2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16434), .B(n16433), .ZN(n16436) );
  OAI211_X1 U19483 ( .C1(n16722), .C2(n16438), .A(n16437), .B(n16436), .ZN(
        n16439) );
  AOI21_X1 U19484 ( .B1(n19726), .B2(n16440), .A(n16439), .ZN(n16441) );
  OAI21_X1 U19485 ( .B1(n16710), .B2(n16442), .A(n16441), .ZN(P2_U3017) );
  NAND2_X1 U19486 ( .A1(n16443), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16445) );
  OAI211_X1 U19487 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n16446), .A(
        n16445), .B(n16444), .ZN(n16449) );
  NOR2_X1 U19488 ( .A1(n16447), .A2(n19728), .ZN(n16448) );
  AOI211_X1 U19489 ( .C1(n16731), .C2(n10453), .A(n16449), .B(n16448), .ZN(
        n16453) );
  NAND3_X1 U19490 ( .A1(n16451), .A2(n19721), .A3(n16450), .ZN(n16452) );
  OAI211_X1 U19491 ( .C1(n16454), .C2(n19706), .A(n16453), .B(n16452), .ZN(
        P2_U3019) );
  XNOR2_X1 U19492 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16457) );
  NAND3_X1 U19493 ( .A1(n16482), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n16713), .ZN(n16456) );
  OAI211_X1 U19494 ( .C1(n16458), .C2(n16457), .A(n16456), .B(n16455), .ZN(
        n16461) );
  NOR2_X1 U19495 ( .A1(n16459), .A2(n19728), .ZN(n16460) );
  AOI211_X1 U19496 ( .C1(n16731), .C2(n10457), .A(n16461), .B(n16460), .ZN(
        n16464) );
  NAND2_X1 U19497 ( .A1(n16462), .A2(n19721), .ZN(n16463) );
  OAI211_X1 U19498 ( .C1(n16465), .C2(n19706), .A(n16464), .B(n16463), .ZN(
        P2_U3020) );
  INV_X1 U19499 ( .A(n16466), .ZN(n16472) );
  AOI21_X1 U19500 ( .B1(n16469), .B2(n16468), .A(n16467), .ZN(n16471) );
  NAND3_X1 U19501 ( .A1(n16482), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n16713), .ZN(n16470) );
  OAI211_X1 U19502 ( .C1(n16472), .C2(n16722), .A(n16471), .B(n16470), .ZN(
        n16473) );
  AOI21_X1 U19503 ( .B1(n16474), .B2(n19712), .A(n16473), .ZN(n16477) );
  NAND3_X1 U19504 ( .A1(n16475), .A2(n19721), .A3(n16184), .ZN(n16476) );
  OAI211_X1 U19505 ( .C1(n16478), .C2(n19706), .A(n16477), .B(n16476), .ZN(
        P2_U3021) );
  OAI21_X1 U19506 ( .B1(n16491), .B2(n16492), .A(n16479), .ZN(n16481) );
  AOI21_X1 U19507 ( .B1(n16482), .B2(n16481), .A(n16480), .ZN(n16485) );
  NAND2_X1 U19508 ( .A1(n16483), .A2(n16731), .ZN(n16484) );
  OAI211_X1 U19509 ( .C1(n16486), .C2(n19728), .A(n16485), .B(n16484), .ZN(
        n16487) );
  AOI21_X1 U19510 ( .B1(n19726), .B2(n16488), .A(n16487), .ZN(n16489) );
  OAI21_X1 U19511 ( .B1(n16710), .B2(n16490), .A(n16489), .ZN(P2_U3022) );
  INV_X1 U19512 ( .A(n16491), .ZN(n16505) );
  OAI211_X1 U19513 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16505), .B(n16492), .ZN(
        n16494) );
  OAI211_X1 U19514 ( .C1(n16509), .C2(n16495), .A(n16494), .B(n16493), .ZN(
        n16498) );
  NOR2_X1 U19515 ( .A1(n16496), .A2(n19728), .ZN(n16497) );
  AOI211_X1 U19516 ( .C1(n19724), .C2(n16499), .A(n16498), .B(n16497), .ZN(
        n16503) );
  NAND3_X1 U19517 ( .A1(n16501), .A2(n19726), .A3(n16500), .ZN(n16502) );
  OAI211_X1 U19518 ( .C1(n16504), .C2(n16710), .A(n16503), .B(n16502), .ZN(
        P2_U3023) );
  NAND2_X1 U19519 ( .A1(n16505), .A2(n16508), .ZN(n16507) );
  OAI211_X1 U19520 ( .C1(n16509), .C2(n16508), .A(n16507), .B(n16506), .ZN(
        n16512) );
  NOR2_X1 U19521 ( .A1(n16510), .A2(n19728), .ZN(n16511) );
  AOI211_X1 U19522 ( .C1(n16731), .C2(n16513), .A(n16512), .B(n16511), .ZN(
        n16517) );
  NAND3_X1 U19523 ( .A1(n16515), .A2(n19721), .A3(n16514), .ZN(n16516) );
  OAI211_X1 U19524 ( .C1(n16518), .C2(n19706), .A(n16517), .B(n16516), .ZN(
        P2_U3024) );
  NOR2_X1 U19525 ( .A1(n16519), .A2(n19728), .ZN(n16529) );
  NOR2_X1 U19526 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n16662), .ZN(
        n16521) );
  AOI21_X1 U19527 ( .B1(n16522), .B2(n16521), .A(n16520), .ZN(n16526) );
  OAI21_X1 U19528 ( .B1(n16523), .B2(n17413), .A(n16635), .ZN(n16548) );
  NOR3_X1 U19529 ( .A1(n16524), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n16662), .ZN(n16534) );
  OAI21_X1 U19530 ( .B1(n16548), .B2(n16534), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16525) );
  OAI211_X1 U19531 ( .C1(n16527), .C2(n16722), .A(n16526), .B(n16525), .ZN(
        n16528) );
  AOI211_X1 U19532 ( .C1(n16530), .C2(n19721), .A(n16529), .B(n16528), .ZN(
        n16531) );
  OAI21_X1 U19533 ( .B1(n16532), .B2(n19706), .A(n16531), .ZN(P2_U3026) );
  AOI211_X1 U19534 ( .C1(n16548), .C2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n16534), .B(n16533), .ZN(n16537) );
  NAND2_X1 U19535 ( .A1(n16535), .A2(n19724), .ZN(n16536) );
  OAI211_X1 U19536 ( .C1(n16538), .C2(n19728), .A(n16537), .B(n16536), .ZN(
        n16539) );
  AOI21_X1 U19537 ( .B1(n16540), .B2(n19721), .A(n16539), .ZN(n16541) );
  OAI21_X1 U19538 ( .B1(n16542), .B2(n19706), .A(n16541), .ZN(P2_U3027) );
  AND4_X1 U19539 ( .A1(n16545), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n16544), .A4(n16543), .ZN(n16546) );
  AOI211_X1 U19540 ( .C1(n16548), .C2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16547), .B(n16546), .ZN(n16551) );
  NAND2_X1 U19541 ( .A1(n16549), .A2(n19724), .ZN(n16550) );
  OAI211_X1 U19542 ( .C1(n16552), .C2(n19728), .A(n16551), .B(n16550), .ZN(
        n16553) );
  INV_X1 U19543 ( .A(n16556), .ZN(n16565) );
  NAND3_X1 U19544 ( .A1(n16558), .A2(n16557), .A3(n19726), .ZN(n16562) );
  AOI21_X1 U19545 ( .B1(n16560), .B2(n19724), .A(n16559), .ZN(n16561) );
  OAI211_X1 U19546 ( .C1(n16563), .C2(n19728), .A(n16562), .B(n16561), .ZN(
        n16564) );
  AOI21_X1 U19547 ( .B1(n16565), .B2(n16567), .A(n16564), .ZN(n16566) );
  OAI21_X1 U19548 ( .B1(n16568), .B2(n16567), .A(n16566), .ZN(P2_U3030) );
  NOR2_X1 U19549 ( .A1(n16569), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16570) );
  AOI211_X1 U19550 ( .C1(n16572), .C2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16571), .B(n16570), .ZN(n16575) );
  NAND2_X1 U19551 ( .A1(n16573), .A2(n16731), .ZN(n16574) );
  OAI211_X1 U19552 ( .C1(n16576), .C2(n19728), .A(n16575), .B(n16574), .ZN(
        n16577) );
  AOI21_X1 U19553 ( .B1(n16578), .B2(n19726), .A(n16577), .ZN(n16579) );
  OAI21_X1 U19554 ( .B1(n16580), .B2(n16710), .A(n16579), .ZN(P2_U3031) );
  INV_X1 U19555 ( .A(n16581), .ZN(n16593) );
  NAND3_X1 U19556 ( .A1(n16582), .A2(n16637), .A3(n16590), .ZN(n16583) );
  OAI211_X1 U19557 ( .C1(n16585), .C2(n16722), .A(n16584), .B(n16583), .ZN(
        n16592) );
  NOR2_X1 U19558 ( .A1(n16589), .A2(n16662), .ZN(n16586) );
  NAND2_X1 U19559 ( .A1(n16586), .A2(n16602), .ZN(n16605) );
  NAND2_X1 U19560 ( .A1(n16733), .A2(n16589), .ZN(n16587) );
  NAND2_X1 U19561 ( .A1(n16635), .A2(n16587), .ZN(n16621) );
  NAND2_X1 U19562 ( .A1(n16604), .A2(n16637), .ZN(n16588) );
  NOR2_X1 U19563 ( .A1(n16589), .A2(n16588), .ZN(n16620) );
  NOR2_X1 U19564 ( .A1(n16621), .A2(n16620), .ZN(n16603) );
  AOI21_X1 U19565 ( .B1(n16605), .B2(n16603), .A(n16590), .ZN(n16591) );
  AOI211_X1 U19566 ( .C1(n16593), .C2(n19712), .A(n16592), .B(n16591), .ZN(
        n16596) );
  NAND2_X1 U19567 ( .A1(n16594), .A2(n19726), .ZN(n16595) );
  OAI211_X1 U19568 ( .C1(n16597), .C2(n16710), .A(n16596), .B(n16595), .ZN(
        P2_U3032) );
  NAND2_X1 U19569 ( .A1(n16598), .A2(n19724), .ZN(n16601) );
  INV_X1 U19570 ( .A(n16599), .ZN(n16600) );
  OAI211_X1 U19571 ( .C1(n16603), .C2(n16602), .A(n16601), .B(n16600), .ZN(
        n16607) );
  NOR2_X1 U19572 ( .A1(n16605), .A2(n16604), .ZN(n16606) );
  NOR2_X1 U19573 ( .A1(n16607), .A2(n16606), .ZN(n16610) );
  NAND2_X1 U19574 ( .A1(n16608), .A2(n19712), .ZN(n16609) );
  OAI211_X1 U19575 ( .C1(n16611), .C2(n19706), .A(n16610), .B(n16609), .ZN(
        n16612) );
  INV_X1 U19576 ( .A(n16612), .ZN(n16613) );
  OAI21_X1 U19577 ( .B1(n16614), .B2(n16710), .A(n16613), .ZN(P2_U3033) );
  NAND3_X1 U19578 ( .A1(n16616), .A2(n19721), .A3(n16615), .ZN(n16627) );
  INV_X1 U19579 ( .A(n16617), .ZN(n16625) );
  INV_X1 U19580 ( .A(n16618), .ZN(n16619) );
  AOI211_X1 U19581 ( .C1(n16621), .C2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n16620), .B(n16619), .ZN(n16622) );
  OAI21_X1 U19582 ( .B1(n16722), .B2(n16623), .A(n16622), .ZN(n16624) );
  AOI21_X1 U19583 ( .B1(n19712), .B2(n16625), .A(n16624), .ZN(n16626) );
  OAI211_X1 U19584 ( .C1(n16628), .C2(n19706), .A(n16627), .B(n16626), .ZN(
        P2_U3034) );
  NAND2_X1 U19585 ( .A1(n16629), .A2(n19721), .ZN(n16643) );
  INV_X1 U19586 ( .A(n16630), .ZN(n16633) );
  NAND3_X1 U19587 ( .A1(n16631), .A2(n16637), .A3(n16638), .ZN(n16632) );
  OAI211_X1 U19588 ( .C1(n16634), .C2(n16722), .A(n16633), .B(n16632), .ZN(
        n16640) );
  INV_X1 U19589 ( .A(n16635), .ZN(n16665) );
  AOI21_X1 U19590 ( .B1(n16636), .B2(n16733), .A(n16665), .ZN(n16649) );
  NAND3_X1 U19591 ( .A1(n16648), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n16637), .ZN(n16645) );
  AOI21_X1 U19592 ( .B1(n16649), .B2(n16645), .A(n16638), .ZN(n16639) );
  AOI211_X1 U19593 ( .C1(n16641), .C2(n19712), .A(n16640), .B(n16639), .ZN(
        n16642) );
  OAI211_X1 U19594 ( .C1(n16644), .C2(n19706), .A(n16643), .B(n16642), .ZN(
        P2_U3035) );
  OAI211_X1 U19595 ( .C1(n16647), .C2(n16722), .A(n16646), .B(n16645), .ZN(
        n16651) );
  NOR2_X1 U19596 ( .A1(n16649), .A2(n16648), .ZN(n16650) );
  AOI211_X1 U19597 ( .C1(n16652), .C2(n19712), .A(n16651), .B(n16650), .ZN(
        n16655) );
  NAND2_X1 U19598 ( .A1(n16653), .A2(n19726), .ZN(n16654) );
  OAI211_X1 U19599 ( .C1(n16656), .C2(n16710), .A(n16655), .B(n16654), .ZN(
        P2_U3036) );
  NAND2_X1 U19600 ( .A1(n16657), .A2(n19721), .ZN(n16667) );
  NOR2_X1 U19601 ( .A1(n16658), .A2(n19728), .ZN(n16664) );
  NAND2_X1 U19602 ( .A1(n16659), .A2(n19724), .ZN(n16661) );
  OAI211_X1 U19603 ( .C1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n16662), .A(
        n16661), .B(n16660), .ZN(n16663) );
  AOI211_X1 U19604 ( .C1(n16665), .C2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16664), .B(n16663), .ZN(n16666) );
  OAI211_X1 U19605 ( .C1(n16668), .C2(n19706), .A(n16667), .B(n16666), .ZN(
        P2_U3037) );
  NAND3_X1 U19606 ( .A1(n16670), .A2(n16669), .A3(n19721), .ZN(n16681) );
  OAI21_X1 U19607 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16683), .ZN(n16672) );
  OAI21_X1 U19608 ( .B1(n16673), .B2(n16672), .A(n16671), .ZN(n16674) );
  AOI21_X1 U19609 ( .B1(n16675), .B2(n19724), .A(n16674), .ZN(n16676) );
  OAI21_X1 U19610 ( .B1(n16688), .B2(n16677), .A(n16676), .ZN(n16678) );
  AOI21_X1 U19611 ( .B1(n19712), .B2(n16679), .A(n16678), .ZN(n16680) );
  OAI211_X1 U19612 ( .C1(n16682), .C2(n19706), .A(n16681), .B(n16680), .ZN(
        P2_U3038) );
  NAND2_X1 U19613 ( .A1(n16687), .A2(n16683), .ZN(n16684) );
  OAI211_X1 U19614 ( .C1(n16686), .C2(n16722), .A(n16685), .B(n16684), .ZN(
        n16690) );
  NOR2_X1 U19615 ( .A1(n16688), .A2(n16687), .ZN(n16689) );
  AOI211_X1 U19616 ( .C1(n16691), .C2(n19712), .A(n16690), .B(n16689), .ZN(
        n16694) );
  OR2_X1 U19617 ( .A1(n16692), .A2(n19706), .ZN(n16693) );
  OAI211_X1 U19618 ( .C1(n16695), .C2(n16710), .A(n16694), .B(n16693), .ZN(
        P2_U3039) );
  INV_X1 U19619 ( .A(n16714), .ZN(n16696) );
  OAI21_X1 U19620 ( .B1(n17413), .B2(n16698), .A(n16696), .ZN(n16706) );
  NAND3_X1 U19621 ( .A1(n16716), .A2(n16698), .A3(n16697), .ZN(n16703) );
  INV_X1 U19622 ( .A(n16699), .ZN(n16700) );
  AOI21_X1 U19623 ( .B1(n16701), .B2(n19724), .A(n16700), .ZN(n16702) );
  OAI211_X1 U19624 ( .C1(n19728), .C2(n16704), .A(n16703), .B(n16702), .ZN(
        n16705) );
  AOI21_X1 U19625 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16706), .A(
        n16705), .ZN(n16709) );
  NAND2_X1 U19626 ( .A1(n16707), .A2(n19726), .ZN(n16708) );
  OAI211_X1 U19627 ( .C1(n16711), .C2(n16710), .A(n16709), .B(n16708), .ZN(
        P2_U3040) );
  NAND2_X1 U19628 ( .A1(n16712), .A2(n19721), .ZN(n16725) );
  OAI21_X1 U19629 ( .B1(n16715), .B2(n16714), .A(n16713), .ZN(n19716) );
  INV_X1 U19630 ( .A(n19716), .ZN(n16719) );
  NAND2_X1 U19631 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16716), .ZN(
        n19704) );
  AOI221_X1 U19632 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n19717), .C2(n16717), .A(
        n19704), .ZN(n16718) );
  AOI21_X1 U19633 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16719), .A(
        n16718), .ZN(n16721) );
  OAI211_X1 U19634 ( .C1(n16722), .C2(n19612), .A(n16721), .B(n16720), .ZN(
        n16723) );
  AOI21_X1 U19635 ( .B1(n19622), .B2(n19712), .A(n16723), .ZN(n16724) );
  OAI211_X1 U19636 ( .C1(n16726), .C2(n19706), .A(n16725), .B(n16724), .ZN(
        P2_U3041) );
  AOI22_X1 U19637 ( .A1(n19721), .A2(n16728), .B1(n19726), .B2(n16727), .ZN(
        n16737) );
  INV_X1 U19638 ( .A(n16729), .ZN(n17404) );
  AOI21_X1 U19639 ( .B1(n17404), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n16730), .ZN(n16736) );
  AOI22_X1 U19640 ( .A1(n19712), .A2(n16732), .B1(n16731), .B2(n19640), .ZN(
        n16735) );
  OAI211_X1 U19641 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n16733), .B(n19729), .ZN(n16734) );
  NAND4_X1 U19642 ( .A1(n16737), .A2(n16736), .A3(n16735), .A4(n16734), .ZN(
        P2_U3045) );
  INV_X1 U19643 ( .A(n16749), .ZN(n16741) );
  INV_X1 U19644 ( .A(n16738), .ZN(n16739) );
  AOI22_X1 U19645 ( .A1(n16739), .A2(n16742), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20248), .ZN(n16740) );
  OAI21_X1 U19646 ( .B1(n16799), .B2(n16741), .A(n16740), .ZN(n16746) );
  OAI21_X1 U19647 ( .B1(n17415), .B2(P2_FLUSH_REG_SCAN_IN), .A(n17419), .ZN(
        n16744) );
  INV_X1 U19648 ( .A(n16744), .ZN(n16745) );
  NOR2_X1 U19649 ( .A1(n20128), .A2(n16745), .ZN(n20481) );
  INV_X1 U19650 ( .A(n20481), .ZN(n20478) );
  MUX2_X1 U19651 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16746), .S(
        n20478), .Z(P2_U3605) );
  INV_X1 U19652 ( .A(n19640), .ZN(n16752) );
  AND2_X1 U19653 ( .A1(n20463), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20459) );
  INV_X1 U19654 ( .A(n20459), .ZN(n20457) );
  INV_X1 U19655 ( .A(n16747), .ZN(n16748) );
  NAND2_X1 U19656 ( .A1(n16749), .A2(n16748), .ZN(n16750) );
  MUX2_X1 U19657 ( .A(n20457), .B(n16750), .S(n20461), .Z(n16751) );
  OAI21_X1 U19658 ( .B1(n16752), .B2(n20304), .A(n16751), .ZN(n16753) );
  MUX2_X1 U19659 ( .A(n16753), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        n20481), .Z(P2_U3604) );
  INV_X1 U19660 ( .A(n16754), .ZN(n16761) );
  OAI222_X1 U19661 ( .A1(n16765), .A2(n16758), .B1(n16757), .B2(n16761), .C1(
        n16756), .C2(n16755), .ZN(n16759) );
  MUX2_X1 U19662 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n16759), .S(
        n17344), .Z(P2_U3601) );
  NAND3_X1 U19663 ( .A1(n16761), .A2(P2_STATE2_REG_1__SCAN_IN), .A3(n16760), 
        .ZN(n16764) );
  NAND2_X1 U19664 ( .A1(n16762), .A2(n20462), .ZN(n16763) );
  OAI211_X1 U19665 ( .C1(n16765), .C2(n20472), .A(n16764), .B(n16763), .ZN(
        n16766) );
  MUX2_X1 U19666 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16766), .S(
        n17344), .Z(P2_U3599) );
  OR2_X1 U19667 ( .A1(n20465), .A2(n20122), .ZN(n20010) );
  OAI21_X1 U19668 ( .B1(n20010), .B2(n20219), .A(n20463), .ZN(n16781) );
  NOR2_X1 U19669 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n16767) );
  NAND2_X1 U19670 ( .A1(n16767), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19912) );
  OR2_X1 U19671 ( .A1(n19912), .A2(n20248), .ZN(n19978) );
  OAI21_X1 U19672 ( .B1(n9802), .B2(n10120), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16768) );
  INV_X1 U19673 ( .A(n19971), .ZN(n16792) );
  NAND2_X1 U19674 ( .A1(n20253), .A2(n16769), .ZN(n19747) );
  OR2_X2 U19675 ( .A1(n19844), .A2(n20219), .ZN(n19975) );
  NAND2_X1 U19676 ( .A1(n19802), .A2(BUF2_REG_24__SCAN_IN), .ZN(n16775) );
  NOR2_X1 U19677 ( .A1(n16772), .A2(n20457), .ZN(n16773) );
  NAND2_X1 U19678 ( .A1(n19803), .A2(BUF1_REG_24__SCAN_IN), .ZN(n16774) );
  NAND2_X1 U19679 ( .A1(n19802), .A2(BUF2_REG_16__SCAN_IN), .ZN(n16777) );
  NAND2_X1 U19680 ( .A1(n19803), .A2(BUF1_REG_16__SCAN_IN), .ZN(n16776) );
  NAND2_X1 U19681 ( .A1(n19807), .A2(n10323), .ZN(n20249) );
  OAI22_X1 U19682 ( .A1(n20008), .A2(n20318), .B1(n19978), .B2(n20249), .ZN(
        n16778) );
  AOI21_X1 U19683 ( .B1(n19915), .B2(n20315), .A(n16778), .ZN(n16783) );
  INV_X1 U19684 ( .A(n19912), .ZN(n16780) );
  NAND2_X1 U19685 ( .A1(n19972), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n16782) );
  OAI211_X1 U19686 ( .C1(n16792), .C2(n19747), .A(n16783), .B(n16782), .ZN(
        P2_U3088) );
  NAND2_X1 U19687 ( .A1(n20253), .A2(n16784), .ZN(n16803) );
  NAND2_X1 U19688 ( .A1(n19802), .A2(BUF2_REG_25__SCAN_IN), .ZN(n16786) );
  NAND2_X1 U19689 ( .A1(n19803), .A2(BUF1_REG_25__SCAN_IN), .ZN(n16785) );
  NAND2_X1 U19690 ( .A1(n19802), .A2(BUF2_REG_17__SCAN_IN), .ZN(n16788) );
  NAND2_X1 U19691 ( .A1(n19803), .A2(BUF1_REG_17__SCAN_IN), .ZN(n16787) );
  INV_X1 U19692 ( .A(n20319), .ZN(n20263) );
  OAI22_X1 U19693 ( .A1(n20008), .A2(n20264), .B1(n20263), .B2(n19978), .ZN(
        n16789) );
  AOI21_X1 U19694 ( .B1(n19915), .B2(n20226), .A(n16789), .ZN(n16791) );
  NAND2_X1 U19695 ( .A1(n19972), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n16790) );
  OAI211_X1 U19696 ( .C1(n16792), .C2(n16803), .A(n16791), .B(n16790), .ZN(
        P2_U3089) );
  AND2_X1 U19697 ( .A1(n20465), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20312) );
  INV_X1 U19698 ( .A(n19875), .ZN(n20460) );
  NAND2_X1 U19699 ( .A1(n20312), .A2(n20460), .ZN(n16793) );
  NAND2_X1 U19700 ( .A1(n20480), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20121) );
  INV_X1 U19701 ( .A(n20121), .ZN(n20117) );
  NAND2_X1 U19702 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20117), .ZN(
        n16800) );
  NAND2_X1 U19703 ( .A1(n16793), .A2(n16800), .ZN(n16798) );
  NAND2_X1 U19704 ( .A1(n19873), .A2(n20117), .ZN(n20169) );
  INV_X1 U19705 ( .A(n20169), .ZN(n20165) );
  AND2_X1 U19706 ( .A1(n20169), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16794) );
  NAND2_X1 U19707 ( .A1(n16795), .A2(n16794), .ZN(n16802) );
  OAI211_X1 U19708 ( .C1(n20165), .C2(n20304), .A(n16802), .B(n20253), .ZN(
        n16796) );
  INV_X1 U19709 ( .A(n16796), .ZN(n16797) );
  INV_X1 U19710 ( .A(n20172), .ZN(n20154) );
  INV_X1 U19711 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16806) );
  NOR2_X2 U19712 ( .A1(n20246), .A2(n19875), .ZN(n20166) );
  AOI22_X1 U19713 ( .A1(n20184), .A2(n20321), .B1(n20166), .B2(n20226), .ZN(
        n16805) );
  OAI21_X1 U19714 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n16800), .A(n20302), 
        .ZN(n16801) );
  AOI22_X1 U19715 ( .A1(n20171), .A2(n20320), .B1(n20165), .B2(n20319), .ZN(
        n16804) );
  OAI211_X1 U19716 ( .C1(n20154), .C2(n16806), .A(n16805), .B(n16804), .ZN(
        P2_U3137) );
  INV_X1 U19717 ( .A(n16807), .ZN(n16809) );
  NAND2_X1 U19718 ( .A1(n19565), .A2(n19554), .ZN(n19574) );
  INV_X1 U19719 ( .A(n17518), .ZN(n19440) );
  NAND2_X1 U19720 ( .A1(n19555), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19438) );
  INV_X1 U19721 ( .A(n19565), .ZN(n19572) );
  NAND3_X1 U19722 ( .A1(n19555), .A2(n19558), .A3(n17521), .ZN(n19446) );
  NOR2_X1 U19723 ( .A1(n19444), .A2(n19446), .ZN(n17909) );
  NAND3_X1 U19724 ( .A1(n18840), .A2(n19572), .A3(n19443), .ZN(n16810) );
  OR2_X1 U19725 ( .A1(n19553), .A2(n18985), .ZN(n16812) );
  NAND2_X1 U19726 ( .A1(n19386), .A2(n17521), .ZN(n16823) );
  INV_X1 U19727 ( .A(n16823), .ZN(n16811) );
  NAND2_X1 U19728 ( .A1(n16812), .A2(n16811), .ZN(n19389) );
  NAND3_X1 U19729 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n17885) );
  NOR2_X1 U19730 ( .A1(n17929), .A2(n17885), .ZN(n16813) );
  NOR2_X1 U19731 ( .A1(n17699), .A2(n16813), .ZN(n17891) );
  NAND2_X1 U19732 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17901) );
  INV_X1 U19733 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19472) );
  OAI21_X1 U19734 ( .B1(n17917), .B2(n17901), .A(n19472), .ZN(n16822) );
  NOR2_X1 U19735 ( .A1(n18684), .A2(n18673), .ZN(n16814) );
  NAND2_X1 U19736 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18642), .ZN(
        n17874) );
  OAI21_X1 U19737 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16814), .A(
        n17874), .ZN(n18663) );
  INV_X1 U19738 ( .A(n16814), .ZN(n17895) );
  NAND2_X1 U19739 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18589) );
  NAND3_X1 U19740 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16815) );
  NAND2_X1 U19741 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18520) );
  NAND2_X1 U19742 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17079) );
  INV_X1 U19743 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18458) );
  NOR2_X1 U19744 ( .A1(n18458), .A2(n18441), .ZN(n18445) );
  INV_X1 U19745 ( .A(n18445), .ZN(n17064) );
  NAND2_X1 U19746 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18406) );
  NAND2_X1 U19747 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18373) );
  NAND2_X1 U19748 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17043) );
  INV_X1 U19749 ( .A(n17043), .ZN(n16816) );
  INV_X1 U19750 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17576) );
  NAND2_X1 U19751 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16956), .ZN(
        n17017) );
  INV_X2 U19752 ( .A(n17017), .ZN(n17000) );
  OAI21_X1 U19753 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17895), .A(
        n17744), .ZN(n17907) );
  INV_X1 U19754 ( .A(n19443), .ZN(n17829) );
  OAI21_X1 U19755 ( .B1(n18663), .B2(n17907), .A(n17829), .ZN(n16817) );
  AOI21_X1 U19756 ( .B1(n18663), .B2(n17907), .A(n16817), .ZN(n16821) );
  NAND2_X1 U19757 ( .A1(n18985), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16818) );
  NAND2_X1 U19758 ( .A1(n19389), .A2(n16818), .ZN(n16819) );
  INV_X1 U19759 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18138) );
  OAI22_X1 U19760 ( .A1(n18657), .A2(n17880), .B1(n17927), .B2(n18138), .ZN(
        n16820) );
  AOI211_X1 U19761 ( .C1(n17891), .C2(n16822), .A(n16821), .B(n16820), .ZN(
        n16827) );
  NAND3_X1 U19762 ( .A1(n18985), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n16823), 
        .ZN(n16824) );
  NAND2_X1 U19763 ( .A1(n17896), .A2(n18138), .ZN(n17879) );
  OAI211_X1 U19764 ( .C1(n17896), .C2(n18138), .A(n17866), .B(n17879), .ZN(
        n16826) );
  OAI211_X1 U19765 ( .C1(n19574), .C2(n16828), .A(n16827), .B(n16826), .ZN(
        P3_U2668) );
  INV_X1 U19766 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17970) );
  INV_X1 U19767 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17626) );
  INV_X1 U19768 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17676) );
  INV_X1 U19769 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n17232) );
  INV_X1 U19770 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17987) );
  NOR2_X1 U19771 ( .A1(n17232), .A2(n17987), .ZN(n16829) );
  AND2_X1 U19772 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17971) );
  NAND4_X1 U19773 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n16829), .A4(n17971), .ZN(n16830) );
  NOR4_X1 U19774 ( .A1(n17970), .A2(n17626), .A3(n17231), .A4(n16830), .ZN(
        n17963) );
  NAND2_X1 U19775 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17963), .ZN(n16832) );
  NAND2_X1 U19776 ( .A1(n16832), .A2(n18148), .ZN(n17964) );
  INV_X1 U19777 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n17544) );
  NAND2_X1 U19778 ( .A1(n18157), .A2(n17544), .ZN(n16831) );
  OAI22_X1 U19779 ( .A1(n17964), .A2(n17544), .B1(n16832), .B2(n16831), .ZN(
        P3_U2672) );
  OR2_X1 U19780 ( .A1(n18251), .A2(n19001), .ZN(n18229) );
  INV_X1 U19781 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18303) );
  INV_X1 U19782 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18300) );
  NAND4_X1 U19783 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n16834)
         );
  NAND2_X1 U19784 ( .A1(n18157), .A2(n18156), .ZN(n16842) );
  INV_X1 U19785 ( .A(n16842), .ZN(n16835) );
  INV_X1 U19786 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n16836) );
  NOR2_X1 U19787 ( .A1(n18241), .A2(n16836), .ZN(n16837) );
  NAND2_X1 U19788 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18224), .ZN(n18215) );
  OAI21_X1 U19789 ( .B1(n18224), .B2(n16837), .A(n18215), .ZN(n16841) );
  AOI22_X1 U19790 ( .A1(n18223), .A2(BUF2_REG_19__SCAN_IN), .B1(n18249), .B2(
        n16839), .ZN(n16840) );
  OAI211_X1 U19791 ( .C1(n18993), .C2(n18229), .A(n16841), .B(n16840), .ZN(
        P3_U2716) );
  AOI22_X1 U19792 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n18223), .B1(n18214), .B2(
        BUF2_REG_1__SCAN_IN), .ZN(n16846) );
  AND2_X1 U19793 ( .A1(n16842), .A2(P3_EAX_REG_17__SCAN_IN), .ZN(n16844) );
  NOR2_X1 U19794 ( .A1(n16842), .A2(P3_EAX_REG_17__SCAN_IN), .ZN(n16843) );
  AOI21_X1 U19795 ( .B1(n18251), .B2(n16844), .A(n16843), .ZN(n16845) );
  OAI211_X1 U19796 ( .C1(n16847), .C2(n18197), .A(n16846), .B(n16845), .ZN(
        P3_U2718) );
  INV_X1 U19797 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n16849) );
  OAI22_X1 U19798 ( .A1(n16849), .A2(n18221), .B1(n18197), .B2(n16848), .ZN(
        n16851) );
  AOI211_X1 U19799 ( .C1(n18231), .C2(n18300), .A(n18241), .B(n18156), .ZN(
        n16850) );
  AOI211_X1 U19800 ( .C1(n18214), .C2(BUF2_REG_0__SCAN_IN), .A(n16851), .B(
        n16850), .ZN(n16852) );
  INV_X1 U19801 ( .A(n16852), .ZN(P3_U2719) );
  INV_X1 U19802 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17491) );
  INV_X1 U19803 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18348) );
  INV_X1 U19804 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18344) );
  NAND2_X1 U19805 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n18240), .ZN(n16856) );
  AOI21_X1 U19806 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n18251), .A(n16859), .ZN(
        n16854) );
  NAND2_X1 U19807 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n16859), .ZN(n18239) );
  INV_X1 U19808 ( .A(n18239), .ZN(n16853) );
  OAI222_X1 U19809 ( .A1(n18255), .A2(n17491), .B1(n18197), .B2(n16855), .C1(
        n16854), .C2(n16853), .ZN(P3_U2722) );
  INV_X1 U19810 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18174) );
  INV_X1 U19811 ( .A(n16856), .ZN(n16863) );
  AOI21_X1 U19812 ( .B1(n18251), .B2(P3_EAX_REG_12__SCAN_IN), .A(n16863), .ZN(
        n16858) );
  OAI222_X1 U19813 ( .A1(n18255), .A2(n18174), .B1(n16859), .B2(n16858), .C1(
        n18197), .C2(n16857), .ZN(P3_U2723) );
  INV_X1 U19814 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17488) );
  AOI21_X1 U19815 ( .B1(n18251), .B2(P3_EAX_REG_11__SCAN_IN), .A(n18240), .ZN(
        n16862) );
  INV_X1 U19816 ( .A(n16860), .ZN(n16861) );
  OAI222_X1 U19817 ( .A1(n18255), .A2(n17488), .B1(n16863), .B2(n16862), .C1(
        n18197), .C2(n16861), .ZN(P3_U2724) );
  AOI22_X1 U19818 ( .A1(n18061), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16871) );
  AOI22_X1 U19819 ( .A1(n18008), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16870) );
  INV_X1 U19820 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16866) );
  NAND2_X1 U19821 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n16865) );
  NAND2_X1 U19822 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n16864) );
  OAI211_X1 U19823 ( .C1(n18112), .C2(n16866), .A(n16865), .B(n16864), .ZN(
        n16867) );
  INV_X1 U19824 ( .A(n16867), .ZN(n16869) );
  NAND2_X1 U19825 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n16868) );
  NAND4_X1 U19826 ( .A1(n16871), .A2(n16870), .A3(n16869), .A4(n16868), .ZN(
        n16877) );
  AOI22_X1 U19827 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18099), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16875) );
  AOI22_X1 U19828 ( .A1(n13361), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16874) );
  AOI22_X1 U19829 ( .A1(n13053), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16873) );
  AOI22_X1 U19830 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16872) );
  NAND4_X1 U19831 ( .A1(n16875), .A2(n16874), .A3(n16873), .A4(n16872), .ZN(
        n16876) );
  INV_X1 U19832 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n19012) );
  INV_X1 U19833 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18336) );
  NOR2_X1 U19834 ( .A1(n18336), .A2(n16878), .ZN(n16895) );
  AOI21_X1 U19835 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n18251), .A(n16895), .ZN(
        n16879) );
  OAI222_X1 U19836 ( .A1(n18197), .A2(n17151), .B1(n18255), .B2(n19012), .C1(
        n16879), .C2(n18247), .ZN(P3_U2728) );
  NAND2_X1 U19837 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n16881) );
  NAND2_X1 U19838 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n16880) );
  OAI211_X1 U19839 ( .C1(n18006), .C2(n16882), .A(n16881), .B(n16880), .ZN(
        n16883) );
  INV_X1 U19840 ( .A(n16883), .ZN(n16887) );
  AOI22_X1 U19841 ( .A1(n18008), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16886) );
  AOI22_X1 U19842 ( .A1(n18061), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16885) );
  NAND2_X1 U19843 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n16884) );
  NAND4_X1 U19844 ( .A1(n16887), .A2(n16886), .A3(n16885), .A4(n16884), .ZN(
        n16893) );
  AOI22_X1 U19845 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16891) );
  AOI22_X1 U19846 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16890) );
  AOI22_X1 U19847 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16889) );
  AOI22_X1 U19848 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16888) );
  NAND4_X1 U19849 ( .A1(n16891), .A2(n16890), .A3(n16889), .A4(n16888), .ZN(
        n16892) );
  INV_X1 U19850 ( .A(n16979), .ZN(n16897) );
  INV_X1 U19851 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n21479) );
  AOI21_X1 U19852 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18251), .A(n16894), .ZN(
        n16896) );
  OAI222_X1 U19853 ( .A1(n18197), .A2(n16897), .B1(n18255), .B2(n21479), .C1(
        n16896), .C2(n16895), .ZN(P3_U2729) );
  INV_X1 U19854 ( .A(n16908), .ZN(n16898) );
  NAND2_X1 U19855 ( .A1(n16898), .A2(n16960), .ZN(n16912) );
  INV_X1 U19856 ( .A(n16912), .ZN(n16900) );
  NAND2_X1 U19857 ( .A1(n16900), .A2(n16899), .ZN(n16916) );
  INV_X1 U19858 ( .A(n16923), .ZN(n16901) );
  NAND2_X1 U19859 ( .A1(n16901), .A2(n16979), .ZN(n16926) );
  OR2_X2 U19860 ( .A1(n16926), .A2(n17151), .ZN(n18583) );
  NAND2_X1 U19861 ( .A1(n16903), .A2(n16902), .ZN(n16907) );
  INV_X1 U19862 ( .A(n16904), .ZN(n16905) );
  NAND2_X1 U19863 ( .A1(n16905), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n16906) );
  XNOR2_X1 U19864 ( .A(n16908), .B(n16960), .ZN(n16910) );
  INV_X1 U19865 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16909) );
  XNOR2_X1 U19866 ( .A(n16910), .B(n16909), .ZN(n18651) );
  NAND2_X1 U19867 ( .A1(n18652), .A2(n18651), .ZN(n18650) );
  NAND2_X1 U19868 ( .A1(n16910), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16911) );
  NAND2_X1 U19869 ( .A1(n18650), .A2(n16911), .ZN(n18645) );
  XNOR2_X1 U19870 ( .A(n16912), .B(n16964), .ZN(n16913) );
  XNOR2_X1 U19871 ( .A(n16913), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18644) );
  NAND2_X1 U19872 ( .A1(n18645), .A2(n18644), .ZN(n18643) );
  INV_X1 U19873 ( .A(n16913), .ZN(n16914) );
  NAND2_X1 U19874 ( .A1(n16914), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n16915) );
  NAND2_X1 U19875 ( .A1(n18643), .A2(n16915), .ZN(n16920) );
  NAND2_X1 U19876 ( .A1(n16916), .A2(n16962), .ZN(n16917) );
  NAND2_X1 U19877 ( .A1(n16923), .A2(n16917), .ZN(n16918) );
  INV_X1 U19878 ( .A(n16918), .ZN(n16919) );
  NAND2_X1 U19879 ( .A1(n16920), .A2(n16919), .ZN(n16921) );
  XNOR2_X1 U19880 ( .A(n16979), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18611) );
  INV_X1 U19881 ( .A(n18611), .ZN(n16922) );
  XNOR2_X1 U19882 ( .A(n16923), .B(n16922), .ZN(n18617) );
  XNOR2_X1 U19883 ( .A(n16923), .B(n16979), .ZN(n16924) );
  NAND2_X1 U19884 ( .A1(n16924), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16925) );
  NAND2_X1 U19885 ( .A1(n16926), .A2(n17151), .ZN(n16927) );
  NAND2_X1 U19886 ( .A1(n18583), .A2(n16927), .ZN(n16928) );
  XNOR2_X1 U19887 ( .A(n17085), .B(n16928), .ZN(n18601) );
  INV_X1 U19888 ( .A(n16928), .ZN(n16929) );
  NAND2_X1 U19889 ( .A1(n17085), .A2(n16929), .ZN(n16930) );
  NOR2_X1 U19890 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18578) );
  INV_X1 U19891 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18489) );
  NOR2_X1 U19892 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17088) );
  INV_X1 U19893 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18760) );
  NAND2_X1 U19894 ( .A1(n17088), .A2(n18760), .ZN(n16934) );
  INV_X1 U19895 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16931) );
  NOR2_X1 U19896 ( .A1(n18882), .A2(n16931), .ZN(n18869) );
  NAND2_X1 U19897 ( .A1(n18831), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18508) );
  NAND2_X1 U19898 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16932) );
  INV_X1 U19899 ( .A(n18814), .ZN(n18487) );
  INV_X1 U19900 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18811) );
  INV_X1 U19901 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18773) );
  AND2_X1 U19902 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18461) );
  INV_X1 U19903 ( .A(n18461), .ZN(n18765) );
  OR2_X1 U19904 ( .A1(n18708), .A2(n18765), .ZN(n16935) );
  NAND2_X1 U19905 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18718) );
  NAND3_X1 U19906 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16936) );
  NOR2_X1 U19907 ( .A1(n18718), .A2(n16936), .ZN(n18687) );
  AND2_X1 U19908 ( .A1(n18687), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16937) );
  AND2_X1 U19909 ( .A1(n18464), .A2(n16937), .ZN(n16941) );
  INV_X1 U19910 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18702) );
  INV_X1 U19911 ( .A(n18718), .ZN(n18734) );
  AND2_X1 U19912 ( .A1(n18461), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18737) );
  NAND3_X1 U19913 ( .A1(n18734), .A2(n18737), .A3(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18713) );
  INV_X1 U19914 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18717) );
  NOR2_X1 U19915 ( .A1(n18713), .A2(n18717), .ZN(n17209) );
  INV_X1 U19916 ( .A(n17209), .ZN(n17169) );
  INV_X1 U19917 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21475) );
  INV_X1 U19918 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18756) );
  NAND2_X1 U19919 ( .A1(n18462), .A2(n18756), .ZN(n16938) );
  NOR2_X1 U19920 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n16938), .ZN(
        n18418) );
  INV_X1 U19921 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18716) );
  NAND3_X1 U19922 ( .A1(n18401), .A2(n18702), .A3(n18717), .ZN(n16939) );
  NAND2_X1 U19923 ( .A1(n17203), .A2(n16939), .ZN(n16940) );
  OR2_X2 U19924 ( .A1(n17198), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18377) );
  NAND2_X1 U19925 ( .A1(n16941), .A2(n18377), .ZN(n18378) );
  INV_X1 U19926 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18361) );
  AND2_X1 U19927 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17180) );
  INV_X1 U19928 ( .A(n17180), .ZN(n16942) );
  OAI21_X1 U19929 ( .B1(n18378), .B2(n16942), .A(n10114), .ZN(n16943) );
  AND2_X1 U19930 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17022) );
  NAND2_X1 U19931 ( .A1(n17022), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17114) );
  NOR2_X1 U19932 ( .A1(n17160), .A2(n17114), .ZN(n16994) );
  INV_X1 U19933 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17142) );
  AOI21_X1 U19934 ( .B1(n9654), .B2(n17142), .A(n10114), .ZN(n16945) );
  AND2_X1 U19935 ( .A1(n16954), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17116) );
  NOR3_X1 U19936 ( .A1(n16994), .A2(n16945), .A3(n17116), .ZN(n16951) );
  NAND2_X1 U19937 ( .A1(n10114), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16946) );
  MUX2_X1 U19938 ( .A(n10114), .B(n16946), .S(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .Z(n16950) );
  AND2_X1 U19939 ( .A1(n16994), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16949) );
  INV_X1 U19940 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17006) );
  AND2_X1 U19941 ( .A1(n17006), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16952) );
  MUX2_X1 U19942 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n16947), .S(
        n18583), .Z(n16948) );
  INV_X1 U19943 ( .A(n18586), .ZN(n18512) );
  INV_X1 U19944 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18389) );
  NOR2_X1 U19945 ( .A1(n17203), .A2(n18389), .ZN(n18376) );
  NAND2_X1 U19946 ( .A1(n18376), .A2(n17180), .ZN(n17182) );
  NOR2_X1 U19947 ( .A1(n17182), .A2(n17114), .ZN(n17133) );
  INV_X1 U19948 ( .A(n16952), .ZN(n17119) );
  NAND2_X1 U19949 ( .A1(n17133), .A2(n17116), .ZN(n16953) );
  OAI211_X1 U19950 ( .C1(n17133), .C2(n16954), .A(n17119), .B(n16953), .ZN(
        n17123) );
  INV_X1 U19951 ( .A(n18439), .ZN(n18516) );
  NAND2_X2 U19952 ( .A1(n18672), .A2(n18516), .ZN(n18426) );
  NOR2_X1 U19953 ( .A1(n18426), .A2(n18684), .ZN(n16955) );
  OR2_X2 U19954 ( .A1(n16955), .A2(n19336), .ZN(n17077) );
  NAND2_X1 U19955 ( .A1(n17077), .A2(n16956), .ZN(n17002) );
  INV_X1 U19956 ( .A(n17002), .ZN(n16957) );
  NOR2_X1 U19957 ( .A1(n18426), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17016) );
  NOR2_X1 U19958 ( .A1(n18684), .A2(n9735), .ZN(n17036) );
  OR2_X1 U19959 ( .A1(n19015), .A2(n16956), .ZN(n17015) );
  OAI211_X1 U19960 ( .C1(n18439), .C2(n17036), .A(n18672), .B(n17015), .ZN(
        n17021) );
  NAND2_X1 U19961 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17209), .ZN(
        n16988) );
  INV_X1 U19962 ( .A(n17176), .ZN(n18689) );
  NAND2_X1 U19963 ( .A1(n16967), .A2(n16960), .ZN(n16965) );
  INV_X1 U19964 ( .A(n16962), .ZN(n16961) );
  NAND2_X1 U19965 ( .A1(n18609), .A2(n16979), .ZN(n16978) );
  NOR2_X1 U19966 ( .A1(n16978), .A2(n17151), .ZN(n16986) );
  XNOR2_X1 U19967 ( .A(n16978), .B(n17153), .ZN(n16982) );
  XNOR2_X1 U19968 ( .A(n16963), .B(n16962), .ZN(n16976) );
  AND2_X1 U19969 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16976), .ZN(
        n16977) );
  XNOR2_X1 U19970 ( .A(n16965), .B(n16964), .ZN(n16973) );
  INV_X1 U19971 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18939) );
  NOR2_X1 U19972 ( .A1(n16973), .A2(n18939), .ZN(n16975) );
  XNOR2_X1 U19973 ( .A(n16967), .B(n16966), .ZN(n16971) );
  NOR2_X1 U19974 ( .A1(n16972), .A2(n18654), .ZN(n18638) );
  AOI21_X1 U19975 ( .B1(n16973), .B2(n18939), .A(n16975), .ZN(n16974) );
  INV_X1 U19976 ( .A(n16974), .ZN(n18637) );
  NOR2_X1 U19977 ( .A1(n18638), .A2(n18637), .ZN(n18636) );
  NOR2_X1 U19978 ( .A1(n16975), .A2(n18636), .ZN(n18628) );
  INV_X1 U19979 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18928) );
  XOR2_X1 U19980 ( .A(n18928), .B(n16976), .Z(n18627) );
  INV_X1 U19981 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17102) );
  OAI21_X1 U19982 ( .B1(n18609), .B2(n16979), .A(n16978), .ZN(n16980) );
  NOR2_X1 U19983 ( .A1(n18598), .A2(n9998), .ZN(n16981) );
  NAND2_X1 U19984 ( .A1(n16986), .A2(n16981), .ZN(n16987) );
  INV_X1 U19985 ( .A(n16981), .ZN(n16985) );
  AND2_X1 U19986 ( .A1(n16983), .A2(n16982), .ZN(n18599) );
  AOI21_X1 U19987 ( .B1(n16986), .B2(n16985), .A(n18599), .ZN(n16984) );
  OAI21_X1 U19988 ( .B1(n16986), .B2(n16985), .A(n16984), .ZN(n18585) );
  NAND2_X1 U19989 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18585), .ZN(
        n18584) );
  INV_X1 U19990 ( .A(n18370), .ZN(n16989) );
  NOR2_X1 U19991 ( .A1(n17181), .A2(n17114), .ZN(n17132) );
  NOR2_X2 U19992 ( .A1(n18658), .A2(n18579), .ZN(n18685) );
  NAND2_X1 U19993 ( .A1(n18953), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n17117) );
  OAI21_X1 U19994 ( .B1(n17862), .B2(n18530), .A(n17117), .ZN(n16991) );
  NOR3_X1 U19995 ( .A1(n17002), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A3(
        n10160), .ZN(n16990) );
  AOI21_X1 U19996 ( .B1(n18512), .B2(n17123), .A(n16992), .ZN(n16993) );
  OAI21_X1 U19997 ( .B1(n17126), .B2(n18556), .A(n16993), .ZN(P3_U2799) );
  NOR2_X1 U19998 ( .A1(n10114), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16995) );
  AOI21_X1 U19999 ( .B1(n9654), .B2(n16995), .A(n16994), .ZN(n16996) );
  XOR2_X1 U20000 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n16996), .Z(
        n17137) );
  NOR2_X1 U20001 ( .A1(n17114), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17130) );
  NAND2_X1 U20002 ( .A1(n18498), .A2(n18675), .ZN(n16998) );
  NAND2_X1 U20003 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18691) );
  INV_X1 U20004 ( .A(n18691), .ZN(n18686) );
  NAND2_X1 U20005 ( .A1(n17180), .A2(n18686), .ZN(n17177) );
  NOR2_X1 U20006 ( .A1(n18359), .A2(n17177), .ZN(n17059) );
  NAND2_X1 U20007 ( .A1(n18612), .A2(n18586), .ZN(n18424) );
  INV_X1 U20008 ( .A(n17181), .ZN(n17128) );
  INV_X1 U20009 ( .A(n17182), .ZN(n17023) );
  OAI22_X1 U20010 ( .A1(n17128), .A2(n18612), .B1(n18586), .B2(n17023), .ZN(
        n17028) );
  AOI21_X1 U20011 ( .B1(n17114), .B2(n18424), .A(n17028), .ZN(n17007) );
  OAI21_X1 U20012 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n17000), .A(
        n16999), .ZN(n17567) );
  INV_X1 U20013 ( .A(n17567), .ZN(n17004) );
  AND2_X1 U20014 ( .A1(n13496), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n17129) );
  AOI21_X1 U20015 ( .B1(n10160), .B2(n17002), .A(n17001), .ZN(n17003) );
  AOI211_X1 U20016 ( .C1(n18432), .C2(n17004), .A(n17129), .B(n17003), .ZN(
        n17005) );
  OAI21_X1 U20017 ( .B1(n17007), .B2(n17006), .A(n17005), .ZN(n17008) );
  AOI21_X1 U20018 ( .B1(n17130), .B2(n17059), .A(n17008), .ZN(n17009) );
  OAI21_X1 U20019 ( .B1(n17137), .B2(n18556), .A(n17009), .ZN(P3_U2800) );
  INV_X1 U20020 ( .A(n17160), .ZN(n17152) );
  OAI22_X1 U20021 ( .A1(n17152), .A2(n9654), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18583), .ZN(n17010) );
  XNOR2_X1 U20022 ( .A(n17010), .B(n17142), .ZN(n17150) );
  INV_X1 U20023 ( .A(n17132), .ZN(n17012) );
  INV_X1 U20024 ( .A(n17022), .ZN(n17138) );
  OAI21_X1 U20025 ( .B1(n17181), .B2(n17138), .A(n17142), .ZN(n17011) );
  NAND3_X1 U20026 ( .A1(n18675), .A2(n17012), .A3(n17011), .ZN(n17014) );
  INV_X1 U20027 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19520) );
  NOR2_X1 U20028 ( .A1(n18840), .A2(n19520), .ZN(n17141) );
  INV_X1 U20029 ( .A(n17141), .ZN(n17013) );
  OAI211_X1 U20030 ( .C1(n17015), .C2(n9735), .A(n17014), .B(n17013), .ZN(
        n17020) );
  INV_X1 U20031 ( .A(n17016), .ZN(n17018) );
  OAI21_X1 U20032 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n17036), .A(
        n17017), .ZN(n17582) );
  AOI21_X1 U20033 ( .B1(n17018), .B2(n18530), .A(n17582), .ZN(n17019) );
  AOI211_X1 U20034 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n17021), .A(
        n17020), .B(n17019), .ZN(n17026) );
  NAND2_X1 U20035 ( .A1(n17023), .A2(n17022), .ZN(n17140) );
  INV_X1 U20036 ( .A(n17140), .ZN(n17157) );
  INV_X1 U20037 ( .A(n17133), .ZN(n17024) );
  OAI211_X1 U20038 ( .C1(n17157), .C2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n18512), .B(n17024), .ZN(n17025) );
  OAI211_X1 U20039 ( .C1(n17150), .C2(n18556), .A(n17026), .B(n17025), .ZN(
        P3_U2801) );
  INV_X1 U20040 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17030) );
  XNOR2_X1 U20041 ( .A(n18583), .B(n17030), .ZN(n17161) );
  AOI211_X1 U20042 ( .C1(n17027), .C2(n17161), .A(n18556), .B(n9619), .ZN(
        n17048) );
  INV_X1 U20043 ( .A(n17028), .ZN(n18362) );
  INV_X1 U20044 ( .A(n18424), .ZN(n17029) );
  AOI211_X1 U20045 ( .C1(n18362), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17030), .B(n17029), .ZN(n17047) );
  INV_X1 U20046 ( .A(n17177), .ZN(n17107) );
  AND2_X1 U20047 ( .A1(n17030), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17031) );
  NAND2_X1 U20048 ( .A1(n17107), .A2(n17031), .ZN(n17168) );
  INV_X1 U20049 ( .A(n17055), .ZN(n17033) );
  AOI21_X1 U20050 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18357), .A(
        n18439), .ZN(n17032) );
  AOI21_X1 U20051 ( .B1(n17033), .B2(n18579), .A(n17032), .ZN(n17034) );
  AND2_X1 U20052 ( .A1(n18672), .A2(n17034), .ZN(n18369) );
  OAI21_X1 U20053 ( .B1(n18426), .B2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n18369), .ZN(n17054) );
  AND2_X1 U20054 ( .A1(n17055), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17554) );
  OR2_X1 U20055 ( .A1(n17554), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17039) );
  INV_X1 U20056 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17598) );
  INV_X1 U20057 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17035) );
  NAND2_X1 U20058 ( .A1(n17598), .A2(n17035), .ZN(n17042) );
  INV_X1 U20059 ( .A(n17036), .ZN(n17037) );
  AND2_X1 U20060 ( .A1(n17042), .A2(n17037), .ZN(n17038) );
  NAND2_X1 U20061 ( .A1(n17039), .A2(n17038), .ZN(n17591) );
  AND2_X1 U20062 ( .A1(n13496), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17171) );
  INV_X1 U20063 ( .A(n17171), .ZN(n17040) );
  OAI21_X1 U20064 ( .B1(n17591), .B2(n18530), .A(n17040), .ZN(n17041) );
  AOI21_X1 U20065 ( .B1(n17054), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n17041), .ZN(n17045) );
  NAND4_X1 U20066 ( .A1(n17077), .A2(n17043), .A3(n17055), .A4(n17042), .ZN(
        n17044) );
  OAI211_X1 U20067 ( .C1(n18359), .C2(n17168), .A(n17045), .B(n17044), .ZN(
        n17046) );
  OR3_X1 U20068 ( .A1(n17048), .A2(n17047), .A3(n17046), .ZN(P3_U2802) );
  NAND2_X1 U20069 ( .A1(n17049), .A2(n17162), .ZN(n17050) );
  MUX2_X1 U20070 ( .A(n17162), .B(n17050), .S(n18583), .Z(n17051) );
  NAND2_X1 U20071 ( .A1(n17051), .A2(n17160), .ZN(n17190) );
  INV_X1 U20072 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n17052) );
  NOR2_X1 U20073 ( .A1(n18840), .A2(n17052), .ZN(n17187) );
  XNOR2_X1 U20074 ( .A(n17554), .B(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17605) );
  NOR2_X1 U20075 ( .A1(n17605), .A2(n18530), .ZN(n17053) );
  AOI211_X1 U20076 ( .C1(n17054), .C2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n17187), .B(n17053), .ZN(n17057) );
  NAND3_X1 U20077 ( .A1(n17077), .A2(n17055), .A3(n17598), .ZN(n17056) );
  OAI211_X1 U20078 ( .C1(n18362), .C2(n17154), .A(n17057), .B(n17056), .ZN(
        n17058) );
  AOI21_X1 U20079 ( .B1(n17059), .B2(n17154), .A(n17058), .ZN(n17060) );
  OAI21_X1 U20080 ( .B1(n17190), .B2(n18556), .A(n17060), .ZN(P3_U2803) );
  INV_X1 U20081 ( .A(n18399), .ZN(n18435) );
  AOI21_X1 U20082 ( .B1(n18464), .B2(n18687), .A(n18401), .ZN(n17061) );
  AOI211_X1 U20083 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18583), .A(
        n18435), .B(n17061), .ZN(n17062) );
  XNOR2_X1 U20084 ( .A(n17062), .B(n18702), .ZN(n18706) );
  INV_X1 U20085 ( .A(n18706), .ZN(n17075) );
  INV_X1 U20086 ( .A(n17203), .ZN(n17063) );
  OAI22_X1 U20087 ( .A1(n17200), .A2(n18612), .B1(n17063), .B2(n18586), .ZN(
        n18387) );
  INV_X1 U20088 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19511) );
  INV_X1 U20089 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18416) );
  NOR2_X1 U20090 ( .A1(n18684), .A2(n18454), .ZN(n18440) );
  INV_X1 U20091 ( .A(n18440), .ZN(n17710) );
  NAND2_X1 U20092 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18403), .ZN(
        n17561) );
  NOR2_X1 U20093 ( .A1(n18416), .A2(n17561), .ZN(n17560) );
  NAND2_X1 U20094 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17560), .ZN(
        n17559) );
  INV_X1 U20095 ( .A(n17559), .ZN(n17065) );
  OAI22_X1 U20096 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17065), .B1(
        n18684), .B2(n18372), .ZN(n17650) );
  OAI22_X1 U20097 ( .A1(n18840), .A2(n19511), .B1(n18530), .B2(n17650), .ZN(
        n17071) );
  OAI21_X1 U20098 ( .B1(n17065), .B2(n18439), .A(n18672), .ZN(n17066) );
  AOI21_X1 U20099 ( .B1(n19336), .B2(n18372), .A(n17066), .ZN(n18371) );
  INV_X1 U20100 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17069) );
  NAND3_X1 U20101 ( .A1(n17067), .A2(n17077), .A3(n17069), .ZN(n17068) );
  OAI21_X1 U20102 ( .B1(n18371), .B2(n17069), .A(n17068), .ZN(n17070) );
  NOR2_X1 U20103 ( .A1(n17071), .A2(n17070), .ZN(n17072) );
  OAI21_X1 U20104 ( .B1(n18359), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n17072), .ZN(n17073) );
  AOI21_X1 U20105 ( .B1(n18387), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n17073), .ZN(n17074) );
  OAI21_X1 U20106 ( .B1(n17075), .B2(n18556), .A(n17074), .ZN(P3_U2807) );
  OR2_X1 U20107 ( .A1(n18709), .A2(n18612), .ZN(n18486) );
  OR2_X1 U20108 ( .A1(n18586), .A2(n10105), .ZN(n18492) );
  NAND2_X1 U20109 ( .A1(n18486), .A2(n18492), .ZN(n18423) );
  INV_X1 U20110 ( .A(n18423), .ZN(n18460) );
  INV_X1 U20111 ( .A(n18481), .ZN(n18398) );
  INV_X1 U20112 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19497) );
  NOR2_X1 U20113 ( .A1(n18684), .A2(n17078), .ZN(n17746) );
  AOI21_X1 U20114 ( .B1(n18579), .B2(n17078), .A(n18658), .ZN(n18500) );
  OAI21_X1 U20115 ( .B1(n17746), .B2(n18439), .A(n18500), .ZN(n18483) );
  INV_X1 U20116 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17076) );
  NAND2_X1 U20117 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17746), .ZN(
        n17732) );
  AND2_X1 U20118 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18471), .ZN(
        n17711) );
  AOI21_X1 U20119 ( .B1(n17076), .B2(n17732), .A(n17711), .ZN(n17725) );
  AOI22_X1 U20120 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18483), .B1(
        n18432), .B2(n17725), .ZN(n17081) );
  NOR2_X1 U20121 ( .A1(n18519), .A2(n17078), .ZN(n18485) );
  OAI211_X1 U20122 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18485), .B(n17079), .ZN(n17080) );
  OAI211_X1 U20123 ( .C1(n19497), .C2(n18840), .A(n17081), .B(n17080), .ZN(
        n17082) );
  AOI21_X1 U20124 ( .B1(n18398), .B2(n18760), .A(n17082), .ZN(n17091) );
  NAND2_X1 U20125 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17083) );
  NOR2_X1 U20126 ( .A1(n18583), .A2(n17083), .ZN(n17084) );
  AND2_X1 U20127 ( .A1(n17085), .A2(n17084), .ZN(n18563) );
  NAND2_X1 U20128 ( .A1(n18563), .A2(n18831), .ZN(n18535) );
  NAND3_X1 U20129 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17086) );
  NOR3_X1 U20130 ( .A1(n18535), .A2(n17086), .A3(n18811), .ZN(n17087) );
  AOI21_X1 U20131 ( .B1(n9880), .B2(n17088), .A(n17087), .ZN(n17089) );
  XNOR2_X1 U20132 ( .A(n17089), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n18793) );
  NAND2_X1 U20133 ( .A1(n18793), .A2(n18588), .ZN(n17090) );
  OAI211_X1 U20134 ( .C1(n18460), .C2(n18760), .A(n17091), .B(n17090), .ZN(
        P3_U2814) );
  NOR3_X1 U20135 ( .A1(n18594), .A2(n18589), .A3(n19015), .ZN(n17092) );
  NAND2_X1 U20136 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17092), .ZN(
        n18559) );
  INV_X1 U20137 ( .A(n18559), .ZN(n17094) );
  INV_X1 U20138 ( .A(n18685), .ZN(n18546) );
  AOI21_X1 U20139 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18546), .A(
        n17092), .ZN(n17093) );
  NAND3_X1 U20140 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(n18615), .ZN(n17835) );
  NOR2_X1 U20141 ( .A1(n18589), .A2(n17835), .ZN(n17827) );
  NAND2_X1 U20142 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17827), .ZN(
        n17799) );
  OAI21_X1 U20143 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17827), .A(
        n17799), .ZN(n17813) );
  OAI22_X1 U20144 ( .A1(n17094), .A2(n17093), .B1(n18667), .B2(n17813), .ZN(
        n17100) );
  INV_X1 U20145 ( .A(n18581), .ZN(n18864) );
  OAI22_X1 U20146 ( .A1(n18498), .A2(n18612), .B1(n18864), .B2(n18586), .ZN(
        n18574) );
  INV_X1 U20147 ( .A(n18574), .ZN(n18551) );
  INV_X1 U20148 ( .A(n18563), .ZN(n17095) );
  NAND2_X1 U20149 ( .A1(n17096), .A2(n17095), .ZN(n18571) );
  NOR2_X1 U20150 ( .A1(n17096), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18566) );
  AOI21_X1 U20151 ( .B1(n18882), .B2(n18563), .A(n18566), .ZN(n17097) );
  OAI21_X1 U20152 ( .B1(n18882), .B2(n18571), .A(n17097), .ZN(n18886) );
  INV_X1 U20153 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19483) );
  NOR2_X1 U20154 ( .A1(n18840), .A2(n19483), .ZN(n18885) );
  AOI21_X1 U20155 ( .B1(n18588), .B2(n18886), .A(n18885), .ZN(n17098) );
  OAI21_X1 U20156 ( .B1(n18551), .B2(n18882), .A(n17098), .ZN(n17099) );
  AOI211_X1 U20157 ( .C1(n18882), .C2(n18554), .A(n17100), .B(n17099), .ZN(
        n17101) );
  INV_X1 U20158 ( .A(n17101), .ZN(P3_U2821) );
  NAND3_X1 U20159 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18919) );
  NOR2_X1 U20160 ( .A1(n17102), .A2(n18919), .ZN(n18911) );
  AND2_X1 U20161 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18911), .ZN(
        n18900) );
  NAND2_X1 U20162 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18900), .ZN(
        n17164) );
  NOR2_X1 U20163 ( .A1(n17164), .A2(n18786), .ZN(n18858) );
  NOR2_X1 U20164 ( .A1(n18689), .A2(n18713), .ZN(n18721) );
  NAND2_X1 U20165 ( .A1(n18858), .A2(n18721), .ZN(n18715) );
  NOR2_X1 U20166 ( .A1(n18717), .A2(n18715), .ZN(n17108) );
  NAND3_X1 U20167 ( .A1(n17108), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17107), .ZN(n17105) );
  INV_X1 U20168 ( .A(n17164), .ZN(n18783) );
  NAND2_X1 U20169 ( .A1(n17176), .A2(n18783), .ZN(n18785) );
  INV_X1 U20170 ( .A(n18785), .ZN(n17103) );
  NAND2_X1 U20171 ( .A1(n18782), .A2(n17103), .ZN(n18711) );
  OR2_X1 U20172 ( .A1(n17169), .A2(n18711), .ZN(n17178) );
  NOR2_X1 U20173 ( .A1(n17178), .A2(n17177), .ZN(n17109) );
  NOR2_X1 U20174 ( .A1(n17109), .A2(n18784), .ZN(n17104) );
  NAND2_X1 U20175 ( .A1(n18783), .A2(n18895), .ZN(n18780) );
  NOR3_X1 U20176 ( .A1(n18765), .A2(n18689), .A3(n18780), .ZN(n18762) );
  NAND2_X1 U20177 ( .A1(n18762), .A2(n18687), .ZN(n18692) );
  NOR2_X1 U20178 ( .A1(n18692), .A2(n17177), .ZN(n17110) );
  NOR2_X1 U20179 ( .A1(n17110), .A2(n18896), .ZN(n17184) );
  AOI211_X1 U20180 ( .C1(n18861), .C2(n17105), .A(n17104), .B(n17184), .ZN(
        n17144) );
  OR2_X1 U20181 ( .A1(n18792), .A2(n18899), .ZN(n18916) );
  INV_X1 U20182 ( .A(n18916), .ZN(n18957) );
  NAND2_X1 U20183 ( .A1(n18957), .A2(n17114), .ZN(n17106) );
  OAI211_X1 U20184 ( .C1(n17144), .C2(n18899), .A(n18855), .B(n17106), .ZN(
        n17134) );
  NAND2_X1 U20185 ( .A1(n17108), .A2(n17107), .ZN(n17112) );
  AOI22_X1 U20186 ( .A1(n19406), .A2(n17110), .B1(n17109), .B2(n18958), .ZN(
        n17111) );
  OAI21_X1 U20187 ( .B1(n18868), .B2(n17112), .A(n17111), .ZN(n17113) );
  AND2_X1 U20188 ( .A1(n17113), .A2(n18944), .ZN(n17127) );
  INV_X1 U20189 ( .A(n17114), .ZN(n17115) );
  NAND3_X1 U20190 ( .A1(n17127), .A2(n17116), .A3(n17115), .ZN(n17118) );
  OAI211_X1 U20191 ( .C1(n18916), .C2(n17119), .A(n17118), .B(n17117), .ZN(
        n17122) );
  AND2_X1 U20192 ( .A1(n18952), .A2(n17120), .ZN(n17121) );
  AOI211_X1 U20193 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n17134), .A(
        n17122), .B(n17121), .ZN(n17125) );
  OR2_X1 U20194 ( .A1(n18906), .A2(n17153), .ZN(n18890) );
  INV_X1 U20195 ( .A(n18890), .ZN(n18823) );
  NAND2_X1 U20196 ( .A1(n17123), .A2(n18823), .ZN(n17124) );
  OAI211_X1 U20197 ( .C1(n17126), .C2(n18873), .A(n17125), .B(n17124), .ZN(
        P3_U2831) );
  AOI21_X1 U20198 ( .B1(n18952), .B2(n17128), .A(n17127), .ZN(n17139) );
  OAI21_X1 U20199 ( .B1(n17182), .B2(n18890), .A(n17139), .ZN(n17131) );
  AOI21_X1 U20200 ( .B1(n17131), .B2(n17130), .A(n17129), .ZN(n17136) );
  OAI22_X1 U20201 ( .A1(n17133), .A2(n18890), .B1(n17132), .B2(n18923), .ZN(
        n17147) );
  OAI21_X1 U20202 ( .B1(n17147), .B2(n17134), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17135) );
  OAI211_X1 U20203 ( .C1(n17137), .C2(n18873), .A(n17136), .B(n17135), .ZN(
        P3_U2832) );
  OAI22_X1 U20204 ( .A1(n17140), .A2(n18890), .B1(n17139), .B2(n17138), .ZN(
        n17143) );
  AOI21_X1 U20205 ( .B1(n17143), .B2(n17142), .A(n17141), .ZN(n17149) );
  INV_X1 U20206 ( .A(n17144), .ZN(n17145) );
  AOI211_X1 U20207 ( .C1(n17154), .C2(n18875), .A(n18955), .B(n17145), .ZN(
        n17156) );
  OAI22_X1 U20208 ( .A1(n17156), .A2(n18953), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18916), .ZN(n17146) );
  OAI21_X1 U20209 ( .B1(n17147), .B2(n17146), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17148) );
  OAI211_X1 U20210 ( .C1(n17150), .C2(n18873), .A(n17149), .B(n17148), .ZN(
        P3_U2833) );
  OR2_X1 U20211 ( .A1(n19399), .A2(n17151), .ZN(n18804) );
  NOR3_X1 U20212 ( .A1(n9619), .A2(n17152), .A3(n18804), .ZN(n17159) );
  OR2_X1 U20213 ( .A1(n19399), .A2(n17153), .ZN(n18863) );
  OAI21_X1 U20214 ( .B1(n17154), .B2(n17181), .A(n19404), .ZN(n17155) );
  OAI211_X1 U20215 ( .C1(n17157), .C2(n18863), .A(n17156), .B(n17155), .ZN(
        n17158) );
  OAI211_X1 U20216 ( .C1(n17159), .C2(n17158), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18840), .ZN(n17175) );
  NOR3_X1 U20217 ( .A1(n17160), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n18906), .ZN(n17173) );
  NOR3_X1 U20218 ( .A1(n17162), .A2(n9882), .A3(n18873), .ZN(n17172) );
  NAND2_X1 U20219 ( .A1(n18498), .A2(n19404), .ZN(n17167) );
  AOI22_X1 U20220 ( .A1(n19406), .A2(n18895), .B1(n18782), .B2(n17163), .ZN(
        n18909) );
  NOR2_X1 U20221 ( .A1(n18909), .A2(n17164), .ZN(n18812) );
  NOR2_X1 U20222 ( .A1(n18863), .A2(n18581), .ZN(n17165) );
  NOR2_X1 U20223 ( .A1(n18812), .A2(n17165), .ZN(n17166) );
  NAND2_X1 U20224 ( .A1(n17167), .A2(n17166), .ZN(n18722) );
  NOR3_X1 U20225 ( .A1(n18797), .A2(n17169), .A3(n17168), .ZN(n17170) );
  NOR4_X1 U20226 ( .A1(n17173), .A2(n17172), .A3(n17171), .A4(n17170), .ZN(
        n17174) );
  NAND2_X1 U20227 ( .A1(n17175), .A2(n17174), .ZN(P3_U2834) );
  NAND3_X1 U20228 ( .A1(n18722), .A2(n17176), .A3(n17209), .ZN(n18703) );
  NOR2_X1 U20229 ( .A1(n18703), .A2(n17177), .ZN(n17186) );
  INV_X1 U20230 ( .A(n18758), .ZN(n17179) );
  OAI21_X1 U20231 ( .B1(n17179), .B2(n17178), .A(n18759), .ZN(n17201) );
  OAI21_X1 U20232 ( .B1(n18686), .B2(n18766), .A(n17201), .ZN(n18690) );
  OAI22_X1 U20233 ( .A1(n18784), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18868), .B2(n17180), .ZN(n17183) );
  OAI211_X1 U20234 ( .C1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n18784), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17193), .ZN(n17185) );
  OAI211_X1 U20235 ( .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n17186), .A(
        n17185), .B(n18944), .ZN(n17189) );
  AOI21_X1 U20236 ( .B1(n18955), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17187), .ZN(n17188) );
  OAI211_X1 U20237 ( .C1(n17190), .C2(n18873), .A(n17189), .B(n17188), .ZN(
        P3_U2835) );
  OAI21_X1 U20238 ( .B1(n9699), .B2(n18361), .A(n17191), .ZN(n17192) );
  INV_X1 U20239 ( .A(n17192), .ZN(n18363) );
  NAND3_X1 U20240 ( .A1(n18361), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n18686), .ZN(n18360) );
  OAI22_X1 U20241 ( .A1(n17193), .A2(n18361), .B1(n18703), .B2(n18360), .ZN(
        n17196) );
  INV_X1 U20242 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n17194) );
  OAI22_X1 U20243 ( .A1(n18855), .A2(n18361), .B1(n18840), .B2(n17194), .ZN(
        n17195) );
  AOI21_X1 U20244 ( .B1(n17196), .B2(n18944), .A(n17195), .ZN(n17197) );
  OAI21_X1 U20245 ( .B1(n18363), .B2(n18873), .A(n17197), .ZN(P3_U2836) );
  NAND2_X1 U20246 ( .A1(n17198), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17199) );
  AND2_X1 U20247 ( .A1(n18377), .A2(n17199), .ZN(n18388) );
  INV_X1 U20248 ( .A(n18792), .ZN(n17208) );
  INV_X1 U20249 ( .A(n19404), .ZN(n18829) );
  OR2_X1 U20250 ( .A1(n17200), .A2(n18829), .ZN(n17205) );
  NAND2_X1 U20251 ( .A1(n17201), .A2(n18855), .ZN(n17202) );
  AOI21_X1 U20252 ( .B1(n17203), .B2(n18712), .A(n17202), .ZN(n17204) );
  NAND2_X1 U20253 ( .A1(n17205), .A2(n17204), .ZN(n17207) );
  AOI211_X1 U20254 ( .C1(n19406), .C2(n18692), .A(n18702), .B(n17207), .ZN(
        n17206) );
  NOR2_X1 U20255 ( .A1(n17206), .A2(n18953), .ZN(n18705) );
  OAI211_X1 U20256 ( .C1(n17208), .C2(n17207), .A(n18705), .B(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17214) );
  NOR2_X1 U20257 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18702), .ZN(
        n18392) );
  NAND2_X1 U20258 ( .A1(n17209), .A2(n18392), .ZN(n17211) );
  INV_X1 U20259 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19513) );
  NOR2_X1 U20260 ( .A1(n18840), .A2(n19513), .ZN(n18383) );
  INV_X1 U20261 ( .A(n18383), .ZN(n17210) );
  OAI21_X1 U20262 ( .B1(n18797), .B2(n17211), .A(n17210), .ZN(n17212) );
  INV_X1 U20263 ( .A(n17212), .ZN(n17213) );
  OAI211_X1 U20264 ( .C1(n18388), .C2(n18873), .A(n17214), .B(n17213), .ZN(
        P3_U2838) );
  NAND2_X1 U20265 ( .A1(n18868), .A2(n17215), .ZN(n17224) );
  MUX2_X1 U20266 ( .A(n18958), .B(n17224), .S(n17217), .Z(n19408) );
  INV_X1 U20267 ( .A(n19408), .ZN(n19409) );
  AOI22_X1 U20268 ( .A1(n17227), .A2(n17217), .B1(n17216), .B2(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n17218) );
  OAI21_X1 U20269 ( .B1(n19409), .B2(n19570), .A(n17218), .ZN(n17219) );
  MUX2_X1 U20270 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n17219), .S(
        n17229), .Z(P3_U3290) );
  NOR2_X1 U20271 ( .A1(n17221), .A2(n17220), .ZN(n17918) );
  AOI22_X1 U20272 ( .A1(n17224), .A2(n17918), .B1(n17223), .B2(n17222), .ZN(
        n19410) );
  AOI22_X1 U20273 ( .A1(n17918), .A2(n17227), .B1(n17226), .B2(n17225), .ZN(
        n17228) );
  OAI21_X1 U20274 ( .B1(n19410), .B2(n19570), .A(n17228), .ZN(n17230) );
  MUX2_X1 U20275 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n17230), .S(
        n17229), .Z(P3_U3289) );
  INV_X1 U20276 ( .A(n17977), .ZN(n17972) );
  NAND2_X1 U20277 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17972), .ZN(n17340) );
  OAI21_X1 U20278 ( .B1(n17971), .B2(n17233), .A(n17982), .ZN(n17969) );
  INV_X1 U20279 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U20280 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18057), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17235) );
  AOI22_X1 U20281 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17234) );
  OAI211_X1 U20282 ( .C1(n13034), .C2(n17236), .A(n17235), .B(n17234), .ZN(
        n17246) );
  INV_X1 U20283 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17238) );
  AOI22_X1 U20284 ( .A1(n18008), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17312), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17237) );
  OAI21_X1 U20285 ( .B1(n17239), .B2(n17238), .A(n17237), .ZN(n17245) );
  AOI22_X1 U20286 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17243) );
  AOI22_X1 U20287 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U20288 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17241) );
  AOI22_X1 U20289 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17240) );
  NAND4_X1 U20290 ( .A1(n17243), .A2(n17242), .A3(n17241), .A4(n17240), .ZN(
        n17244) );
  NOR3_X1 U20291 ( .A1(n17246), .A2(n17245), .A3(n17244), .ZN(n17338) );
  INV_X1 U20292 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18086) );
  INV_X1 U20293 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18080) );
  OAI22_X1 U20294 ( .A1(n18077), .A2(n18086), .B1(n9640), .B2(n18080), .ZN(
        n17251) );
  INV_X1 U20295 ( .A(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17249) );
  AOI22_X1 U20296 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17322), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U20297 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17247) );
  OAI211_X1 U20298 ( .C1(n18112), .C2(n17249), .A(n17248), .B(n17247), .ZN(
        n17250) );
  AOI211_X1 U20299 ( .C1(n17293), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n17251), .B(n17250), .ZN(n17259) );
  AOI22_X1 U20300 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17258) );
  AOI22_X1 U20301 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17257) );
  INV_X1 U20302 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17252) );
  NOR2_X1 U20303 ( .A1(n18085), .A2(n17252), .ZN(n17255) );
  INV_X1 U20304 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17253) );
  INV_X1 U20305 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18076) );
  OAI22_X1 U20306 ( .A1(n10446), .A2(n17253), .B1(n13229), .B2(n18076), .ZN(
        n17254) );
  AOI211_X1 U20307 ( .C1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .C2(n17266), .A(
        n17255), .B(n17254), .ZN(n17256) );
  NAND4_X1 U20308 ( .A1(n17259), .A2(n17258), .A3(n17257), .A4(n17256), .ZN(
        n17984) );
  AOI22_X1 U20309 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18108), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17261) );
  NAND2_X1 U20310 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n17260) );
  AND2_X1 U20311 ( .A1(n17261), .A2(n17260), .ZN(n17265) );
  AOI22_X1 U20312 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17264) );
  AOI22_X1 U20313 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17322), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17263) );
  NAND2_X1 U20314 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n17262) );
  NAND4_X1 U20315 ( .A1(n17265), .A2(n17264), .A3(n17263), .A4(n17262), .ZN(
        n17272) );
  AOI22_X1 U20316 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17270) );
  AOI22_X1 U20317 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17312), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17269) );
  AOI22_X1 U20318 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17268) );
  AOI22_X1 U20319 ( .A1(n17266), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17267) );
  NAND4_X1 U20320 ( .A1(n17270), .A2(n17269), .A3(n17268), .A4(n17267), .ZN(
        n17271) );
  OR2_X1 U20321 ( .A1(n17272), .A2(n17271), .ZN(n17998) );
  NAND2_X1 U20322 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n17274) );
  NAND2_X1 U20323 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n17273) );
  OAI211_X1 U20324 ( .C1(n17276), .C2(n17275), .A(n17274), .B(n17273), .ZN(
        n17277) );
  INV_X1 U20325 ( .A(n17277), .ZN(n17282) );
  AOI22_X1 U20326 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17281) );
  AOI22_X1 U20327 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17322), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17280) );
  NAND2_X1 U20328 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n17279) );
  NAND4_X1 U20329 ( .A1(n17282), .A2(n17281), .A3(n17280), .A4(n17279), .ZN(
        n17288) );
  AOI22_X1 U20330 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20331 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17312), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17285) );
  AOI22_X1 U20332 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17284) );
  AOI22_X1 U20333 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17283) );
  NAND4_X1 U20334 ( .A1(n17286), .A2(n17285), .A3(n17284), .A4(n17283), .ZN(
        n17287) );
  OR2_X1 U20335 ( .A1(n17288), .A2(n17287), .ZN(n17997) );
  AND2_X1 U20336 ( .A1(n17998), .A2(n17997), .ZN(n17995) );
  NAND2_X1 U20337 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n17290) );
  NAND2_X1 U20338 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n17289) );
  OAI211_X1 U20339 ( .C1(n17276), .C2(n17291), .A(n17290), .B(n17289), .ZN(
        n17292) );
  INV_X1 U20340 ( .A(n17292), .ZN(n17297) );
  AOI22_X1 U20341 ( .A1(n18008), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17296) );
  AOI22_X1 U20342 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17322), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17295) );
  NAND2_X1 U20343 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n17294) );
  NAND4_X1 U20344 ( .A1(n17297), .A2(n17296), .A3(n17295), .A4(n17294), .ZN(
        n17306) );
  AOI22_X1 U20345 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17304) );
  AOI22_X1 U20346 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17303) );
  AOI22_X1 U20347 ( .A1(n17299), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18100), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17302) );
  AOI22_X1 U20348 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17301) );
  NAND4_X1 U20349 ( .A1(n17304), .A2(n17303), .A3(n17302), .A4(n17301), .ZN(
        n17305) );
  OR2_X1 U20350 ( .A1(n17306), .A2(n17305), .ZN(n17988) );
  AND2_X1 U20351 ( .A1(n17995), .A2(n17988), .ZN(n17990) );
  NAND2_X1 U20352 ( .A1(n17984), .A2(n17990), .ZN(n17983) );
  INV_X1 U20353 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17309) );
  AOI22_X1 U20354 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17322), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17308) );
  AOI22_X1 U20355 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17307) );
  OAI211_X1 U20356 ( .C1(n18112), .C2(n17309), .A(n17308), .B(n17307), .ZN(
        n17319) );
  AOI22_X1 U20357 ( .A1(n18008), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17310) );
  OAI21_X1 U20358 ( .B1(n17239), .B2(n17311), .A(n17310), .ZN(n17318) );
  AOI22_X1 U20359 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17316) );
  AOI22_X1 U20360 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17312), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17315) );
  AOI22_X1 U20361 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17314) );
  AOI22_X1 U20362 ( .A1(n17266), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17313) );
  NAND4_X1 U20363 ( .A1(n17316), .A2(n17315), .A3(n17314), .A4(n17313), .ZN(
        n17317) );
  NOR3_X1 U20364 ( .A1(n17319), .A2(n17318), .A3(n17317), .ZN(n17979) );
  NOR2_X1 U20365 ( .A1(n17983), .A2(n17979), .ZN(n17978) );
  INV_X1 U20366 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17321) );
  OAI22_X1 U20367 ( .A1(n18077), .A2(n17321), .B1(n9640), .B2(n17320), .ZN(
        n17328) );
  INV_X1 U20368 ( .A(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17326) );
  AOI22_X1 U20369 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17322), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17325) );
  AOI22_X1 U20370 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17324) );
  OAI211_X1 U20371 ( .C1(n18112), .C2(n17326), .A(n17325), .B(n17324), .ZN(
        n17327) );
  AOI211_X1 U20372 ( .C1(n17293), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n17328), .B(n17327), .ZN(n17337) );
  AOI22_X1 U20373 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17336) );
  AOI22_X1 U20374 ( .A1(n13053), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17335) );
  NOR2_X1 U20375 ( .A1(n10444), .A2(n18135), .ZN(n17333) );
  INV_X1 U20376 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17331) );
  INV_X1 U20377 ( .A(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18040) );
  OAI22_X1 U20378 ( .A1(n10446), .A2(n17331), .B1(n13229), .B2(n18040), .ZN(
        n17332) );
  AOI211_X1 U20379 ( .C1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .C2(n17300), .A(
        n17333), .B(n17332), .ZN(n17334) );
  NAND4_X1 U20380 ( .A1(n17337), .A2(n17336), .A3(n17335), .A4(n17334), .ZN(
        n17975) );
  NAND2_X1 U20381 ( .A1(n17978), .A2(n17975), .ZN(n17974) );
  NOR2_X1 U20382 ( .A1(n17974), .A2(n17338), .ZN(n17968) );
  AOI21_X1 U20383 ( .B1(n17338), .B2(n17974), .A(n17968), .ZN(n18170) );
  AOI22_X1 U20384 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17969), .B1(n18170), 
        .B2(n18151), .ZN(n17339) );
  OAI21_X1 U20385 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17340), .A(n17339), .ZN(
        P3_U2675) );
  NAND3_X1 U20386 ( .A1(n17344), .A2(n20462), .A3(n17341), .ZN(n17342) );
  OAI21_X1 U20387 ( .B1(n17344), .B2(n17343), .A(n17342), .ZN(P2_U3595) );
  AND2_X1 U20388 ( .A1(n20615), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U20389 ( .A1(n17345), .A2(n20478), .ZN(P2_U3047) );
  INV_X1 U20390 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17348) );
  AOI22_X1 U20391 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(n20541), .B1(n20532), 
        .B2(n17346), .ZN(n17347) );
  OAI211_X1 U20392 ( .C1(n20565), .C2(n17348), .A(n17347), .B(n20667), .ZN(
        n17353) );
  NAND3_X1 U20393 ( .A1(n20505), .A2(P1_REIP_REG_9__SCAN_IN), .A3(n17356), 
        .ZN(n17349) );
  OAI21_X1 U20394 ( .B1(n17351), .B2(n17350), .A(n17349), .ZN(n17352) );
  AOI211_X1 U20395 ( .C1(n17354), .C2(n20575), .A(n17353), .B(n17352), .ZN(
        n17355) );
  OAI21_X1 U20396 ( .B1(n17357), .B2(n17356), .A(n17355), .ZN(P1_U2830) );
  AOI22_X1 U20397 ( .A1(n20641), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20683), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n17364) );
  NAND2_X1 U20398 ( .A1(n17359), .A2(n17358), .ZN(n17360) );
  XNOR2_X1 U20399 ( .A(n17361), .B(n17360), .ZN(n17391) );
  INV_X1 U20400 ( .A(n17362), .ZN(n20528) );
  AOI22_X1 U20401 ( .A1(n17391), .A2(n20650), .B1(n20528), .B2(n20649), .ZN(
        n17363) );
  OAI211_X1 U20402 ( .C1(n20654), .C2(n20521), .A(n17364), .B(n17363), .ZN(
        P1_U2992) );
  INV_X1 U20403 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n17365) );
  NOR2_X1 U20404 ( .A1(n20667), .A2(n17365), .ZN(n17398) );
  AOI21_X1 U20405 ( .B1(n20641), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n17398), .ZN(n17370) );
  XNOR2_X1 U20406 ( .A(n17366), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17367) );
  XNOR2_X1 U20407 ( .A(n17368), .B(n17367), .ZN(n17400) );
  AOI22_X1 U20408 ( .A1(n20591), .A2(n20649), .B1(n17400), .B2(n20650), .ZN(
        n17369) );
  OAI211_X1 U20409 ( .C1(n20654), .C2(n20534), .A(n17370), .B(n17369), .ZN(
        P1_U2993) );
  AOI21_X1 U20410 ( .B1(n20641), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n17371), .ZN(n17376) );
  INV_X1 U20411 ( .A(n17372), .ZN(n17374) );
  INV_X1 U20412 ( .A(n17373), .ZN(n20546) );
  AOI22_X1 U20413 ( .A1(n17374), .A2(n20650), .B1(n20649), .B2(n20546), .ZN(
        n17375) );
  OAI211_X1 U20414 ( .C1(n20654), .C2(n20543), .A(n17376), .B(n17375), .ZN(
        P1_U2994) );
  INV_X1 U20415 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17389) );
  OAI21_X1 U20416 ( .B1(n17379), .B2(n17378), .A(n17377), .ZN(n17399) );
  AOI21_X1 U20417 ( .B1(n17389), .B2(n20702), .A(n17399), .ZN(n17393) );
  INV_X1 U20418 ( .A(n17380), .ZN(n17381) );
  AOI21_X1 U20419 ( .B1(n17382), .B2(n20696), .A(n17381), .ZN(n17387) );
  NAND2_X1 U20420 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17384) );
  INV_X1 U20421 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17394) );
  AOI211_X1 U20422 ( .C1(n17388), .C2(n17394), .A(n17389), .B(n17403), .ZN(
        n17383) );
  AOI22_X1 U20423 ( .A1(n17385), .A2(n20699), .B1(n17384), .B2(n17383), .ZN(
        n17386) );
  OAI211_X1 U20424 ( .C1(n17393), .C2(n17388), .A(n17387), .B(n17386), .ZN(
        P1_U3023) );
  OR2_X1 U20425 ( .A1(n17389), .A2(n17403), .ZN(n17395) );
  INV_X1 U20426 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21438) );
  OAI22_X1 U20427 ( .A1(n20668), .A2(n20526), .B1(n21438), .B2(n20667), .ZN(
        n17390) );
  AOI21_X1 U20428 ( .B1(n17391), .B2(n20699), .A(n17390), .ZN(n17392) );
  OAI221_X1 U20429 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17395), .C1(
        n17394), .C2(n17393), .A(n17392), .ZN(P1_U3024) );
  AND2_X1 U20430 ( .A1(n14193), .A2(n17396), .ZN(n17397) );
  AOI21_X1 U20431 ( .B1(n20696), .B2(n10449), .A(n17398), .ZN(n17402) );
  AOI22_X1 U20432 ( .A1(n17400), .A2(n20699), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17399), .ZN(n17401) );
  OAI211_X1 U20433 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n17403), .A(
        n17402), .B(n17401), .ZN(P1_U3025) );
  AOI22_X1 U20434 ( .A1(n19724), .A2(n19651), .B1(n17404), .B2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17412) );
  AOI21_X1 U20435 ( .B1(n19712), .B2(n17406), .A(n17405), .ZN(n17407) );
  OAI21_X1 U20436 ( .B1(n19706), .B2(n17408), .A(n17407), .ZN(n17409) );
  AOI21_X1 U20437 ( .B1(n19721), .B2(n17410), .A(n17409), .ZN(n17411) );
  OAI211_X1 U20438 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n17413), .A(
        n17412), .B(n17411), .ZN(P2_U3046) );
  INV_X1 U20439 ( .A(n17414), .ZN(n17429) );
  INV_X1 U20440 ( .A(n17415), .ZN(n17420) );
  INV_X1 U20441 ( .A(n17416), .ZN(n17417) );
  AOI211_X1 U20442 ( .C1(n17420), .C2(n17419), .A(n17418), .B(n17417), .ZN(
        n17427) );
  OAI21_X1 U20443 ( .B1(n17422), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n17421), 
        .ZN(n17424) );
  NAND2_X1 U20444 ( .A1(n17425), .A2(n20381), .ZN(n17423) );
  AOI22_X1 U20445 ( .A1(n17425), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n17424), 
        .B2(n17423), .ZN(n17426) );
  OAI211_X1 U20446 ( .C1(n17429), .C2(n17428), .A(n17427), .B(n17426), .ZN(
        P2_U3176) );
  NOR3_X1 U20447 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n17431) );
  NOR4_X1 U20448 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17430) );
  NAND4_X1 U20449 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17431), .A3(n17430), .A4(
        U215), .ZN(U213) );
  INV_X1 U20450 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19657) );
  INV_X2 U20451 ( .A(U214), .ZN(n17473) );
  NOR2_X2 U20452 ( .A1(n17473), .A2(n17432), .ZN(n17475) );
  INV_X1 U20453 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17511) );
  OAI222_X1 U20454 ( .A1(U212), .A2(n19657), .B1(n17472), .B2(n17433), .C1(
        U214), .C2(n17511), .ZN(U216) );
  AOI222_X1 U20455 ( .A1(n17470), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n17475), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n17473), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n17434) );
  INV_X1 U20456 ( .A(n17434), .ZN(U217) );
  AOI22_X1 U20457 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17470), .ZN(n17435) );
  OAI21_X1 U20458 ( .B1(n16049), .B2(n17472), .A(n17435), .ZN(U218) );
  INV_X1 U20459 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n17437) );
  AOI22_X1 U20460 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17470), .ZN(n17436) );
  OAI21_X1 U20461 ( .B1(n17437), .B2(n17472), .A(n17436), .ZN(U219) );
  AOI22_X1 U20462 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17470), .ZN(n17438) );
  OAI21_X1 U20463 ( .B1(n16065), .B2(n17472), .A(n17438), .ZN(U220) );
  AOI22_X1 U20464 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17470), .ZN(n17439) );
  OAI21_X1 U20465 ( .B1(n17440), .B2(n17472), .A(n17439), .ZN(U221) );
  AOI22_X1 U20466 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n17470), .ZN(n17441) );
  OAI21_X1 U20467 ( .B1(n16079), .B2(n17472), .A(n17441), .ZN(U222) );
  INV_X1 U20468 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n17443) );
  AOI22_X1 U20469 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n17470), .ZN(n17442) );
  OAI21_X1 U20470 ( .B1(n17443), .B2(n17472), .A(n17442), .ZN(U223) );
  AOI22_X1 U20471 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17470), .ZN(n17444) );
  OAI21_X1 U20472 ( .B1(n16091), .B2(n17472), .A(n17444), .ZN(U224) );
  AOI22_X1 U20473 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n17470), .ZN(n17445) );
  OAI21_X1 U20474 ( .B1(n16097), .B2(n17472), .A(n17445), .ZN(U225) );
  AOI22_X1 U20475 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n17470), .ZN(n17446) );
  OAI21_X1 U20476 ( .B1(n16103), .B2(n17472), .A(n17446), .ZN(U226) );
  AOI22_X1 U20477 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17470), .ZN(n17447) );
  OAI21_X1 U20478 ( .B1(n16110), .B2(n17472), .A(n17447), .ZN(U227) );
  AOI22_X1 U20479 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17470), .ZN(n17448) );
  OAI21_X1 U20480 ( .B1(n16118), .B2(n17472), .A(n17448), .ZN(U228) );
  AOI22_X1 U20481 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n17470), .ZN(n17449) );
  OAI21_X1 U20482 ( .B1(n17450), .B2(n17472), .A(n17449), .ZN(U229) );
  AOI22_X1 U20483 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n17470), .ZN(n17451) );
  OAI21_X1 U20484 ( .B1(n16130), .B2(n17472), .A(n17451), .ZN(U230) );
  INV_X1 U20485 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n21452) );
  AOI22_X1 U20486 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n17475), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n17473), .ZN(n17452) );
  OAI21_X1 U20487 ( .B1(n21452), .B2(U212), .A(n17452), .ZN(U231) );
  INV_X1 U20488 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n17454) );
  AOI22_X1 U20489 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n17475), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n17473), .ZN(n17453) );
  OAI21_X1 U20490 ( .B1(n17454), .B2(U212), .A(n17453), .ZN(U232) );
  INV_X1 U20491 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n21493) );
  AOI22_X1 U20492 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n17475), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n17473), .ZN(n17455) );
  OAI21_X1 U20493 ( .B1(n21493), .B2(U212), .A(n17455), .ZN(U233) );
  INV_X1 U20494 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n17492) );
  AOI22_X1 U20495 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n17475), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n17473), .ZN(n17456) );
  OAI21_X1 U20496 ( .B1(n17492), .B2(U212), .A(n17456), .ZN(U234) );
  AOI22_X1 U20497 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n17470), .ZN(n17457) );
  OAI21_X1 U20498 ( .B1(n17458), .B2(n17472), .A(n17457), .ZN(U235) );
  INV_X1 U20499 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n17489) );
  AOI22_X1 U20500 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n17475), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n17473), .ZN(n17459) );
  OAI21_X1 U20501 ( .B1(n17489), .B2(U212), .A(n17459), .ZN(U236) );
  AOI22_X1 U20502 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n17470), .ZN(n17460) );
  OAI21_X1 U20503 ( .B1(n17461), .B2(n17472), .A(n17460), .ZN(U237) );
  INV_X1 U20504 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n17486) );
  AOI22_X1 U20505 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n17475), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n17473), .ZN(n17462) );
  OAI21_X1 U20506 ( .B1(n17486), .B2(U212), .A(n17462), .ZN(U238) );
  AOI222_X1 U20507 ( .A1(n17470), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n17475), 
        .B2(BUF1_REG_8__SCAN_IN), .C1(n17473), .C2(P1_DATAO_REG_8__SCAN_IN), 
        .ZN(n17463) );
  INV_X1 U20508 ( .A(n17463), .ZN(U239) );
  INV_X1 U20509 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n17484) );
  AOI22_X1 U20510 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n17475), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n17473), .ZN(n17464) );
  OAI21_X1 U20511 ( .B1(n17484), .B2(U212), .A(n17464), .ZN(U240) );
  AOI22_X1 U20512 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n17470), .ZN(n17465) );
  OAI21_X1 U20513 ( .B1(n13257), .B2(n17472), .A(n17465), .ZN(U241) );
  INV_X1 U20514 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n17482) );
  AOI22_X1 U20515 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n17475), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n17473), .ZN(n17466) );
  OAI21_X1 U20516 ( .B1(n17482), .B2(U212), .A(n17466), .ZN(U242) );
  INV_X1 U20517 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n17468) );
  AOI22_X1 U20518 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n17470), .ZN(n17467) );
  OAI21_X1 U20519 ( .B1(n17468), .B2(n17472), .A(n17467), .ZN(U243) );
  INV_X1 U20520 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n17480) );
  AOI22_X1 U20521 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n17475), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n17473), .ZN(n17469) );
  OAI21_X1 U20522 ( .B1(n17480), .B2(U212), .A(n17469), .ZN(U244) );
  AOI22_X1 U20523 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n17473), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n17470), .ZN(n17471) );
  OAI21_X1 U20524 ( .B1(n13855), .B2(n17472), .A(n17471), .ZN(U245) );
  INV_X1 U20525 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n17478) );
  AOI22_X1 U20526 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n17475), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n17473), .ZN(n17474) );
  OAI21_X1 U20527 ( .B1(n17478), .B2(U212), .A(n17474), .ZN(U246) );
  INV_X1 U20528 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n17477) );
  AOI22_X1 U20529 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n17475), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n17473), .ZN(n17476) );
  OAI21_X1 U20530 ( .B1(n17477), .B2(U212), .A(n17476), .ZN(U247) );
  AOI22_X1 U20531 ( .A1(n17509), .A2(n17477), .B1(n13222), .B2(U215), .ZN(U251) );
  INV_X1 U20532 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18986) );
  AOI22_X1 U20533 ( .A1(n17509), .A2(n17478), .B1(n18986), .B2(U215), .ZN(U252) );
  OAI22_X1 U20534 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n17509), .ZN(n17479) );
  INV_X1 U20535 ( .A(n17479), .ZN(U253) );
  AOI22_X1 U20536 ( .A1(n17509), .A2(n17480), .B1(n18993), .B2(U215), .ZN(U254) );
  OAI22_X1 U20537 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n17509), .ZN(n17481) );
  INV_X1 U20538 ( .A(n17481), .ZN(U255) );
  AOI22_X1 U20539 ( .A1(n17497), .A2(n17482), .B1(n19002), .B2(U215), .ZN(U256) );
  OAI22_X1 U20540 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n17509), .ZN(n17483) );
  INV_X1 U20541 ( .A(n17483), .ZN(U257) );
  AOI22_X1 U20542 ( .A1(n17509), .A2(n17484), .B1(n19012), .B2(U215), .ZN(U258) );
  INV_X1 U20543 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n21420) );
  INV_X1 U20544 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n18254) );
  AOI22_X1 U20545 ( .A1(n17509), .A2(n21420), .B1(n18254), .B2(U215), .ZN(U259) );
  AOI22_X1 U20546 ( .A1(n17497), .A2(n17486), .B1(n17485), .B2(U215), .ZN(U260) );
  OAI22_X1 U20547 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n17497), .ZN(n17487) );
  INV_X1 U20548 ( .A(n17487), .ZN(U261) );
  AOI22_X1 U20549 ( .A1(n17509), .A2(n17489), .B1(n17488), .B2(U215), .ZN(U262) );
  OAI22_X1 U20550 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n17497), .ZN(n17490) );
  INV_X1 U20551 ( .A(n17490), .ZN(U263) );
  AOI22_X1 U20552 ( .A1(n17497), .A2(n17492), .B1(n17491), .B2(U215), .ZN(U264) );
  OAI22_X1 U20553 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17497), .ZN(n17493) );
  INV_X1 U20554 ( .A(n17493), .ZN(U265) );
  OAI22_X1 U20555 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n17497), .ZN(n17494) );
  INV_X1 U20556 ( .A(n17494), .ZN(U266) );
  AOI22_X1 U20557 ( .A1(n17497), .A2(n21452), .B1(n16849), .B2(U215), .ZN(U267) );
  OAI22_X1 U20558 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17497), .ZN(n17495) );
  INV_X1 U20559 ( .A(n17495), .ZN(U268) );
  OAI22_X1 U20560 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17509), .ZN(n17496) );
  INV_X1 U20561 ( .A(n17496), .ZN(U269) );
  OAI22_X1 U20562 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17497), .ZN(n17498) );
  INV_X1 U20563 ( .A(n17498), .ZN(U270) );
  OAI22_X1 U20564 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17509), .ZN(n17499) );
  INV_X1 U20565 ( .A(n17499), .ZN(U271) );
  OAI22_X1 U20566 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17509), .ZN(n17500) );
  INV_X1 U20567 ( .A(n17500), .ZN(U272) );
  OAI22_X1 U20568 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n17509), .ZN(n17501) );
  INV_X1 U20569 ( .A(n17501), .ZN(U273) );
  OAI22_X1 U20570 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17509), .ZN(n17502) );
  INV_X1 U20571 ( .A(n17502), .ZN(U274) );
  OAI22_X1 U20572 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17509), .ZN(n17503) );
  INV_X1 U20573 ( .A(n17503), .ZN(U275) );
  OAI22_X1 U20574 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17509), .ZN(n17504) );
  INV_X1 U20575 ( .A(n17504), .ZN(U276) );
  OAI22_X1 U20576 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17509), .ZN(n17505) );
  INV_X1 U20577 ( .A(n17505), .ZN(U277) );
  OAI22_X1 U20578 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17509), .ZN(n17506) );
  INV_X1 U20579 ( .A(n17506), .ZN(U278) );
  OAI22_X1 U20580 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17509), .ZN(n17507) );
  INV_X1 U20581 ( .A(n17507), .ZN(U279) );
  OAI22_X1 U20582 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17509), .ZN(n17508) );
  INV_X1 U20583 ( .A(n17508), .ZN(U280) );
  INV_X1 U20584 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19661) );
  INV_X1 U20585 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19006) );
  AOI22_X1 U20586 ( .A1(n17509), .A2(n19661), .B1(n19006), .B2(U215), .ZN(U281) );
  INV_X1 U20587 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19014) );
  AOI22_X1 U20588 ( .A1(n17509), .A2(n19657), .B1(n19014), .B2(U215), .ZN(U282) );
  INV_X1 U20589 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17510) );
  AOI222_X1 U20590 ( .A1(n17511), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19657), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17510), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n17512) );
  INV_X2 U20591 ( .A(n17514), .ZN(n17513) );
  INV_X1 U20592 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19485) );
  INV_X1 U20593 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20408) );
  AOI22_X1 U20594 ( .A1(n17513), .A2(n19485), .B1(n20408), .B2(n17514), .ZN(
        U347) );
  INV_X1 U20595 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19484) );
  INV_X1 U20596 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20407) );
  AOI22_X1 U20597 ( .A1(n17513), .A2(n19484), .B1(n20407), .B2(n17514), .ZN(
        U348) );
  INV_X1 U20598 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19481) );
  INV_X1 U20599 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20405) );
  AOI22_X1 U20600 ( .A1(n17513), .A2(n19481), .B1(n20405), .B2(n17514), .ZN(
        U349) );
  INV_X1 U20601 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19480) );
  INV_X1 U20602 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20403) );
  AOI22_X1 U20603 ( .A1(n17513), .A2(n19480), .B1(n20403), .B2(n17514), .ZN(
        U350) );
  INV_X1 U20604 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19478) );
  INV_X1 U20605 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20401) );
  AOI22_X1 U20606 ( .A1(n17513), .A2(n19478), .B1(n20401), .B2(n17514), .ZN(
        U351) );
  INV_X1 U20607 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19476) );
  INV_X1 U20608 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20399) );
  AOI22_X1 U20609 ( .A1(n17513), .A2(n19476), .B1(n20399), .B2(n17514), .ZN(
        U352) );
  INV_X1 U20610 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19474) );
  INV_X1 U20611 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20397) );
  AOI22_X1 U20612 ( .A1(n17513), .A2(n19474), .B1(n20397), .B2(n17514), .ZN(
        U353) );
  INV_X1 U20613 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19471) );
  AOI22_X1 U20614 ( .A1(n17513), .A2(n19471), .B1(n20395), .B2(n17514), .ZN(
        U354) );
  INV_X1 U20615 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19525) );
  INV_X1 U20616 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20447) );
  AOI22_X1 U20617 ( .A1(n17513), .A2(n19525), .B1(n20447), .B2(n17514), .ZN(
        U355) );
  INV_X1 U20618 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19521) );
  INV_X1 U20619 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20442) );
  AOI22_X1 U20620 ( .A1(n17513), .A2(n19521), .B1(n20442), .B2(n17514), .ZN(
        U356) );
  INV_X1 U20621 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19518) );
  INV_X1 U20622 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20440) );
  AOI22_X1 U20623 ( .A1(n17513), .A2(n19518), .B1(n20440), .B2(n17514), .ZN(
        U357) );
  INV_X1 U20624 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19517) );
  INV_X1 U20625 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20437) );
  AOI22_X1 U20626 ( .A1(n17513), .A2(n19517), .B1(n20437), .B2(n17514), .ZN(
        U358) );
  INV_X1 U20627 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n21507) );
  INV_X1 U20628 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20436) );
  AOI22_X1 U20629 ( .A1(n17513), .A2(n21507), .B1(n20436), .B2(n17514), .ZN(
        U359) );
  INV_X1 U20630 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19516) );
  INV_X1 U20631 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20434) );
  AOI22_X1 U20632 ( .A1(n17513), .A2(n19516), .B1(n20434), .B2(n17514), .ZN(
        U360) );
  INV_X1 U20633 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19514) );
  INV_X1 U20634 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20432) );
  AOI22_X1 U20635 ( .A1(n17513), .A2(n19514), .B1(n20432), .B2(n17514), .ZN(
        U361) );
  INV_X1 U20636 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19512) );
  INV_X1 U20637 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20430) );
  AOI22_X1 U20638 ( .A1(n17513), .A2(n19512), .B1(n20430), .B2(n17514), .ZN(
        U362) );
  INV_X1 U20639 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19510) );
  INV_X1 U20640 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20428) );
  AOI22_X1 U20641 ( .A1(n17513), .A2(n19510), .B1(n20428), .B2(n17514), .ZN(
        U363) );
  INV_X1 U20642 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19508) );
  INV_X1 U20643 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20427) );
  AOI22_X1 U20644 ( .A1(n17513), .A2(n19508), .B1(n20427), .B2(n17514), .ZN(
        U364) );
  INV_X1 U20645 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19470) );
  INV_X1 U20646 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20393) );
  AOI22_X1 U20647 ( .A1(n17513), .A2(n19470), .B1(n20393), .B2(n17514), .ZN(
        U365) );
  INV_X1 U20648 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19505) );
  INV_X1 U20649 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20425) );
  AOI22_X1 U20650 ( .A1(n17513), .A2(n19505), .B1(n20425), .B2(n17514), .ZN(
        U366) );
  INV_X1 U20651 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19503) );
  INV_X1 U20652 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20424) );
  AOI22_X1 U20653 ( .A1(n17513), .A2(n19503), .B1(n20424), .B2(n17514), .ZN(
        U367) );
  INV_X1 U20654 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19502) );
  INV_X1 U20655 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20422) );
  AOI22_X1 U20656 ( .A1(n17513), .A2(n19502), .B1(n20422), .B2(n17514), .ZN(
        U368) );
  INV_X1 U20657 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19499) );
  INV_X1 U20658 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20421) );
  AOI22_X1 U20659 ( .A1(n17513), .A2(n19499), .B1(n20421), .B2(n17514), .ZN(
        U369) );
  INV_X1 U20660 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19498) );
  INV_X1 U20661 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20419) );
  AOI22_X1 U20662 ( .A1(n17513), .A2(n19498), .B1(n20419), .B2(n17514), .ZN(
        U370) );
  INV_X1 U20663 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19496) );
  INV_X1 U20664 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20417) );
  AOI22_X1 U20665 ( .A1(n17513), .A2(n19496), .B1(n20417), .B2(n17514), .ZN(
        U371) );
  INV_X1 U20666 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19493) );
  INV_X1 U20667 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20415) );
  AOI22_X1 U20668 ( .A1(n17513), .A2(n19493), .B1(n20415), .B2(n17514), .ZN(
        U372) );
  INV_X1 U20669 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19492) );
  INV_X1 U20670 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20414) );
  AOI22_X1 U20671 ( .A1(n17513), .A2(n19492), .B1(n20414), .B2(n17514), .ZN(
        U373) );
  INV_X1 U20672 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19490) );
  INV_X1 U20673 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20412) );
  AOI22_X1 U20674 ( .A1(n17513), .A2(n19490), .B1(n20412), .B2(n17514), .ZN(
        U374) );
  INV_X1 U20675 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19488) );
  INV_X1 U20676 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20410) );
  AOI22_X1 U20677 ( .A1(n17513), .A2(n19488), .B1(n20410), .B2(n17514), .ZN(
        U375) );
  INV_X1 U20678 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19467) );
  INV_X1 U20679 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20392) );
  AOI22_X1 U20680 ( .A1(n17513), .A2(n19467), .B1(n20392), .B2(n17514), .ZN(
        U376) );
  INV_X1 U20681 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19464) );
  NOR2_X1 U20682 ( .A1(n19452), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19454) );
  OAI22_X1 U20683 ( .A1(n19464), .A2(n19454), .B1(n19452), .B2(
        P3_STATE_REG_0__SCAN_IN), .ZN(n19448) );
  INV_X1 U20684 ( .A(n19448), .ZN(n19536) );
  AOI21_X1 U20685 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19536), .ZN(n17515) );
  INV_X1 U20686 ( .A(n17515), .ZN(P3_U2633) );
  NOR2_X1 U20687 ( .A1(n18295), .A2(n17523), .ZN(n17516) );
  OAI21_X1 U20688 ( .B1(n17516), .B2(n18293), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17517) );
  OAI21_X1 U20689 ( .B1(n17519), .B2(n17518), .A(n17517), .ZN(P3_U2634) );
  INV_X1 U20690 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19466) );
  AOI21_X1 U20691 ( .B1(n19464), .B2(n19466), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17520) );
  AOI22_X1 U20692 ( .A1(n19531), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17520), 
        .B2(n19568), .ZN(P3_U2635) );
  OAI21_X1 U20693 ( .B1(n19450), .B2(BS16), .A(n19536), .ZN(n19534) );
  OAI21_X1 U20694 ( .B1(n19536), .B2(n17521), .A(n19534), .ZN(P3_U2636) );
  OAI211_X1 U20695 ( .C1(n18295), .C2(n17523), .A(n17522), .B(n19401), .ZN(
        n19422) );
  NAND2_X1 U20696 ( .A1(n19561), .A2(n19422), .ZN(n19550) );
  INV_X1 U20697 ( .A(n19550), .ZN(n19552) );
  OAI21_X1 U20698 ( .B1(n19552), .B2(n17525), .A(n17524), .ZN(P3_U2637) );
  NOR4_X1 U20699 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n17529) );
  NOR4_X1 U20700 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n17528) );
  NOR4_X1 U20701 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17527) );
  NOR4_X1 U20702 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n17526) );
  NAND4_X1 U20703 ( .A1(n17529), .A2(n17528), .A3(n17527), .A4(n17526), .ZN(
        n17535) );
  NOR4_X1 U20704 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17533) );
  AOI211_X1 U20705 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_8__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17532) );
  NOR4_X1 U20706 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n17531) );
  NOR4_X1 U20707 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n17530) );
  NAND4_X1 U20708 ( .A1(n17533), .A2(n17532), .A3(n17531), .A4(n17530), .ZN(
        n17534) );
  NOR2_X1 U20709 ( .A1(n17535), .A2(n17534), .ZN(n19548) );
  INV_X1 U20710 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17537) );
  NOR3_X1 U20711 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A3(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n17538) );
  OAI21_X1 U20712 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17538), .A(n19548), .ZN(
        n17536) );
  OAI21_X1 U20713 ( .B1(n19548), .B2(n17537), .A(n17536), .ZN(P3_U2638) );
  INV_X1 U20714 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19541) );
  INV_X1 U20715 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19535) );
  AOI21_X1 U20716 ( .B1(n19541), .B2(n19535), .A(n17538), .ZN(n17540) );
  INV_X1 U20717 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17539) );
  INV_X1 U20718 ( .A(n19548), .ZN(n19543) );
  AOI22_X1 U20719 ( .A1(n19548), .A2(n17540), .B1(n17539), .B2(n19543), .ZN(
        P3_U2639) );
  INV_X1 U20720 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17867) );
  NAND2_X1 U20721 ( .A1(n17878), .A2(n17867), .ZN(n17865) );
  INV_X1 U20722 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17848) );
  NAND2_X1 U20723 ( .A1(n17852), .A2(n17848), .ZN(n17845) );
  NAND2_X1 U20724 ( .A1(n17823), .A2(n17816), .ZN(n17815) );
  INV_X1 U20725 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17792) );
  NAND2_X1 U20726 ( .A1(n17802), .A2(n17792), .ZN(n17791) );
  NAND2_X1 U20727 ( .A1(n17772), .A2(n17767), .ZN(n17766) );
  NOR2_X2 U20728 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17766), .ZN(n17748) );
  NAND2_X1 U20729 ( .A1(n17748), .A2(n17736), .ZN(n17735) );
  NOR2_X2 U20730 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17735), .ZN(n17727) );
  NAND2_X1 U20731 ( .A1(n17727), .A2(n17717), .ZN(n17716) );
  INV_X1 U20732 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n21434) );
  NAND2_X1 U20733 ( .A1(n17696), .A2(n21434), .ZN(n17693) );
  INV_X1 U20734 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17667) );
  NAND2_X1 U20735 ( .A1(n17678), .A2(n17667), .ZN(n17666) );
  NAND2_X1 U20736 ( .A1(n17654), .A2(n17987), .ZN(n17647) );
  NAND2_X1 U20737 ( .A1(n17627), .A2(n17626), .ZN(n17611) );
  INV_X1 U20738 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17602) );
  NAND2_X1 U20739 ( .A1(n17610), .A2(n17602), .ZN(n17601) );
  NAND2_X1 U20740 ( .A1(n17587), .A2(n17970), .ZN(n17566) );
  NOR2_X1 U20741 ( .A1(n17926), .A2(n17566), .ZN(n17573) );
  INV_X1 U20742 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17547) );
  INV_X1 U20743 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19526) );
  NAND2_X1 U20744 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n17593) );
  INV_X1 U20745 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19509) );
  INV_X1 U20746 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19507) );
  NOR4_X1 U20747 ( .A1(n19513), .A2(n19511), .A3(n19509), .A4(n19507), .ZN(
        n17553) );
  INV_X1 U20748 ( .A(n17553), .ZN(n17543) );
  INV_X1 U20749 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19489) );
  NAND3_X1 U20750 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .ZN(n17797) );
  INV_X1 U20751 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19486) );
  NOR2_X1 U20752 ( .A1(n19486), .A2(n19483), .ZN(n17785) );
  INV_X1 U20753 ( .A(n17785), .ZN(n17807) );
  NOR3_X1 U20754 ( .A1(n17885), .A2(n17797), .A3(n17807), .ZN(n17541) );
  NAND4_X1 U20755 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(P3_REIP_REG_5__SCAN_IN), 
        .A3(P3_REIP_REG_4__SCAN_IN), .A4(n17541), .ZN(n17771) );
  NOR2_X1 U20756 ( .A1(n19489), .A2(n17771), .ZN(n17749) );
  NAND2_X1 U20757 ( .A1(n17902), .A2(n17623), .ZN(n17741) );
  INV_X1 U20758 ( .A(n17741), .ZN(n17542) );
  INV_X1 U20759 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19506) );
  INV_X1 U20760 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19500) );
  NAND2_X1 U20761 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n17708) );
  NOR2_X1 U20762 ( .A1(n19500), .A2(n17708), .ZN(n17549) );
  NAND3_X1 U20763 ( .A1(n17549), .A2(P3_REIP_REG_19__SCAN_IN), .A3(
        P3_REIP_REG_18__SCAN_IN), .ZN(n17551) );
  NOR2_X1 U20764 ( .A1(n19506), .A2(n17551), .ZN(n17621) );
  NAND2_X1 U20765 ( .A1(n17542), .A2(n17621), .ZN(n17673) );
  NOR2_X1 U20766 ( .A1(n17543), .A2(n17673), .ZN(n17625) );
  NAND3_X1 U20767 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n17625), .ZN(n17592) );
  NOR2_X1 U20768 ( .A1(n17593), .A2(n17592), .ZN(n17579) );
  NAND2_X1 U20769 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17579), .ZN(n17548) );
  NOR3_X1 U20770 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19526), .A3(n17548), 
        .ZN(n17546) );
  OAI22_X1 U20771 ( .A1(n10163), .A2(n17880), .B1(n17544), .B2(n17927), .ZN(
        n17545) );
  AOI211_X1 U20772 ( .C1(n17573), .C2(n17547), .A(n17546), .B(n17545), .ZN(
        n17565) );
  NOR2_X1 U20773 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n17548), .ZN(n17571) );
  INV_X1 U20774 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19515) );
  NOR2_X1 U20775 ( .A1(n17194), .A2(n19515), .ZN(n17552) );
  NAND2_X1 U20776 ( .A1(n17623), .A2(n17899), .ZN(n17750) );
  INV_X1 U20777 ( .A(n17549), .ZN(n17685) );
  NOR2_X1 U20778 ( .A1(n17750), .A2(n17685), .ZN(n17698) );
  INV_X1 U20779 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19504) );
  INV_X1 U20780 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19501) );
  NOR2_X1 U20781 ( .A1(n19504), .A2(n19501), .ZN(n17550) );
  AOI21_X1 U20782 ( .B1(n17698), .B2(n17550), .A(n17699), .ZN(n17674) );
  NOR3_X1 U20783 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n17741), .A3(n17551), 
        .ZN(n17680) );
  NOR2_X1 U20784 ( .A1(n17674), .A2(n17680), .ZN(n17672) );
  OAI221_X1 U20785 ( .B1(n17699), .B2(n17553), .C1(n17699), .C2(n17552), .A(
        n17672), .ZN(n17609) );
  AOI221_X1 U20786 ( .B1(n19520), .B2(n17902), .C1(n17593), .C2(n17902), .A(
        n17609), .ZN(n17569) );
  INV_X1 U20787 ( .A(n17569), .ZN(n17578) );
  OAI21_X1 U20788 ( .B1(n17571), .B2(n17578), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n17564) );
  NOR2_X1 U20789 ( .A1(n17862), .A2(n19443), .ZN(n17915) );
  NAND2_X1 U20790 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18357), .ZN(
        n17555) );
  AOI21_X1 U20791 ( .B1(n10167), .B2(n17555), .A(n17554), .ZN(n18358) );
  INV_X1 U20792 ( .A(n18358), .ZN(n17616) );
  INV_X1 U20793 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18385) );
  NOR3_X1 U20794 ( .A1(n18684), .A2(n18372), .A3(n18385), .ZN(n17556) );
  OAI21_X1 U20795 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17556), .A(
        n17555), .ZN(n18375) );
  NOR2_X1 U20796 ( .A1(n18684), .A2(n18372), .ZN(n17558) );
  INV_X1 U20797 ( .A(n17556), .ZN(n17557) );
  OAI21_X1 U20798 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17558), .A(
        n17557), .ZN(n18396) );
  OAI21_X1 U20799 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17560), .A(
        n17559), .ZN(n18409) );
  INV_X1 U20800 ( .A(n18403), .ZN(n17686) );
  NOR2_X1 U20801 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17732), .ZN(
        n17712) );
  OAI21_X1 U20802 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18403), .A(
        n17561), .ZN(n18425) );
  NAND2_X1 U20803 ( .A1(n17682), .A2(n18425), .ZN(n17681) );
  AOI21_X1 U20804 ( .B1(n18416), .B2(n17561), .A(n17560), .ZN(n17562) );
  INV_X1 U20805 ( .A(n17562), .ZN(n18413) );
  NAND2_X1 U20806 ( .A1(n17744), .A2(n17664), .ZN(n17661) );
  NAND2_X1 U20807 ( .A1(n18409), .A2(n17661), .ZN(n17660) );
  NAND2_X1 U20808 ( .A1(n17744), .A2(n17660), .ZN(n17649) );
  NAND2_X1 U20809 ( .A1(n17650), .A2(n17649), .ZN(n17648) );
  NAND2_X1 U20810 ( .A1(n17744), .A2(n17648), .ZN(n17641) );
  NAND2_X1 U20811 ( .A1(n18396), .A2(n17641), .ZN(n17640) );
  NAND2_X1 U20812 ( .A1(n17744), .A2(n17640), .ZN(n17629) );
  NAND2_X1 U20813 ( .A1(n18375), .A2(n17629), .ZN(n17628) );
  NAND2_X1 U20814 ( .A1(n17744), .A2(n17628), .ZN(n17615) );
  NAND2_X1 U20815 ( .A1(n17616), .A2(n17615), .ZN(n17614) );
  NAND2_X1 U20816 ( .A1(n17744), .A2(n17614), .ZN(n17604) );
  NAND2_X1 U20817 ( .A1(n17605), .A2(n17604), .ZN(n17603) );
  NAND2_X1 U20818 ( .A1(n17744), .A2(n17603), .ZN(n17590) );
  NAND2_X1 U20819 ( .A1(n17591), .A2(n17590), .ZN(n17589) );
  NAND2_X1 U20820 ( .A1(n17744), .A2(n17589), .ZN(n17581) );
  NAND2_X1 U20821 ( .A1(n17582), .A2(n17581), .ZN(n17580) );
  NAND3_X1 U20822 ( .A1(n17915), .A2(n17567), .A3(n17568), .ZN(n17563) );
  NAND3_X1 U20823 ( .A1(n17565), .A2(n17564), .A3(n17563), .ZN(P3_U2640) );
  NAND2_X1 U20824 ( .A1(n17866), .A2(n17566), .ZN(n17585) );
  OAI22_X1 U20825 ( .A1(n17569), .A2(n19526), .B1(n10160), .B2(n17880), .ZN(
        n17570) );
  AOI211_X1 U20826 ( .C1(n17572), .C2(n17829), .A(n17571), .B(n17570), .ZN(
        n17575) );
  OAI21_X1 U20827 ( .B1(n17884), .B2(n17573), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n17574) );
  OAI211_X1 U20828 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n17585), .A(n17575), .B(
        n17574), .ZN(P3_U2641) );
  NOR2_X1 U20829 ( .A1(n17587), .A2(n17970), .ZN(n17586) );
  OAI22_X1 U20830 ( .A1(n17576), .A2(n17880), .B1(n17927), .B2(n17970), .ZN(
        n17577) );
  AOI221_X1 U20831 ( .B1(n17579), .B2(n19520), .C1(n17578), .C2(
        P3_REIP_REG_29__SCAN_IN), .A(n17577), .ZN(n17584) );
  OAI211_X1 U20832 ( .C1(n17582), .C2(n17581), .A(n17909), .B(n17580), .ZN(
        n17583) );
  OAI211_X1 U20833 ( .C1(n17586), .C2(n17585), .A(n17584), .B(n17583), .ZN(
        P3_U2642) );
  AOI22_X1 U20834 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17914), .B1(
        n17884), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17597) );
  AOI211_X1 U20835 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17601), .A(n17587), .B(
        n17926), .ZN(n17588) );
  AOI21_X1 U20836 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(n17609), .A(n17588), 
        .ZN(n17596) );
  OAI211_X1 U20837 ( .C1(n17591), .C2(n17590), .A(n17909), .B(n17589), .ZN(
        n17595) );
  INV_X1 U20838 ( .A(n17592), .ZN(n17600) );
  OAI211_X1 U20839 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n17600), .B(n17593), .ZN(n17594) );
  NAND4_X1 U20840 ( .A1(n17597), .A2(n17596), .A3(n17595), .A4(n17594), .ZN(
        P3_U2643) );
  OAI22_X1 U20841 ( .A1(n17598), .A2(n17880), .B1(n17927), .B2(n17602), .ZN(
        n17599) );
  AOI221_X1 U20842 ( .B1(n17600), .B2(n17052), .C1(n17609), .C2(
        P3_REIP_REG_27__SCAN_IN), .A(n17599), .ZN(n17608) );
  OAI211_X1 U20843 ( .C1(n17610), .C2(n17602), .A(n17866), .B(n17601), .ZN(
        n17607) );
  OAI211_X1 U20844 ( .C1(n17605), .C2(n17604), .A(n17829), .B(n17603), .ZN(
        n17606) );
  NAND3_X1 U20845 ( .A1(n17608), .A2(n17607), .A3(n17606), .ZN(P3_U2644) );
  INV_X1 U20846 ( .A(n17609), .ZN(n17620) );
  AOI21_X1 U20847 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n17625), .A(
        P3_REIP_REG_26__SCAN_IN), .ZN(n17619) );
  AOI211_X1 U20848 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17611), .A(n17610), .B(
        n17926), .ZN(n17613) );
  NOR2_X1 U20849 ( .A1(n10167), .A2(n17880), .ZN(n17612) );
  AOI211_X1 U20850 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17884), .A(n17613), .B(
        n17612), .ZN(n17618) );
  OAI211_X1 U20851 ( .C1(n17616), .C2(n17615), .A(n17909), .B(n17614), .ZN(
        n17617) );
  OAI211_X1 U20852 ( .C1(n17620), .C2(n17619), .A(n17618), .B(n17617), .ZN(
        P3_U2645) );
  NAND2_X1 U20853 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n17658) );
  NOR2_X1 U20854 ( .A1(n19511), .A2(n17658), .ZN(n17622) );
  NAND3_X1 U20855 ( .A1(n17623), .A2(n17622), .A3(n17621), .ZN(n17637) );
  AOI21_X1 U20856 ( .B1(n17902), .B2(n17637), .A(n17929), .ZN(n17644) );
  OAI21_X1 U20857 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n17917), .A(n17644), 
        .ZN(n17624) );
  AOI22_X1 U20858 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17914), .B1(
        P3_REIP_REG_25__SCAN_IN), .B2(n17624), .ZN(n17633) );
  NOR2_X1 U20859 ( .A1(n17627), .A2(n17926), .ZN(n17634) );
  AOI22_X1 U20860 ( .A1(n17634), .A2(n17626), .B1(n17625), .B2(n19515), .ZN(
        n17632) );
  OAI221_X1 U20861 ( .B1(n17884), .B2(n17866), .C1(n17884), .C2(n17627), .A(
        P3_EBX_REG_25__SCAN_IN), .ZN(n17631) );
  OAI211_X1 U20862 ( .C1(n18375), .C2(n17629), .A(n17909), .B(n17628), .ZN(
        n17630) );
  NAND4_X1 U20863 ( .A1(n17633), .A2(n17632), .A3(n17631), .A4(n17630), .ZN(
        P3_U2646) );
  INV_X1 U20864 ( .A(n17634), .ZN(n17635) );
  AOI21_X1 U20865 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17647), .A(n17635), .ZN(
        n17639) );
  NAND2_X1 U20866 ( .A1(n17902), .A2(n19513), .ZN(n17636) );
  OAI22_X1 U20867 ( .A1(n18385), .A2(n17880), .B1(n17637), .B2(n17636), .ZN(
        n17638) );
  AOI211_X1 U20868 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17884), .A(n17639), .B(
        n17638), .ZN(n17643) );
  OAI211_X1 U20869 ( .C1(n18396), .C2(n17641), .A(n17909), .B(n17640), .ZN(
        n17642) );
  OAI211_X1 U20870 ( .C1(n17644), .C2(n19513), .A(n17643), .B(n17642), .ZN(
        P3_U2647) );
  NOR3_X1 U20871 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n17658), .A3(n17673), 
        .ZN(n17646) );
  OAI22_X1 U20872 ( .A1(n17644), .A2(n19511), .B1(n17927), .B2(n17987), .ZN(
        n17645) );
  AOI211_X1 U20873 ( .C1(n17914), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n17646), .B(n17645), .ZN(n17653) );
  OAI211_X1 U20874 ( .C1(n17654), .C2(n17987), .A(n17866), .B(n17647), .ZN(
        n17652) );
  OAI211_X1 U20875 ( .C1(n17650), .C2(n17649), .A(n17829), .B(n17648), .ZN(
        n17651) );
  NAND3_X1 U20876 ( .A1(n17653), .A2(n17652), .A3(n17651), .ZN(P3_U2648) );
  AOI21_X1 U20877 ( .B1(n19509), .B2(n19507), .A(n17673), .ZN(n17659) );
  AOI211_X1 U20878 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17666), .A(n17654), .B(
        n17926), .ZN(n17657) );
  AOI22_X1 U20879 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17914), .B1(
        n17884), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n17655) );
  INV_X1 U20880 ( .A(n17655), .ZN(n17656) );
  AOI211_X1 U20881 ( .C1(n17659), .C2(n17658), .A(n17657), .B(n17656), .ZN(
        n17663) );
  OAI211_X1 U20882 ( .C1(n18409), .C2(n17661), .A(n17829), .B(n17660), .ZN(
        n17662) );
  OAI211_X1 U20883 ( .C1(n17672), .C2(n19509), .A(n17663), .B(n17662), .ZN(
        P3_U2649) );
  AOI22_X1 U20884 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17914), .B1(
        n17884), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n17670) );
  OAI211_X1 U20885 ( .C1(n18413), .C2(n17665), .A(n17829), .B(n17664), .ZN(
        n17669) );
  OAI211_X1 U20886 ( .C1(n17678), .C2(n17667), .A(n17866), .B(n17666), .ZN(
        n17668) );
  AND3_X1 U20887 ( .A1(n17670), .A2(n17669), .A3(n17668), .ZN(n17671) );
  OAI221_X1 U20888 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n17673), .C1(n19507), 
        .C2(n17672), .A(n17671), .ZN(P3_U2650) );
  INV_X1 U20889 ( .A(n17674), .ZN(n17690) );
  AOI21_X1 U20890 ( .B1(n17693), .B2(P3_EBX_REG_20__SCAN_IN), .A(n17926), .ZN(
        n17675) );
  INV_X1 U20891 ( .A(n17675), .ZN(n17677) );
  OAI22_X1 U20892 ( .A1(n17678), .A2(n17677), .B1(n17927), .B2(n17676), .ZN(
        n17679) );
  AOI211_X1 U20893 ( .C1(n17914), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n17680), .B(n17679), .ZN(n17684) );
  OAI211_X1 U20894 ( .C1(n17682), .C2(n18425), .A(n17829), .B(n17681), .ZN(
        n17683) );
  OAI211_X1 U20895 ( .C1(n19506), .C2(n17690), .A(n17684), .B(n17683), .ZN(
        P3_U2651) );
  NOR2_X1 U20896 ( .A1(n17685), .A2(n17741), .ZN(n17705) );
  AOI21_X1 U20897 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n17705), .A(
        P3_REIP_REG_19__SCAN_IN), .ZN(n17691) );
  NAND2_X1 U20898 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18440), .ZN(
        n17700) );
  INV_X1 U20899 ( .A(n17700), .ZN(n17687) );
  AOI21_X1 U20900 ( .B1(n17712), .B2(n17687), .A(n17862), .ZN(n17688) );
  OAI21_X1 U20901 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17687), .A(
        n17686), .ZN(n18443) );
  XOR2_X1 U20902 ( .A(n17688), .B(n18443), .Z(n17689) );
  OAI22_X1 U20903 ( .A1(n17691), .A2(n17690), .B1(n19443), .B2(n17689), .ZN(
        n17692) );
  AOI211_X1 U20904 ( .C1(n17884), .C2(P3_EBX_REG_19__SCAN_IN), .A(n13496), .B(
        n17692), .ZN(n17695) );
  OAI211_X1 U20905 ( .C1(n17696), .C2(n21434), .A(n17866), .B(n17693), .ZN(
        n17694) );
  OAI211_X1 U20906 ( .C1(n17880), .C2(n18441), .A(n17695), .B(n17694), .ZN(
        P3_U2652) );
  INV_X1 U20907 ( .A(n18840), .ZN(n18953) );
  AOI211_X1 U20908 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17716), .A(n17696), .B(
        n17926), .ZN(n17697) );
  AOI211_X1 U20909 ( .C1(n17884), .C2(P3_EBX_REG_18__SCAN_IN), .A(n18953), .B(
        n17697), .ZN(n17707) );
  NOR2_X1 U20910 ( .A1(n17699), .A2(n17698), .ZN(n17714) );
  OAI21_X1 U20911 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18440), .A(
        n17700), .ZN(n18455) );
  NOR2_X1 U20912 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18684), .ZN(
        n17910) );
  INV_X1 U20913 ( .A(n17910), .ZN(n17701) );
  OAI21_X1 U20914 ( .B1(n18454), .B2(n17701), .A(n17744), .ZN(n17703) );
  OAI21_X1 U20915 ( .B1(n18455), .B2(n17703), .A(n17829), .ZN(n17702) );
  AOI21_X1 U20916 ( .B1(n18455), .B2(n17703), .A(n17702), .ZN(n17704) );
  AOI221_X1 U20917 ( .B1(n17714), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n17705), 
        .C2(n19501), .A(n17704), .ZN(n17706) );
  OAI211_X1 U20918 ( .C1(n18458), .C2(n17880), .A(n17707), .B(n17706), .ZN(
        P3_U2653) );
  NOR3_X1 U20919 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n17708), .A3(n17741), 
        .ZN(n17709) );
  AOI211_X1 U20920 ( .C1(n17884), .C2(P3_EBX_REG_17__SCAN_IN), .A(n18953), .B(
        n17709), .ZN(n17721) );
  OAI21_X1 U20921 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17711), .A(
        n17710), .ZN(n18472) );
  AOI21_X1 U20922 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17712), .A(
        n17862), .ZN(n17713) );
  XNOR2_X1 U20923 ( .A(n18472), .B(n17713), .ZN(n17715) );
  AOI22_X1 U20924 ( .A1(n17829), .A2(n17715), .B1(P3_REIP_REG_17__SCAN_IN), 
        .B2(n17714), .ZN(n17720) );
  OAI211_X1 U20925 ( .C1(n17727), .C2(n17717), .A(n17866), .B(n17716), .ZN(
        n17719) );
  NAND2_X1 U20926 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17914), .ZN(
        n17718) );
  NAND4_X1 U20927 ( .A1(n17721), .A2(n17720), .A3(n17719), .A4(n17718), .ZN(
        P3_U2654) );
  INV_X1 U20928 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19495) );
  OAI21_X1 U20929 ( .B1(n17750), .B2(n19495), .A(n17933), .ZN(n17742) );
  NOR3_X1 U20930 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n19495), .A3(n17741), 
        .ZN(n17722) );
  AOI211_X1 U20931 ( .C1(n17884), .C2(P3_EBX_REG_16__SCAN_IN), .A(n18953), .B(
        n17722), .ZN(n17731) );
  INV_X1 U20932 ( .A(n17726), .ZN(n17724) );
  INV_X1 U20933 ( .A(n17725), .ZN(n17723) );
  AOI221_X1 U20934 ( .B1(n17726), .B2(n17725), .C1(n17724), .C2(n17723), .A(
        n19443), .ZN(n17729) );
  AOI211_X1 U20935 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17735), .A(n17727), .B(
        n17926), .ZN(n17728) );
  AOI211_X1 U20936 ( .C1(n17914), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n17729), .B(n17728), .ZN(n17730) );
  OAI211_X1 U20937 ( .C1(n19497), .C2(n17742), .A(n17731), .B(n17730), .ZN(
        P3_U2655) );
  INV_X1 U20938 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18484) );
  OAI21_X1 U20939 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17746), .A(
        n17732), .ZN(n18497) );
  INV_X1 U20940 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18501) );
  INV_X1 U20941 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18533) );
  INV_X1 U20942 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18558) );
  NOR2_X1 U20943 ( .A1(n18558), .A2(n17799), .ZN(n17798) );
  NAND2_X1 U20944 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17798), .ZN(
        n18515) );
  NOR2_X1 U20945 ( .A1(n18533), .A2(n18515), .ZN(n17777) );
  INV_X1 U20946 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17928) );
  NAND2_X1 U20947 ( .A1(n17777), .A2(n17928), .ZN(n17758) );
  INV_X1 U20948 ( .A(n17758), .ZN(n17760) );
  NAND2_X1 U20949 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17760), .ZN(
        n17743) );
  OAI21_X1 U20950 ( .B1(n18501), .B2(n17743), .A(n17744), .ZN(n17734) );
  AOI21_X1 U20951 ( .B1(n18497), .B2(n17734), .A(n19443), .ZN(n17733) );
  OAI21_X1 U20952 ( .B1(n18497), .B2(n17734), .A(n17733), .ZN(n17738) );
  OAI211_X1 U20953 ( .C1(n17748), .C2(n17736), .A(n17866), .B(n17735), .ZN(
        n17737) );
  OAI211_X1 U20954 ( .C1(n17880), .C2(n18484), .A(n17738), .B(n17737), .ZN(
        n17739) );
  AOI211_X1 U20955 ( .C1(n17884), .C2(P3_EBX_REG_15__SCAN_IN), .A(n18953), .B(
        n17739), .ZN(n17740) );
  OAI221_X1 U20956 ( .B1(n17742), .B2(n19495), .C1(n17742), .C2(n17741), .A(
        n17740), .ZN(P3_U2656) );
  NAND2_X1 U20957 ( .A1(n17744), .A2(n17743), .ZN(n17747) );
  NAND2_X1 U20958 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17745), .ZN(
        n17757) );
  AOI21_X1 U20959 ( .B1(n18501), .B2(n17757), .A(n17746), .ZN(n18503) );
  XOR2_X1 U20960 ( .A(n17747), .B(n18503), .Z(n17756) );
  AOI211_X1 U20961 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17766), .A(n17748), .B(
        n17926), .ZN(n17754) );
  INV_X1 U20962 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19491) );
  NAND2_X1 U20963 ( .A1(n17902), .A2(n17749), .ZN(n17762) );
  NOR2_X1 U20964 ( .A1(n19491), .A2(n17762), .ZN(n17751) );
  OAI211_X1 U20965 ( .C1(n17751), .C2(P3_REIP_REG_14__SCAN_IN), .A(n17933), 
        .B(n17750), .ZN(n17752) );
  OAI211_X1 U20966 ( .C1(n18501), .C2(n17880), .A(n17752), .B(n18840), .ZN(
        n17753) );
  AOI211_X1 U20967 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17884), .A(n17754), .B(
        n17753), .ZN(n17755) );
  OAI21_X1 U20968 ( .B1(n17756), .B2(n19443), .A(n17755), .ZN(P3_U2657) );
  OAI21_X1 U20969 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17777), .A(
        n17757), .ZN(n18523) );
  INV_X1 U20970 ( .A(n18523), .ZN(n17770) );
  NAND2_X1 U20971 ( .A1(n17915), .A2(n17758), .ZN(n17776) );
  AOI21_X1 U20972 ( .B1(n17902), .B2(n17771), .A(n17929), .ZN(n17788) );
  OAI21_X1 U20973 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n17917), .A(n17788), 
        .ZN(n17765) );
  AOI22_X1 U20974 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17914), .B1(
        n17884), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n17759) );
  INV_X1 U20975 ( .A(n17759), .ZN(n17764) );
  OAI211_X1 U20976 ( .C1(n17760), .C2(n17862), .A(n17909), .B(n17770), .ZN(
        n17761) );
  OAI211_X1 U20977 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n17762), .A(n18840), 
        .B(n17761), .ZN(n17763) );
  AOI211_X1 U20978 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n17765), .A(n17764), 
        .B(n17763), .ZN(n17769) );
  OAI211_X1 U20979 ( .C1(n17772), .C2(n17767), .A(n17866), .B(n17766), .ZN(
        n17768) );
  OAI211_X1 U20980 ( .C1(n17770), .C2(n17776), .A(n17769), .B(n17768), .ZN(
        P3_U2658) );
  INV_X1 U20981 ( .A(n17771), .ZN(n17775) );
  NOR2_X1 U20982 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17917), .ZN(n17774) );
  AOI211_X1 U20983 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17791), .A(n17772), .B(
        n17926), .ZN(n17773) );
  AOI211_X1 U20984 ( .C1(n17775), .C2(n17774), .A(n13496), .B(n17773), .ZN(
        n17784) );
  INV_X1 U20985 ( .A(n17776), .ZN(n17782) );
  AOI21_X1 U20986 ( .B1(n18533), .B2(n18515), .A(n17777), .ZN(n17778) );
  INV_X1 U20987 ( .A(n17778), .ZN(n18529) );
  OAI21_X1 U20988 ( .B1(n17862), .B2(n17928), .A(n17909), .ZN(n17925) );
  AOI211_X1 U20989 ( .C1(n17744), .C2(n18515), .A(n18529), .B(n17925), .ZN(
        n17781) );
  OAI22_X1 U20990 ( .A1(n18533), .A2(n17880), .B1(n17927), .B2(n17779), .ZN(
        n17780) );
  AOI211_X1 U20991 ( .C1(n17782), .C2(n18529), .A(n17781), .B(n17780), .ZN(
        n17783) );
  OAI211_X1 U20992 ( .C1(n19489), .C2(n17788), .A(n17784), .B(n17783), .ZN(
        P3_U2659) );
  INV_X1 U20993 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17795) );
  INV_X1 U20994 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19473) );
  NOR3_X1 U20995 ( .A1(n17917), .A2(n17885), .A3(n19473), .ZN(n17864) );
  NAND2_X1 U20996 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n17864), .ZN(n17860) );
  NOR2_X1 U20997 ( .A1(n17797), .A2(n17860), .ZN(n17821) );
  AOI21_X1 U20998 ( .B1(n17785), .B2(n17821), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n17789) );
  NAND2_X1 U20999 ( .A1(n10144), .A2(n17910), .ZN(n17851) );
  NOR2_X1 U21000 ( .A1(n18589), .A2(n17851), .ZN(n17810) );
  AOI21_X1 U21001 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17810), .A(
        n17862), .ZN(n17801) );
  AOI21_X1 U21002 ( .B1(n17744), .B2(n18558), .A(n17801), .ZN(n17786) );
  OAI21_X1 U21003 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17798), .A(
        n18515), .ZN(n18549) );
  XNOR2_X1 U21004 ( .A(n17786), .B(n18549), .ZN(n17787) );
  OAI22_X1 U21005 ( .A1(n17789), .A2(n17788), .B1(n19443), .B2(n17787), .ZN(
        n17790) );
  AOI211_X1 U21006 ( .C1(n17884), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18953), .B(
        n17790), .ZN(n17794) );
  OAI211_X1 U21007 ( .C1(n17802), .C2(n17792), .A(n17866), .B(n17791), .ZN(
        n17793) );
  OAI211_X1 U21008 ( .C1(n17880), .C2(n17795), .A(n17794), .B(n17793), .ZN(
        P3_U2660) );
  NAND2_X1 U21009 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .ZN(n17796) );
  AOI221_X1 U21010 ( .B1(n17885), .B2(n17902), .C1(n17796), .C2(n17902), .A(
        n17929), .ZN(n17859) );
  INV_X1 U21011 ( .A(n17859), .ZN(n17863) );
  AOI21_X1 U21012 ( .B1(n17933), .B2(n17797), .A(n17863), .ZN(n17834) );
  AOI21_X1 U21013 ( .B1(n18558), .B2(n17799), .A(n17798), .ZN(n18562) );
  INV_X1 U21014 ( .A(n18562), .ZN(n17800) );
  INV_X1 U21015 ( .A(n17801), .ZN(n17812) );
  AOI221_X1 U21016 ( .B1(n18562), .B2(n17801), .C1(n17800), .C2(n17812), .A(
        n19443), .ZN(n17806) );
  AOI211_X1 U21017 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17815), .A(n17802), .B(
        n17926), .ZN(n17805) );
  AOI22_X1 U21018 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17914), .B1(
        n17884), .B2(P3_EBX_REG_10__SCAN_IN), .ZN(n17803) );
  INV_X1 U21019 ( .A(n17803), .ZN(n17804) );
  NOR4_X1 U21020 ( .A1(n18953), .A2(n17806), .A3(n17805), .A4(n17804), .ZN(
        n17809) );
  OAI211_X1 U21021 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n17821), .B(n17807), .ZN(n17808) );
  OAI211_X1 U21022 ( .C1(n17834), .C2(n19486), .A(n17809), .B(n17808), .ZN(
        P3_U2661) );
  INV_X1 U21023 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17819) );
  NAND2_X1 U21024 ( .A1(n17862), .A2(n17829), .ZN(n17913) );
  OAI21_X1 U21025 ( .B1(n17810), .B2(n17813), .A(n17829), .ZN(n17811) );
  AOI22_X1 U21026 ( .A1(n17813), .A2(n17812), .B1(n17913), .B2(n17811), .ZN(
        n17814) );
  AOI211_X1 U21027 ( .C1(n17884), .C2(P3_EBX_REG_9__SCAN_IN), .A(n18953), .B(
        n17814), .ZN(n17818) );
  OAI211_X1 U21028 ( .C1(n17823), .C2(n17816), .A(n17866), .B(n17815), .ZN(
        n17817) );
  OAI211_X1 U21029 ( .C1(n17880), .C2(n17819), .A(n17818), .B(n17817), .ZN(
        n17820) );
  AOI21_X1 U21030 ( .B1(n17821), .B2(n19483), .A(n17820), .ZN(n17822) );
  OAI21_X1 U21031 ( .B1(n17834), .B2(n19483), .A(n17822), .ZN(P3_U2662) );
  INV_X1 U21032 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19482) );
  INV_X1 U21033 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19479) );
  INV_X1 U21034 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19477) );
  NOR4_X1 U21035 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n19479), .A3(n19477), .A4(
        n17860), .ZN(n17826) );
  AOI211_X1 U21036 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17845), .A(n17823), .B(
        n17926), .ZN(n17825) );
  INV_X1 U21037 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17828) );
  OAI22_X1 U21038 ( .A1(n17828), .A2(n17880), .B1(n17927), .B2(n18119), .ZN(
        n17824) );
  NOR4_X1 U21039 ( .A1(n18953), .A2(n17826), .A3(n17825), .A4(n17824), .ZN(
        n17833) );
  INV_X1 U21040 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18596) );
  NOR2_X1 U21041 ( .A1(n18594), .A2(n18596), .ZN(n18590) );
  NAND2_X1 U21042 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18590), .ZN(
        n17836) );
  AOI21_X1 U21043 ( .B1(n17828), .B2(n17836), .A(n17827), .ZN(n18580) );
  AOI21_X1 U21044 ( .B1(n18590), .B2(n17910), .A(n17862), .ZN(n17839) );
  INV_X1 U21045 ( .A(n18580), .ZN(n17831) );
  INV_X1 U21046 ( .A(n17839), .ZN(n17830) );
  OAI221_X1 U21047 ( .B1(n18580), .B2(n17839), .C1(n17831), .C2(n17830), .A(
        n17829), .ZN(n17832) );
  OAI211_X1 U21048 ( .C1(n17834), .C2(n19482), .A(n17833), .B(n17832), .ZN(
        P3_U2663) );
  NOR2_X1 U21049 ( .A1(n19477), .A2(n17860), .ZN(n17844) );
  OAI21_X1 U21050 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n17860), .A(n17859), .ZN(
        n17843) );
  INV_X1 U21051 ( .A(n17835), .ZN(n17849) );
  OAI21_X1 U21052 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17849), .A(
        n17836), .ZN(n18606) );
  INV_X1 U21053 ( .A(n18606), .ZN(n17840) );
  INV_X1 U21054 ( .A(n17913), .ZN(n17838) );
  AOI21_X1 U21055 ( .B1(n17840), .B2(n17851), .A(n19443), .ZN(n17837) );
  OAI22_X1 U21056 ( .A1(n17840), .A2(n17839), .B1(n17838), .B2(n17837), .ZN(
        n17841) );
  OAI211_X1 U21057 ( .C1(n18596), .C2(n17880), .A(n18840), .B(n17841), .ZN(
        n17842) );
  AOI221_X1 U21058 ( .B1(n17844), .B2(n19479), .C1(n17843), .C2(
        P3_REIP_REG_7__SCAN_IN), .A(n17842), .ZN(n17847) );
  OAI211_X1 U21059 ( .C1(n17852), .C2(n17848), .A(n17866), .B(n17845), .ZN(
        n17846) );
  OAI211_X1 U21060 ( .C1(n17848), .C2(n17927), .A(n17847), .B(n17846), .ZN(
        P3_U2664) );
  INV_X1 U21061 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n21483) );
  NAND2_X1 U21062 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18615), .ZN(
        n17861) );
  AOI21_X1 U21063 ( .B1(n21483), .B2(n17861), .A(n17849), .ZN(n17850) );
  INV_X1 U21064 ( .A(n17850), .ZN(n18622) );
  AOI211_X1 U21065 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n17744), .A(
        n18622), .B(n17925), .ZN(n17857) );
  NAND3_X1 U21066 ( .A1(n17851), .A2(n17915), .A3(n18622), .ZN(n17855) );
  AOI211_X1 U21067 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17865), .A(n17852), .B(
        n17926), .ZN(n17853) );
  AOI211_X1 U21068 ( .C1(n17884), .C2(P3_EBX_REG_6__SCAN_IN), .A(n13496), .B(
        n17853), .ZN(n17854) );
  NAND2_X1 U21069 ( .A1(n17855), .A2(n17854), .ZN(n17856) );
  AOI211_X1 U21070 ( .C1(n17914), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n17857), .B(n17856), .ZN(n17858) );
  OAI221_X1 U21071 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n17860), .C1(n19477), 
        .C2(n17859), .A(n17858), .ZN(P3_U2665) );
  NOR2_X1 U21072 ( .A1(n18684), .A2(n18630), .ZN(n17873) );
  OAI21_X1 U21073 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17873), .A(
        n17861), .ZN(n18635) );
  AOI21_X1 U21074 ( .B1(n17873), .B2(n17928), .A(n17862), .ZN(n17876) );
  XOR2_X1 U21075 ( .A(n18635), .B(n17876), .Z(n17872) );
  OAI21_X1 U21076 ( .B1(P3_REIP_REG_5__SCAN_IN), .B2(n17864), .A(n17863), .ZN(
        n17869) );
  OAI211_X1 U21077 ( .C1(n17878), .C2(n17867), .A(n17866), .B(n17865), .ZN(
        n17868) );
  OAI211_X1 U21078 ( .C1(n17880), .C2(n18629), .A(n17869), .B(n17868), .ZN(
        n17870) );
  AOI211_X1 U21079 ( .C1(n17884), .C2(P3_EBX_REG_5__SCAN_IN), .A(n13496), .B(
        n17870), .ZN(n17871) );
  OAI21_X1 U21080 ( .B1(n19443), .B2(n17872), .A(n17871), .ZN(P3_U2666) );
  INV_X1 U21081 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17881) );
  NAND2_X1 U21082 ( .A1(n18642), .A2(n17881), .ZN(n18639) );
  INV_X1 U21083 ( .A(n18639), .ZN(n17877) );
  AOI21_X1 U21084 ( .B1(n17881), .B2(n17874), .A(n17873), .ZN(n17875) );
  INV_X1 U21085 ( .A(n17875), .ZN(n18649) );
  AOI22_X1 U21086 ( .A1(n17910), .A2(n17877), .B1(n17876), .B2(n18649), .ZN(
        n17894) );
  AOI211_X1 U21087 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17879), .A(n17878), .B(
        n17926), .ZN(n17883) );
  OAI22_X1 U21088 ( .A1(n17881), .A2(n17880), .B1(n18649), .B2(n17913), .ZN(
        n17882) );
  AOI211_X1 U21089 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17884), .A(n17883), .B(
        n17882), .ZN(n17893) );
  NOR2_X1 U21090 ( .A1(n17917), .A2(n17885), .ZN(n17888) );
  AOI21_X1 U21091 ( .B1(n17886), .B2(n10445), .A(n19574), .ZN(n17887) );
  AOI211_X1 U21092 ( .C1(n17888), .C2(n19473), .A(n18953), .B(n17887), .ZN(
        n17889) );
  INV_X1 U21093 ( .A(n17889), .ZN(n17890) );
  AOI21_X1 U21094 ( .B1(n17891), .B2(P3_REIP_REG_4__SCAN_IN), .A(n17890), .ZN(
        n17892) );
  OAI211_X1 U21095 ( .C1(n17894), .C2(n19443), .A(n17893), .B(n17892), .ZN(
        P3_U2667) );
  OAI21_X1 U21096 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17895), .ZN(n18666) );
  INV_X1 U21097 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n18153) );
  NAND2_X1 U21098 ( .A1(n18153), .A2(n17916), .ZN(n17897) );
  AOI211_X1 U21099 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17897), .A(n17896), .B(
        n17926), .ZN(n17906) );
  OAI22_X1 U21100 ( .A1(n17899), .A2(n19469), .B1(n17898), .B2(n19574), .ZN(
        n17900) );
  INV_X1 U21101 ( .A(n17900), .ZN(n17904) );
  OAI211_X1 U21102 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17902), .B(n17901), .ZN(n17903) );
  OAI211_X1 U21103 ( .C1(n18143), .C2(n17927), .A(n17904), .B(n17903), .ZN(
        n17905) );
  AOI211_X1 U21104 ( .C1(n17914), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n17906), .B(n17905), .ZN(n17912) );
  INV_X1 U21105 ( .A(n17907), .ZN(n17908) );
  OAI211_X1 U21106 ( .C1(n17910), .C2(n18666), .A(n17909), .B(n17908), .ZN(
        n17911) );
  OAI211_X1 U21107 ( .C1(n17913), .C2(n18666), .A(n17912), .B(n17911), .ZN(
        P3_U2669) );
  AOI21_X1 U21108 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17915), .A(
        n17914), .ZN(n17924) );
  OAI22_X1 U21109 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17917), .B1(n17927), 
        .B2(n17916), .ZN(n17922) );
  INV_X1 U21110 ( .A(n17918), .ZN(n17919) );
  OAI22_X1 U21111 ( .A1(n17926), .A2(n17920), .B1(n19574), .B2(n17919), .ZN(
        n17921) );
  AOI211_X1 U21112 ( .C1(n17929), .C2(P3_REIP_REG_1__SCAN_IN), .A(n17922), .B(
        n17921), .ZN(n17923) );
  OAI221_X1 U21113 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17925), .C1(
        n18684), .C2(n17924), .A(n17923), .ZN(P3_U2670) );
  AOI21_X1 U21114 ( .B1(n17927), .B2(n17926), .A(n18153), .ZN(n17932) );
  NOR3_X1 U21115 ( .A1(n17930), .A2(n17929), .A3(n17928), .ZN(n17931) );
  AOI211_X1 U21116 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(n17933), .A(n17932), .B(
        n17931), .ZN(n17934) );
  OAI21_X1 U21117 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19574), .A(
        n17934), .ZN(P3_U2671) );
  INV_X1 U21118 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17935) );
  INV_X1 U21119 ( .A(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18005) );
  OAI22_X1 U21120 ( .A1(n18077), .A2(n17935), .B1(n9640), .B2(n18005), .ZN(
        n17940) );
  INV_X1 U21121 ( .A(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17938) );
  AOI22_X1 U21122 ( .A1(n18061), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17937) );
  AOI22_X1 U21123 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17936) );
  OAI211_X1 U21124 ( .C1(n18112), .C2(n17938), .A(n17937), .B(n17936), .ZN(
        n17939) );
  AOI211_X1 U21125 ( .C1(n17293), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n17940), .B(n17939), .ZN(n17948) );
  AOI22_X1 U21126 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17947) );
  AOI22_X1 U21127 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17946) );
  INV_X1 U21128 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17941) );
  NOR2_X1 U21129 ( .A1(n13229), .A2(n17941), .ZN(n17944) );
  INV_X1 U21130 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17942) );
  OAI22_X1 U21131 ( .A1(n10444), .A2(n18127), .B1(n18085), .B2(n17942), .ZN(
        n17943) );
  AOI211_X1 U21132 ( .C1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .C2(n18099), .A(
        n17944), .B(n17943), .ZN(n17945) );
  NAND4_X1 U21133 ( .A1(n17948), .A2(n17947), .A3(n17946), .A4(n17945), .ZN(
        n17967) );
  NAND2_X1 U21134 ( .A1(n17968), .A2(n17967), .ZN(n17966) );
  AOI22_X1 U21135 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17952) );
  AOI22_X1 U21136 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17951) );
  AOI22_X1 U21137 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17950) );
  AOI22_X1 U21138 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18101), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17949) );
  NAND4_X1 U21139 ( .A1(n17952), .A2(n17951), .A3(n17950), .A4(n17949), .ZN(
        n17961) );
  INV_X1 U21140 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17956) );
  AOI22_X1 U21141 ( .A1(n18061), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17955) );
  AOI22_X1 U21142 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18108), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17954) );
  OAI211_X1 U21143 ( .C1(n17956), .C2(n18112), .A(n17955), .B(n17954), .ZN(
        n17960) );
  INV_X1 U21144 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17958) );
  AOI22_X1 U21145 ( .A1(n18008), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17957) );
  OAI21_X1 U21146 ( .B1(n17239), .B2(n17958), .A(n17957), .ZN(n17959) );
  OR3_X1 U21147 ( .A1(n17961), .A2(n17960), .A3(n17959), .ZN(n17962) );
  XOR2_X1 U21148 ( .A(n17966), .B(n17962), .Z(n18161) );
  NOR2_X1 U21149 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17963), .ZN(n17965) );
  OAI22_X1 U21150 ( .A1(n18161), .A2(n18148), .B1(n17965), .B2(n17964), .ZN(
        P3_U2673) );
  OAI21_X1 U21151 ( .B1(n17968), .B2(n17967), .A(n17966), .ZN(n18169) );
  OAI222_X1 U21152 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17972), .B1(
        P3_EBX_REG_29__SCAN_IN), .B2(n17971), .C1(n17970), .C2(n17969), .ZN(
        n17973) );
  OAI21_X1 U21153 ( .B1(n18169), .B2(n18148), .A(n17973), .ZN(P3_U2674) );
  OAI21_X1 U21154 ( .B1(n17978), .B2(n17975), .A(n17974), .ZN(n18179) );
  NAND3_X1 U21155 ( .A1(n17977), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n18148), 
        .ZN(n17976) );
  OAI221_X1 U21156 ( .B1(n17977), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n18148), 
        .C2(n18179), .A(n17976), .ZN(P3_U2676) );
  INV_X1 U21157 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n21530) );
  AOI21_X1 U21158 ( .B1(n17979), .B2(n17983), .A(n17978), .ZN(n18180) );
  NAND2_X1 U21159 ( .A1(n18180), .A2(n18151), .ZN(n17980) );
  OAI221_X1 U21160 ( .B1(n17982), .B2(n21530), .C1(n17982), .C2(n17981), .A(
        n17980), .ZN(P3_U2677) );
  AOI21_X1 U21161 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18148), .A(n17993), .ZN(
        n17985) );
  OAI21_X1 U21162 ( .B1(n17990), .B2(n17984), .A(n17983), .ZN(n18187) );
  OAI22_X1 U21163 ( .A1(n17986), .A2(n17985), .B1(n18148), .B2(n18187), .ZN(
        P3_U2678) );
  NOR2_X1 U21164 ( .A1(n17987), .A2(n17994), .ZN(n18000) );
  AOI21_X1 U21165 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18148), .A(n18000), .ZN(
        n17992) );
  NOR2_X1 U21166 ( .A1(n17995), .A2(n17988), .ZN(n17989) );
  NOR2_X1 U21167 ( .A1(n17990), .A2(n17989), .ZN(n18188) );
  INV_X1 U21168 ( .A(n18188), .ZN(n17991) );
  OAI22_X1 U21169 ( .A1(n17993), .A2(n17992), .B1(n18148), .B2(n17991), .ZN(
        P3_U2679) );
  INV_X1 U21170 ( .A(n17994), .ZN(n18020) );
  AOI21_X1 U21171 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18148), .A(n18020), .ZN(
        n17999) );
  INV_X1 U21172 ( .A(n17995), .ZN(n17996) );
  OAI21_X1 U21173 ( .B1(n17998), .B2(n17997), .A(n17996), .ZN(n18196) );
  OAI22_X1 U21174 ( .A1(n18000), .A2(n17999), .B1(n18148), .B2(n18196), .ZN(
        P3_U2680) );
  AOI21_X1 U21175 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18148), .A(n18001), .ZN(
        n18019) );
  NAND2_X1 U21176 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n18004) );
  NAND2_X1 U21177 ( .A1(n18002), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n18003) );
  OAI211_X1 U21178 ( .C1(n18006), .C2(n18005), .A(n18004), .B(n18003), .ZN(
        n18007) );
  INV_X1 U21179 ( .A(n18007), .ZN(n18012) );
  AOI22_X1 U21180 ( .A1(n18008), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18011) );
  AOI22_X1 U21181 ( .A1(n18061), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18010) );
  NAND2_X1 U21182 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n18009) );
  NAND4_X1 U21183 ( .A1(n18012), .A2(n18011), .A3(n18010), .A4(n18009), .ZN(
        n18018) );
  AOI22_X1 U21184 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18016) );
  AOI22_X1 U21185 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18015) );
  AOI22_X1 U21186 ( .A1(n13053), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18014) );
  AOI22_X1 U21187 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18013) );
  NAND4_X1 U21188 ( .A1(n18016), .A2(n18015), .A3(n18014), .A4(n18013), .ZN(
        n18017) );
  NOR2_X1 U21189 ( .A1(n18018), .A2(n18017), .ZN(n18201) );
  OAI22_X1 U21190 ( .A1(n18020), .A2(n18019), .B1(n18201), .B2(n18148), .ZN(
        P3_U2681) );
  NOR2_X1 U21191 ( .A1(n18021), .A2(n19010), .ZN(n18054) );
  NAND2_X1 U21192 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18054), .ZN(n18037) );
  AOI22_X1 U21193 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18107), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18023) );
  NAND2_X1 U21194 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n18022) );
  AND2_X1 U21195 ( .A1(n18023), .A2(n18022), .ZN(n18027) );
  AOI22_X1 U21196 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18026) );
  AOI22_X1 U21197 ( .A1(n18061), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18025) );
  NAND2_X1 U21198 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n18024) );
  NAND4_X1 U21199 ( .A1(n18027), .A2(n18026), .A3(n18025), .A4(n18024), .ZN(
        n18034) );
  AOI22_X1 U21200 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18032) );
  AOI22_X1 U21201 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18031) );
  AOI22_X1 U21202 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18030) );
  AOI22_X1 U21203 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18029) );
  NAND4_X1 U21204 ( .A1(n18032), .A2(n18031), .A3(n18030), .A4(n18029), .ZN(
        n18033) );
  OR2_X1 U21205 ( .A1(n18034), .A2(n18033), .ZN(n18208) );
  OAI21_X1 U21206 ( .B1(n18052), .B2(n17667), .A(n18148), .ZN(n18035) );
  OAI21_X1 U21207 ( .B1(n18148), .B2(n18208), .A(n18035), .ZN(n18036) );
  OAI21_X1 U21208 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n18037), .A(n18036), .ZN(
        P3_U2682) );
  NAND2_X1 U21209 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n18039) );
  NAND2_X1 U21210 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n18038) );
  OAI211_X1 U21211 ( .C1(n17276), .C2(n18040), .A(n18039), .B(n18038), .ZN(
        n18041) );
  INV_X1 U21212 ( .A(n18041), .ZN(n18045) );
  AOI22_X1 U21213 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18044) );
  AOI22_X1 U21214 ( .A1(n18061), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18043) );
  NAND2_X1 U21215 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n18042) );
  NAND4_X1 U21216 ( .A1(n18045), .A2(n18044), .A3(n18043), .A4(n18042), .ZN(
        n18051) );
  AOI22_X1 U21217 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18049) );
  AOI22_X1 U21218 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18048) );
  AOI22_X1 U21219 ( .A1(n18101), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18047) );
  AOI22_X1 U21220 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18046) );
  NAND4_X1 U21221 ( .A1(n18049), .A2(n18048), .A3(n18047), .A4(n18046), .ZN(
        n18050) );
  NOR2_X1 U21222 ( .A1(n18051), .A2(n18050), .ZN(n18212) );
  NOR2_X1 U21223 ( .A1(n18052), .A2(n18151), .ZN(n18053) );
  OAI21_X1 U21224 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18054), .A(n18053), .ZN(
        n18055) );
  OAI21_X1 U21225 ( .B1(n18212), .B2(n18148), .A(n18055), .ZN(P3_U2683) );
  NAND3_X1 U21226 ( .A1(n18148), .A2(P3_EBX_REG_18__SCAN_IN), .A3(n18056), 
        .ZN(n18074) );
  NAND2_X1 U21227 ( .A1(n18057), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n18059) );
  NAND2_X1 U21228 ( .A1(n13507), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n18058) );
  OAI211_X1 U21229 ( .C1(n17276), .C2(n18076), .A(n18059), .B(n18058), .ZN(
        n18060) );
  INV_X1 U21230 ( .A(n18060), .ZN(n18065) );
  AOI22_X1 U21231 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18064) );
  AOI22_X1 U21232 ( .A1(n18061), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18063) );
  NAND2_X1 U21233 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n18062) );
  NAND4_X1 U21234 ( .A1(n18065), .A2(n18064), .A3(n18063), .A4(n18062), .ZN(
        n18071) );
  AOI22_X1 U21235 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18069) );
  AOI22_X1 U21236 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18068) );
  AOI22_X1 U21237 ( .A1(n13053), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18067) );
  AOI22_X1 U21238 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18066) );
  NAND4_X1 U21239 ( .A1(n18069), .A2(n18068), .A3(n18067), .A4(n18066), .ZN(
        n18070) );
  OR2_X1 U21240 ( .A1(n18071), .A2(n18070), .ZN(n18222) );
  AOI22_X1 U21241 ( .A1(n18072), .A2(n21491), .B1(n18151), .B2(n18222), .ZN(
        n18073) );
  NAND2_X1 U21242 ( .A1(n18074), .A2(n18073), .ZN(P3_U2685) );
  NAND2_X1 U21243 ( .A1(n18094), .A2(n18157), .ZN(n18097) );
  OAI22_X1 U21244 ( .A1(n18077), .A2(n18076), .B1(n9640), .B2(n18075), .ZN(
        n18082) );
  AOI22_X1 U21245 ( .A1(n18061), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18079) );
  AOI22_X1 U21246 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18107), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18078) );
  OAI211_X1 U21247 ( .C1(n18112), .C2(n18080), .A(n18079), .B(n18078), .ZN(
        n18081) );
  AOI211_X1 U21248 ( .C1(n17293), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n18082), .B(n18081), .ZN(n18092) );
  AOI22_X1 U21249 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13361), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18091) );
  AOI22_X1 U21250 ( .A1(n13053), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18090) );
  INV_X1 U21251 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18083) );
  NOR2_X1 U21252 ( .A1(n13229), .A2(n18083), .ZN(n18088) );
  INV_X1 U21253 ( .A(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18084) );
  OAI22_X1 U21254 ( .A1(n10444), .A2(n18086), .B1(n18085), .B2(n18084), .ZN(
        n18087) );
  AOI211_X1 U21255 ( .C1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .C2(n18099), .A(
        n18088), .B(n18087), .ZN(n18089) );
  NAND4_X1 U21256 ( .A1(n18092), .A2(n18091), .A3(n18090), .A4(n18089), .ZN(
        n18244) );
  INV_X1 U21257 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n18093) );
  OAI21_X1 U21258 ( .B1(n18094), .B2(n18093), .A(n18148), .ZN(n18095) );
  OAI21_X1 U21259 ( .B1(n18244), .B2(n18148), .A(n18095), .ZN(n18096) );
  OAI21_X1 U21260 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n18097), .A(n18096), .ZN(
        P3_U2693) );
  AOI22_X1 U21261 ( .A1(n18098), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9568), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18105) );
  AOI22_X1 U21262 ( .A1(n18099), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18104) );
  AOI22_X1 U21263 ( .A1(n18100), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18103) );
  AOI22_X1 U21264 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18101), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18102) );
  NAND4_X1 U21265 ( .A1(n18105), .A2(n18104), .A3(n18103), .A4(n18102), .ZN(
        n18117) );
  INV_X1 U21266 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18111) );
  AOI22_X1 U21267 ( .A1(n18061), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18110) );
  AOI22_X1 U21268 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18107), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18109) );
  OAI211_X1 U21269 ( .C1(n18112), .C2(n18111), .A(n18110), .B(n18109), .ZN(
        n18116) );
  INV_X1 U21270 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18114) );
  AOI22_X1 U21271 ( .A1(n17278), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14312), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18113) );
  OAI21_X1 U21272 ( .B1(n17239), .B2(n18114), .A(n18113), .ZN(n18115) );
  OR3_X1 U21273 ( .A1(n18117), .A2(n18116), .A3(n18115), .ZN(n18248) );
  INV_X1 U21274 ( .A(n18118), .ZN(n18125) );
  OAI21_X1 U21275 ( .B1(n18119), .B2(n18125), .A(n18148), .ZN(n18120) );
  OAI21_X1 U21276 ( .B1(n18148), .B2(n18248), .A(n18120), .ZN(n18121) );
  OAI21_X1 U21277 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n18122), .A(n18121), .ZN(
        P3_U2695) );
  NAND2_X1 U21278 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n18137), .ZN(n18130) );
  INV_X1 U21279 ( .A(n18130), .ZN(n18126) );
  AND2_X1 U21280 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18126), .ZN(n18129) );
  AOI21_X1 U21281 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n18148), .A(n18129), .ZN(
        n18124) );
  INV_X1 U21282 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18123) );
  OAI22_X1 U21283 ( .A1(n18125), .A2(n18124), .B1(n18123), .B2(n18148), .ZN(
        P3_U2696) );
  AOI21_X1 U21284 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n18148), .A(n18126), .ZN(
        n18128) );
  OAI22_X1 U21285 ( .A1(n18129), .A2(n18128), .B1(n18127), .B2(n18148), .ZN(
        P3_U2697) );
  OAI21_X1 U21286 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n18131), .A(n18130), .ZN(
        n18132) );
  AOI22_X1 U21287 ( .A1(n18151), .A2(n18133), .B1(n18132), .B2(n18148), .ZN(
        P3_U2698) );
  NAND2_X1 U21288 ( .A1(n18134), .A2(n18150), .ZN(n18146) );
  NOR2_X1 U21289 ( .A1(n18138), .A2(n18146), .ZN(n18142) );
  AOI21_X1 U21290 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18148), .A(n18142), .ZN(
        n18136) );
  OAI22_X1 U21291 ( .A1(n18137), .A2(n18136), .B1(n18135), .B2(n18148), .ZN(
        P3_U2699) );
  OAI21_X1 U21292 ( .B1(n18138), .B2(n18151), .A(n18146), .ZN(n18139) );
  INV_X1 U21293 ( .A(n18139), .ZN(n18141) );
  INV_X1 U21294 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18140) );
  OAI22_X1 U21295 ( .A1(n18142), .A2(n18141), .B1(n18140), .B2(n18148), .ZN(
        P3_U2700) );
  OAI211_X1 U21296 ( .C1(n18145), .C2(n18144), .A(n18143), .B(n18148), .ZN(
        n18147) );
  OAI211_X1 U21297 ( .C1(n18148), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n18147), .B(n18146), .ZN(n18149) );
  INV_X1 U21298 ( .A(n18149), .ZN(P3_U2701) );
  AOI22_X1 U21299 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18151), .B1(
        n18150), .B2(n18153), .ZN(n18152) );
  OAI21_X1 U21300 ( .B1(n18154), .B2(n18153), .A(n18152), .ZN(P3_U2703) );
  INV_X1 U21301 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18318) );
  INV_X1 U21302 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n18315) );
  INV_X1 U21303 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n21429) );
  INV_X1 U21304 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18312) );
  INV_X1 U21305 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n21415) );
  INV_X1 U21306 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18310) );
  INV_X1 U21307 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18308) );
  NOR4_X1 U21308 ( .A1(n21415), .A2(n18310), .A3(n18308), .A4(n18303), .ZN(
        n18155) );
  NAND4_X1 U21309 ( .A1(n18156), .A2(P3_EAX_REG_20__SCAN_IN), .A3(
        P3_EAX_REG_19__SCAN_IN), .A4(n18155), .ZN(n18195) );
  NOR2_X2 U21310 ( .A1(n18312), .A2(n18195), .ZN(n18194) );
  NAND2_X1 U21311 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18175), .ZN(n18171) );
  NAND2_X1 U21312 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18166), .ZN(n18165) );
  NOR2_X1 U21313 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n18165), .ZN(n18159) );
  NAND2_X1 U21314 ( .A1(n18251), .A2(n18165), .ZN(n18164) );
  OAI21_X1 U21315 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n18203), .A(n18164), .ZN(
        n18158) );
  AOI22_X1 U21316 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n18159), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n18158), .ZN(n18160) );
  OAI21_X1 U21317 ( .B1(n19014), .B2(n18221), .A(n18160), .ZN(P3_U2704) );
  INV_X1 U21318 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18324) );
  OAI22_X1 U21319 ( .A1(n18161), .A2(n18197), .B1(n19006), .B2(n18221), .ZN(
        n18162) );
  AOI21_X1 U21320 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n18214), .A(n18162), .ZN(
        n18163) );
  OAI221_X1 U21321 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n18165), .C1(n18324), 
        .C2(n18164), .A(n18163), .ZN(P3_U2705) );
  AOI22_X1 U21322 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18214), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18223), .ZN(n18168) );
  OAI211_X1 U21323 ( .C1(n18166), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18251), .B(
        n18165), .ZN(n18167) );
  OAI211_X1 U21324 ( .C1(n18169), .C2(n18197), .A(n18168), .B(n18167), .ZN(
        P3_U2706) );
  AOI22_X1 U21325 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18223), .B1(n18249), .B2(
        n18170), .ZN(n18173) );
  OAI211_X1 U21326 ( .C1(n18175), .C2(P3_EAX_REG_28__SCAN_IN), .A(n18251), .B(
        n18171), .ZN(n18172) );
  OAI211_X1 U21327 ( .C1(n18229), .C2(n18174), .A(n18173), .B(n18172), .ZN(
        P3_U2707) );
  AOI22_X1 U21328 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18214), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18223), .ZN(n18178) );
  AOI211_X1 U21329 ( .C1(n18318), .C2(n18181), .A(n18175), .B(n18241), .ZN(
        n18176) );
  INV_X1 U21330 ( .A(n18176), .ZN(n18177) );
  OAI211_X1 U21331 ( .C1(n18179), .C2(n18197), .A(n18178), .B(n18177), .ZN(
        P3_U2708) );
  INV_X1 U21332 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18246) );
  AOI22_X1 U21333 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18223), .B1(n18249), .B2(
        n18180), .ZN(n18183) );
  OAI211_X1 U21334 ( .C1(n9644), .C2(P3_EAX_REG_26__SCAN_IN), .A(n18251), .B(
        n18181), .ZN(n18182) );
  OAI211_X1 U21335 ( .C1(n18229), .C2(n18246), .A(n18183), .B(n18182), .ZN(
        P3_U2709) );
  AOI22_X1 U21336 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18214), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18223), .ZN(n18186) );
  AOI211_X1 U21337 ( .C1(n18315), .C2(n18190), .A(n9644), .B(n18241), .ZN(
        n18184) );
  INV_X1 U21338 ( .A(n18184), .ZN(n18185) );
  OAI211_X1 U21339 ( .C1(n18187), .C2(n18197), .A(n18186), .B(n18185), .ZN(
        P3_U2710) );
  AOI22_X1 U21340 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18223), .B1(n18249), .B2(
        n18188), .ZN(n18193) );
  OAI21_X1 U21341 ( .B1(n21429), .B2(n18241), .A(n18189), .ZN(n18191) );
  NAND2_X1 U21342 ( .A1(n18191), .A2(n18190), .ZN(n18192) );
  OAI211_X1 U21343 ( .C1(n18229), .C2(n18254), .A(n18193), .B(n18192), .ZN(
        P3_U2711) );
  AOI211_X1 U21344 ( .C1(n18312), .C2(n18195), .A(n18241), .B(n18194), .ZN(
        n18199) );
  OAI22_X1 U21345 ( .A1(n19012), .A2(n18229), .B1(n18197), .B2(n18196), .ZN(
        n18198) );
  AOI211_X1 U21346 ( .C1(n18223), .C2(BUF2_REG_23__SCAN_IN), .A(n18199), .B(
        n18198), .ZN(n18200) );
  INV_X1 U21347 ( .A(n18200), .ZN(P3_U2712) );
  INV_X1 U21348 ( .A(n18201), .ZN(n18202) );
  AOI22_X1 U21349 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18223), .B1(n18249), .B2(
        n18202), .ZN(n18207) );
  NAND3_X1 U21350 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(n18224), .ZN(n18216) );
  NAND2_X1 U21351 ( .A1(n18251), .A2(n18216), .ZN(n18209) );
  OAI21_X1 U21352 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18203), .A(n18209), .ZN(
        n18205) );
  NOR2_X1 U21353 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18216), .ZN(n18204) );
  AOI22_X1 U21354 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18205), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n18204), .ZN(n18206) );
  OAI211_X1 U21355 ( .C1(n21479), .C2(n18229), .A(n18207), .B(n18206), .ZN(
        P3_U2713) );
  AOI22_X1 U21356 ( .A1(n18223), .A2(BUF2_REG_21__SCAN_IN), .B1(n18249), .B2(
        n18208), .ZN(n18211) );
  INV_X1 U21357 ( .A(n18209), .ZN(n18218) );
  AOI22_X1 U21358 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18214), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n18218), .ZN(n18210) );
  OAI211_X1 U21359 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n18216), .A(n18211), .B(
        n18210), .ZN(P3_U2714) );
  INV_X1 U21360 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18998) );
  INV_X1 U21361 ( .A(n18212), .ZN(n18213) );
  AOI22_X1 U21362 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18214), .B1(n18249), .B2(
        n18213), .ZN(n18220) );
  INV_X1 U21363 ( .A(n18215), .ZN(n18217) );
  AOI22_X1 U21364 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18218), .B1(n18217), 
        .B2(n18216), .ZN(n18219) );
  OAI211_X1 U21365 ( .C1(n18998), .C2(n18221), .A(n18220), .B(n18219), .ZN(
        P3_U2715) );
  AOI22_X1 U21366 ( .A1(n18223), .A2(BUF2_REG_18__SCAN_IN), .B1(n18249), .B2(
        n18222), .ZN(n18228) );
  AOI211_X1 U21367 ( .C1(n18303), .C2(n18225), .A(n18224), .B(n18241), .ZN(
        n18226) );
  INV_X1 U21368 ( .A(n18226), .ZN(n18227) );
  OAI211_X1 U21369 ( .C1(n18229), .C2(n21444), .A(n18228), .B(n18227), .ZN(
        P3_U2717) );
  AOI22_X1 U21370 ( .A1(n18249), .A2(n18230), .B1(BUF2_REG_15__SCAN_IN), .B2(
        n18236), .ZN(n18233) );
  OAI211_X1 U21371 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n9650), .A(n18251), .B(
        n18231), .ZN(n18232) );
  NAND2_X1 U21372 ( .A1(n18233), .A2(n18232), .ZN(P3_U2720) );
  INV_X1 U21373 ( .A(n18234), .ZN(n18235) );
  AOI22_X1 U21374 ( .A1(n18236), .A2(BUF2_REG_14__SCAN_IN), .B1(n18249), .B2(
        n18235), .ZN(n18238) );
  INV_X1 U21375 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n18352) );
  OR3_X1 U21376 ( .A1(n18352), .A2(n18241), .A3(n9650), .ZN(n18237) );
  OAI211_X1 U21377 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n18239), .A(n18238), .B(
        n18237), .ZN(P3_U2721) );
  AOI211_X1 U21378 ( .C1(n18242), .C2(n18344), .A(n18241), .B(n18240), .ZN(
        n18243) );
  AOI21_X1 U21379 ( .B1(n18249), .B2(n18244), .A(n18243), .ZN(n18245) );
  OAI21_X1 U21380 ( .B1(n18246), .B2(n18255), .A(n18245), .ZN(P3_U2725) );
  INV_X1 U21381 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18340) );
  AOI22_X1 U21382 ( .A1(n18249), .A2(n18248), .B1(n18247), .B2(n18340), .ZN(
        n18253) );
  NAND3_X1 U21383 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18251), .A3(n18250), .ZN(
        n18252) );
  OAI211_X1 U21384 ( .C1(n18255), .C2(n18254), .A(n18253), .B(n18252), .ZN(
        P3_U2727) );
  OR2_X1 U21385 ( .A1(n19444), .A2(n18439), .ZN(n19562) );
  NOR2_X4 U21386 ( .A1(n18290), .A2(n18273), .ZN(n18283) );
  AND2_X1 U21387 ( .A1(n18283), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U21388 ( .A1(n18273), .A2(n18978), .ZN(n18272) );
  AOI22_X1 U21389 ( .A1(n18290), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18257) );
  OAI21_X1 U21390 ( .B1(n18324), .B2(n18272), .A(n18257), .ZN(P3_U2737) );
  INV_X1 U21391 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18322) );
  AOI22_X1 U21392 ( .A1(n18290), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18258) );
  OAI21_X1 U21393 ( .B1(n18322), .B2(n18272), .A(n18258), .ZN(P3_U2738) );
  INV_X1 U21394 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18320) );
  AOI22_X1 U21395 ( .A1(n18290), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18259) );
  OAI21_X1 U21396 ( .B1(n18320), .B2(n18272), .A(n18259), .ZN(P3_U2739) );
  AOI22_X1 U21397 ( .A1(n18290), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18260) );
  OAI21_X1 U21398 ( .B1(n18318), .B2(n18272), .A(n18260), .ZN(P3_U2740) );
  AOI22_X1 U21399 ( .A1(n18290), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18261) );
  OAI21_X1 U21400 ( .B1(n10174), .B2(n18272), .A(n18261), .ZN(P3_U2741) );
  AOI22_X1 U21401 ( .A1(n18290), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18262) );
  OAI21_X1 U21402 ( .B1(n18315), .B2(n18272), .A(n18262), .ZN(P3_U2742) );
  AOI22_X1 U21403 ( .A1(n18290), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18263) );
  OAI21_X1 U21404 ( .B1(n21429), .B2(n18272), .A(n18263), .ZN(P3_U2743) );
  INV_X2 U21405 ( .A(n19562), .ZN(n18290) );
  AOI22_X1 U21406 ( .A1(n18290), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18264) );
  OAI21_X1 U21407 ( .B1(n18312), .B2(n18272), .A(n18264), .ZN(P3_U2744) );
  AOI22_X1 U21408 ( .A1(n18290), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18265) );
  OAI21_X1 U21409 ( .B1(n18310), .B2(n18272), .A(n18265), .ZN(P3_U2745) );
  AOI22_X1 U21410 ( .A1(n18290), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18266) );
  OAI21_X1 U21411 ( .B1(n18308), .B2(n18272), .A(n18266), .ZN(P3_U2746) );
  INV_X1 U21412 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18306) );
  AOI22_X1 U21413 ( .A1(n18290), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18267) );
  OAI21_X1 U21414 ( .B1(n18306), .B2(n18272), .A(n18267), .ZN(P3_U2747) );
  AOI22_X1 U21415 ( .A1(n18290), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18268) );
  OAI21_X1 U21416 ( .B1(n16836), .B2(n18272), .A(n18268), .ZN(P3_U2748) );
  AOI22_X1 U21417 ( .A1(n18290), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18269) );
  OAI21_X1 U21418 ( .B1(n18303), .B2(n18272), .A(n18269), .ZN(P3_U2749) );
  AOI22_X1 U21419 ( .A1(n18290), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18270) );
  OAI21_X1 U21420 ( .B1(n21415), .B2(n18272), .A(n18270), .ZN(P3_U2750) );
  AOI22_X1 U21421 ( .A1(n18290), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18271) );
  OAI21_X1 U21422 ( .B1(n18300), .B2(n18272), .A(n18271), .ZN(P3_U2751) );
  INV_X1 U21423 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18356) );
  AOI22_X1 U21424 ( .A1(n18290), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18274) );
  OAI21_X1 U21425 ( .B1(n18356), .B2(n18292), .A(n18274), .ZN(P3_U2752) );
  AOI22_X1 U21426 ( .A1(n18290), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18275) );
  OAI21_X1 U21427 ( .B1(n18352), .B2(n18292), .A(n18275), .ZN(P3_U2753) );
  INV_X1 U21428 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18350) );
  AOI22_X1 U21429 ( .A1(n18290), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18276) );
  OAI21_X1 U21430 ( .B1(n18350), .B2(n18292), .A(n18276), .ZN(P3_U2754) );
  AOI22_X1 U21431 ( .A1(n18290), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18277) );
  OAI21_X1 U21432 ( .B1(n18348), .B2(n18292), .A(n18277), .ZN(P3_U2755) );
  INV_X1 U21433 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18346) );
  AOI22_X1 U21434 ( .A1(n18290), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18278) );
  OAI21_X1 U21435 ( .B1(n18346), .B2(n18292), .A(n18278), .ZN(P3_U2756) );
  AOI22_X1 U21436 ( .A1(n18290), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18279) );
  OAI21_X1 U21437 ( .B1(n18344), .B2(n18292), .A(n18279), .ZN(P3_U2757) );
  INV_X1 U21438 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18342) );
  AOI22_X1 U21439 ( .A1(n18290), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18280) );
  OAI21_X1 U21440 ( .B1(n18342), .B2(n18292), .A(n18280), .ZN(P3_U2758) );
  AOI22_X1 U21441 ( .A1(n18290), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18281) );
  OAI21_X1 U21442 ( .B1(n18340), .B2(n18292), .A(n18281), .ZN(P3_U2759) );
  INV_X1 U21443 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18338) );
  AOI22_X1 U21444 ( .A1(n18290), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18282) );
  OAI21_X1 U21445 ( .B1(n18338), .B2(n18292), .A(n18282), .ZN(P3_U2760) );
  AOI22_X1 U21446 ( .A1(n18290), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18284) );
  OAI21_X1 U21447 ( .B1(n18336), .B2(n18292), .A(n18284), .ZN(P3_U2761) );
  INV_X1 U21448 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18334) );
  AOI22_X1 U21449 ( .A1(n18290), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18285) );
  OAI21_X1 U21450 ( .B1(n18334), .B2(n18292), .A(n18285), .ZN(P3_U2762) );
  AOI22_X1 U21451 ( .A1(n18290), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18286) );
  OAI21_X1 U21452 ( .B1(n18332), .B2(n18292), .A(n18286), .ZN(P3_U2763) );
  INV_X1 U21453 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18330) );
  AOI22_X1 U21454 ( .A1(n18290), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18287) );
  OAI21_X1 U21455 ( .B1(n18330), .B2(n18292), .A(n18287), .ZN(P3_U2764) );
  INV_X1 U21456 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18328) );
  AOI22_X1 U21457 ( .A1(n18290), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18288) );
  OAI21_X1 U21458 ( .B1(n18328), .B2(n18292), .A(n18288), .ZN(P3_U2765) );
  INV_X1 U21459 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n21435) );
  AOI22_X1 U21460 ( .A1(n18290), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18289) );
  OAI21_X1 U21461 ( .B1(n21435), .B2(n18292), .A(n18289), .ZN(P3_U2766) );
  AOI22_X1 U21462 ( .A1(n18290), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18283), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18291) );
  OAI21_X1 U21463 ( .B1(n21512), .B2(n18292), .A(n18291), .ZN(P3_U2767) );
  INV_X1 U21464 ( .A(n18293), .ZN(n18297) );
  INV_X1 U21465 ( .A(n19386), .ZN(n19563) );
  NAND2_X1 U21466 ( .A1(n18985), .A2(n19563), .ZN(n18294) );
  AOI22_X1 U21467 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n10447), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18353), .ZN(n18299) );
  OAI21_X1 U21468 ( .B1(n18300), .B2(n18355), .A(n18299), .ZN(P3_U2768) );
  AOI22_X1 U21469 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n10447), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18353), .ZN(n18301) );
  OAI21_X1 U21470 ( .B1(n21415), .B2(n18355), .A(n18301), .ZN(P3_U2769) );
  AOI22_X1 U21471 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n10447), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18353), .ZN(n18302) );
  OAI21_X1 U21472 ( .B1(n18303), .B2(n18355), .A(n18302), .ZN(P3_U2770) );
  AOI22_X1 U21473 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n10447), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18353), .ZN(n18304) );
  OAI21_X1 U21474 ( .B1(n16836), .B2(n18355), .A(n18304), .ZN(P3_U2771) );
  AOI22_X1 U21475 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n10447), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18353), .ZN(n18305) );
  OAI21_X1 U21476 ( .B1(n18306), .B2(n18355), .A(n18305), .ZN(P3_U2772) );
  AOI22_X1 U21477 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n10447), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18353), .ZN(n18307) );
  OAI21_X1 U21478 ( .B1(n18308), .B2(n18355), .A(n18307), .ZN(P3_U2773) );
  AOI22_X1 U21479 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n10447), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18353), .ZN(n18309) );
  OAI21_X1 U21480 ( .B1(n18310), .B2(n18355), .A(n18309), .ZN(P3_U2774) );
  AOI22_X1 U21481 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n10447), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18353), .ZN(n18311) );
  OAI21_X1 U21482 ( .B1(n18312), .B2(n18355), .A(n18311), .ZN(P3_U2775) );
  AOI22_X1 U21483 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n10447), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18353), .ZN(n18313) );
  OAI21_X1 U21484 ( .B1(n21429), .B2(n18355), .A(n18313), .ZN(P3_U2776) );
  AOI22_X1 U21485 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n10447), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18353), .ZN(n18314) );
  OAI21_X1 U21486 ( .B1(n18315), .B2(n18355), .A(n18314), .ZN(P3_U2777) );
  AOI22_X1 U21487 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n10447), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18353), .ZN(n18316) );
  OAI21_X1 U21488 ( .B1(n10174), .B2(n18355), .A(n18316), .ZN(P3_U2778) );
  AOI22_X1 U21489 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n10447), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18353), .ZN(n18317) );
  OAI21_X1 U21490 ( .B1(n18318), .B2(n18355), .A(n18317), .ZN(P3_U2779) );
  AOI22_X1 U21491 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n10447), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18353), .ZN(n18319) );
  OAI21_X1 U21492 ( .B1(n18320), .B2(n18355), .A(n18319), .ZN(P3_U2780) );
  AOI22_X1 U21493 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n10447), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18353), .ZN(n18321) );
  OAI21_X1 U21494 ( .B1(n18322), .B2(n18355), .A(n18321), .ZN(P3_U2781) );
  AOI22_X1 U21495 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n10447), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18353), .ZN(n18323) );
  OAI21_X1 U21496 ( .B1(n18324), .B2(n18355), .A(n18323), .ZN(P3_U2782) );
  AOI22_X1 U21497 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n10447), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18353), .ZN(n18325) );
  OAI21_X1 U21498 ( .B1(n21512), .B2(n18355), .A(n18325), .ZN(P3_U2783) );
  AOI22_X1 U21499 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n10447), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18353), .ZN(n18326) );
  OAI21_X1 U21500 ( .B1(n21435), .B2(n18355), .A(n18326), .ZN(P3_U2784) );
  AOI22_X1 U21501 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n10447), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18353), .ZN(n18327) );
  OAI21_X1 U21502 ( .B1(n18328), .B2(n18355), .A(n18327), .ZN(P3_U2785) );
  AOI22_X1 U21503 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n10447), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18353), .ZN(n18329) );
  OAI21_X1 U21504 ( .B1(n18330), .B2(n18355), .A(n18329), .ZN(P3_U2786) );
  AOI22_X1 U21505 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n10447), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18353), .ZN(n18331) );
  OAI21_X1 U21506 ( .B1(n18332), .B2(n18355), .A(n18331), .ZN(P3_U2787) );
  AOI22_X1 U21507 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n10447), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18353), .ZN(n18333) );
  OAI21_X1 U21508 ( .B1(n18334), .B2(n18355), .A(n18333), .ZN(P3_U2788) );
  AOI22_X1 U21509 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n10447), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18353), .ZN(n18335) );
  OAI21_X1 U21510 ( .B1(n18336), .B2(n18355), .A(n18335), .ZN(P3_U2789) );
  AOI22_X1 U21511 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n10447), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18353), .ZN(n18337) );
  OAI21_X1 U21512 ( .B1(n18338), .B2(n18355), .A(n18337), .ZN(P3_U2790) );
  AOI22_X1 U21513 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n10447), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18353), .ZN(n18339) );
  OAI21_X1 U21514 ( .B1(n18340), .B2(n18355), .A(n18339), .ZN(P3_U2791) );
  AOI22_X1 U21515 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n10447), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18353), .ZN(n18341) );
  OAI21_X1 U21516 ( .B1(n18342), .B2(n18355), .A(n18341), .ZN(P3_U2792) );
  AOI22_X1 U21517 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n10447), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18353), .ZN(n18343) );
  OAI21_X1 U21518 ( .B1(n18344), .B2(n18355), .A(n18343), .ZN(P3_U2793) );
  AOI22_X1 U21519 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n10447), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18353), .ZN(n18345) );
  OAI21_X1 U21520 ( .B1(n18346), .B2(n18355), .A(n18345), .ZN(P3_U2794) );
  AOI22_X1 U21521 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n10447), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18353), .ZN(n18347) );
  OAI21_X1 U21522 ( .B1(n18348), .B2(n18355), .A(n18347), .ZN(P3_U2795) );
  AOI22_X1 U21523 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n10447), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18353), .ZN(n18349) );
  OAI21_X1 U21524 ( .B1(n18350), .B2(n18355), .A(n18349), .ZN(P3_U2796) );
  AOI22_X1 U21525 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n10447), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18353), .ZN(n18351) );
  OAI21_X1 U21526 ( .B1(n18352), .B2(n18355), .A(n18351), .ZN(P3_U2797) );
  AOI22_X1 U21527 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n10447), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18353), .ZN(n18354) );
  OAI21_X1 U21528 ( .B1(n18356), .B2(n18355), .A(n18354), .ZN(P3_U2798) );
  AOI21_X1 U21529 ( .B1(n18357), .B2(n19336), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18368) );
  AOI22_X1 U21530 ( .A1(n13496), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n18358), 
        .B2(n18681), .ZN(n18367) );
  INV_X1 U21531 ( .A(n18359), .ZN(n18393) );
  INV_X1 U21532 ( .A(n18360), .ZN(n18365) );
  OAI22_X1 U21533 ( .A1(n18363), .A2(n18556), .B1(n18362), .B2(n18361), .ZN(
        n18364) );
  AOI21_X1 U21534 ( .B1(n18393), .B2(n18365), .A(n18364), .ZN(n18366) );
  OAI211_X1 U21535 ( .C1(n18369), .C2(n18368), .A(n18367), .B(n18366), .ZN(
        P3_U2804) );
  XOR2_X1 U21536 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n18370), .Z(
        n18693) );
  OAI21_X1 U21537 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18439), .A(
        n18371), .ZN(n18384) );
  NOR2_X1 U21538 ( .A1(n18519), .A2(n18372), .ZN(n18386) );
  OAI211_X1 U21539 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n18386), .B(n18373), .ZN(n18374) );
  NAND2_X1 U21540 ( .A1(n18953), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18700) );
  OAI211_X1 U21541 ( .C1(n18530), .C2(n18375), .A(n18374), .B(n18700), .ZN(
        n18381) );
  XNOR2_X1 U21542 ( .A(n18376), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18696) );
  MUX2_X1 U21543 ( .A(n18378), .B(n18377), .S(n18583), .Z(n18379) );
  XOR2_X1 U21544 ( .A(n18379), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18695) );
  OAI22_X1 U21545 ( .A1(n18586), .A2(n18696), .B1(n18556), .B2(n18695), .ZN(
        n18380) );
  AOI211_X1 U21546 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n18384), .A(
        n18381), .B(n18380), .ZN(n18382) );
  OAI21_X1 U21547 ( .B1(n18612), .B2(n18693), .A(n18382), .ZN(P3_U2805) );
  AOI221_X1 U21548 ( .B1(n18386), .B2(n18385), .C1(n18384), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18383), .ZN(n18395) );
  INV_X1 U21549 ( .A(n18387), .ZN(n18390) );
  OAI22_X1 U21550 ( .A1(n18390), .A2(n18389), .B1(n18388), .B2(n18556), .ZN(
        n18391) );
  AOI21_X1 U21551 ( .B1(n18393), .B2(n18392), .A(n18391), .ZN(n18394) );
  OAI211_X1 U21552 ( .C1(n18530), .C2(n18396), .A(n18395), .B(n18394), .ZN(
        P3_U2806) );
  INV_X1 U21553 ( .A(n18713), .ZN(n18397) );
  NAND2_X1 U21554 ( .A1(n18398), .A2(n18397), .ZN(n18412) );
  AOI21_X1 U21555 ( .B1(n18713), .B2(n18424), .A(n18423), .ZN(n18422) );
  NOR2_X1 U21556 ( .A1(n18708), .A2(n18713), .ZN(n18400) );
  OAI21_X1 U21557 ( .B1(n18401), .B2(n18400), .A(n18399), .ZN(n18402) );
  XNOR2_X1 U21558 ( .A(n18402), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18725) );
  OAI21_X1 U21559 ( .B1(n18403), .B2(n18439), .A(n18672), .ZN(n18404) );
  AOI21_X1 U21560 ( .B1(n18579), .B2(n18405), .A(n18404), .ZN(n18428) );
  OAI21_X1 U21561 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18426), .A(
        n18428), .ZN(n18415) );
  AOI22_X1 U21562 ( .A1(n13496), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18415), .ZN(n18408) );
  NOR2_X1 U21563 ( .A1(n18519), .A2(n18405), .ZN(n18417) );
  OAI211_X1 U21564 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n18417), .B(n18406), .ZN(n18407) );
  OAI211_X1 U21565 ( .C1(n18409), .C2(n18530), .A(n18408), .B(n18407), .ZN(
        n18410) );
  AOI21_X1 U21566 ( .B1(n18588), .B2(n18725), .A(n18410), .ZN(n18411) );
  OAI221_X1 U21567 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18412), 
        .C1(n18717), .C2(n18422), .A(n18411), .ZN(P3_U2808) );
  OAI22_X1 U21568 ( .A1(n18840), .A2(n19507), .B1(n18530), .B2(n18413), .ZN(
        n18414) );
  AOI221_X1 U21569 ( .B1(n18417), .B2(n18416), .C1(n18415), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18414), .ZN(n18421) );
  INV_X1 U21570 ( .A(n18464), .ZN(n18447) );
  NAND3_X1 U21571 ( .A1(n10105), .A2(n10114), .A3(n18737), .ZN(n18448) );
  INV_X1 U21572 ( .A(n18448), .ZN(n18433) );
  AOI22_X1 U21573 ( .A1(n18447), .A2(n18418), .B1(n18433), .B2(n18734), .ZN(
        n18419) );
  XNOR2_X1 U21574 ( .A(n18419), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n18739) );
  NOR2_X1 U21575 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18718), .ZN(
        n18738) );
  INV_X1 U21576 ( .A(n18737), .ZN(n18729) );
  NOR2_X1 U21577 ( .A1(n18729), .A2(n18481), .ZN(n18450) );
  AOI22_X1 U21578 ( .A1(n18588), .A2(n18739), .B1(n18738), .B2(n18450), .ZN(
        n18420) );
  OAI211_X1 U21579 ( .C1(n18422), .C2(n18716), .A(n18421), .B(n18420), .ZN(
        P3_U2809) );
  NAND2_X1 U21580 ( .A1(n18737), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18745) );
  AOI21_X1 U21581 ( .B1(n18745), .B2(n18424), .A(n18423), .ZN(n18453) );
  INV_X1 U21582 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18714) );
  INV_X1 U21583 ( .A(n18425), .ZN(n18431) );
  INV_X1 U21584 ( .A(n18426), .ZN(n18430) );
  AOI21_X1 U21585 ( .B1(n9769), .B2(n19336), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18427) );
  OAI22_X1 U21586 ( .A1(n18428), .A2(n18427), .B1(n18840), .B2(n19506), .ZN(
        n18429) );
  AOI221_X1 U21587 ( .B1(n18432), .B2(n18431), .C1(n18430), .C2(n18431), .A(
        n18429), .ZN(n18438) );
  OAI22_X1 U21588 ( .A1(n18433), .A2(n18756), .B1(n18462), .B2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18434) );
  NOR2_X1 U21589 ( .A1(n18435), .A2(n18434), .ZN(n18436) );
  XNOR2_X1 U21590 ( .A(n18436), .B(n18714), .ZN(n18744) );
  NOR2_X1 U21591 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18756), .ZN(
        n18742) );
  AOI22_X1 U21592 ( .A1(n18588), .A2(n18744), .B1(n18450), .B2(n18742), .ZN(
        n18437) );
  OAI211_X1 U21593 ( .C1(n18453), .C2(n18714), .A(n18438), .B(n18437), .ZN(
        P3_U2810) );
  AOI21_X1 U21594 ( .B1(n18579), .B2(n18454), .A(n18658), .ZN(n18473) );
  OAI21_X1 U21595 ( .B1(n18440), .B2(n18439), .A(n18473), .ZN(n18457) );
  NOR2_X1 U21596 ( .A1(n18840), .A2(n19504), .ZN(n18752) );
  AOI211_X1 U21597 ( .C1(n18458), .C2(n18441), .A(n18454), .B(n18519), .ZN(
        n18442) );
  INV_X1 U21598 ( .A(n18442), .ZN(n18444) );
  OAI22_X1 U21599 ( .A1(n18445), .A2(n18444), .B1(n18443), .B2(n18530), .ZN(
        n18446) );
  AOI211_X1 U21600 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n18457), .A(
        n18752), .B(n18446), .ZN(n18452) );
  NAND2_X1 U21601 ( .A1(n18447), .A2(n18462), .ZN(n18467) );
  NAND2_X1 U21602 ( .A1(n18467), .A2(n18448), .ZN(n18449) );
  XNOR2_X1 U21603 ( .A(n18449), .B(n18756), .ZN(n18753) );
  AOI22_X1 U21604 ( .A1(n18588), .A2(n18753), .B1(n18450), .B2(n18756), .ZN(
        n18451) );
  OAI211_X1 U21605 ( .C1(n18453), .C2(n18756), .A(n18452), .B(n18451), .ZN(
        P3_U2811) );
  NAND2_X1 U21606 ( .A1(n18461), .A2(n21475), .ZN(n18772) );
  NOR2_X1 U21607 ( .A1(n18519), .A2(n18454), .ZN(n18459) );
  OAI22_X1 U21608 ( .A1(n18840), .A2(n19501), .B1(n18530), .B2(n18455), .ZN(
        n18456) );
  AOI221_X1 U21609 ( .B1(n18459), .B2(n18458), .C1(n18457), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18456), .ZN(n18470) );
  OAI21_X1 U21610 ( .B1(n18461), .B2(n18481), .A(n18460), .ZN(n18478) );
  NAND2_X1 U21611 ( .A1(n10114), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18466) );
  INV_X1 U21612 ( .A(n18462), .ZN(n18463) );
  NAND2_X1 U21613 ( .A1(n18463), .A2(n18466), .ZN(n18465) );
  MUX2_X1 U21614 ( .A(n18466), .B(n18465), .S(n18464), .Z(n18468) );
  NAND2_X1 U21615 ( .A1(n18468), .A2(n18467), .ZN(n18767) );
  AOI22_X1 U21616 ( .A1(n18478), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n18588), .B2(n18767), .ZN(n18469) );
  OAI211_X1 U21617 ( .C1(n18481), .C2(n18772), .A(n18470), .B(n18469), .ZN(
        P3_U2812) );
  NAND2_X1 U21618 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18773), .ZN(
        n18779) );
  AOI21_X1 U21619 ( .B1(n18471), .B2(n19336), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18474) );
  OAI22_X1 U21620 ( .A1(n18474), .A2(n18473), .B1(n18667), .B2(n18472), .ZN(
        n18475) );
  AOI21_X1 U21621 ( .B1(n13496), .B2(P3_REIP_REG_17__SCAN_IN), .A(n18475), 
        .ZN(n18480) );
  XNOR2_X1 U21622 ( .A(n18476), .B(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18775) );
  INV_X1 U21623 ( .A(n18775), .ZN(n18477) );
  AOI22_X1 U21624 ( .A1(n18478), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n18588), .B2(n18477), .ZN(n18479) );
  OAI211_X1 U21625 ( .C1(n18481), .C2(n18779), .A(n18480), .B(n18479), .ZN(
        P3_U2813) );
  NOR2_X1 U21626 ( .A1(n18840), .A2(n19495), .ZN(n18482) );
  AOI221_X1 U21627 ( .B1(n18485), .B2(n18484), .C1(n18483), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18482), .ZN(n18496) );
  INV_X1 U21628 ( .A(n18486), .ZN(n18494) );
  OAI21_X1 U21629 ( .B1(n18866), .B2(n18487), .A(n18811), .ZN(n18807) );
  INV_X1 U21630 ( .A(n18508), .ZN(n18813) );
  NAND2_X1 U21631 ( .A1(n18563), .A2(n18813), .ZN(n18504) );
  OAI21_X1 U21632 ( .B1(n18489), .B2(n18504), .A(n18488), .ZN(n18490) );
  INV_X1 U21633 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18817) );
  NAND2_X1 U21634 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18817), .ZN(
        n18844) );
  NAND2_X1 U21635 ( .A1(n18490), .A2(n18844), .ZN(n18491) );
  XNOR2_X1 U21636 ( .A(n18491), .B(n18811), .ZN(n18805) );
  AND2_X1 U21637 ( .A1(n18509), .A2(n18811), .ZN(n18799) );
  OAI22_X1 U21638 ( .A1(n18805), .A2(n18556), .B1(n18799), .B2(n18492), .ZN(
        n18493) );
  AOI21_X1 U21639 ( .B1(n18494), .B2(n18807), .A(n18493), .ZN(n18495) );
  OAI211_X1 U21640 ( .C1(n18530), .C2(n18497), .A(n18496), .B(n18495), .ZN(
        P3_U2815) );
  NOR2_X1 U21641 ( .A1(n18866), .A2(n18508), .ZN(n18830) );
  NAND2_X1 U21642 ( .A1(n18814), .A2(n18498), .ZN(n18499) );
  OAI221_X1 U21643 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18830), .A(n18499), .ZN(
        n18827) );
  OR2_X1 U21644 ( .A1(n18518), .A2(n19015), .ZN(n18545) );
  AOI221_X1 U21645 ( .B1(n18520), .B2(n18501), .C1(n18545), .C2(n18501), .A(
        n18500), .ZN(n18502) );
  INV_X1 U21646 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19494) );
  NOR2_X1 U21647 ( .A1(n18840), .A2(n19494), .ZN(n18821) );
  AOI211_X1 U21648 ( .C1(n18503), .C2(n18681), .A(n18502), .B(n18821), .ZN(
        n18514) );
  INV_X1 U21649 ( .A(n18504), .ZN(n18505) );
  OAI21_X1 U21650 ( .B1(n18506), .B2(n18505), .A(n18844), .ZN(n18507) );
  XOR2_X1 U21651 ( .A(n18489), .B(n18507), .Z(n18824) );
  NOR2_X1 U21652 ( .A1(n18581), .A2(n18508), .ZN(n18834) );
  NAND2_X1 U21653 ( .A1(n18834), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18511) );
  INV_X1 U21654 ( .A(n18509), .ZN(n18510) );
  AOI21_X1 U21655 ( .B1(n18511), .B2(n18489), .A(n18510), .ZN(n18822) );
  AOI22_X1 U21656 ( .A1(n18824), .A2(n18588), .B1(n18512), .B2(n18822), .ZN(
        n18513) );
  OAI211_X1 U21657 ( .C1(n18612), .C2(n18827), .A(n18514), .B(n18513), .ZN(
        P3_U2816) );
  NAND2_X1 U21658 ( .A1(n18554), .A2(n18831), .ZN(n18541) );
  AOI22_X1 U21659 ( .A1(n18516), .A2(n18515), .B1(n18579), .B2(n18518), .ZN(
        n18517) );
  NAND2_X1 U21660 ( .A1(n18517), .A2(n18672), .ZN(n18532) );
  NOR2_X1 U21661 ( .A1(n18519), .A2(n18518), .ZN(n18534) );
  OAI211_X1 U21662 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18534), .B(n18520), .ZN(n18522) );
  NAND2_X1 U21663 ( .A1(n18953), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n18521) );
  OAI211_X1 U21664 ( .C1(n18530), .C2(n18523), .A(n18522), .B(n18521), .ZN(
        n18524) );
  AOI21_X1 U21665 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18532), .A(
        n18524), .ZN(n18528) );
  OAI22_X1 U21666 ( .A1(n18830), .A2(n18612), .B1(n18834), .B2(n18586), .ZN(
        n18538) );
  INV_X1 U21667 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18854) );
  AOI21_X1 U21668 ( .B1(n18583), .B2(n18854), .A(n18834), .ZN(n18525) );
  AOI21_X1 U21669 ( .B1(n18583), .B2(n18536), .A(n18525), .ZN(n18526) );
  XOR2_X1 U21670 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18526), .Z(
        n18828) );
  AOI22_X1 U21671 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18538), .B1(
        n18588), .B2(n18828), .ZN(n18527) );
  OAI211_X1 U21672 ( .C1(n18844), .C2(n18541), .A(n18528), .B(n18527), .ZN(
        P3_U2817) );
  NAND2_X1 U21673 ( .A1(n18953), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18852) );
  OAI21_X1 U21674 ( .B1(n18530), .B2(n18529), .A(n18852), .ZN(n18531) );
  AOI221_X1 U21675 ( .B1(n18534), .B2(n18533), .C1(n18532), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n18531), .ZN(n18540) );
  NAND2_X1 U21676 ( .A1(n18536), .A2(n18535), .ZN(n18537) );
  XNOR2_X1 U21677 ( .A(n18537), .B(n18854), .ZN(n18851) );
  AOI22_X1 U21678 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18538), .B1(
        n18588), .B2(n18851), .ZN(n18539) );
  OAI211_X1 U21679 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18541), .A(
        n18540), .B(n18539), .ZN(P3_U2818) );
  AND2_X1 U21680 ( .A1(n18563), .A2(n18869), .ZN(n18569) );
  INV_X1 U21681 ( .A(n18569), .ZN(n18542) );
  NAND2_X1 U21682 ( .A1(n18543), .A2(n18542), .ZN(n18544) );
  XNOR2_X1 U21683 ( .A(n18544), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18874) );
  INV_X1 U21684 ( .A(n18869), .ZN(n18550) );
  NOR2_X1 U21685 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18550), .ZN(
        n18856) );
  NOR2_X1 U21686 ( .A1(n18558), .A2(n18559), .ZN(n18557) );
  OAI211_X1 U21687 ( .C1(n18557), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n18546), .B(n18545), .ZN(n18548) );
  NAND2_X1 U21688 ( .A1(n18953), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n18547) );
  OAI211_X1 U21689 ( .C1(n18667), .C2(n18549), .A(n18548), .B(n18547), .ZN(
        n18553) );
  NAND2_X1 U21690 ( .A1(n18554), .A2(n18550), .ZN(n18577) );
  AOI21_X1 U21691 ( .B1(n18551), .B2(n18577), .A(n9875), .ZN(n18552) );
  AOI211_X1 U21692 ( .C1(n18856), .C2(n18554), .A(n18553), .B(n18552), .ZN(
        n18555) );
  OAI21_X1 U21693 ( .B1(n18874), .B2(n18556), .A(n18555), .ZN(P3_U2819) );
  AOI211_X1 U21694 ( .C1(n18559), .C2(n18558), .A(n18685), .B(n18557), .ZN(
        n18561) );
  NOR2_X1 U21695 ( .A1(n18840), .A2(n19486), .ZN(n18560) );
  AOI211_X1 U21696 ( .C1(n18562), .C2(n18681), .A(n18561), .B(n18560), .ZN(
        n18576) );
  NAND2_X1 U21697 ( .A1(n18563), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18564) );
  NAND2_X1 U21698 ( .A1(n18564), .A2(n16931), .ZN(n18565) );
  OR2_X1 U21699 ( .A1(n18566), .A2(n18565), .ZN(n18573) );
  NAND2_X1 U21700 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18882), .ZN(
        n18567) );
  NOR2_X1 U21701 ( .A1(n18568), .A2(n18567), .ZN(n18570) );
  AOI21_X1 U21702 ( .B1(n18571), .B2(n18570), .A(n18569), .ZN(n18572) );
  AND2_X1 U21703 ( .A1(n18573), .A2(n18572), .ZN(n18877) );
  AOI22_X1 U21704 ( .A1(n18574), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n18588), .B2(n18877), .ZN(n18575) );
  OAI211_X1 U21705 ( .C1(n18578), .C2(n18577), .A(n18576), .B(n18575), .ZN(
        P3_U2820) );
  INV_X1 U21706 ( .A(n18579), .ZN(n18641) );
  OAI21_X1 U21707 ( .B1(n10144), .B2(n18641), .A(n18672), .ZN(n18595) );
  AOI22_X1 U21708 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18595), .B1(
        n18580), .B2(n18681), .ZN(n18593) );
  NAND2_X1 U21709 ( .A1(n18582), .A2(n18581), .ZN(n18889) );
  XNOR2_X1 U21710 ( .A(n18889), .B(n18583), .ZN(n18893) );
  OAI21_X1 U21711 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18585), .A(
        n18584), .ZN(n18891) );
  OAI22_X1 U21712 ( .A1(n18891), .A2(n18612), .B1(n18586), .B2(n18889), .ZN(
        n18587) );
  AOI21_X1 U21713 ( .B1(n18588), .B2(n18893), .A(n18587), .ZN(n18592) );
  NAND2_X1 U21714 ( .A1(n18953), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18903) );
  OAI211_X1 U21715 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18590), .A(
        n19336), .B(n18589), .ZN(n18591) );
  NAND4_X1 U21716 ( .A1(n18593), .A2(n18592), .A3(n18903), .A4(n18591), .ZN(
        P3_U2822) );
  NOR2_X1 U21717 ( .A1(n18594), .A2(n19015), .ZN(n18597) );
  NOR2_X1 U21718 ( .A1(n18840), .A2(n19479), .ZN(n18905) );
  AOI221_X1 U21719 ( .B1(n18597), .B2(n18596), .C1(n18595), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18905), .ZN(n18605) );
  NOR2_X1 U21720 ( .A1(n18599), .A2(n18598), .ZN(n18600) );
  XOR2_X1 U21721 ( .A(n18600), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18908) );
  OR2_X1 U21722 ( .A1(n18601), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18602) );
  AND2_X1 U21723 ( .A1(n18603), .A2(n18602), .ZN(n18907) );
  AOI22_X1 U21724 ( .A1(n18908), .A2(n18675), .B1(n18680), .B2(n18907), .ZN(
        n18604) );
  OAI211_X1 U21725 ( .C1(n18667), .C2(n18606), .A(n18605), .B(n18604), .ZN(
        P3_U2823) );
  NAND2_X1 U21726 ( .A1(n18615), .A2(n19336), .ZN(n18613) );
  INV_X1 U21727 ( .A(n18609), .ZN(n18607) );
  AOI22_X1 U21728 ( .A1(n18609), .A2(n18626), .B1(n18608), .B2(n18607), .ZN(
        n18610) );
  XOR2_X1 U21729 ( .A(n18611), .B(n18610), .Z(n18924) );
  OAI22_X1 U21730 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18613), .B1(
        n18924), .B2(n18612), .ZN(n18614) );
  AOI21_X1 U21731 ( .B1(n13496), .B2(P3_REIP_REG_6__SCAN_IN), .A(n18614), .ZN(
        n18621) );
  AOI21_X1 U21732 ( .B1(n19336), .B2(n18615), .A(n18685), .ZN(n18632) );
  OAI21_X1 U21733 ( .B1(n18618), .B2(n18617), .A(n18616), .ZN(n18619) );
  INV_X1 U21734 ( .A(n18619), .ZN(n18915) );
  AOI22_X1 U21735 ( .A1(n18632), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n18680), .B2(n18915), .ZN(n18620) );
  OAI211_X1 U21736 ( .C1(n18667), .C2(n18622), .A(n18621), .B(n18620), .ZN(
        P3_U2824) );
  OR2_X1 U21737 ( .A1(n18623), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18624) );
  AND2_X1 U21738 ( .A1(n18625), .A2(n18624), .ZN(n18926) );
  AOI22_X1 U21739 ( .A1(n18680), .A2(n18926), .B1(n18953), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n18634) );
  AOI21_X1 U21740 ( .B1(n18628), .B2(n18627), .A(n18626), .ZN(n18925) );
  OAI21_X1 U21741 ( .B1(n18658), .B2(n18630), .A(n18629), .ZN(n18631) );
  AOI22_X1 U21742 ( .A1(n18675), .A2(n18925), .B1(n18632), .B2(n18631), .ZN(
        n18633) );
  OAI211_X1 U21743 ( .C1(n18667), .C2(n18635), .A(n18634), .B(n18633), .ZN(
        P3_U2825) );
  AOI21_X1 U21744 ( .B1(n18638), .B2(n18637), .A(n18636), .ZN(n18933) );
  OAI22_X1 U21745 ( .A1(n18840), .A2(n19473), .B1(n19015), .B2(n18639), .ZN(
        n18640) );
  AOI21_X1 U21746 ( .B1(n18675), .B2(n18933), .A(n18640), .ZN(n18648) );
  OAI21_X1 U21747 ( .B1(n18642), .B2(n18641), .A(n18672), .ZN(n18660) );
  OAI21_X1 U21748 ( .B1(n18645), .B2(n18644), .A(n18643), .ZN(n18646) );
  INV_X1 U21749 ( .A(n18646), .ZN(n18935) );
  AOI22_X1 U21750 ( .A1(n18660), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n18680), .B2(n18935), .ZN(n18647) );
  OAI211_X1 U21751 ( .C1(n18667), .C2(n18649), .A(n18648), .B(n18647), .ZN(
        P3_U2826) );
  OAI21_X1 U21752 ( .B1(n18652), .B2(n18651), .A(n18650), .ZN(n18653) );
  INV_X1 U21753 ( .A(n18653), .ZN(n18941) );
  AOI22_X1 U21754 ( .A1(n18680), .A2(n18941), .B1(n13496), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n18662) );
  AOI21_X1 U21755 ( .B1(n18656), .B2(n18655), .A(n18654), .ZN(n18942) );
  OAI21_X1 U21756 ( .B1(n18658), .B2(n18673), .A(n18657), .ZN(n18659) );
  AOI22_X1 U21757 ( .A1(n18675), .A2(n18942), .B1(n18660), .B2(n18659), .ZN(
        n18661) );
  OAI211_X1 U21758 ( .C1(n18667), .C2(n18663), .A(n18662), .B(n18661), .ZN(
        P3_U2827) );
  INV_X1 U21759 ( .A(n18680), .ZN(n18664) );
  OAI22_X1 U21760 ( .A1(n18667), .A2(n18666), .B1(n18665), .B2(n18664), .ZN(
        n18668) );
  AOI211_X1 U21761 ( .C1(n18675), .C2(n18670), .A(n18669), .B(n18668), .ZN(
        n18671) );
  OAI221_X1 U21762 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19015), .C1(
        n18673), .C2(n18672), .A(n18671), .ZN(P3_U2828) );
  XOR2_X1 U21763 ( .A(n18674), .B(n18678), .Z(n18951) );
  AOI22_X1 U21764 ( .A1(n18675), .A2(n18951), .B1(n13496), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18683) );
  OAI21_X1 U21765 ( .B1(n18678), .B2(n18677), .A(n18676), .ZN(n18679) );
  INV_X1 U21766 ( .A(n18679), .ZN(n18949) );
  AOI22_X1 U21767 ( .A1(n18681), .A2(n18684), .B1(n18680), .B2(n18949), .ZN(
        n18682) );
  OAI211_X1 U21768 ( .C1(n18685), .C2(n18684), .A(n18683), .B(n18682), .ZN(
        P3_U2829) );
  NAND4_X1 U21769 ( .A1(n18687), .A2(n18686), .A3(n18812), .A4(n10359), .ZN(
        n18688) );
  NOR3_X1 U21770 ( .A1(n18765), .A2(n18689), .A3(n18688), .ZN(n18699) );
  AOI221_X1 U21771 ( .B1(n18692), .B2(n19406), .C1(n18691), .C2(n19406), .A(
        n18690), .ZN(n18694) );
  OAI22_X1 U21772 ( .A1(n18694), .A2(n10359), .B1(n18829), .B2(n18693), .ZN(
        n18698) );
  OAI22_X1 U21773 ( .A1(n18890), .A2(n18696), .B1(n18873), .B2(n18695), .ZN(
        n18697) );
  AOI221_X1 U21774 ( .B1(n18699), .B2(n18944), .C1(n18698), .C2(n18944), .A(
        n18697), .ZN(n18701) );
  OAI211_X1 U21775 ( .C1(n18855), .C2(n10359), .A(n18701), .B(n18700), .ZN(
        P3_U2837) );
  OAI21_X1 U21776 ( .B1(n18955), .B2(n18703), .A(n18702), .ZN(n18704) );
  AOI22_X1 U21777 ( .A1(n18894), .A2(n18706), .B1(n18705), .B2(n18704), .ZN(
        n18707) );
  OAI21_X1 U21778 ( .B1(n18840), .B2(n19511), .A(n18707), .ZN(P3_U2839) );
  NAND2_X1 U21779 ( .A1(n18712), .A2(n18708), .ZN(n18798) );
  OAI21_X1 U21780 ( .B1(n18709), .B2(n18829), .A(n18798), .ZN(n18730) );
  AOI21_X1 U21781 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18762), .A(
        n18896), .ZN(n18710) );
  AOI221_X1 U21782 ( .B1(n18711), .B2(n18958), .C1(n18745), .C2(n18958), .A(
        n18710), .ZN(n18731) );
  NOR2_X1 U21783 ( .A1(n19404), .A2(n18712), .ZN(n18867) );
  INV_X1 U21784 ( .A(n18867), .ZN(n18764) );
  AOI22_X1 U21785 ( .A1(n18958), .A2(n18714), .B1(n18713), .B2(n18764), .ZN(
        n18733) );
  AOI22_X1 U21786 ( .A1(n18875), .A2(n18716), .B1(n18861), .B2(n18715), .ZN(
        n18720) );
  AOI21_X1 U21787 ( .B1(n19406), .B2(n18718), .A(n18717), .ZN(n18719) );
  NAND4_X1 U21788 ( .A1(n18731), .A2(n18733), .A3(n18720), .A4(n18719), .ZN(
        n18724) );
  AND2_X1 U21789 ( .A1(n18722), .A2(n18721), .ZN(n18723) );
  OAI22_X1 U21790 ( .A1(n18730), .A2(n18724), .B1(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18723), .ZN(n18728) );
  AOI22_X1 U21791 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18955), .B1(
        n18894), .B2(n18725), .ZN(n18727) );
  NAND2_X1 U21792 ( .A1(n18953), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18726) );
  OAI211_X1 U21793 ( .C1(n18899), .C2(n18728), .A(n18727), .B(n18726), .ZN(
        P3_U2840) );
  NOR3_X1 U21794 ( .A1(n18729), .A2(n18786), .A3(n18785), .ZN(n18732) );
  NOR2_X1 U21795 ( .A1(n18730), .A2(n18899), .ZN(n18791) );
  OAI211_X1 U21796 ( .C1(n18868), .C2(n18732), .A(n18791), .B(n18731), .ZN(
        n18746) );
  OAI21_X1 U21797 ( .B1(n18734), .B2(n18747), .A(n18733), .ZN(n18735) );
  OAI21_X1 U21798 ( .B1(n18746), .B2(n18735), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18741) );
  INV_X1 U21799 ( .A(n18797), .ZN(n18736) );
  NAND2_X1 U21800 ( .A1(n18737), .A2(n18736), .ZN(n18757) );
  INV_X1 U21801 ( .A(n18757), .ZN(n18743) );
  AOI22_X1 U21802 ( .A1(n18894), .A2(n18739), .B1(n18738), .B2(n18743), .ZN(
        n18740) );
  OAI221_X1 U21803 ( .B1(n13496), .B2(n18741), .C1(n18840), .C2(n19507), .A(
        n18740), .ZN(P3_U2841) );
  AOI22_X1 U21804 ( .A1(n18894), .A2(n18744), .B1(n18743), .B2(n18742), .ZN(
        n18751) );
  OAI221_X1 U21805 ( .B1(n18746), .B2(n18745), .C1(n18746), .C2(n18764), .A(
        n18840), .ZN(n18755) );
  INV_X1 U21806 ( .A(n18755), .ZN(n18749) );
  NOR3_X1 U21807 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18747), .A3(
        n19555), .ZN(n18748) );
  OAI21_X1 U21808 ( .B1(n18749), .B2(n18748), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18750) );
  OAI211_X1 U21809 ( .C1(n19506), .C2(n18840), .A(n18751), .B(n18750), .ZN(
        P3_U2842) );
  AOI21_X1 U21810 ( .B1(n18894), .B2(n18753), .A(n18752), .ZN(n18754) );
  OAI221_X1 U21811 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18757), 
        .C1(n18756), .C2(n18755), .A(n18754), .ZN(P3_U2843) );
  OAI21_X1 U21812 ( .B1(n18782), .B2(n18766), .A(n18758), .ZN(n18897) );
  OAI21_X1 U21813 ( .B1(n18785), .B2(n18760), .A(n18759), .ZN(n18761) );
  OAI211_X1 U21814 ( .C1(n18762), .C2(n18896), .A(n18791), .B(n18761), .ZN(
        n18763) );
  AOI211_X1 U21815 ( .C1(n18765), .C2(n18764), .A(n18897), .B(n18763), .ZN(
        n18774) );
  OAI21_X1 U21816 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18766), .A(
        n18774), .ZN(n18769) );
  NOR2_X1 U21817 ( .A1(n13496), .A2(n21475), .ZN(n18768) );
  AOI22_X1 U21818 ( .A1(n18769), .A2(n18768), .B1(n18894), .B2(n18767), .ZN(
        n18771) );
  NAND2_X1 U21819 ( .A1(n18953), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18770) );
  OAI211_X1 U21820 ( .C1(n18772), .C2(n18797), .A(n18771), .B(n18770), .ZN(
        P3_U2844) );
  NOR3_X1 U21821 ( .A1(n18774), .A2(n18953), .A3(n18773), .ZN(n18777) );
  OAI22_X1 U21822 ( .A1(n18775), .A2(n18873), .B1(n19500), .B2(n18840), .ZN(
        n18776) );
  NOR2_X1 U21823 ( .A1(n18777), .A2(n18776), .ZN(n18778) );
  OAI21_X1 U21824 ( .B1(n18797), .B2(n18779), .A(n18778), .ZN(P3_U2845) );
  NAND2_X1 U21825 ( .A1(n19406), .A2(n18780), .ZN(n18781) );
  OAI221_X1 U21826 ( .B1(n18784), .B2(n18783), .C1(n18784), .C2(n18782), .A(
        n18781), .ZN(n18859) );
  NOR2_X1 U21827 ( .A1(n18786), .A2(n18785), .ZN(n18787) );
  AOI21_X1 U21828 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18868), .A(
        n18787), .ZN(n18788) );
  INV_X1 U21829 ( .A(n18788), .ZN(n18789) );
  OAI21_X1 U21830 ( .B1(n18814), .B2(n18839), .A(n18789), .ZN(n18790) );
  NOR2_X1 U21831 ( .A1(n18859), .A2(n18790), .ZN(n18800) );
  AOI221_X1 U21832 ( .B1(n18792), .B2(n18791), .C1(n18800), .C2(n18791), .A(
        n13496), .ZN(n18794) );
  AOI22_X1 U21833 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18794), .B1(
        n18894), .B2(n18793), .ZN(n18796) );
  NAND2_X1 U21834 ( .A1(n18953), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n18795) );
  OAI211_X1 U21835 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n18797), .A(
        n18796), .B(n18795), .ZN(P3_U2846) );
  AOI21_X1 U21836 ( .B1(n18812), .B2(n18814), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18801) );
  OAI22_X1 U21837 ( .A1(n18801), .A2(n18800), .B1(n18799), .B2(n18798), .ZN(
        n18802) );
  INV_X1 U21838 ( .A(n18802), .ZN(n18803) );
  OAI21_X1 U21839 ( .B1(n18805), .B2(n18804), .A(n18803), .ZN(n18806) );
  AOI22_X1 U21840 ( .A1(n13496), .A2(P3_REIP_REG_15__SCAN_IN), .B1(n18944), 
        .B2(n18806), .ZN(n18810) );
  NAND3_X1 U21841 ( .A1(n18952), .A2(n18808), .A3(n18807), .ZN(n18809) );
  OAI211_X1 U21842 ( .C1(n18855), .C2(n18811), .A(n18810), .B(n18809), .ZN(
        P3_U2847) );
  NAND4_X1 U21843 ( .A1(n18831), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(n18812), .ZN(n18819) );
  NAND2_X1 U21844 ( .A1(n18858), .A2(n18813), .ZN(n18845) );
  NAND2_X1 U21845 ( .A1(n18861), .A2(n18845), .ZN(n18838) );
  OAI211_X1 U21846 ( .C1(n18814), .C2(n18839), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18838), .ZN(n18815) );
  AOI211_X1 U21847 ( .C1(n18817), .C2(n18816), .A(n18859), .B(n18815), .ZN(
        n18818) );
  AOI211_X1 U21848 ( .C1(n18489), .C2(n18819), .A(n18818), .B(n18899), .ZN(
        n18820) );
  AOI211_X1 U21849 ( .C1(n18955), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18821), .B(n18820), .ZN(n18826) );
  AOI22_X1 U21850 ( .A1(n18824), .A2(n18894), .B1(n18823), .B2(n18822), .ZN(
        n18825) );
  OAI211_X1 U21851 ( .C1(n18923), .C2(n18827), .A(n18826), .B(n18825), .ZN(
        P3_U2848) );
  NAND2_X1 U21852 ( .A1(n18831), .A2(n18881), .ZN(n18848) );
  AOI22_X1 U21853 ( .A1(n13496), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18894), 
        .B2(n18828), .ZN(n18843) );
  OR2_X1 U21854 ( .A1(n18830), .A2(n18829), .ZN(n18837) );
  INV_X1 U21855 ( .A(n18859), .ZN(n18833) );
  INV_X1 U21856 ( .A(n18831), .ZN(n18832) );
  NAND2_X1 U21857 ( .A1(n18875), .A2(n18832), .ZN(n18857) );
  OAI211_X1 U21858 ( .C1(n18834), .C2(n18863), .A(n18833), .B(n18857), .ZN(
        n18835) );
  INV_X1 U21859 ( .A(n18835), .ZN(n18836) );
  AND2_X1 U21860 ( .A1(n18837), .A2(n18836), .ZN(n18846) );
  OAI211_X1 U21861 ( .C1(n18839), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18846), .B(n18838), .ZN(n18841) );
  OAI211_X1 U21862 ( .C1(n18899), .C2(n18841), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18840), .ZN(n18842) );
  OAI211_X1 U21863 ( .C1(n18848), .C2(n18844), .A(n18843), .B(n18842), .ZN(
        P3_U2849) );
  OAI21_X1 U21864 ( .B1(n18861), .B2(n18854), .A(n18845), .ZN(n18847) );
  NAND2_X1 U21865 ( .A1(n18847), .A2(n18846), .ZN(n18850) );
  OAI21_X1 U21866 ( .B1(n18899), .B2(n18854), .A(n18848), .ZN(n18849) );
  AOI22_X1 U21867 ( .A1(n18894), .A2(n18851), .B1(n18850), .B2(n18849), .ZN(
        n18853) );
  OAI211_X1 U21868 ( .C1(n18855), .C2(n18854), .A(n18853), .B(n18852), .ZN(
        P3_U2850) );
  AOI22_X1 U21869 ( .A1(n13496), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18881), 
        .B2(n18856), .ZN(n18872) );
  INV_X1 U21870 ( .A(n18857), .ZN(n18870) );
  INV_X1 U21871 ( .A(n18858), .ZN(n18860) );
  AOI211_X1 U21872 ( .C1(n18861), .C2(n18860), .A(n18899), .B(n18859), .ZN(
        n18862) );
  OAI21_X1 U21873 ( .B1(n18864), .B2(n18863), .A(n18862), .ZN(n18865) );
  AOI21_X1 U21874 ( .B1(n19404), .B2(n18866), .A(n18865), .ZN(n18883) );
  OAI221_X1 U21875 ( .B1(n18869), .B2(n18868), .C1(n18869), .C2(n18867), .A(
        n18883), .ZN(n18876) );
  OAI211_X1 U21876 ( .C1(n18870), .C2(n18876), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18840), .ZN(n18871) );
  OAI211_X1 U21877 ( .C1(n18874), .C2(n18873), .A(n18872), .B(n18871), .ZN(
        P3_U2851) );
  OAI221_X1 U21878 ( .B1(n18876), .B2(n18875), .C1(n18876), .C2(n18882), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18880) );
  NOR2_X1 U21879 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18882), .ZN(
        n18878) );
  AOI22_X1 U21880 ( .A1(n18881), .A2(n18878), .B1(n18894), .B2(n18877), .ZN(
        n18879) );
  OAI221_X1 U21881 ( .B1(n13496), .B2(n18880), .C1(n18840), .C2(n19486), .A(
        n18879), .ZN(P3_U2852) );
  INV_X1 U21882 ( .A(n18881), .ZN(n18888) );
  NOR3_X1 U21883 ( .A1(n13496), .A2(n18883), .A3(n18882), .ZN(n18884) );
  AOI211_X1 U21884 ( .C1(n18894), .C2(n18886), .A(n18885), .B(n18884), .ZN(
        n18887) );
  OAI21_X1 U21885 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18888), .A(
        n18887), .ZN(P3_U2853) );
  OAI22_X1 U21886 ( .A1(n18891), .A2(n18923), .B1(n18890), .B2(n18889), .ZN(
        n18892) );
  AOI21_X1 U21887 ( .B1(n18894), .B2(n18893), .A(n18892), .ZN(n18904) );
  NOR2_X1 U21888 ( .A1(n18896), .A2(n18895), .ZN(n18898) );
  NOR2_X1 U21889 ( .A1(n18898), .A2(n18897), .ZN(n18932) );
  AOI21_X1 U21890 ( .B1(n18900), .B2(n18932), .A(n18916), .ZN(n18910) );
  OAI21_X1 U21891 ( .B1(n18955), .B2(n18910), .A(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18902) );
  NOR2_X1 U21892 ( .A1(n18909), .A2(n18899), .ZN(n18934) );
  NAND3_X1 U21893 ( .A1(n18900), .A2(n18934), .A3(n10350), .ZN(n18901) );
  NAND4_X1 U21894 ( .A1(n18904), .A2(n18903), .A3(n18902), .A4(n18901), .ZN(
        P3_U2854) );
  AOI21_X1 U21895 ( .B1(n18955), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18905), .ZN(n18914) );
  INV_X1 U21896 ( .A(n18906), .ZN(n18950) );
  AOI22_X1 U21897 ( .A1(n18908), .A2(n18952), .B1(n18950), .B2(n18907), .ZN(
        n18913) );
  INV_X1 U21898 ( .A(n18909), .ZN(n18945) );
  OAI221_X1 U21899 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18911), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18945), .A(n18910), .ZN(
        n18912) );
  NAND3_X1 U21900 ( .A1(n18914), .A2(n18913), .A3(n18912), .ZN(P3_U2855) );
  AOI22_X1 U21901 ( .A1(n18950), .A2(n18915), .B1(n13496), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n18922) );
  INV_X1 U21902 ( .A(n18919), .ZN(n18917) );
  AOI21_X1 U21903 ( .B1(n18932), .B2(n18917), .A(n18916), .ZN(n18918) );
  OR2_X1 U21904 ( .A1(n18918), .A2(n18955), .ZN(n18927) );
  NOR2_X1 U21905 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18919), .ZN(
        n18920) );
  AOI22_X1 U21906 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18927), .B1(
        n18934), .B2(n18920), .ZN(n18921) );
  OAI211_X1 U21907 ( .C1(n18924), .C2(n18923), .A(n18922), .B(n18921), .ZN(
        P3_U2856) );
  AOI22_X1 U21908 ( .A1(n13496), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18952), 
        .B2(n18925), .ZN(n18931) );
  AOI22_X1 U21909 ( .A1(n18927), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n18950), .B2(n18926), .ZN(n18930) );
  NAND4_X1 U21910 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n18934), .A4(n18928), .ZN(
        n18929) );
  NAND3_X1 U21911 ( .A1(n18931), .A2(n18930), .A3(n18929), .ZN(P3_U2857) );
  NAND2_X1 U21912 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18932), .ZN(
        n18943) );
  AOI21_X1 U21913 ( .B1(n18957), .B2(n18943), .A(n18955), .ZN(n18940) );
  AOI22_X1 U21914 ( .A1(n13496), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18952), 
        .B2(n18933), .ZN(n18938) );
  AND2_X1 U21915 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18934), .ZN(
        n18936) );
  AOI22_X1 U21916 ( .A1(n18936), .A2(n18939), .B1(n18950), .B2(n18935), .ZN(
        n18937) );
  OAI211_X1 U21917 ( .C1(n18940), .C2(n18939), .A(n18938), .B(n18937), .ZN(
        P3_U2858) );
  AOI22_X1 U21918 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18955), .B1(
        n18953), .B2(P3_REIP_REG_3__SCAN_IN), .ZN(n18948) );
  AOI22_X1 U21919 ( .A1(n18952), .A2(n18942), .B1(n18950), .B2(n18941), .ZN(
        n18947) );
  OAI211_X1 U21920 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18945), .A(
        n18944), .B(n18943), .ZN(n18946) );
  NAND3_X1 U21921 ( .A1(n18948), .A2(n18947), .A3(n18946), .ZN(P3_U2859) );
  AOI22_X1 U21922 ( .A1(n18952), .A2(n18951), .B1(n18950), .B2(n18949), .ZN(
        n18962) );
  NAND2_X1 U21923 ( .A1(n18953), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18961) );
  OAI21_X1 U21924 ( .B1(n18955), .B2(n18954), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18960) );
  OAI211_X1 U21925 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18958), .A(
        n18957), .B(n18956), .ZN(n18959) );
  NAND4_X1 U21926 ( .A1(n18962), .A2(n18961), .A3(n18960), .A4(n18959), .ZN(
        P3_U2861) );
  INV_X1 U21927 ( .A(n18963), .ZN(n18964) );
  OAI211_X1 U21928 ( .C1(n18964), .C2(P3_FLUSH_REG_SCAN_IN), .A(
        P3_STATE2_REG_1__SCAN_IN), .B(P3_STATE2_REG_2__SCAN_IN), .ZN(n19433)
         );
  OAI21_X1 U21929 ( .B1(n18967), .B2(n18965), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18966) );
  OAI221_X1 U21930 ( .B1(n18967), .B2(n19433), .C1(n18967), .C2(n19019), .A(
        n18966), .ZN(P3_U2863) );
  NAND2_X1 U21931 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19146) );
  AOI221_X1 U21932 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19146), .C1(n18969), 
        .C2(n19146), .A(n18968), .ZN(n18974) );
  NOR2_X1 U21933 ( .A1(n18970), .A2(n13074), .ZN(n18971) );
  OAI21_X1 U21934 ( .B1(n18971), .B2(n19309), .A(n18975), .ZN(n18972) );
  AOI22_X1 U21935 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18974), .B1(
        n18972), .B2(n13077), .ZN(P3_U2865) );
  INV_X1 U21936 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19394) );
  NAND2_X1 U21937 ( .A1(n13077), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19236) );
  INV_X1 U21938 ( .A(n19236), .ZN(n19258) );
  NOR2_X1 U21939 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13077), .ZN(
        n19148) );
  NOR2_X1 U21940 ( .A1(n19258), .A2(n19148), .ZN(n18973) );
  OAI22_X1 U21941 ( .A1(n18974), .A2(n19394), .B1(n18973), .B2(n18972), .ZN(
        P3_U2866) );
  NOR2_X1 U21942 ( .A1(n19395), .A2(n18975), .ZN(P3_U2867) );
  NOR2_X1 U21943 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19084) );
  NOR2_X1 U21944 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19064) );
  NAND2_X1 U21945 ( .A1(n19084), .A2(n19064), .ZN(n19041) );
  NOR2_X1 U21946 ( .A1(n18977), .A2(n18976), .ZN(n19009) );
  NAND2_X1 U21947 ( .A1(n18978), .A2(n19009), .ZN(n19340) );
  NOR2_X2 U21948 ( .A1(n19015), .A2(n16849), .ZN(n19337) );
  NAND2_X1 U21949 ( .A1(n19407), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19213) );
  INV_X1 U21950 ( .A(n19213), .ZN(n18979) );
  NOR2_X1 U21951 ( .A1(n13077), .A2(n19394), .ZN(n18980) );
  NAND2_X1 U21952 ( .A1(n18979), .A2(n18980), .ZN(n19330) );
  NOR2_X2 U21953 ( .A1(n19011), .A2(n13222), .ZN(n19332) );
  NOR2_X1 U21954 ( .A1(n19394), .A2(n19146), .ZN(n19333) );
  NAND2_X1 U21955 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19333), .ZN(
        n19384) );
  NAND2_X1 U21956 ( .A1(n19384), .A2(n19041), .ZN(n18981) );
  INV_X1 U21957 ( .A(n18981), .ZN(n19039) );
  NOR2_X1 U21958 ( .A1(n19385), .A2(n19039), .ZN(n19013) );
  AOI22_X1 U21959 ( .A1(n19337), .A2(n19035), .B1(n19332), .B2(n19013), .ZN(
        n18984) );
  NOR2_X1 U21960 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19407), .ZN(
        n19189) );
  NOR2_X1 U21961 ( .A1(n19189), .A2(n18979), .ZN(n19261) );
  INV_X1 U21962 ( .A(n18980), .ZN(n18982) );
  NOR2_X1 U21963 ( .A1(n19261), .A2(n18982), .ZN(n19310) );
  AOI21_X1 U21964 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n19011), .ZN(n19307) );
  AOI22_X1 U21965 ( .A1(n19336), .A2(n19310), .B1(n19307), .B2(n18981), .ZN(
        n19016) );
  AND2_X1 U21966 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19336), .ZN(n19331) );
  NOR2_X1 U21967 ( .A1(n18982), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19335) );
  NAND2_X1 U21968 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19335), .ZN(
        n19306) );
  INV_X1 U21969 ( .A(n19306), .ZN(n19379) );
  AOI22_X1 U21970 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19016), .B1(
        n19331), .B2(n19379), .ZN(n18983) );
  OAI211_X1 U21971 ( .C1(n19041), .C2(n19340), .A(n18984), .B(n18983), .ZN(
        P3_U2868) );
  NAND2_X1 U21972 ( .A1(n18985), .A2(n19009), .ZN(n19346) );
  NOR2_X2 U21973 ( .A1(n19011), .A2(n18986), .ZN(n19342) );
  AOI22_X1 U21974 ( .A1(n19342), .A2(n19013), .B1(n19341), .B2(n19379), .ZN(
        n18988) );
  AND2_X1 U21975 ( .A1(n19336), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19343) );
  AOI22_X1 U21976 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19016), .B1(
        n19343), .B2(n19035), .ZN(n18987) );
  OAI211_X1 U21977 ( .C1(n19041), .C2(n19346), .A(n18988), .B(n18987), .ZN(
        P3_U2869) );
  NAND2_X1 U21978 ( .A1(n18989), .A2(n19009), .ZN(n19352) );
  AND2_X1 U21979 ( .A1(n19336), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19348) );
  NOR2_X2 U21980 ( .A1(n19011), .A2(n21444), .ZN(n19347) );
  AOI22_X1 U21981 ( .A1(n19348), .A2(n19035), .B1(n19347), .B2(n19013), .ZN(
        n18991) );
  AND2_X1 U21982 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19336), .ZN(n19349) );
  AOI22_X1 U21983 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19016), .B1(
        n19349), .B2(n19379), .ZN(n18990) );
  OAI211_X1 U21984 ( .C1(n19041), .C2(n19352), .A(n18991), .B(n18990), .ZN(
        P3_U2870) );
  NAND2_X1 U21985 ( .A1(n18992), .A2(n19009), .ZN(n19358) );
  NOR2_X2 U21986 ( .A1(n19011), .A2(n18993), .ZN(n19354) );
  AND2_X1 U21987 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19336), .ZN(n19353) );
  AOI22_X1 U21988 ( .A1(n19354), .A2(n19013), .B1(n19353), .B2(n19379), .ZN(
        n18995) );
  AND2_X1 U21989 ( .A1(n19336), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19355) );
  AOI22_X1 U21990 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19016), .B1(
        n19355), .B2(n19035), .ZN(n18994) );
  OAI211_X1 U21991 ( .C1(n19041), .C2(n19358), .A(n18995), .B(n18994), .ZN(
        P3_U2871) );
  NAND2_X1 U21992 ( .A1(n18996), .A2(n19009), .ZN(n19364) );
  NOR2_X2 U21993 ( .A1(n19011), .A2(n18997), .ZN(n19360) );
  NOR2_X2 U21994 ( .A1(n19015), .A2(n18998), .ZN(n19359) );
  AOI22_X1 U21995 ( .A1(n19360), .A2(n19013), .B1(n19359), .B2(n19035), .ZN(
        n19000) );
  AND2_X1 U21996 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19336), .ZN(n19361) );
  AOI22_X1 U21997 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19016), .B1(
        n19361), .B2(n19379), .ZN(n18999) );
  OAI211_X1 U21998 ( .C1(n19041), .C2(n19364), .A(n19000), .B(n18999), .ZN(
        P3_U2872) );
  NAND2_X1 U21999 ( .A1(n19001), .A2(n19009), .ZN(n19370) );
  AND2_X1 U22000 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19336), .ZN(n19366) );
  NOR2_X2 U22001 ( .A1(n19011), .A2(n19002), .ZN(n19365) );
  AOI22_X1 U22002 ( .A1(n19366), .A2(n19379), .B1(n19365), .B2(n19013), .ZN(
        n19004) );
  AND2_X1 U22003 ( .A1(n19336), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19367) );
  AOI22_X1 U22004 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19016), .B1(
        n19367), .B2(n19035), .ZN(n19003) );
  OAI211_X1 U22005 ( .C1(n19041), .C2(n19370), .A(n19004), .B(n19003), .ZN(
        P3_U2873) );
  NAND2_X1 U22006 ( .A1(n19005), .A2(n19009), .ZN(n19376) );
  AND2_X1 U22007 ( .A1(n19336), .A2(BUF2_REG_22__SCAN_IN), .ZN(n19372) );
  NOR2_X2 U22008 ( .A1(n19011), .A2(n21479), .ZN(n19371) );
  AOI22_X1 U22009 ( .A1(n19372), .A2(n19035), .B1(n19371), .B2(n19013), .ZN(
        n19008) );
  NOR2_X2 U22010 ( .A1(n19006), .A2(n19015), .ZN(n19373) );
  AOI22_X1 U22011 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19016), .B1(
        n19373), .B2(n19379), .ZN(n19007) );
  OAI211_X1 U22012 ( .C1(n19041), .C2(n19376), .A(n19008), .B(n19007), .ZN(
        P3_U2874) );
  NAND2_X1 U22013 ( .A1(n19010), .A2(n19009), .ZN(n21549) );
  NAND2_X1 U22014 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19336), .ZN(n21551) );
  INV_X1 U22015 ( .A(n21551), .ZN(n19380) );
  NOR2_X2 U22016 ( .A1(n19012), .A2(n19011), .ZN(n21544) );
  AOI22_X1 U22017 ( .A1(n19380), .A2(n19035), .B1(n21544), .B2(n19013), .ZN(
        n19018) );
  NOR2_X2 U22018 ( .A1(n19015), .A2(n19014), .ZN(n21546) );
  AOI22_X1 U22019 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19016), .B1(
        n21546), .B2(n19379), .ZN(n19017) );
  OAI211_X1 U22020 ( .C1(n21549), .C2(n19041), .A(n19018), .B(n19017), .ZN(
        P3_U2875) );
  NAND2_X1 U22021 ( .A1(n19064), .A2(n19189), .ZN(n19063) );
  INV_X1 U22022 ( .A(n19064), .ZN(n19062) );
  NAND2_X1 U22023 ( .A1(n13074), .A2(n19438), .ZN(n19191) );
  NOR2_X1 U22024 ( .A1(n19062), .A2(n19191), .ZN(n19034) );
  AOI22_X1 U22025 ( .A1(n19332), .A2(n19034), .B1(n19331), .B2(n19035), .ZN(
        n19021) );
  NAND2_X1 U22026 ( .A1(n19263), .A2(n19019), .ZN(n19192) );
  NOR2_X1 U22027 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19192), .ZN(
        n19107) );
  AOI22_X1 U22028 ( .A1(n19336), .A2(n19333), .B1(n19107), .B2(n19064), .ZN(
        n19036) );
  AOI22_X1 U22029 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19036), .B1(
        n19057), .B2(n19337), .ZN(n19020) );
  OAI211_X1 U22030 ( .C1(n19063), .C2(n19340), .A(n19021), .B(n19020), .ZN(
        P3_U2876) );
  AOI22_X1 U22031 ( .A1(n19057), .A2(n19343), .B1(n19342), .B2(n19034), .ZN(
        n19023) );
  AOI22_X1 U22032 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19036), .B1(
        n19341), .B2(n19035), .ZN(n19022) );
  OAI211_X1 U22033 ( .C1(n19063), .C2(n19346), .A(n19023), .B(n19022), .ZN(
        P3_U2877) );
  AOI22_X1 U22034 ( .A1(n19057), .A2(n19348), .B1(n19347), .B2(n19034), .ZN(
        n19025) );
  AOI22_X1 U22035 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19036), .B1(
        n19349), .B2(n19035), .ZN(n19024) );
  OAI211_X1 U22036 ( .C1(n19063), .C2(n19352), .A(n19025), .B(n19024), .ZN(
        P3_U2878) );
  AOI22_X1 U22037 ( .A1(n19354), .A2(n19034), .B1(n19353), .B2(n19035), .ZN(
        n19027) );
  AOI22_X1 U22038 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19036), .B1(
        n19057), .B2(n19355), .ZN(n19026) );
  OAI211_X1 U22039 ( .C1(n19063), .C2(n19358), .A(n19027), .B(n19026), .ZN(
        P3_U2879) );
  AOI22_X1 U22040 ( .A1(n19057), .A2(n19359), .B1(n19360), .B2(n19034), .ZN(
        n19029) );
  AOI22_X1 U22041 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19036), .B1(
        n19361), .B2(n19035), .ZN(n19028) );
  OAI211_X1 U22042 ( .C1(n19063), .C2(n19364), .A(n19029), .B(n19028), .ZN(
        P3_U2880) );
  AOI22_X1 U22043 ( .A1(n19057), .A2(n19367), .B1(n19365), .B2(n19034), .ZN(
        n19031) );
  AOI22_X1 U22044 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19036), .B1(
        n19366), .B2(n19035), .ZN(n19030) );
  OAI211_X1 U22045 ( .C1(n19063), .C2(n19370), .A(n19031), .B(n19030), .ZN(
        P3_U2881) );
  AOI22_X1 U22046 ( .A1(n19057), .A2(n19372), .B1(n19371), .B2(n19034), .ZN(
        n19033) );
  AOI22_X1 U22047 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19036), .B1(
        n19373), .B2(n19035), .ZN(n19032) );
  OAI211_X1 U22048 ( .C1(n19063), .C2(n19376), .A(n19033), .B(n19032), .ZN(
        P3_U2882) );
  AOI22_X1 U22049 ( .A1(n19380), .A2(n19057), .B1(n21544), .B2(n19034), .ZN(
        n19038) );
  AOI22_X1 U22050 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19036), .B1(
        n21546), .B2(n19035), .ZN(n19037) );
  OAI211_X1 U22051 ( .C1(n21549), .C2(n19063), .A(n19038), .B(n19037), .ZN(
        P3_U2883) );
  NOR2_X2 U22052 ( .A1(n19062), .A2(n19213), .ZN(n21547) );
  INV_X1 U22053 ( .A(n21547), .ZN(n19061) );
  AOI21_X1 U22054 ( .B1(n19061), .B2(n19063), .A(n19385), .ZN(n19056) );
  AOI22_X1 U22055 ( .A1(n19057), .A2(n19331), .B1(n19332), .B2(n19056), .ZN(
        n19043) );
  AOI221_X1 U22056 ( .B1(n19039), .B2(n19063), .C1(n19085), .C2(n19063), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19040) );
  OAI21_X1 U22057 ( .B1(n21547), .B2(n19040), .A(n19263), .ZN(n19058) );
  INV_X1 U22058 ( .A(n19041), .ZN(n19080) );
  AOI22_X1 U22059 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19058), .B1(
        n19080), .B2(n19337), .ZN(n19042) );
  OAI211_X1 U22060 ( .C1(n19061), .C2(n19340), .A(n19043), .B(n19042), .ZN(
        P3_U2884) );
  AOI22_X1 U22061 ( .A1(n19057), .A2(n19341), .B1(n19056), .B2(n19342), .ZN(
        n19045) );
  AOI22_X1 U22062 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19058), .B1(
        n19080), .B2(n19343), .ZN(n19044) );
  OAI211_X1 U22063 ( .C1(n19061), .C2(n19346), .A(n19045), .B(n19044), .ZN(
        P3_U2885) );
  AOI22_X1 U22064 ( .A1(n19057), .A2(n19349), .B1(n19056), .B2(n19347), .ZN(
        n19047) );
  AOI22_X1 U22065 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19058), .B1(
        n19080), .B2(n19348), .ZN(n19046) );
  OAI211_X1 U22066 ( .C1(n19061), .C2(n19352), .A(n19047), .B(n19046), .ZN(
        P3_U2886) );
  AOI22_X1 U22067 ( .A1(n19057), .A2(n19353), .B1(n19056), .B2(n19354), .ZN(
        n19049) );
  AOI22_X1 U22068 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19058), .B1(
        n19080), .B2(n19355), .ZN(n19048) );
  OAI211_X1 U22069 ( .C1(n19061), .C2(n19358), .A(n19049), .B(n19048), .ZN(
        P3_U2887) );
  AOI22_X1 U22070 ( .A1(n19080), .A2(n19359), .B1(n19056), .B2(n19360), .ZN(
        n19051) );
  AOI22_X1 U22071 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19058), .B1(
        n19057), .B2(n19361), .ZN(n19050) );
  OAI211_X1 U22072 ( .C1(n19061), .C2(n19364), .A(n19051), .B(n19050), .ZN(
        P3_U2888) );
  AOI22_X1 U22073 ( .A1(n19080), .A2(n19367), .B1(n19056), .B2(n19365), .ZN(
        n19053) );
  AOI22_X1 U22074 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19058), .B1(
        n19057), .B2(n19366), .ZN(n19052) );
  OAI211_X1 U22075 ( .C1(n19061), .C2(n19370), .A(n19053), .B(n19052), .ZN(
        P3_U2889) );
  AOI22_X1 U22076 ( .A1(n19057), .A2(n19373), .B1(n19056), .B2(n19371), .ZN(
        n19055) );
  AOI22_X1 U22077 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19058), .B1(
        n19080), .B2(n19372), .ZN(n19054) );
  OAI211_X1 U22078 ( .C1(n19061), .C2(n19376), .A(n19055), .B(n19054), .ZN(
        P3_U2890) );
  AOI22_X1 U22079 ( .A1(n19380), .A2(n19080), .B1(n21544), .B2(n19056), .ZN(
        n19060) );
  AOI22_X1 U22080 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19058), .B1(
        n21546), .B2(n19057), .ZN(n19059) );
  OAI211_X1 U22081 ( .C1(n21549), .C2(n19061), .A(n19060), .B(n19059), .ZN(
        P3_U2891) );
  NOR2_X1 U22082 ( .A1(n13074), .A2(n19062), .ZN(n19108) );
  NAND2_X1 U22083 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19108), .ZN(
        n21552) );
  AND2_X1 U22084 ( .A1(n19438), .A2(n19108), .ZN(n19079) );
  AOI22_X1 U22085 ( .A1(n19103), .A2(n19337), .B1(n19332), .B2(n19079), .ZN(
        n19066) );
  AOI21_X1 U22086 ( .B1(n13074), .B2(n19085), .A(n19192), .ZN(n19147) );
  NAND2_X1 U22087 ( .A1(n19064), .A2(n19147), .ZN(n19081) );
  AOI22_X1 U22088 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19081), .B1(
        n19080), .B2(n19331), .ZN(n19065) );
  OAI211_X1 U22089 ( .C1(n21552), .C2(n19340), .A(n19066), .B(n19065), .ZN(
        P3_U2892) );
  AOI22_X1 U22090 ( .A1(n19080), .A2(n19341), .B1(n19342), .B2(n19079), .ZN(
        n19068) );
  AOI22_X1 U22091 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19081), .B1(
        n19103), .B2(n19343), .ZN(n19067) );
  OAI211_X1 U22092 ( .C1(n21552), .C2(n19346), .A(n19068), .B(n19067), .ZN(
        P3_U2893) );
  AOI22_X1 U22093 ( .A1(n19103), .A2(n19348), .B1(n19347), .B2(n19079), .ZN(
        n19070) );
  AOI22_X1 U22094 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19081), .B1(
        n19080), .B2(n19349), .ZN(n19069) );
  OAI211_X1 U22095 ( .C1(n21552), .C2(n19352), .A(n19070), .B(n19069), .ZN(
        P3_U2894) );
  AOI22_X1 U22096 ( .A1(n19080), .A2(n19353), .B1(n19354), .B2(n19079), .ZN(
        n19072) );
  AOI22_X1 U22097 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19081), .B1(
        n19103), .B2(n19355), .ZN(n19071) );
  OAI211_X1 U22098 ( .C1(n21552), .C2(n19358), .A(n19072), .B(n19071), .ZN(
        P3_U2895) );
  AOI22_X1 U22099 ( .A1(n19103), .A2(n19359), .B1(n19360), .B2(n19079), .ZN(
        n19074) );
  AOI22_X1 U22100 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19081), .B1(
        n19080), .B2(n19361), .ZN(n19073) );
  OAI211_X1 U22101 ( .C1(n21552), .C2(n19364), .A(n19074), .B(n19073), .ZN(
        P3_U2896) );
  AOI22_X1 U22102 ( .A1(n19103), .A2(n19367), .B1(n19365), .B2(n19079), .ZN(
        n19076) );
  AOI22_X1 U22103 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19081), .B1(
        n19080), .B2(n19366), .ZN(n19075) );
  OAI211_X1 U22104 ( .C1(n21552), .C2(n19370), .A(n19076), .B(n19075), .ZN(
        P3_U2897) );
  AOI22_X1 U22105 ( .A1(n19080), .A2(n19373), .B1(n19371), .B2(n19079), .ZN(
        n19078) );
  AOI22_X1 U22106 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19081), .B1(
        n19103), .B2(n19372), .ZN(n19077) );
  OAI211_X1 U22107 ( .C1(n21552), .C2(n19376), .A(n19078), .B(n19077), .ZN(
        P3_U2898) );
  AOI22_X1 U22108 ( .A1(n21546), .A2(n19080), .B1(n21544), .B2(n19079), .ZN(
        n19083) );
  AOI22_X1 U22109 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19081), .B1(
        n19380), .B2(n19103), .ZN(n19082) );
  OAI211_X1 U22110 ( .C1(n21552), .C2(n21549), .A(n19083), .B(n19082), .ZN(
        P3_U2899) );
  INV_X1 U22111 ( .A(n19084), .ZN(n19414) );
  INV_X1 U22112 ( .A(n19148), .ZN(n19123) );
  NOR2_X2 U22113 ( .A1(n19414), .A2(n19123), .ZN(n19164) );
  AOI21_X1 U22114 ( .B1(n21552), .B2(n19124), .A(n19385), .ZN(n19102) );
  AOI22_X1 U22115 ( .A1(n19103), .A2(n19331), .B1(n19332), .B2(n19102), .ZN(
        n19089) );
  NOR2_X1 U22116 ( .A1(n21547), .A2(n19103), .ZN(n19086) );
  AOI221_X1 U22117 ( .B1(n19086), .B2(n21552), .C1(n19085), .C2(n21552), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19087) );
  OAI21_X1 U22118 ( .B1(n19164), .B2(n19087), .A(n19263), .ZN(n19104) );
  AOI22_X1 U22119 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19104), .B1(
        n21547), .B2(n19337), .ZN(n19088) );
  OAI211_X1 U22120 ( .C1(n19340), .C2(n19124), .A(n19089), .B(n19088), .ZN(
        P3_U2900) );
  AOI22_X1 U22121 ( .A1(n21547), .A2(n19343), .B1(n19342), .B2(n19102), .ZN(
        n19091) );
  AOI22_X1 U22122 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19104), .B1(
        n19103), .B2(n19341), .ZN(n19090) );
  OAI211_X1 U22123 ( .C1(n19346), .C2(n19124), .A(n19091), .B(n19090), .ZN(
        P3_U2901) );
  AOI22_X1 U22124 ( .A1(n21547), .A2(n19348), .B1(n19347), .B2(n19102), .ZN(
        n19093) );
  AOI22_X1 U22125 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19104), .B1(
        n19103), .B2(n19349), .ZN(n19092) );
  OAI211_X1 U22126 ( .C1(n19352), .C2(n19124), .A(n19093), .B(n19092), .ZN(
        P3_U2902) );
  AOI22_X1 U22127 ( .A1(n19103), .A2(n19353), .B1(n19354), .B2(n19102), .ZN(
        n19095) );
  AOI22_X1 U22128 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19104), .B1(
        n21547), .B2(n19355), .ZN(n19094) );
  OAI211_X1 U22129 ( .C1(n19358), .C2(n19124), .A(n19095), .B(n19094), .ZN(
        P3_U2903) );
  AOI22_X1 U22130 ( .A1(n19103), .A2(n19361), .B1(n19360), .B2(n19102), .ZN(
        n19097) );
  AOI22_X1 U22131 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19104), .B1(
        n21547), .B2(n19359), .ZN(n19096) );
  OAI211_X1 U22132 ( .C1(n19364), .C2(n19124), .A(n19097), .B(n19096), .ZN(
        P3_U2904) );
  AOI22_X1 U22133 ( .A1(n19103), .A2(n19366), .B1(n19365), .B2(n19102), .ZN(
        n19099) );
  AOI22_X1 U22134 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19104), .B1(
        n21547), .B2(n19367), .ZN(n19098) );
  OAI211_X1 U22135 ( .C1(n19370), .C2(n19124), .A(n19099), .B(n19098), .ZN(
        P3_U2905) );
  AOI22_X1 U22136 ( .A1(n19103), .A2(n19373), .B1(n19371), .B2(n19102), .ZN(
        n19101) );
  AOI22_X1 U22137 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19104), .B1(
        n21547), .B2(n19372), .ZN(n19100) );
  OAI211_X1 U22138 ( .C1(n19376), .C2(n19124), .A(n19101), .B(n19100), .ZN(
        P3_U2906) );
  AOI22_X1 U22139 ( .A1(n19380), .A2(n21547), .B1(n21544), .B2(n19102), .ZN(
        n19106) );
  AOI22_X1 U22140 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19104), .B1(
        n21546), .B2(n19103), .ZN(n19105) );
  OAI211_X1 U22141 ( .C1(n21549), .C2(n19124), .A(n19106), .B(n19105), .ZN(
        P3_U2907) );
  NAND2_X1 U22142 ( .A1(n19148), .A2(n19189), .ZN(n21550) );
  NOR2_X1 U22143 ( .A1(n19123), .A2(n19191), .ZN(n21545) );
  AOI22_X1 U22144 ( .A1(n21547), .A2(n19331), .B1(n21545), .B2(n19332), .ZN(
        n19110) );
  AOI22_X1 U22145 ( .A1(n19336), .A2(n19108), .B1(n19107), .B2(n19148), .ZN(
        n21555) );
  AOI22_X1 U22146 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n21555), .B1(
        n19141), .B2(n19337), .ZN(n19109) );
  OAI211_X1 U22147 ( .C1(n21550), .C2(n19340), .A(n19110), .B(n19109), .ZN(
        P3_U2908) );
  AOI22_X1 U22148 ( .A1(n21547), .A2(n19341), .B1(n21545), .B2(n19342), .ZN(
        n19112) );
  AOI22_X1 U22149 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n21555), .B1(
        n19141), .B2(n19343), .ZN(n19111) );
  OAI211_X1 U22150 ( .C1(n21550), .C2(n19346), .A(n19112), .B(n19111), .ZN(
        P3_U2909) );
  AOI22_X1 U22151 ( .A1(n19141), .A2(n19348), .B1(n21545), .B2(n19347), .ZN(
        n19114) );
  AOI22_X1 U22152 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n21555), .B1(
        n21547), .B2(n19349), .ZN(n19113) );
  OAI211_X1 U22153 ( .C1(n21550), .C2(n19352), .A(n19114), .B(n19113), .ZN(
        P3_U2910) );
  AOI22_X1 U22154 ( .A1(n21547), .A2(n19353), .B1(n21545), .B2(n19354), .ZN(
        n19116) );
  AOI22_X1 U22155 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n21555), .B1(
        n19141), .B2(n19355), .ZN(n19115) );
  OAI211_X1 U22156 ( .C1(n21550), .C2(n19358), .A(n19116), .B(n19115), .ZN(
        P3_U2911) );
  AOI22_X1 U22157 ( .A1(n19141), .A2(n19359), .B1(n21545), .B2(n19360), .ZN(
        n19118) );
  AOI22_X1 U22158 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n21555), .B1(
        n21547), .B2(n19361), .ZN(n19117) );
  OAI211_X1 U22159 ( .C1(n21550), .C2(n19364), .A(n19118), .B(n19117), .ZN(
        P3_U2912) );
  AOI22_X1 U22160 ( .A1(n21547), .A2(n19366), .B1(n21545), .B2(n19365), .ZN(
        n19120) );
  AOI22_X1 U22161 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n21555), .B1(
        n19141), .B2(n19367), .ZN(n19119) );
  OAI211_X1 U22162 ( .C1(n21550), .C2(n19370), .A(n19120), .B(n19119), .ZN(
        P3_U2913) );
  AOI22_X1 U22163 ( .A1(n19141), .A2(n19372), .B1(n21545), .B2(n19371), .ZN(
        n19122) );
  AOI22_X1 U22164 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n21555), .B1(
        n21547), .B2(n19373), .ZN(n19121) );
  OAI211_X1 U22165 ( .C1(n21550), .C2(n19376), .A(n19122), .B(n19121), .ZN(
        P3_U2914) );
  NOR2_X2 U22166 ( .A1(n19123), .A2(n19213), .ZN(n19209) );
  NAND2_X1 U22167 ( .A1(n21550), .A2(n19145), .ZN(n19168) );
  AND2_X1 U22168 ( .A1(n19438), .A2(n19168), .ZN(n19140) );
  AOI22_X1 U22169 ( .A1(n19337), .A2(n19164), .B1(n19332), .B2(n19140), .ZN(
        n19127) );
  NAND2_X1 U22170 ( .A1(n21552), .A2(n19124), .ZN(n19125) );
  OAI221_X1 U22171 ( .B1(n19168), .B2(n19309), .C1(n19168), .C2(n19125), .A(
        n19307), .ZN(n19142) );
  AOI22_X1 U22172 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19142), .B1(
        n19141), .B2(n19331), .ZN(n19126) );
  OAI211_X1 U22173 ( .C1(n19340), .C2(n19145), .A(n19127), .B(n19126), .ZN(
        P3_U2916) );
  AOI22_X1 U22174 ( .A1(n19343), .A2(n19164), .B1(n19342), .B2(n19140), .ZN(
        n19129) );
  AOI22_X1 U22175 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19142), .B1(
        n19141), .B2(n19341), .ZN(n19128) );
  OAI211_X1 U22176 ( .C1(n19346), .C2(n19145), .A(n19129), .B(n19128), .ZN(
        P3_U2917) );
  AOI22_X1 U22177 ( .A1(n19348), .A2(n19164), .B1(n19347), .B2(n19140), .ZN(
        n19131) );
  AOI22_X1 U22178 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19142), .B1(
        n19141), .B2(n19349), .ZN(n19130) );
  OAI211_X1 U22179 ( .C1(n19352), .C2(n19145), .A(n19131), .B(n19130), .ZN(
        P3_U2918) );
  AOI22_X1 U22180 ( .A1(n19355), .A2(n19164), .B1(n19354), .B2(n19140), .ZN(
        n19133) );
  AOI22_X1 U22181 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19142), .B1(
        n19141), .B2(n19353), .ZN(n19132) );
  OAI211_X1 U22182 ( .C1(n19358), .C2(n19145), .A(n19133), .B(n19132), .ZN(
        P3_U2919) );
  AOI22_X1 U22183 ( .A1(n19141), .A2(n19361), .B1(n19360), .B2(n19140), .ZN(
        n19135) );
  AOI22_X1 U22184 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19142), .B1(
        n19359), .B2(n19164), .ZN(n19134) );
  OAI211_X1 U22185 ( .C1(n19364), .C2(n19145), .A(n19135), .B(n19134), .ZN(
        P3_U2920) );
  AOI22_X1 U22186 ( .A1(n19141), .A2(n19366), .B1(n19365), .B2(n19140), .ZN(
        n19137) );
  AOI22_X1 U22187 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19142), .B1(
        n19367), .B2(n19164), .ZN(n19136) );
  OAI211_X1 U22188 ( .C1(n19370), .C2(n19145), .A(n19137), .B(n19136), .ZN(
        P3_U2921) );
  AOI22_X1 U22189 ( .A1(n19141), .A2(n19373), .B1(n19371), .B2(n19140), .ZN(
        n19139) );
  AOI22_X1 U22190 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19142), .B1(
        n19372), .B2(n19164), .ZN(n19138) );
  OAI211_X1 U22191 ( .C1(n19376), .C2(n19145), .A(n19139), .B(n19138), .ZN(
        P3_U2922) );
  AOI22_X1 U22192 ( .A1(n19380), .A2(n19164), .B1(n21544), .B2(n19140), .ZN(
        n19144) );
  AOI22_X1 U22193 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19142), .B1(
        n19141), .B2(n21546), .ZN(n19143) );
  OAI211_X1 U22194 ( .C1(n21549), .C2(n19145), .A(n19144), .B(n19143), .ZN(
        P3_U2923) );
  NOR2_X1 U22195 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19146), .ZN(
        n19193) );
  NAND2_X1 U22196 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19193), .ZN(
        n19190) );
  AND2_X1 U22197 ( .A1(n19438), .A2(n19193), .ZN(n19163) );
  AOI22_X1 U22198 ( .A1(n19332), .A2(n19163), .B1(n19331), .B2(n19164), .ZN(
        n19150) );
  NAND2_X1 U22199 ( .A1(n19148), .A2(n19147), .ZN(n19165) );
  AOI22_X1 U22200 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19165), .B1(
        n19184), .B2(n19337), .ZN(n19149) );
  OAI211_X1 U22201 ( .C1(n19340), .C2(n19190), .A(n19150), .B(n19149), .ZN(
        P3_U2924) );
  AOI22_X1 U22202 ( .A1(n19342), .A2(n19163), .B1(n19341), .B2(n19164), .ZN(
        n19152) );
  AOI22_X1 U22203 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19165), .B1(
        n19184), .B2(n19343), .ZN(n19151) );
  OAI211_X1 U22204 ( .C1(n19346), .C2(n19190), .A(n19152), .B(n19151), .ZN(
        P3_U2925) );
  AOI22_X1 U22205 ( .A1(n19184), .A2(n19348), .B1(n19347), .B2(n19163), .ZN(
        n19154) );
  AOI22_X1 U22206 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19165), .B1(
        n19349), .B2(n19164), .ZN(n19153) );
  OAI211_X1 U22207 ( .C1(n19352), .C2(n19190), .A(n19154), .B(n19153), .ZN(
        P3_U2926) );
  AOI22_X1 U22208 ( .A1(n19354), .A2(n19163), .B1(n19353), .B2(n19164), .ZN(
        n19156) );
  AOI22_X1 U22209 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19165), .B1(
        n19184), .B2(n19355), .ZN(n19155) );
  OAI211_X1 U22210 ( .C1(n19358), .C2(n19190), .A(n19156), .B(n19155), .ZN(
        P3_U2927) );
  AOI22_X1 U22211 ( .A1(n19184), .A2(n19359), .B1(n19360), .B2(n19163), .ZN(
        n19158) );
  AOI22_X1 U22212 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19165), .B1(
        n19361), .B2(n19164), .ZN(n19157) );
  OAI211_X1 U22213 ( .C1(n19364), .C2(n19190), .A(n19158), .B(n19157), .ZN(
        P3_U2928) );
  AOI22_X1 U22214 ( .A1(n19366), .A2(n19164), .B1(n19365), .B2(n19163), .ZN(
        n19160) );
  AOI22_X1 U22215 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19165), .B1(
        n19184), .B2(n19367), .ZN(n19159) );
  OAI211_X1 U22216 ( .C1(n19370), .C2(n19190), .A(n19160), .B(n19159), .ZN(
        P3_U2929) );
  AOI22_X1 U22217 ( .A1(n19371), .A2(n19163), .B1(n19373), .B2(n19164), .ZN(
        n19162) );
  AOI22_X1 U22218 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19165), .B1(
        n19184), .B2(n19372), .ZN(n19161) );
  OAI211_X1 U22219 ( .C1(n19376), .C2(n19190), .A(n19162), .B(n19161), .ZN(
        P3_U2930) );
  AOI22_X1 U22220 ( .A1(n19380), .A2(n19184), .B1(n21544), .B2(n19163), .ZN(
        n19167) );
  AOI22_X1 U22221 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19165), .B1(
        n21546), .B2(n19164), .ZN(n19166) );
  OAI211_X1 U22222 ( .C1(n21549), .C2(n19190), .A(n19167), .B(n19166), .ZN(
        P3_U2931) );
  NOR2_X2 U22223 ( .A1(n19414), .A2(n19236), .ZN(n19254) );
  NAND2_X1 U22224 ( .A1(n19190), .A2(n19188), .ZN(n19214) );
  AND2_X1 U22225 ( .A1(n19438), .A2(n19214), .ZN(n19183) );
  AOI22_X1 U22226 ( .A1(n19337), .A2(n19209), .B1(n19332), .B2(n19183), .ZN(
        n19170) );
  OAI221_X1 U22227 ( .B1(n19214), .B2(n19309), .C1(n19214), .C2(n19168), .A(
        n19307), .ZN(n19185) );
  AOI22_X1 U22228 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19185), .B1(
        n19184), .B2(n19331), .ZN(n19169) );
  OAI211_X1 U22229 ( .C1(n19340), .C2(n19188), .A(n19170), .B(n19169), .ZN(
        P3_U2932) );
  AOI22_X1 U22230 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19185), .B1(
        n19342), .B2(n19183), .ZN(n19172) );
  AOI22_X1 U22231 ( .A1(n19184), .A2(n19341), .B1(n19343), .B2(n19209), .ZN(
        n19171) );
  OAI211_X1 U22232 ( .C1(n19346), .C2(n19188), .A(n19172), .B(n19171), .ZN(
        P3_U2933) );
  AOI22_X1 U22233 ( .A1(n19348), .A2(n19209), .B1(n19347), .B2(n19183), .ZN(
        n19174) );
  AOI22_X1 U22234 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19185), .B1(
        n19184), .B2(n19349), .ZN(n19173) );
  OAI211_X1 U22235 ( .C1(n19352), .C2(n19188), .A(n19174), .B(n19173), .ZN(
        P3_U2934) );
  AOI22_X1 U22236 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19185), .B1(
        n19354), .B2(n19183), .ZN(n19176) );
  AOI22_X1 U22237 ( .A1(n19184), .A2(n19353), .B1(n19355), .B2(n19209), .ZN(
        n19175) );
  OAI211_X1 U22238 ( .C1(n19358), .C2(n19188), .A(n19176), .B(n19175), .ZN(
        P3_U2935) );
  AOI22_X1 U22239 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19185), .B1(
        n19360), .B2(n19183), .ZN(n19178) );
  AOI22_X1 U22240 ( .A1(n19184), .A2(n19361), .B1(n19359), .B2(n19209), .ZN(
        n19177) );
  OAI211_X1 U22241 ( .C1(n19364), .C2(n19188), .A(n19178), .B(n19177), .ZN(
        P3_U2936) );
  AOI22_X1 U22242 ( .A1(n19365), .A2(n19183), .B1(n19367), .B2(n19209), .ZN(
        n19180) );
  AOI22_X1 U22243 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19185), .B1(
        n19184), .B2(n19366), .ZN(n19179) );
  OAI211_X1 U22244 ( .C1(n19370), .C2(n19188), .A(n19180), .B(n19179), .ZN(
        P3_U2937) );
  AOI22_X1 U22245 ( .A1(n19372), .A2(n19209), .B1(n19371), .B2(n19183), .ZN(
        n19182) );
  AOI22_X1 U22246 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19185), .B1(
        n19184), .B2(n19373), .ZN(n19181) );
  OAI211_X1 U22247 ( .C1(n19376), .C2(n19188), .A(n19182), .B(n19181), .ZN(
        P3_U2938) );
  AOI22_X1 U22248 ( .A1(n19380), .A2(n19209), .B1(n21544), .B2(n19183), .ZN(
        n19187) );
  AOI22_X1 U22249 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19185), .B1(
        n19184), .B2(n21546), .ZN(n19186) );
  OAI211_X1 U22250 ( .C1(n21549), .C2(n19188), .A(n19187), .B(n19186), .ZN(
        P3_U2939) );
  NAND2_X1 U22251 ( .A1(n19189), .A2(n19258), .ZN(n19238) );
  NOR2_X1 U22252 ( .A1(n19191), .A2(n19236), .ZN(n19208) );
  AOI22_X1 U22253 ( .A1(n19337), .A2(n19231), .B1(n19332), .B2(n19208), .ZN(
        n19195) );
  INV_X1 U22254 ( .A(n19192), .ZN(n19334) );
  NOR2_X1 U22255 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19236), .ZN(
        n19237) );
  AOI22_X1 U22256 ( .A1(n19336), .A2(n19193), .B1(n19334), .B2(n19237), .ZN(
        n19210) );
  AOI22_X1 U22257 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19210), .B1(
        n19331), .B2(n19209), .ZN(n19194) );
  OAI211_X1 U22258 ( .C1(n19340), .C2(n19238), .A(n19195), .B(n19194), .ZN(
        P3_U2940) );
  AOI22_X1 U22259 ( .A1(n19342), .A2(n19208), .B1(n19341), .B2(n19209), .ZN(
        n19197) );
  AOI22_X1 U22260 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19210), .B1(
        n19343), .B2(n19231), .ZN(n19196) );
  OAI211_X1 U22261 ( .C1(n19346), .C2(n19238), .A(n19197), .B(n19196), .ZN(
        P3_U2941) );
  AOI22_X1 U22262 ( .A1(n19348), .A2(n19231), .B1(n19347), .B2(n19208), .ZN(
        n19199) );
  AOI22_X1 U22263 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19210), .B1(
        n19349), .B2(n19209), .ZN(n19198) );
  OAI211_X1 U22264 ( .C1(n19352), .C2(n19238), .A(n19199), .B(n19198), .ZN(
        P3_U2942) );
  AOI22_X1 U22265 ( .A1(n19355), .A2(n19231), .B1(n19354), .B2(n19208), .ZN(
        n19201) );
  AOI22_X1 U22266 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19210), .B1(
        n19353), .B2(n19209), .ZN(n19200) );
  OAI211_X1 U22267 ( .C1(n19358), .C2(n19238), .A(n19201), .B(n19200), .ZN(
        P3_U2943) );
  AOI22_X1 U22268 ( .A1(n19361), .A2(n19209), .B1(n19360), .B2(n19208), .ZN(
        n19203) );
  AOI22_X1 U22269 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19210), .B1(
        n19359), .B2(n19231), .ZN(n19202) );
  OAI211_X1 U22270 ( .C1(n19364), .C2(n19238), .A(n19203), .B(n19202), .ZN(
        P3_U2944) );
  AOI22_X1 U22271 ( .A1(n19365), .A2(n19208), .B1(n19367), .B2(n19231), .ZN(
        n19205) );
  AOI22_X1 U22272 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19210), .B1(
        n19366), .B2(n19209), .ZN(n19204) );
  OAI211_X1 U22273 ( .C1(n19370), .C2(n19238), .A(n19205), .B(n19204), .ZN(
        P3_U2945) );
  AOI22_X1 U22274 ( .A1(n19371), .A2(n19208), .B1(n19373), .B2(n19209), .ZN(
        n19207) );
  AOI22_X1 U22275 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19210), .B1(
        n19372), .B2(n19231), .ZN(n19206) );
  OAI211_X1 U22276 ( .C1(n19376), .C2(n19238), .A(n19207), .B(n19206), .ZN(
        P3_U2946) );
  AOI22_X1 U22277 ( .A1(n21546), .A2(n19209), .B1(n21544), .B2(n19208), .ZN(
        n19212) );
  AOI22_X1 U22278 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19210), .B1(
        n19380), .B2(n19231), .ZN(n19211) );
  OAI211_X1 U22279 ( .C1(n21549), .C2(n19238), .A(n19212), .B(n19211), .ZN(
        P3_U2947) );
  NOR2_X2 U22280 ( .A1(n19213), .A2(n19236), .ZN(n19302) );
  AOI21_X1 U22281 ( .B1(n19238), .B2(n19235), .A(n19385), .ZN(n19230) );
  AOI22_X1 U22282 ( .A1(n19332), .A2(n19230), .B1(n19331), .B2(n19231), .ZN(
        n19217) );
  NAND2_X1 U22283 ( .A1(n19238), .A2(n19235), .ZN(n19215) );
  OAI221_X1 U22284 ( .B1(n19215), .B2(n19309), .C1(n19215), .C2(n19214), .A(
        n19307), .ZN(n19232) );
  AOI22_X1 U22285 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19232), .B1(
        n19337), .B2(n19254), .ZN(n19216) );
  OAI211_X1 U22286 ( .C1(n19340), .C2(n19235), .A(n19217), .B(n19216), .ZN(
        P3_U2948) );
  AOI22_X1 U22287 ( .A1(n19342), .A2(n19230), .B1(n19341), .B2(n19231), .ZN(
        n19219) );
  AOI22_X1 U22288 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19232), .B1(
        n19343), .B2(n19254), .ZN(n19218) );
  OAI211_X1 U22289 ( .C1(n19346), .C2(n19235), .A(n19219), .B(n19218), .ZN(
        P3_U2949) );
  AOI22_X1 U22290 ( .A1(n19349), .A2(n19231), .B1(n19347), .B2(n19230), .ZN(
        n19221) );
  AOI22_X1 U22291 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19232), .B1(
        n19348), .B2(n19254), .ZN(n19220) );
  OAI211_X1 U22292 ( .C1(n19352), .C2(n19235), .A(n19221), .B(n19220), .ZN(
        P3_U2950) );
  AOI22_X1 U22293 ( .A1(n19354), .A2(n19230), .B1(n19353), .B2(n19231), .ZN(
        n19223) );
  AOI22_X1 U22294 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19232), .B1(
        n19355), .B2(n19254), .ZN(n19222) );
  OAI211_X1 U22295 ( .C1(n19358), .C2(n19235), .A(n19223), .B(n19222), .ZN(
        P3_U2951) );
  AOI22_X1 U22296 ( .A1(n19360), .A2(n19230), .B1(n19359), .B2(n19254), .ZN(
        n19225) );
  AOI22_X1 U22297 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19232), .B1(
        n19361), .B2(n19231), .ZN(n19224) );
  OAI211_X1 U22298 ( .C1(n19364), .C2(n19235), .A(n19225), .B(n19224), .ZN(
        P3_U2952) );
  AOI22_X1 U22299 ( .A1(n19365), .A2(n19230), .B1(n19367), .B2(n19254), .ZN(
        n19227) );
  AOI22_X1 U22300 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19232), .B1(
        n19366), .B2(n19231), .ZN(n19226) );
  OAI211_X1 U22301 ( .C1(n19370), .C2(n19235), .A(n19227), .B(n19226), .ZN(
        P3_U2953) );
  AOI22_X1 U22302 ( .A1(n19372), .A2(n19254), .B1(n19371), .B2(n19230), .ZN(
        n19229) );
  AOI22_X1 U22303 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19232), .B1(
        n19373), .B2(n19231), .ZN(n19228) );
  OAI211_X1 U22304 ( .C1(n19376), .C2(n19235), .A(n19229), .B(n19228), .ZN(
        P3_U2954) );
  AOI22_X1 U22305 ( .A1(n19380), .A2(n19254), .B1(n21544), .B2(n19230), .ZN(
        n19234) );
  AOI22_X1 U22306 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19232), .B1(
        n21546), .B2(n19231), .ZN(n19233) );
  OAI211_X1 U22307 ( .C1(n21549), .C2(n19235), .A(n19234), .B(n19233), .ZN(
        P3_U2955) );
  NOR2_X1 U22308 ( .A1(n13074), .A2(n19236), .ZN(n19286) );
  NAND2_X1 U22309 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19286), .ZN(
        n19284) );
  AND2_X1 U22310 ( .A1(n19438), .A2(n19286), .ZN(n19253) );
  AOI22_X1 U22311 ( .A1(n19332), .A2(n19253), .B1(n19331), .B2(n19254), .ZN(
        n19240) );
  AOI22_X1 U22312 ( .A1(n19336), .A2(n19237), .B1(n19334), .B2(n19286), .ZN(
        n19255) );
  AOI22_X1 U22313 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19255), .B1(
        n19337), .B2(n19279), .ZN(n19239) );
  OAI211_X1 U22314 ( .C1(n19340), .C2(n19284), .A(n19240), .B(n19239), .ZN(
        P3_U2956) );
  AOI22_X1 U22315 ( .A1(n19342), .A2(n19253), .B1(n19341), .B2(n19254), .ZN(
        n19242) );
  AOI22_X1 U22316 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19255), .B1(
        n19343), .B2(n19279), .ZN(n19241) );
  OAI211_X1 U22317 ( .C1(n19346), .C2(n19284), .A(n19242), .B(n19241), .ZN(
        P3_U2957) );
  AOI22_X1 U22318 ( .A1(n19348), .A2(n19279), .B1(n19347), .B2(n19253), .ZN(
        n19244) );
  AOI22_X1 U22319 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19255), .B1(
        n19349), .B2(n19254), .ZN(n19243) );
  OAI211_X1 U22320 ( .C1(n19352), .C2(n19284), .A(n19244), .B(n19243), .ZN(
        P3_U2958) );
  AOI22_X1 U22321 ( .A1(n19354), .A2(n19253), .B1(n19353), .B2(n19254), .ZN(
        n19246) );
  AOI22_X1 U22322 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19255), .B1(
        n19355), .B2(n19279), .ZN(n19245) );
  OAI211_X1 U22323 ( .C1(n19358), .C2(n19284), .A(n19246), .B(n19245), .ZN(
        P3_U2959) );
  AOI22_X1 U22324 ( .A1(n19361), .A2(n19254), .B1(n19360), .B2(n19253), .ZN(
        n19248) );
  AOI22_X1 U22325 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19255), .B1(
        n19359), .B2(n19279), .ZN(n19247) );
  OAI211_X1 U22326 ( .C1(n19364), .C2(n19284), .A(n19248), .B(n19247), .ZN(
        P3_U2960) );
  AOI22_X1 U22327 ( .A1(n19365), .A2(n19253), .B1(n19367), .B2(n19279), .ZN(
        n19250) );
  AOI22_X1 U22328 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19255), .B1(
        n19366), .B2(n19254), .ZN(n19249) );
  OAI211_X1 U22329 ( .C1(n19370), .C2(n19284), .A(n19250), .B(n19249), .ZN(
        P3_U2961) );
  AOI22_X1 U22330 ( .A1(n19371), .A2(n19253), .B1(n19373), .B2(n19254), .ZN(
        n19252) );
  AOI22_X1 U22331 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19255), .B1(
        n19372), .B2(n19279), .ZN(n19251) );
  OAI211_X1 U22332 ( .C1(n19376), .C2(n19284), .A(n19252), .B(n19251), .ZN(
        P3_U2962) );
  AOI22_X1 U22333 ( .A1(n19380), .A2(n19279), .B1(n21544), .B2(n19253), .ZN(
        n19257) );
  AOI22_X1 U22334 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19255), .B1(
        n21546), .B2(n19254), .ZN(n19256) );
  OAI211_X1 U22335 ( .C1(n21549), .C2(n19284), .A(n19257), .B(n19256), .ZN(
        P3_U2963) );
  INV_X1 U22336 ( .A(n19335), .ZN(n19285) );
  NOR2_X2 U22337 ( .A1(n19285), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19378) );
  NAND2_X1 U22338 ( .A1(n19284), .A2(n19283), .ZN(n19308) );
  INV_X1 U22339 ( .A(n19308), .ZN(n19259) );
  NOR2_X1 U22340 ( .A1(n19385), .A2(n19259), .ZN(n19278) );
  AOI22_X1 U22341 ( .A1(n19337), .A2(n19302), .B1(n19332), .B2(n19278), .ZN(
        n19265) );
  NAND2_X1 U22342 ( .A1(n19309), .A2(n19258), .ZN(n19260) );
  OAI21_X1 U22343 ( .B1(n19261), .B2(n19260), .A(n19259), .ZN(n19262) );
  OAI211_X1 U22344 ( .C1(n19378), .C2(n19539), .A(n19263), .B(n19262), .ZN(
        n19280) );
  AOI22_X1 U22345 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19280), .B1(
        n19331), .B2(n19279), .ZN(n19264) );
  OAI211_X1 U22346 ( .C1(n19340), .C2(n19283), .A(n19265), .B(n19264), .ZN(
        P3_U2964) );
  AOI22_X1 U22347 ( .A1(n19342), .A2(n19278), .B1(n19341), .B2(n19279), .ZN(
        n19267) );
  AOI22_X1 U22348 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19280), .B1(
        n19343), .B2(n19302), .ZN(n19266) );
  OAI211_X1 U22349 ( .C1(n19346), .C2(n19283), .A(n19267), .B(n19266), .ZN(
        P3_U2965) );
  AOI22_X1 U22350 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19280), .B1(
        n19347), .B2(n19278), .ZN(n19269) );
  AOI22_X1 U22351 ( .A1(n19348), .A2(n19302), .B1(n19349), .B2(n19279), .ZN(
        n19268) );
  OAI211_X1 U22352 ( .C1(n19352), .C2(n19283), .A(n19269), .B(n19268), .ZN(
        P3_U2966) );
  AOI22_X1 U22353 ( .A1(n19355), .A2(n19302), .B1(n19354), .B2(n19278), .ZN(
        n19271) );
  AOI22_X1 U22354 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19280), .B1(
        n19353), .B2(n19279), .ZN(n19270) );
  OAI211_X1 U22355 ( .C1(n19358), .C2(n19283), .A(n19271), .B(n19270), .ZN(
        P3_U2967) );
  AOI22_X1 U22356 ( .A1(n19360), .A2(n19278), .B1(n19359), .B2(n19302), .ZN(
        n19273) );
  AOI22_X1 U22357 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19280), .B1(
        n19361), .B2(n19279), .ZN(n19272) );
  OAI211_X1 U22358 ( .C1(n19364), .C2(n19283), .A(n19273), .B(n19272), .ZN(
        P3_U2968) );
  AOI22_X1 U22359 ( .A1(n19365), .A2(n19278), .B1(n19367), .B2(n19302), .ZN(
        n19275) );
  AOI22_X1 U22360 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19280), .B1(
        n19366), .B2(n19279), .ZN(n19274) );
  OAI211_X1 U22361 ( .C1(n19370), .C2(n19283), .A(n19275), .B(n19274), .ZN(
        P3_U2969) );
  AOI22_X1 U22362 ( .A1(n19372), .A2(n19302), .B1(n19371), .B2(n19278), .ZN(
        n19277) );
  AOI22_X1 U22363 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19280), .B1(
        n19373), .B2(n19279), .ZN(n19276) );
  OAI211_X1 U22364 ( .C1(n19376), .C2(n19283), .A(n19277), .B(n19276), .ZN(
        P3_U2970) );
  AOI22_X1 U22365 ( .A1(n21546), .A2(n19279), .B1(n21544), .B2(n19278), .ZN(
        n19282) );
  AOI22_X1 U22366 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19280), .B1(
        n19380), .B2(n19302), .ZN(n19281) );
  OAI211_X1 U22367 ( .C1(n21549), .C2(n19283), .A(n19282), .B(n19281), .ZN(
        P3_U2971) );
  NOR2_X1 U22368 ( .A1(n19385), .A2(n19285), .ZN(n19301) );
  AOI22_X1 U22369 ( .A1(n19337), .A2(n19326), .B1(n19332), .B2(n19301), .ZN(
        n19288) );
  AOI22_X1 U22370 ( .A1(n19336), .A2(n19286), .B1(n19334), .B2(n19335), .ZN(
        n19303) );
  AOI22_X1 U22371 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19303), .B1(
        n19331), .B2(n19302), .ZN(n19287) );
  OAI211_X1 U22372 ( .C1(n19340), .C2(n19306), .A(n19288), .B(n19287), .ZN(
        P3_U2972) );
  AOI22_X1 U22373 ( .A1(n19343), .A2(n19326), .B1(n19342), .B2(n19301), .ZN(
        n19290) );
  AOI22_X1 U22374 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19303), .B1(
        n19341), .B2(n19302), .ZN(n19289) );
  OAI211_X1 U22375 ( .C1(n19346), .C2(n19306), .A(n19290), .B(n19289), .ZN(
        P3_U2973) );
  AOI22_X1 U22376 ( .A1(n19349), .A2(n19302), .B1(n19347), .B2(n19301), .ZN(
        n19292) );
  AOI22_X1 U22377 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19303), .B1(
        n19348), .B2(n19326), .ZN(n19291) );
  OAI211_X1 U22378 ( .C1(n19352), .C2(n19306), .A(n19292), .B(n19291), .ZN(
        P3_U2974) );
  AOI22_X1 U22379 ( .A1(n19354), .A2(n19301), .B1(n19353), .B2(n19302), .ZN(
        n19294) );
  AOI22_X1 U22380 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19303), .B1(
        n19355), .B2(n19326), .ZN(n19293) );
  OAI211_X1 U22381 ( .C1(n19358), .C2(n19306), .A(n19294), .B(n19293), .ZN(
        P3_U2975) );
  AOI22_X1 U22382 ( .A1(n19360), .A2(n19301), .B1(n19359), .B2(n19326), .ZN(
        n19296) );
  AOI22_X1 U22383 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19303), .B1(
        n19361), .B2(n19302), .ZN(n19295) );
  OAI211_X1 U22384 ( .C1(n19364), .C2(n19306), .A(n19296), .B(n19295), .ZN(
        P3_U2976) );
  AOI22_X1 U22385 ( .A1(n19365), .A2(n19301), .B1(n19367), .B2(n19326), .ZN(
        n19298) );
  AOI22_X1 U22386 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19303), .B1(
        n19366), .B2(n19302), .ZN(n19297) );
  OAI211_X1 U22387 ( .C1(n19370), .C2(n19306), .A(n19298), .B(n19297), .ZN(
        P3_U2977) );
  AOI22_X1 U22388 ( .A1(n19372), .A2(n19326), .B1(n19371), .B2(n19301), .ZN(
        n19300) );
  AOI22_X1 U22389 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19303), .B1(
        n19373), .B2(n19302), .ZN(n19299) );
  OAI211_X1 U22390 ( .C1(n19376), .C2(n19306), .A(n19300), .B(n19299), .ZN(
        P3_U2978) );
  AOI22_X1 U22391 ( .A1(n19380), .A2(n19326), .B1(n21544), .B2(n19301), .ZN(
        n19305) );
  AOI22_X1 U22392 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19303), .B1(
        n21546), .B2(n19302), .ZN(n19304) );
  OAI211_X1 U22393 ( .C1(n21549), .C2(n19306), .A(n19305), .B(n19304), .ZN(
        P3_U2979) );
  AND2_X1 U22394 ( .A1(n19438), .A2(n19310), .ZN(n19325) );
  AOI22_X1 U22395 ( .A1(n19332), .A2(n19325), .B1(n19331), .B2(n19326), .ZN(
        n19312) );
  OAI221_X1 U22396 ( .B1(n19310), .B2(n19309), .C1(n19310), .C2(n19308), .A(
        n19307), .ZN(n19327) );
  AOI22_X1 U22397 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19327), .B1(
        n19337), .B2(n19378), .ZN(n19311) );
  OAI211_X1 U22398 ( .C1(n19340), .C2(n19330), .A(n19312), .B(n19311), .ZN(
        P3_U2980) );
  AOI22_X1 U22399 ( .A1(n19343), .A2(n19378), .B1(n19342), .B2(n19325), .ZN(
        n19314) );
  AOI22_X1 U22400 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19327), .B1(
        n19341), .B2(n19326), .ZN(n19313) );
  OAI211_X1 U22401 ( .C1(n19346), .C2(n19330), .A(n19314), .B(n19313), .ZN(
        P3_U2981) );
  AOI22_X1 U22402 ( .A1(n19349), .A2(n19326), .B1(n19347), .B2(n19325), .ZN(
        n19316) );
  AOI22_X1 U22403 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19327), .B1(
        n19348), .B2(n19378), .ZN(n19315) );
  OAI211_X1 U22404 ( .C1(n19352), .C2(n19330), .A(n19316), .B(n19315), .ZN(
        P3_U2982) );
  AOI22_X1 U22405 ( .A1(n19355), .A2(n19378), .B1(n19354), .B2(n19325), .ZN(
        n19318) );
  AOI22_X1 U22406 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19327), .B1(
        n19353), .B2(n19326), .ZN(n19317) );
  OAI211_X1 U22407 ( .C1(n19358), .C2(n19330), .A(n19318), .B(n19317), .ZN(
        P3_U2983) );
  AOI22_X1 U22408 ( .A1(n19360), .A2(n19325), .B1(n19359), .B2(n19378), .ZN(
        n19320) );
  AOI22_X1 U22409 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19327), .B1(
        n19361), .B2(n19326), .ZN(n19319) );
  OAI211_X1 U22410 ( .C1(n19364), .C2(n19330), .A(n19320), .B(n19319), .ZN(
        P3_U2984) );
  AOI22_X1 U22411 ( .A1(n19365), .A2(n19325), .B1(n19367), .B2(n19378), .ZN(
        n19322) );
  AOI22_X1 U22412 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19327), .B1(
        n19366), .B2(n19326), .ZN(n19321) );
  OAI211_X1 U22413 ( .C1(n19370), .C2(n19330), .A(n19322), .B(n19321), .ZN(
        P3_U2985) );
  AOI22_X1 U22414 ( .A1(n19371), .A2(n19325), .B1(n19373), .B2(n19326), .ZN(
        n19324) );
  AOI22_X1 U22415 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19327), .B1(
        n19372), .B2(n19378), .ZN(n19323) );
  OAI211_X1 U22416 ( .C1(n19376), .C2(n19330), .A(n19324), .B(n19323), .ZN(
        P3_U2986) );
  AOI22_X1 U22417 ( .A1(n19380), .A2(n19378), .B1(n21544), .B2(n19325), .ZN(
        n19329) );
  AOI22_X1 U22418 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19327), .B1(
        n21546), .B2(n19326), .ZN(n19328) );
  OAI211_X1 U22419 ( .C1(n21549), .C2(n19330), .A(n19329), .B(n19328), .ZN(
        P3_U2987) );
  AND2_X1 U22420 ( .A1(n19438), .A2(n19333), .ZN(n19377) );
  AOI22_X1 U22421 ( .A1(n19332), .A2(n19377), .B1(n19331), .B2(n19378), .ZN(
        n19339) );
  AOI22_X1 U22422 ( .A1(n19336), .A2(n19335), .B1(n19334), .B2(n19333), .ZN(
        n19381) );
  AOI22_X1 U22423 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19381), .B1(
        n19337), .B2(n19379), .ZN(n19338) );
  OAI211_X1 U22424 ( .C1(n19384), .C2(n19340), .A(n19339), .B(n19338), .ZN(
        P3_U2988) );
  AOI22_X1 U22425 ( .A1(n19342), .A2(n19377), .B1(n19341), .B2(n19378), .ZN(
        n19345) );
  AOI22_X1 U22426 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19381), .B1(
        n19343), .B2(n19379), .ZN(n19344) );
  OAI211_X1 U22427 ( .C1(n19384), .C2(n19346), .A(n19345), .B(n19344), .ZN(
        P3_U2989) );
  AOI22_X1 U22428 ( .A1(n19348), .A2(n19379), .B1(n19347), .B2(n19377), .ZN(
        n19351) );
  AOI22_X1 U22429 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19381), .B1(
        n19349), .B2(n19378), .ZN(n19350) );
  OAI211_X1 U22430 ( .C1(n19384), .C2(n19352), .A(n19351), .B(n19350), .ZN(
        P3_U2990) );
  AOI22_X1 U22431 ( .A1(n19354), .A2(n19377), .B1(n19353), .B2(n19378), .ZN(
        n19357) );
  AOI22_X1 U22432 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19381), .B1(
        n19355), .B2(n19379), .ZN(n19356) );
  OAI211_X1 U22433 ( .C1(n19384), .C2(n19358), .A(n19357), .B(n19356), .ZN(
        P3_U2991) );
  AOI22_X1 U22434 ( .A1(n19360), .A2(n19377), .B1(n19359), .B2(n19379), .ZN(
        n19363) );
  AOI22_X1 U22435 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19381), .B1(
        n19361), .B2(n19378), .ZN(n19362) );
  OAI211_X1 U22436 ( .C1(n19384), .C2(n19364), .A(n19363), .B(n19362), .ZN(
        P3_U2992) );
  AOI22_X1 U22437 ( .A1(n19366), .A2(n19378), .B1(n19365), .B2(n19377), .ZN(
        n19369) );
  AOI22_X1 U22438 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19381), .B1(
        n19367), .B2(n19379), .ZN(n19368) );
  OAI211_X1 U22439 ( .C1(n19384), .C2(n19370), .A(n19369), .B(n19368), .ZN(
        P3_U2993) );
  AOI22_X1 U22440 ( .A1(n19372), .A2(n19379), .B1(n19371), .B2(n19377), .ZN(
        n19375) );
  AOI22_X1 U22441 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19381), .B1(
        n19373), .B2(n19378), .ZN(n19374) );
  OAI211_X1 U22442 ( .C1(n19384), .C2(n19376), .A(n19375), .B(n19374), .ZN(
        P3_U2994) );
  AOI22_X1 U22443 ( .A1(n21546), .A2(n19378), .B1(n21544), .B2(n19377), .ZN(
        n19383) );
  AOI22_X1 U22444 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19381), .B1(
        n19380), .B2(n19379), .ZN(n19382) );
  OAI211_X1 U22445 ( .C1(n21549), .C2(n19384), .A(n19383), .B(n19382), .ZN(
        P3_U2995) );
  NAND2_X1 U22446 ( .A1(n19385), .A2(n19444), .ZN(n19387) );
  OAI22_X1 U22447 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19387), .B1(
        n19562), .B2(n19386), .ZN(n19437) );
  AND2_X1 U22448 ( .A1(n19388), .A2(n9649), .ZN(n19432) );
  INV_X1 U22449 ( .A(n19389), .ZN(n19431) );
  INV_X1 U22450 ( .A(n19426), .ZN(n19412) );
  NAND2_X1 U22451 ( .A1(n19412), .A2(n19390), .ZN(n19393) );
  NAND2_X1 U22452 ( .A1(n19426), .A2(n19391), .ZN(n19392) );
  NAND2_X1 U22453 ( .A1(n19393), .A2(n19392), .ZN(n19416) );
  INV_X1 U22454 ( .A(n19416), .ZN(n19418) );
  AOI21_X1 U22455 ( .B1(n19395), .B2(n19394), .A(n19418), .ZN(n19429) );
  OR2_X1 U22456 ( .A1(n19426), .A2(n19396), .ZN(n19397) );
  AOI22_X1 U22457 ( .A1(n19412), .A2(n19398), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19397), .ZN(n19428) );
  OAI22_X1 U22458 ( .A1(n19402), .A2(n19401), .B1(n19400), .B2(n19399), .ZN(
        n19403) );
  AOI221_X1 U22459 ( .B1(n19406), .B2(n19405), .C1(n19404), .C2(n19405), .A(
        n19403), .ZN(n19551) );
  NOR3_X1 U22460 ( .A1(n19408), .A2(n13074), .A3(n19407), .ZN(n19411) );
  OAI22_X1 U22461 ( .A1(n19411), .A2(n19410), .B1(n19409), .B2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19413) );
  NAND2_X1 U22462 ( .A1(n19413), .A2(n19412), .ZN(n19415) );
  OAI211_X1 U22463 ( .C1(n19416), .C2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n19415), .B(n19414), .ZN(n19417) );
  OAI21_X1 U22464 ( .B1(n13077), .B2(n19418), .A(n19417), .ZN(n19419) );
  AOI211_X1 U22465 ( .C1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n19428), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n19419), .ZN(n19425) );
  NOR2_X1 U22466 ( .A1(P3_MORE_REG_SCAN_IN), .A2(P3_FLUSH_REG_SCAN_IN), .ZN(
        n19423) );
  OAI211_X1 U22467 ( .C1(n19423), .C2(n19422), .A(n19421), .B(n19420), .ZN(
        n19424) );
  AOI211_X1 U22468 ( .C1(n19426), .C2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n19425), .B(n19424), .ZN(n19427) );
  OAI211_X1 U22469 ( .C1(n19429), .C2(n19428), .A(n19551), .B(n19427), .ZN(
        n19434) );
  AOI211_X1 U22470 ( .C1(n19432), .C2(n19431), .A(n19430), .B(n19434), .ZN(
        n19537) );
  AOI21_X1 U22471 ( .B1(n19563), .B2(n19555), .A(n19537), .ZN(n19439) );
  OAI211_X1 U22472 ( .C1(P3_STATE2_REG_1__SCAN_IN), .C2(n19438), .A(n19439), 
        .B(n19433), .ZN(n19435) );
  AOI22_X1 U22473 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19435), .B1(n19561), 
        .B2(n19434), .ZN(n19436) );
  OAI21_X1 U22474 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19437), .A(n19436), 
        .ZN(P3_U2996) );
  NAND2_X1 U22475 ( .A1(n19563), .A2(n18290), .ZN(n19442) );
  NAND4_X1 U22476 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n19563), .A4(n19555), .ZN(n19445) );
  NAND3_X1 U22477 ( .A1(n19440), .A2(n19439), .A3(n19438), .ZN(n19441) );
  NAND4_X1 U22478 ( .A1(n19443), .A2(n19442), .A3(n19445), .A4(n19441), .ZN(
        P3_U2997) );
  NAND2_X1 U22479 ( .A1(n19555), .A2(n19444), .ZN(n19447) );
  AND4_X1 U22480 ( .A1(n19447), .A2(n19446), .A3(n19445), .A4(n19538), .ZN(
        P3_U2998) );
  AND2_X1 U22481 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19448), .ZN(
        P3_U2999) );
  AND2_X1 U22482 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19448), .ZN(
        P3_U3000) );
  AND2_X1 U22483 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19448), .ZN(
        P3_U3001) );
  AND2_X1 U22484 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19448), .ZN(
        P3_U3002) );
  AND2_X1 U22485 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19448), .ZN(
        P3_U3003) );
  AND2_X1 U22486 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19448), .ZN(
        P3_U3004) );
  AND2_X1 U22487 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19448), .ZN(
        P3_U3005) );
  AND2_X1 U22488 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19448), .ZN(
        P3_U3006) );
  AND2_X1 U22489 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19448), .ZN(
        P3_U3007) );
  AND2_X1 U22490 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19448), .ZN(
        P3_U3008) );
  AND2_X1 U22491 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19448), .ZN(
        P3_U3009) );
  AND2_X1 U22492 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19449), .ZN(
        P3_U3010) );
  AND2_X1 U22493 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19449), .ZN(
        P3_U3011) );
  AND2_X1 U22494 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19449), .ZN(
        P3_U3012) );
  AND2_X1 U22495 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19449), .ZN(
        P3_U3013) );
  AND2_X1 U22496 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19449), .ZN(
        P3_U3014) );
  AND2_X1 U22497 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19449), .ZN(
        P3_U3015) );
  AND2_X1 U22498 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19449), .ZN(
        P3_U3016) );
  AND2_X1 U22499 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19449), .ZN(
        P3_U3017) );
  AND2_X1 U22500 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19449), .ZN(
        P3_U3018) );
  AND2_X1 U22501 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19449), .ZN(
        P3_U3019) );
  AND2_X1 U22502 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19449), .ZN(
        P3_U3020) );
  AND2_X1 U22503 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19449), .ZN(P3_U3021) );
  INV_X1 U22504 ( .A(P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(n21476) );
  NOR2_X1 U22505 ( .A1(n21476), .A2(n19536), .ZN(P3_U3022) );
  AND2_X1 U22506 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19448), .ZN(P3_U3023) );
  AND2_X1 U22507 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19449), .ZN(P3_U3024) );
  AND2_X1 U22508 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19448), .ZN(P3_U3025) );
  AND2_X1 U22509 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19449), .ZN(P3_U3026) );
  AND2_X1 U22510 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19449), .ZN(P3_U3027) );
  AND2_X1 U22511 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19449), .ZN(P3_U3028) );
  NAND2_X1 U22512 ( .A1(n19563), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19460) );
  INV_X1 U22513 ( .A(n19460), .ZN(n19457) );
  OAI21_X1 U22514 ( .B1(n19450), .B2(n21300), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19451) );
  AOI22_X1 U22515 ( .A1(n19457), .A2(n19466), .B1(n19568), .B2(n19451), .ZN(
        n19453) );
  NAND3_X1 U22516 ( .A1(NA), .A2(n19464), .A3(n19452), .ZN(n19458) );
  OAI211_X1 U22517 ( .C1(P3_STATE_REG_0__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n19453), .B(n19458), .ZN(P3_U3029) );
  NAND2_X1 U22518 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n19459) );
  AOI22_X1 U22519 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n19459), .B1(HOLD), 
        .B2(n19454), .ZN(n19456) );
  INV_X1 U22520 ( .A(n19553), .ZN(n19455) );
  OAI211_X1 U22521 ( .C1(n19456), .C2(n19464), .A(n19460), .B(n19455), .ZN(
        P3_U3030) );
  AOI21_X1 U22522 ( .B1(n19464), .B2(n19458), .A(n19457), .ZN(n19465) );
  INV_X1 U22523 ( .A(n19459), .ZN(n19462) );
  OAI22_X1 U22524 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19460), .ZN(n19461) );
  OAI22_X1 U22525 ( .A1(n19462), .A2(n19461), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19463) );
  OAI22_X1 U22526 ( .A1(n19465), .A2(n19466), .B1(n19464), .B2(n19463), .ZN(
        P3_U3031) );
  INV_X2 U22527 ( .A(n19468), .ZN(n19527) );
  OAI222_X1 U22528 ( .A1(n19541), .A2(n19527), .B1(n19467), .B2(n19524), .C1(
        n19469), .C2(n19522), .ZN(P3_U3032) );
  OAI222_X1 U22529 ( .A1(n19522), .A2(n19472), .B1(n19470), .B2(n19524), .C1(
        n19469), .C2(n19527), .ZN(P3_U3033) );
  OAI222_X1 U22530 ( .A1(n19472), .A2(n19527), .B1(n19471), .B2(n19524), .C1(
        n19473), .C2(n19522), .ZN(P3_U3034) );
  INV_X1 U22531 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19475) );
  OAI222_X1 U22532 ( .A1(n19522), .A2(n19475), .B1(n19474), .B2(n19524), .C1(
        n19473), .C2(n19527), .ZN(P3_U3035) );
  OAI222_X1 U22533 ( .A1(n19522), .A2(n19477), .B1(n19476), .B2(n19524), .C1(
        n19475), .C2(n19527), .ZN(P3_U3036) );
  OAI222_X1 U22534 ( .A1(n19522), .A2(n19479), .B1(n19478), .B2(n19524), .C1(
        n19477), .C2(n19527), .ZN(P3_U3037) );
  OAI222_X1 U22535 ( .A1(n19522), .A2(n19482), .B1(n19480), .B2(n19531), .C1(
        n19479), .C2(n19527), .ZN(P3_U3038) );
  OAI222_X1 U22536 ( .A1(n19482), .A2(n19527), .B1(n19481), .B2(n19524), .C1(
        n19483), .C2(n19522), .ZN(P3_U3039) );
  OAI222_X1 U22537 ( .A1(n19522), .A2(n19486), .B1(n19484), .B2(n19531), .C1(
        n19483), .C2(n19527), .ZN(P3_U3040) );
  INV_X1 U22538 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19487) );
  OAI222_X1 U22539 ( .A1(n19486), .A2(n19527), .B1(n19485), .B2(n19531), .C1(
        n19487), .C2(n19522), .ZN(P3_U3041) );
  OAI222_X1 U22540 ( .A1(n19522), .A2(n19489), .B1(n19488), .B2(n19531), .C1(
        n19487), .C2(n19527), .ZN(P3_U3042) );
  OAI222_X1 U22541 ( .A1(n19522), .A2(n19491), .B1(n19490), .B2(n19531), .C1(
        n19489), .C2(n19527), .ZN(P3_U3043) );
  OAI222_X1 U22542 ( .A1(n19522), .A2(n19494), .B1(n19492), .B2(n19531), .C1(
        n19491), .C2(n19527), .ZN(P3_U3044) );
  OAI222_X1 U22543 ( .A1(n19494), .A2(n19527), .B1(n19493), .B2(n19531), .C1(
        n19495), .C2(n19522), .ZN(P3_U3045) );
  OAI222_X1 U22544 ( .A1(n19522), .A2(n19497), .B1(n19496), .B2(n19531), .C1(
        n19495), .C2(n19527), .ZN(P3_U3046) );
  OAI222_X1 U22545 ( .A1(n19522), .A2(n19500), .B1(n19498), .B2(n19531), .C1(
        n19497), .C2(n19527), .ZN(P3_U3047) );
  OAI222_X1 U22546 ( .A1(n19500), .A2(n19527), .B1(n19499), .B2(n19531), .C1(
        n19501), .C2(n19522), .ZN(P3_U3048) );
  OAI222_X1 U22547 ( .A1(n19522), .A2(n19504), .B1(n19502), .B2(n19531), .C1(
        n19501), .C2(n19527), .ZN(P3_U3049) );
  OAI222_X1 U22548 ( .A1(n19504), .A2(n19527), .B1(n19503), .B2(n19531), .C1(
        n19506), .C2(n19522), .ZN(P3_U3050) );
  OAI222_X1 U22549 ( .A1(n19506), .A2(n19527), .B1(n19505), .B2(n19531), .C1(
        n19507), .C2(n19522), .ZN(P3_U3051) );
  OAI222_X1 U22550 ( .A1(n19522), .A2(n19509), .B1(n19508), .B2(n19531), .C1(
        n19507), .C2(n19527), .ZN(P3_U3052) );
  OAI222_X1 U22551 ( .A1(n19522), .A2(n19511), .B1(n19510), .B2(n19531), .C1(
        n19509), .C2(n19527), .ZN(P3_U3053) );
  OAI222_X1 U22552 ( .A1(n19522), .A2(n19513), .B1(n19512), .B2(n19524), .C1(
        n19511), .C2(n19527), .ZN(P3_U3054) );
  OAI222_X1 U22553 ( .A1(n19522), .A2(n19515), .B1(n19514), .B2(n19524), .C1(
        n19513), .C2(n19527), .ZN(P3_U3055) );
  OAI222_X1 U22554 ( .A1(n19522), .A2(n17194), .B1(n19516), .B2(n19524), .C1(
        n19515), .C2(n19527), .ZN(P3_U3056) );
  OAI222_X1 U22555 ( .A1(n19522), .A2(n17052), .B1(n21507), .B2(n19524), .C1(
        n17194), .C2(n19527), .ZN(P3_U3057) );
  INV_X1 U22556 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19519) );
  OAI222_X1 U22557 ( .A1(n19522), .A2(n19519), .B1(n19517), .B2(n19524), .C1(
        n17052), .C2(n19527), .ZN(P3_U3058) );
  OAI222_X1 U22558 ( .A1(n19519), .A2(n19527), .B1(n19518), .B2(n19524), .C1(
        n19520), .C2(n19522), .ZN(P3_U3059) );
  OAI222_X1 U22559 ( .A1(n19522), .A2(n19526), .B1(n19521), .B2(n19524), .C1(
        n19520), .C2(n19527), .ZN(P3_U3060) );
  INV_X1 U22560 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19523) );
  OAI222_X1 U22561 ( .A1(n19527), .A2(n19526), .B1(n19525), .B2(n19524), .C1(
        n19523), .C2(n19522), .ZN(P3_U3061) );
  OAI22_X1 U22562 ( .A1(n19568), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n19524), .ZN(n19528) );
  INV_X1 U22563 ( .A(n19528), .ZN(P3_U3274) );
  OAI22_X1 U22564 ( .A1(n19568), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n19524), .ZN(n19529) );
  INV_X1 U22565 ( .A(n19529), .ZN(P3_U3275) );
  OAI22_X1 U22566 ( .A1(n19568), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n19524), .ZN(n19530) );
  INV_X1 U22567 ( .A(n19530), .ZN(P3_U3276) );
  OAI22_X1 U22568 ( .A1(n19568), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19531), .ZN(n19532) );
  INV_X1 U22569 ( .A(n19532), .ZN(P3_U3277) );
  OAI21_X1 U22570 ( .B1(n19536), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19534), 
        .ZN(n19533) );
  INV_X1 U22571 ( .A(n19533), .ZN(P3_U3280) );
  OAI21_X1 U22572 ( .B1(n19536), .B2(n19535), .A(n19534), .ZN(P3_U3281) );
  NOR2_X1 U22573 ( .A1(n19537), .A2(n19558), .ZN(n19540) );
  OAI21_X1 U22574 ( .B1(n19540), .B2(n19539), .A(n19538), .ZN(P3_U3282) );
  AOI21_X1 U22575 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19542) );
  AOI22_X1 U22576 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19542), .B2(n19541), .ZN(n19545) );
  INV_X1 U22577 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19544) );
  AOI22_X1 U22578 ( .A1(n19548), .A2(n19545), .B1(n19544), .B2(n19543), .ZN(
        P3_U3292) );
  INV_X1 U22579 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19547) );
  OAI21_X1 U22580 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19548), .ZN(n19546) );
  OAI21_X1 U22581 ( .B1(n19548), .B2(n19547), .A(n19546), .ZN(P3_U3293) );
  INV_X1 U22582 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19549) );
  AOI22_X1 U22583 ( .A1(n19531), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19549), 
        .B2(n19568), .ZN(P3_U3294) );
  INV_X1 U22584 ( .A(P3_MORE_REG_SCAN_IN), .ZN(n21460) );
  AOI22_X1 U22585 ( .A1(n19552), .A2(n19551), .B1(n21460), .B2(n19550), .ZN(
        P3_U3295) );
  OAI21_X1 U22586 ( .B1(n19554), .B2(P3_STATEBS16_REG_SCAN_IN), .A(n19553), 
        .ZN(n19556) );
  AOI211_X1 U22587 ( .C1(n19557), .C2(n19556), .A(n19563), .B(n19555), .ZN(
        n19559) );
  OAI22_X1 U22588 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .B1(n19559), .B2(n19558), .ZN(n19567) );
  OAI22_X1 U22589 ( .A1(n19563), .A2(n19562), .B1(n19561), .B2(n19560), .ZN(
        n19564) );
  NOR2_X1 U22590 ( .A1(n19565), .A2(n19564), .ZN(n19566) );
  MUX2_X1 U22591 ( .A(n19567), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n19566), 
        .Z(P3_U3296) );
  OAI22_X1 U22592 ( .A1(n19568), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n19524), .ZN(n19569) );
  INV_X1 U22593 ( .A(n19569), .ZN(P3_U3297) );
  OAI21_X1 U22594 ( .B1(n19570), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n19572), 
        .ZN(n19575) );
  OAI22_X1 U22595 ( .A1(n19575), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19572), 
        .B2(n19571), .ZN(n19573) );
  INV_X1 U22596 ( .A(n19573), .ZN(P3_U3298) );
  OAI21_X1 U22597 ( .B1(n19575), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n19574), 
        .ZN(n19576) );
  INV_X1 U22598 ( .A(n19576), .ZN(P3_U3299) );
  INV_X1 U22599 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20385) );
  NAND2_X1 U22600 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20391), .ZN(n20378) );
  NAND2_X1 U22601 ( .A1(n20385), .A2(n20370), .ZN(n20374) );
  OAI21_X1 U22602 ( .B1(n20385), .B2(n20378), .A(n20374), .ZN(n20456) );
  AOI21_X1 U22603 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20456), .ZN(n19577) );
  INV_X1 U22604 ( .A(n19577), .ZN(P2_U2815) );
  AOI22_X1 U22605 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(n20483), .B1(n20383), .B2(
        n20385), .ZN(n19578) );
  OAI21_X1 U22606 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n20483), .A(n19578), 
        .ZN(P2_U2817) );
  OAI21_X1 U22607 ( .B1(n20383), .B2(BS16), .A(n20456), .ZN(n20454) );
  OAI21_X1 U22608 ( .B1(n20456), .B2(n20122), .A(n20454), .ZN(P2_U2818) );
  INV_X1 U22609 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n19580) );
  OAI21_X1 U22610 ( .B1(n19581), .B2(n19580), .A(n19579), .ZN(P2_U2819) );
  NOR4_X1 U22611 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19585) );
  NOR4_X1 U22612 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19584) );
  NOR4_X1 U22613 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19583) );
  NOR4_X1 U22614 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19582) );
  NAND4_X1 U22615 ( .A1(n19585), .A2(n19584), .A3(n19583), .A4(n19582), .ZN(
        n19591) );
  NOR4_X1 U22616 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19589) );
  AOI211_X1 U22617 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19588) );
  NOR4_X1 U22618 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19587) );
  NOR4_X1 U22619 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19586) );
  NAND4_X1 U22620 ( .A1(n19589), .A2(n19588), .A3(n19587), .A4(n19586), .ZN(
        n19590) );
  NOR2_X1 U22621 ( .A1(n19591), .A2(n19590), .ZN(n19602) );
  INV_X1 U22622 ( .A(n19602), .ZN(n19600) );
  NOR2_X1 U22623 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19600), .ZN(n19594) );
  INV_X1 U22624 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19592) );
  AOI22_X1 U22625 ( .A1(n19594), .A2(n19595), .B1(n19600), .B2(n19592), .ZN(
        P2_U2820) );
  OR3_X1 U22626 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19599) );
  INV_X1 U22627 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19593) );
  AOI22_X1 U22628 ( .A1(n19594), .A2(n19599), .B1(n19600), .B2(n19593), .ZN(
        P2_U2821) );
  INV_X1 U22629 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20455) );
  NAND2_X1 U22630 ( .A1(n19594), .A2(n20455), .ZN(n19598) );
  OAI21_X1 U22631 ( .B1(n19595), .B2(n10612), .A(n19602), .ZN(n19596) );
  OAI21_X1 U22632 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19602), .A(n19596), 
        .ZN(n19597) );
  OAI221_X1 U22633 ( .B1(n19598), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19598), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19597), .ZN(P2_U2822) );
  INV_X1 U22634 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19601) );
  OAI221_X1 U22635 ( .B1(n19602), .B2(n19601), .C1(n19600), .C2(n19599), .A(
        n19598), .ZN(P2_U2823) );
  INV_X1 U22636 ( .A(n19603), .ZN(n19610) );
  AOI21_X1 U22637 ( .B1(n19605), .B2(P2_REIP_REG_5__SCAN_IN), .A(n19604), .ZN(
        n19606) );
  OAI21_X1 U22638 ( .B1(n19607), .B2(n11071), .A(n19606), .ZN(n19608) );
  AOI21_X1 U22639 ( .B1(n19610), .B2(n19609), .A(n19608), .ZN(n19624) );
  NOR2_X1 U22640 ( .A1(n19612), .A2(n19611), .ZN(n19620) );
  NOR2_X1 U22641 ( .A1(n19613), .A2(n19615), .ZN(n19614) );
  MUX2_X1 U22642 ( .A(n19615), .B(n19614), .S(n9609), .Z(n19618) );
  NOR3_X1 U22643 ( .A1(n19618), .A2(n19617), .A3(n19616), .ZN(n19619) );
  AOI211_X1 U22644 ( .C1(n19622), .C2(n19621), .A(n19620), .B(n19619), .ZN(
        n19623) );
  OAI211_X1 U22645 ( .C1(n12624), .C2(n19625), .A(n19624), .B(n19623), .ZN(
        P2_U2850) );
  INV_X1 U22646 ( .A(n19626), .ZN(n19710) );
  AOI22_X1 U22647 ( .A1(n19710), .A2(n19648), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19647), .ZN(n19631) );
  XNOR2_X1 U22648 ( .A(n19628), .B(n19627), .ZN(n19629) );
  NAND2_X1 U22649 ( .A1(n19629), .A2(n19649), .ZN(n19630) );
  OAI211_X1 U22650 ( .C1(n19632), .C2(n19655), .A(n19631), .B(n19630), .ZN(
        P2_U2915) );
  AOI22_X1 U22651 ( .A1(n20469), .A2(n19648), .B1(n19647), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19638) );
  OAI21_X1 U22652 ( .B1(n19635), .B2(n19634), .A(n19633), .ZN(n19636) );
  NAND2_X1 U22653 ( .A1(n19636), .A2(n19649), .ZN(n19637) );
  OAI211_X1 U22654 ( .C1(n19639), .C2(n19655), .A(n19638), .B(n19637), .ZN(
        P2_U2916) );
  AOI22_X1 U22655 ( .A1(n19648), .A2(n19640), .B1(n19647), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19645) );
  OAI21_X1 U22656 ( .B1(n19642), .B2(n19650), .A(n19641), .ZN(n19643) );
  NAND2_X1 U22657 ( .A1(n19643), .A2(n19649), .ZN(n19644) );
  OAI211_X1 U22658 ( .C1(n19646), .C2(n19655), .A(n19645), .B(n19644), .ZN(
        P2_U2918) );
  AOI22_X1 U22659 ( .A1(n19648), .A2(n19651), .B1(n19647), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n19654) );
  OAI211_X1 U22660 ( .C1(n19652), .C2(n19651), .A(n19650), .B(n19649), .ZN(
        n19653) );
  OAI211_X1 U22661 ( .C1(n19656), .C2(n19655), .A(n19654), .B(n19653), .ZN(
        P2_U2919) );
  NOR2_X1 U22662 ( .A1(n19662), .A2(n19657), .ZN(P2_U2920) );
  INV_X1 U22663 ( .A(n19658), .ZN(n19659) );
  AOI22_X1 U22664 ( .A1(n19659), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n19694), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19660) );
  OAI21_X1 U22665 ( .B1(n19662), .B2(n19661), .A(n19660), .ZN(P2_U2921) );
  AOI22_X1 U22666 ( .A1(n19694), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19663) );
  OAI21_X1 U22667 ( .B1(n19664), .B2(n19696), .A(n19663), .ZN(P2_U2936) );
  INV_X1 U22668 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19666) );
  AOI22_X1 U22669 ( .A1(n19694), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19665) );
  OAI21_X1 U22670 ( .B1(n19666), .B2(n19696), .A(n19665), .ZN(P2_U2937) );
  AOI22_X1 U22671 ( .A1(n19694), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19667) );
  OAI21_X1 U22672 ( .B1(n19668), .B2(n19696), .A(n19667), .ZN(P2_U2938) );
  AOI22_X1 U22673 ( .A1(n19694), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19669) );
  OAI21_X1 U22674 ( .B1(n19670), .B2(n19696), .A(n19669), .ZN(P2_U2939) );
  AOI22_X1 U22675 ( .A1(n19694), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19671) );
  OAI21_X1 U22676 ( .B1(n19672), .B2(n19696), .A(n19671), .ZN(P2_U2940) );
  AOI22_X1 U22677 ( .A1(n19694), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19673) );
  OAI21_X1 U22678 ( .B1(n19674), .B2(n19696), .A(n19673), .ZN(P2_U2941) );
  AOI22_X1 U22679 ( .A1(n19694), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19675) );
  OAI21_X1 U22680 ( .B1(n19676), .B2(n19696), .A(n19675), .ZN(P2_U2942) );
  AOI22_X1 U22681 ( .A1(n19694), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19677) );
  OAI21_X1 U22682 ( .B1(n19678), .B2(n19696), .A(n19677), .ZN(P2_U2943) );
  AOI22_X1 U22683 ( .A1(n19694), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19679) );
  OAI21_X1 U22684 ( .B1(n19680), .B2(n19696), .A(n19679), .ZN(P2_U2944) );
  AOI22_X1 U22685 ( .A1(n19694), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19681) );
  OAI21_X1 U22686 ( .B1(n19682), .B2(n19696), .A(n19681), .ZN(P2_U2945) );
  AOI22_X1 U22687 ( .A1(n19694), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19683) );
  OAI21_X1 U22688 ( .B1(n19684), .B2(n19696), .A(n19683), .ZN(P2_U2946) );
  INV_X1 U22689 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19686) );
  AOI22_X1 U22690 ( .A1(n19694), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19685) );
  OAI21_X1 U22691 ( .B1(n19686), .B2(n19696), .A(n19685), .ZN(P2_U2947) );
  INV_X1 U22692 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19688) );
  AOI22_X1 U22693 ( .A1(n19694), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19687) );
  OAI21_X1 U22694 ( .B1(n19688), .B2(n19696), .A(n19687), .ZN(P2_U2948) );
  INV_X1 U22695 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19690) );
  AOI22_X1 U22696 ( .A1(n19694), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19689) );
  OAI21_X1 U22697 ( .B1(n19690), .B2(n19696), .A(n19689), .ZN(P2_U2949) );
  INV_X1 U22698 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19692) );
  AOI22_X1 U22699 ( .A1(n19694), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19691) );
  OAI21_X1 U22700 ( .B1(n19692), .B2(n19696), .A(n19691), .ZN(P2_U2950) );
  AOI22_X1 U22701 ( .A1(n19694), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19693), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19695) );
  OAI21_X1 U22702 ( .B1(n12274), .B2(n19696), .A(n19695), .ZN(P2_U2951) );
  AOI22_X1 U22703 ( .A1(n19701), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19700), .ZN(n19699) );
  NAND2_X1 U22704 ( .A1(n19698), .A2(n19697), .ZN(n19702) );
  NAND2_X1 U22705 ( .A1(n19699), .A2(n19702), .ZN(P2_U2966) );
  AOI22_X1 U22706 ( .A1(n19701), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n19700), .ZN(n19703) );
  NAND2_X1 U22707 ( .A1(n19703), .A2(n19702), .ZN(P2_U2981) );
  OAI22_X1 U22708 ( .A1(n19705), .A2(n16417), .B1(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19704), .ZN(n19709) );
  NOR2_X1 U22709 ( .A1(n19707), .A2(n19706), .ZN(n19708) );
  AOI211_X1 U22710 ( .C1(n19710), .C2(n19724), .A(n19709), .B(n19708), .ZN(
        n19715) );
  AOI22_X1 U22711 ( .A1(n19713), .A2(n19721), .B1(n19712), .B2(n19711), .ZN(
        n19714) );
  OAI211_X1 U22712 ( .C1(n19717), .C2(n19716), .A(n19715), .B(n19714), .ZN(
        P2_U3042) );
  AOI22_X1 U22713 ( .A1(n19721), .A2(n19720), .B1(n19719), .B2(n19718), .ZN(
        n19738) );
  OR2_X1 U22714 ( .A1(n19723), .A2(n19722), .ZN(n19734) );
  AOI22_X1 U22715 ( .A1(n19726), .A2(n19725), .B1(n19724), .B2(n20477), .ZN(
        n19733) );
  OR2_X1 U22716 ( .A1(n19728), .A2(n19727), .ZN(n19732) );
  OR2_X1 U22717 ( .A1(n19730), .A2(n19729), .ZN(n19731) );
  AND4_X1 U22718 ( .A1(n19734), .A2(n19733), .A3(n19732), .A4(n19731), .ZN(
        n19737) );
  NAND4_X1 U22719 ( .A1(n19738), .A2(n19737), .A3(n19736), .A4(n19735), .ZN(
        P2_U3044) );
  OR2_X2 U22720 ( .A1(n20214), .A2(n20458), .ZN(n20355) );
  NOR2_X1 U22721 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19848), .ZN(
        n19817) );
  AND2_X1 U22722 ( .A1(n19817), .A2(n20248), .ZN(n19745) );
  INV_X1 U22723 ( .A(n19745), .ZN(n19808) );
  OAI22_X1 U22724 ( .A1(n20355), .A2(n20262), .B1(n19808), .B2(n20249), .ZN(
        n19740) );
  INV_X1 U22725 ( .A(n19740), .ZN(n19753) );
  INV_X1 U22726 ( .A(n19843), .ZN(n19741) );
  INV_X2 U22727 ( .A(n20355), .ZN(n20362) );
  OAI21_X1 U22728 ( .B1(n19741), .B2(n20362), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19742) );
  NAND2_X1 U22729 ( .A1(n19742), .A2(n20463), .ZN(n19751) );
  NOR2_X1 U22730 ( .A1(n19743), .A2(n20471), .ZN(n20358) );
  NOR2_X1 U22731 ( .A1(n19751), .A2(n20358), .ZN(n19744) );
  AOI211_X1 U22732 ( .C1(n19749), .C2(n20252), .A(P2_STATE2_REG_3__SCAN_IN), 
        .B(n19744), .ZN(n19746) );
  OAI21_X2 U22733 ( .B1(n19746), .B2(n19745), .A(n20253), .ZN(n19812) );
  INV_X1 U22734 ( .A(n20358), .ZN(n20310) );
  INV_X1 U22735 ( .A(n19751), .ZN(n19748) );
  NOR2_X1 U22736 ( .A1(n19748), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19750) );
  OAI222_X4 U22737 ( .A1(n19751), .A2(n20310), .B1(n19808), .B2(n19750), .C1(
        n20302), .C2(n19749), .ZN(n19811) );
  AOI22_X1 U22738 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19812), .B1(
        n20307), .B2(n19811), .ZN(n19752) );
  OAI211_X1 U22739 ( .C1(n20318), .C2(n19843), .A(n19753), .B(n19752), .ZN(
        P2_U3048) );
  OAI22_X1 U22740 ( .A1(n20355), .A2(n20324), .B1(n20263), .B2(n19808), .ZN(
        n19754) );
  INV_X1 U22741 ( .A(n19754), .ZN(n19756) );
  AOI22_X1 U22742 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19812), .B1(
        n20320), .B2(n19811), .ZN(n19755) );
  OAI211_X1 U22743 ( .C1(n20264), .C2(n19843), .A(n19756), .B(n19755), .ZN(
        P2_U3049) );
  NAND2_X1 U22744 ( .A1(n19802), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19758) );
  NAND2_X1 U22745 ( .A1(n19803), .A2(BUF1_REG_18__SCAN_IN), .ZN(n19757) );
  NAND2_X1 U22746 ( .A1(n19758), .A2(n19757), .ZN(n20194) );
  NAND2_X1 U22747 ( .A1(n19802), .A2(BUF2_REG_26__SCAN_IN), .ZN(n19760) );
  NAND2_X1 U22748 ( .A1(n19803), .A2(BUF1_REG_26__SCAN_IN), .ZN(n19759) );
  NAND2_X1 U22749 ( .A1(n19807), .A2(n10584), .ZN(n20268) );
  OAI22_X1 U22750 ( .A1(n20355), .A2(n20272), .B1(n19808), .B2(n20268), .ZN(
        n19761) );
  INV_X1 U22751 ( .A(n19761), .ZN(n19764) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19812), .B1(
        n20326), .B2(n19811), .ZN(n19763) );
  OAI211_X1 U22753 ( .C1(n20330), .C2(n19843), .A(n19764), .B(n19763), .ZN(
        P2_U3050) );
  NAND2_X1 U22754 ( .A1(n19802), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19766) );
  NAND2_X1 U22755 ( .A1(n19803), .A2(BUF1_REG_19__SCAN_IN), .ZN(n19765) );
  NAND2_X1 U22756 ( .A1(n19802), .A2(BUF2_REG_27__SCAN_IN), .ZN(n19768) );
  NAND2_X1 U22757 ( .A1(n19803), .A2(BUF1_REG_27__SCAN_IN), .ZN(n19767) );
  NAND2_X1 U22758 ( .A1(n19807), .A2(n10585), .ZN(n20273) );
  OAI22_X1 U22759 ( .A1(n20355), .A2(n20336), .B1(n19808), .B2(n20273), .ZN(
        n19769) );
  INV_X1 U22760 ( .A(n19769), .ZN(n19772) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19812), .B1(
        n20332), .B2(n19811), .ZN(n19771) );
  OAI211_X1 U22762 ( .C1(n20274), .C2(n19843), .A(n19772), .B(n19771), .ZN(
        P2_U3051) );
  NAND2_X1 U22763 ( .A1(n19802), .A2(BUF2_REG_20__SCAN_IN), .ZN(n19774) );
  NAND2_X1 U22764 ( .A1(n19803), .A2(BUF1_REG_20__SCAN_IN), .ZN(n19773) );
  NAND2_X1 U22765 ( .A1(n19802), .A2(BUF2_REG_28__SCAN_IN), .ZN(n19776) );
  NAND2_X1 U22766 ( .A1(n19803), .A2(BUF1_REG_28__SCAN_IN), .ZN(n19775) );
  OAI22_X1 U22767 ( .A1(n20355), .A2(n20282), .B1(n19808), .B2(n20278), .ZN(
        n19778) );
  INV_X1 U22768 ( .A(n19778), .ZN(n19781) );
  AOI22_X1 U22769 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19812), .B1(
        n20338), .B2(n19811), .ZN(n19780) );
  OAI211_X1 U22770 ( .C1(n20342), .C2(n19843), .A(n19781), .B(n19780), .ZN(
        P2_U3052) );
  NAND2_X1 U22771 ( .A1(n19802), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19783) );
  NAND2_X1 U22772 ( .A1(n19803), .A2(BUF1_REG_21__SCAN_IN), .ZN(n19782) );
  NAND2_X1 U22773 ( .A1(n19802), .A2(BUF2_REG_29__SCAN_IN), .ZN(n19785) );
  NAND2_X1 U22774 ( .A1(n19803), .A2(BUF1_REG_29__SCAN_IN), .ZN(n19784) );
  OAI22_X1 U22775 ( .A1(n20355), .A2(n20284), .B1(n19808), .B2(n20283), .ZN(
        n19786) );
  INV_X1 U22776 ( .A(n19786), .ZN(n19789) );
  AOI22_X1 U22777 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19812), .B1(
        n20344), .B2(n19811), .ZN(n19788) );
  OAI211_X1 U22778 ( .C1(n20348), .C2(n19843), .A(n19789), .B(n19788), .ZN(
        P2_U3053) );
  NAND2_X1 U22779 ( .A1(n19802), .A2(BUF2_REG_22__SCAN_IN), .ZN(n19791) );
  NAND2_X1 U22780 ( .A1(n19803), .A2(BUF1_REG_22__SCAN_IN), .ZN(n19790) );
  NAND2_X1 U22781 ( .A1(n19802), .A2(BUF2_REG_30__SCAN_IN), .ZN(n19793) );
  NAND2_X1 U22782 ( .A1(n19803), .A2(BUF1_REG_30__SCAN_IN), .ZN(n19792) );
  OAI22_X1 U22783 ( .A1(n20355), .A2(n20289), .B1(n19808), .B2(n20288), .ZN(
        n19796) );
  INV_X1 U22784 ( .A(n19796), .ZN(n19799) );
  AOI22_X1 U22785 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19812), .B1(
        n20350), .B2(n19811), .ZN(n19798) );
  OAI211_X1 U22786 ( .C1(n20356), .C2(n19843), .A(n19799), .B(n19798), .ZN(
        P2_U3054) );
  NAND2_X1 U22787 ( .A1(n19802), .A2(BUF2_REG_23__SCAN_IN), .ZN(n19801) );
  NAND2_X1 U22788 ( .A1(n19803), .A2(BUF1_REG_23__SCAN_IN), .ZN(n19800) );
  NAND2_X1 U22789 ( .A1(n19802), .A2(BUF2_REG_31__SCAN_IN), .ZN(n19805) );
  NAND2_X1 U22790 ( .A1(n19803), .A2(BUF1_REG_31__SCAN_IN), .ZN(n19804) );
  NAND2_X1 U22791 ( .A1(n19807), .A2(n19806), .ZN(n20293) );
  OAI22_X1 U22792 ( .A1(n20355), .A2(n20367), .B1(n19808), .B2(n20293), .ZN(
        n19809) );
  INV_X1 U22793 ( .A(n19809), .ZN(n19814) );
  AOI22_X1 U22794 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19812), .B1(
        n20359), .B2(n19811), .ZN(n19813) );
  OAI211_X1 U22795 ( .C1(n20295), .C2(n19843), .A(n19814), .B(n19813), .ZN(
        P2_U3055) );
  AND2_X1 U22796 ( .A1(n20176), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20080) );
  NAND2_X1 U22797 ( .A1(n20080), .A2(n19876), .ZN(n19820) );
  AND2_X1 U22798 ( .A1(n19820), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19815) );
  NAND2_X1 U22799 ( .A1(n19816), .A2(n19815), .ZN(n19822) );
  INV_X1 U22800 ( .A(n19817), .ZN(n19819) );
  OAI21_X1 U22801 ( .B1(n19819), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20302), 
        .ZN(n19818) );
  INV_X1 U22802 ( .A(n19820), .ZN(n19838) );
  AOI22_X1 U22803 ( .A1(n19839), .A2(n20307), .B1(n20306), .B2(n19838), .ZN(
        n19825) );
  OAI21_X1 U22804 ( .B1(n20010), .B2(n20091), .A(n19819), .ZN(n19823) );
  NAND2_X1 U22805 ( .A1(n19820), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19821) );
  NAND4_X1 U22806 ( .A1(n19823), .A2(n20253), .A3(n19822), .A4(n19821), .ZN(
        n19840) );
  AOI22_X1 U22807 ( .A1(n19840), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n19869), .B2(n20189), .ZN(n19824) );
  OAI211_X1 U22808 ( .C1(n20262), .C2(n19843), .A(n19825), .B(n19824), .ZN(
        P2_U3056) );
  AOI22_X1 U22809 ( .A1(n19839), .A2(n20320), .B1(n20319), .B2(n19838), .ZN(
        n19827) );
  AOI22_X1 U22810 ( .A1(n19840), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n19869), .B2(n20321), .ZN(n19826) );
  OAI211_X1 U22811 ( .C1(n20324), .C2(n19843), .A(n19827), .B(n19826), .ZN(
        P2_U3057) );
  AOI22_X1 U22812 ( .A1(n19839), .A2(n20326), .B1(n19838), .B2(n20325), .ZN(
        n19829) );
  AOI22_X1 U22813 ( .A1(n19840), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n19869), .B2(n20194), .ZN(n19828) );
  OAI211_X1 U22814 ( .C1(n20272), .C2(n19843), .A(n19829), .B(n19828), .ZN(
        P2_U3058) );
  AOI22_X1 U22815 ( .A1(n19839), .A2(n20332), .B1(n19838), .B2(n20331), .ZN(
        n19831) );
  AOI22_X1 U22816 ( .A1(n19840), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n19869), .B2(n20333), .ZN(n19830) );
  OAI211_X1 U22817 ( .C1(n20336), .C2(n19843), .A(n19831), .B(n19830), .ZN(
        P2_U3059) );
  AOI22_X1 U22818 ( .A1(n19839), .A2(n20338), .B1(n19838), .B2(n20337), .ZN(
        n19833) );
  AOI22_X1 U22819 ( .A1(n19840), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n19869), .B2(n20199), .ZN(n19832) );
  OAI211_X1 U22820 ( .C1(n20282), .C2(n19843), .A(n19833), .B(n19832), .ZN(
        P2_U3060) );
  AOI22_X1 U22821 ( .A1(n19839), .A2(n20344), .B1(n19838), .B2(n20343), .ZN(
        n19835) );
  AOI22_X1 U22822 ( .A1(n19840), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n19869), .B2(n20202), .ZN(n19834) );
  OAI211_X1 U22823 ( .C1(n20284), .C2(n19843), .A(n19835), .B(n19834), .ZN(
        P2_U3061) );
  AOI22_X1 U22824 ( .A1(n19839), .A2(n20350), .B1(n19838), .B2(n20349), .ZN(
        n19837) );
  AOI22_X1 U22825 ( .A1(n19840), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n19869), .B2(n20205), .ZN(n19836) );
  OAI211_X1 U22826 ( .C1(n20289), .C2(n19843), .A(n19837), .B(n19836), .ZN(
        P2_U3062) );
  AOI22_X1 U22827 ( .A1(n19839), .A2(n20359), .B1(n19838), .B2(n20357), .ZN(
        n19842) );
  AOI22_X1 U22828 ( .A1(n19840), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n19869), .B2(n20361), .ZN(n19841) );
  OAI211_X1 U22829 ( .C1(n20367), .C2(n19843), .A(n19842), .B(n19841), .ZN(
        P2_U3063) );
  NOR2_X1 U22830 ( .A1(n20176), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20118) );
  NAND2_X1 U22831 ( .A1(n20118), .A2(n19876), .ZN(n19849) );
  INV_X1 U22832 ( .A(n19849), .ZN(n19867) );
  OAI21_X1 U22833 ( .B1(n9731), .B2(n19867), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19845) );
  AOI22_X1 U22834 ( .A1(n19868), .A2(n20307), .B1(n20306), .B2(n19867), .ZN(
        n19854) );
  AOI21_X1 U22835 ( .B1(n19911), .B2(n19846), .A(n20122), .ZN(n19852) );
  INV_X1 U22836 ( .A(n19847), .ZN(n20179) );
  NOR2_X1 U22837 ( .A1(n20179), .A2(n19848), .ZN(n19851) );
  OAI211_X1 U22838 ( .C1(n19852), .C2(n19851), .A(n20128), .B(n19850), .ZN(
        n19870) );
  AOI22_X1 U22839 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19870), .B1(
        n19869), .B2(n20315), .ZN(n19853) );
  OAI211_X1 U22840 ( .C1(n20318), .C2(n19911), .A(n19854), .B(n19853), .ZN(
        P2_U3064) );
  AOI22_X1 U22841 ( .A1(n19868), .A2(n20320), .B1(n20319), .B2(n19867), .ZN(
        n19856) );
  AOI22_X1 U22842 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19870), .B1(
        n19869), .B2(n20226), .ZN(n19855) );
  OAI211_X1 U22843 ( .C1(n20264), .C2(n19911), .A(n19856), .B(n19855), .ZN(
        P2_U3065) );
  AOI22_X1 U22844 ( .A1(n19868), .A2(n20326), .B1(n19867), .B2(n20325), .ZN(
        n19858) );
  AOI22_X1 U22845 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19870), .B1(
        n19869), .B2(n20327), .ZN(n19857) );
  OAI211_X1 U22846 ( .C1(n20330), .C2(n19911), .A(n19858), .B(n19857), .ZN(
        P2_U3066) );
  AOI22_X1 U22847 ( .A1(n19868), .A2(n20332), .B1(n19867), .B2(n20331), .ZN(
        n19860) );
  AOI22_X1 U22848 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19870), .B1(
        n19869), .B2(n20231), .ZN(n19859) );
  OAI211_X1 U22849 ( .C1(n20274), .C2(n19911), .A(n19860), .B(n19859), .ZN(
        P2_U3067) );
  AOI22_X1 U22850 ( .A1(n19868), .A2(n20338), .B1(n19867), .B2(n20337), .ZN(
        n19862) );
  AOI22_X1 U22851 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19870), .B1(
        n19869), .B2(n20339), .ZN(n19861) );
  OAI211_X1 U22852 ( .C1(n20342), .C2(n19911), .A(n19862), .B(n19861), .ZN(
        P2_U3068) );
  AOI22_X1 U22853 ( .A1(n19868), .A2(n20344), .B1(n19867), .B2(n20343), .ZN(
        n19864) );
  AOI22_X1 U22854 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19870), .B1(
        n19869), .B2(n20345), .ZN(n19863) );
  OAI211_X1 U22855 ( .C1(n20348), .C2(n19911), .A(n19864), .B(n19863), .ZN(
        P2_U3069) );
  AOI22_X1 U22856 ( .A1(n19868), .A2(n20350), .B1(n19867), .B2(n20349), .ZN(
        n19866) );
  AOI22_X1 U22857 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19870), .B1(
        n19869), .B2(n20351), .ZN(n19865) );
  OAI211_X1 U22858 ( .C1(n20356), .C2(n19911), .A(n19866), .B(n19865), .ZN(
        P2_U3070) );
  AOI22_X1 U22859 ( .A1(n19868), .A2(n20359), .B1(n19867), .B2(n20357), .ZN(
        n19872) );
  AOI22_X1 U22860 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19870), .B1(
        n19869), .B2(n20241), .ZN(n19871) );
  OAI211_X1 U22861 ( .C1(n20295), .C2(n19911), .A(n19872), .B(n19871), .ZN(
        P2_U3071) );
  OR2_X2 U22862 ( .A1(n20017), .A2(n19875), .ZN(n19949) );
  NAND2_X1 U22863 ( .A1(n19873), .A2(n19876), .ZN(n19905) );
  OAI22_X1 U22864 ( .A1(n19911), .A2(n20262), .B1(n19905), .B2(n20249), .ZN(
        n19874) );
  INV_X1 U22865 ( .A(n19874), .ZN(n19886) );
  OAI21_X1 U22866 ( .B1(n20010), .B2(n19875), .A(n20463), .ZN(n19884) );
  NAND2_X1 U22867 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19876), .ZN(
        n19883) );
  INV_X1 U22868 ( .A(n19883), .ZN(n19878) );
  OAI211_X1 U22869 ( .C1(n19879), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20252), 
        .B(n19905), .ZN(n19877) );
  OAI211_X1 U22870 ( .C1(n19884), .C2(n19878), .A(n20128), .B(n19877), .ZN(
        n19908) );
  INV_X1 U22871 ( .A(n19879), .ZN(n19881) );
  INV_X1 U22872 ( .A(n19905), .ZN(n19880) );
  OAI21_X1 U22873 ( .B1(n19881), .B2(n19880), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19882) );
  AOI22_X1 U22874 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19908), .B1(
        n20307), .B2(n19907), .ZN(n19885) );
  OAI211_X1 U22875 ( .C1(n20318), .C2(n19949), .A(n19886), .B(n19885), .ZN(
        P2_U3072) );
  OAI22_X1 U22876 ( .A1(n19911), .A2(n20324), .B1(n20263), .B2(n19905), .ZN(
        n19887) );
  INV_X1 U22877 ( .A(n19887), .ZN(n19889) );
  AOI22_X1 U22878 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19908), .B1(
        n20320), .B2(n19907), .ZN(n19888) );
  OAI211_X1 U22879 ( .C1(n20264), .C2(n19949), .A(n19889), .B(n19888), .ZN(
        P2_U3073) );
  OAI22_X1 U22880 ( .A1(n19949), .A2(n20330), .B1(n19905), .B2(n20268), .ZN(
        n19890) );
  INV_X1 U22881 ( .A(n19890), .ZN(n19892) );
  AOI22_X1 U22882 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19908), .B1(
        n20326), .B2(n19907), .ZN(n19891) );
  OAI211_X1 U22883 ( .C1(n20272), .C2(n19911), .A(n19892), .B(n19891), .ZN(
        P2_U3074) );
  OAI22_X1 U22884 ( .A1(n19949), .A2(n20274), .B1(n19905), .B2(n20273), .ZN(
        n19893) );
  INV_X1 U22885 ( .A(n19893), .ZN(n19895) );
  AOI22_X1 U22886 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19908), .B1(
        n20332), .B2(n19907), .ZN(n19894) );
  OAI211_X1 U22887 ( .C1(n20336), .C2(n19911), .A(n19895), .B(n19894), .ZN(
        P2_U3075) );
  OAI22_X1 U22888 ( .A1(n19911), .A2(n20282), .B1(n19905), .B2(n20278), .ZN(
        n19896) );
  INV_X1 U22889 ( .A(n19896), .ZN(n19898) );
  AOI22_X1 U22890 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19908), .B1(
        n20338), .B2(n19907), .ZN(n19897) );
  OAI211_X1 U22891 ( .C1(n20342), .C2(n19949), .A(n19898), .B(n19897), .ZN(
        P2_U3076) );
  OAI22_X1 U22892 ( .A1(n19949), .A2(n20348), .B1(n19905), .B2(n20283), .ZN(
        n19899) );
  INV_X1 U22893 ( .A(n19899), .ZN(n19901) );
  AOI22_X1 U22894 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19908), .B1(
        n20344), .B2(n19907), .ZN(n19900) );
  OAI211_X1 U22895 ( .C1(n20284), .C2(n19911), .A(n19901), .B(n19900), .ZN(
        P2_U3077) );
  OAI22_X1 U22896 ( .A1(n19911), .A2(n20289), .B1(n19905), .B2(n20288), .ZN(
        n19902) );
  INV_X1 U22897 ( .A(n19902), .ZN(n19904) );
  AOI22_X1 U22898 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19908), .B1(
        n20350), .B2(n19907), .ZN(n19903) );
  OAI211_X1 U22899 ( .C1(n20356), .C2(n19949), .A(n19904), .B(n19903), .ZN(
        P2_U3078) );
  OAI22_X1 U22900 ( .A1(n19949), .A2(n20295), .B1(n19905), .B2(n20293), .ZN(
        n19906) );
  INV_X1 U22901 ( .A(n19906), .ZN(n19910) );
  AOI22_X1 U22902 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19908), .B1(
        n20359), .B2(n19907), .ZN(n19909) );
  OAI211_X1 U22903 ( .C1(n20367), .C2(n19911), .A(n19910), .B(n19909), .ZN(
        P2_U3079) );
  OR2_X1 U22904 ( .A1(n19912), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19948) );
  OAI22_X1 U22905 ( .A1(n19975), .A2(n20318), .B1(n19948), .B2(n20249), .ZN(
        n19913) );
  INV_X1 U22906 ( .A(n19913), .ZN(n19929) );
  INV_X1 U22907 ( .A(n19949), .ZN(n19914) );
  OAI21_X1 U22908 ( .B1(n19915), .B2(n19914), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19916) );
  NAND2_X1 U22909 ( .A1(n19916), .A2(n20463), .ZN(n19927) );
  INV_X1 U22910 ( .A(n19917), .ZN(n19918) );
  NAND2_X1 U22911 ( .A1(n19918), .A2(n20179), .ZN(n20186) );
  NOR2_X1 U22912 ( .A1(n20186), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19922) );
  INV_X1 U22913 ( .A(n19919), .ZN(n19924) );
  OAI21_X1 U22914 ( .B1(n19924), .B2(n20302), .A(n20304), .ZN(n19920) );
  NAND2_X1 U22915 ( .A1(n19920), .A2(n19948), .ZN(n19921) );
  OAI211_X1 U22916 ( .C1(n19927), .C2(n19922), .A(n20128), .B(n19921), .ZN(
        n19952) );
  INV_X1 U22917 ( .A(n19922), .ZN(n19926) );
  INV_X1 U22918 ( .A(n19948), .ZN(n19923) );
  OAI21_X1 U22919 ( .B1(n19924), .B2(n19923), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19925) );
  AOI22_X1 U22920 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19952), .B1(
        n19951), .B2(n20307), .ZN(n19928) );
  OAI211_X1 U22921 ( .C1(n20262), .C2(n19949), .A(n19929), .B(n19928), .ZN(
        P2_U3080) );
  OAI22_X1 U22922 ( .A1(n19975), .A2(n20264), .B1(n20263), .B2(n19948), .ZN(
        n19930) );
  INV_X1 U22923 ( .A(n19930), .ZN(n19932) );
  AOI22_X1 U22924 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19952), .B1(
        n19951), .B2(n20320), .ZN(n19931) );
  OAI211_X1 U22925 ( .C1(n20324), .C2(n19949), .A(n19932), .B(n19931), .ZN(
        P2_U3081) );
  OAI22_X1 U22926 ( .A1(n19949), .A2(n20272), .B1(n19948), .B2(n20268), .ZN(
        n19933) );
  INV_X1 U22927 ( .A(n19933), .ZN(n19935) );
  AOI22_X1 U22928 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19952), .B1(
        n19951), .B2(n20326), .ZN(n19934) );
  OAI211_X1 U22929 ( .C1(n20330), .C2(n19975), .A(n19935), .B(n19934), .ZN(
        P2_U3082) );
  OAI22_X1 U22930 ( .A1(n19949), .A2(n20336), .B1(n19948), .B2(n20273), .ZN(
        n19936) );
  INV_X1 U22931 ( .A(n19936), .ZN(n19938) );
  AOI22_X1 U22932 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19952), .B1(
        n19951), .B2(n20332), .ZN(n19937) );
  OAI211_X1 U22933 ( .C1(n20274), .C2(n19975), .A(n19938), .B(n19937), .ZN(
        P2_U3083) );
  OAI22_X1 U22934 ( .A1(n19949), .A2(n20282), .B1(n19948), .B2(n20278), .ZN(
        n19939) );
  INV_X1 U22935 ( .A(n19939), .ZN(n19941) );
  AOI22_X1 U22936 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19952), .B1(
        n19951), .B2(n20338), .ZN(n19940) );
  OAI211_X1 U22937 ( .C1(n20342), .C2(n19975), .A(n19941), .B(n19940), .ZN(
        P2_U3084) );
  OAI22_X1 U22938 ( .A1(n19975), .A2(n20348), .B1(n19948), .B2(n20283), .ZN(
        n19942) );
  INV_X1 U22939 ( .A(n19942), .ZN(n19944) );
  AOI22_X1 U22940 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19952), .B1(
        n19951), .B2(n20344), .ZN(n19943) );
  OAI211_X1 U22941 ( .C1(n20284), .C2(n19949), .A(n19944), .B(n19943), .ZN(
        P2_U3085) );
  OAI22_X1 U22942 ( .A1(n19975), .A2(n20356), .B1(n19948), .B2(n20288), .ZN(
        n19945) );
  INV_X1 U22943 ( .A(n19945), .ZN(n19947) );
  AOI22_X1 U22944 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19952), .B1(
        n19951), .B2(n20350), .ZN(n19946) );
  OAI211_X1 U22945 ( .C1(n20289), .C2(n19949), .A(n19947), .B(n19946), .ZN(
        P2_U3086) );
  OAI22_X1 U22946 ( .A1(n19949), .A2(n20367), .B1(n19948), .B2(n20293), .ZN(
        n19950) );
  INV_X1 U22947 ( .A(n19950), .ZN(n19954) );
  AOI22_X1 U22948 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19952), .B1(
        n19951), .B2(n20359), .ZN(n19953) );
  OAI211_X1 U22949 ( .C1(n20295), .C2(n19975), .A(n19954), .B(n19953), .ZN(
        P2_U3087) );
  OAI22_X1 U22950 ( .A1(n20008), .A2(n20330), .B1(n19978), .B2(n20268), .ZN(
        n19955) );
  INV_X1 U22951 ( .A(n19955), .ZN(n19957) );
  AOI22_X1 U22952 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19972), .B1(
        n20326), .B2(n19971), .ZN(n19956) );
  OAI211_X1 U22953 ( .C1(n20272), .C2(n19975), .A(n19957), .B(n19956), .ZN(
        P2_U3090) );
  OAI22_X1 U22954 ( .A1(n19975), .A2(n20336), .B1(n19978), .B2(n20273), .ZN(
        n19958) );
  INV_X1 U22955 ( .A(n19958), .ZN(n19960) );
  AOI22_X1 U22956 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19972), .B1(
        n20332), .B2(n19971), .ZN(n19959) );
  OAI211_X1 U22957 ( .C1(n20274), .C2(n20008), .A(n19960), .B(n19959), .ZN(
        P2_U3091) );
  OAI22_X1 U22958 ( .A1(n19975), .A2(n20282), .B1(n19978), .B2(n20278), .ZN(
        n19961) );
  INV_X1 U22959 ( .A(n19961), .ZN(n19963) );
  AOI22_X1 U22960 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19972), .B1(
        n20338), .B2(n19971), .ZN(n19962) );
  OAI211_X1 U22961 ( .C1(n20342), .C2(n20008), .A(n19963), .B(n19962), .ZN(
        P2_U3092) );
  OAI22_X1 U22962 ( .A1(n20008), .A2(n20348), .B1(n19978), .B2(n20283), .ZN(
        n19964) );
  INV_X1 U22963 ( .A(n19964), .ZN(n19966) );
  AOI22_X1 U22964 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19972), .B1(
        n20344), .B2(n19971), .ZN(n19965) );
  OAI211_X1 U22965 ( .C1(n20284), .C2(n19975), .A(n19966), .B(n19965), .ZN(
        P2_U3093) );
  OAI22_X1 U22966 ( .A1(n20008), .A2(n20356), .B1(n19978), .B2(n20288), .ZN(
        n19967) );
  INV_X1 U22967 ( .A(n19967), .ZN(n19969) );
  AOI22_X1 U22968 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19972), .B1(
        n20350), .B2(n19971), .ZN(n19968) );
  OAI211_X1 U22969 ( .C1(n20289), .C2(n19975), .A(n19969), .B(n19968), .ZN(
        P2_U3094) );
  OAI22_X1 U22970 ( .A1(n20008), .A2(n20295), .B1(n19978), .B2(n20293), .ZN(
        n19970) );
  INV_X1 U22971 ( .A(n19970), .ZN(n19974) );
  AOI22_X1 U22972 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19972), .B1(
        n20359), .B2(n19971), .ZN(n19973) );
  OAI211_X1 U22973 ( .C1(n20367), .C2(n19975), .A(n19974), .B(n19973), .ZN(
        P2_U3095) );
  NAND2_X1 U22974 ( .A1(n20009), .A2(n20248), .ZN(n19981) );
  AND2_X1 U22975 ( .A1(n19981), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19976) );
  NAND2_X1 U22976 ( .A1(n19977), .A2(n19976), .ZN(n19983) );
  INV_X1 U22977 ( .A(n19983), .ZN(n19980) );
  NAND2_X1 U22978 ( .A1(n19981), .A2(n19978), .ZN(n19986) );
  AOI21_X1 U22979 ( .B1(n19986), .B2(n20304), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19979) );
  INV_X1 U22980 ( .A(n19981), .ZN(n20003) );
  AOI22_X1 U22981 ( .A1(n20004), .A2(n20307), .B1(n20003), .B2(n20306), .ZN(
        n19990) );
  NAND2_X1 U22982 ( .A1(n20313), .A2(n19982), .ZN(n19988) );
  AOI21_X1 U22983 ( .B1(n20008), .B2(n19988), .A(n20122), .ZN(n19987) );
  OAI211_X1 U22984 ( .C1(n20003), .C2(n20304), .A(n19983), .B(n20253), .ZN(
        n19984) );
  INV_X1 U22985 ( .A(n19984), .ZN(n19985) );
  AOI22_X1 U22986 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20005), .B1(
        n20036), .B2(n20189), .ZN(n19989) );
  OAI211_X1 U22987 ( .C1(n20262), .C2(n20008), .A(n19990), .B(n19989), .ZN(
        P2_U3096) );
  AOI22_X1 U22988 ( .A1(n20004), .A2(n20320), .B1(n20319), .B2(n20003), .ZN(
        n19992) );
  AOI22_X1 U22989 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20005), .B1(
        n20036), .B2(n20321), .ZN(n19991) );
  OAI211_X1 U22990 ( .C1(n20324), .C2(n20008), .A(n19992), .B(n19991), .ZN(
        P2_U3097) );
  AOI22_X1 U22991 ( .A1(n20004), .A2(n20326), .B1(n20003), .B2(n20325), .ZN(
        n19994) );
  AOI22_X1 U22992 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20005), .B1(
        n20036), .B2(n20194), .ZN(n19993) );
  OAI211_X1 U22993 ( .C1(n20272), .C2(n20008), .A(n19994), .B(n19993), .ZN(
        P2_U3098) );
  AOI22_X1 U22994 ( .A1(n20004), .A2(n20332), .B1(n20003), .B2(n20331), .ZN(
        n19996) );
  AOI22_X1 U22995 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20005), .B1(
        n20036), .B2(n20333), .ZN(n19995) );
  OAI211_X1 U22996 ( .C1(n20336), .C2(n20008), .A(n19996), .B(n19995), .ZN(
        P2_U3099) );
  AOI22_X1 U22997 ( .A1(n20004), .A2(n20338), .B1(n20003), .B2(n20337), .ZN(
        n19998) );
  AOI22_X1 U22998 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20005), .B1(
        n20036), .B2(n20199), .ZN(n19997) );
  OAI211_X1 U22999 ( .C1(n20282), .C2(n20008), .A(n19998), .B(n19997), .ZN(
        P2_U3100) );
  AOI22_X1 U23000 ( .A1(n20004), .A2(n20344), .B1(n20003), .B2(n20343), .ZN(
        n20000) );
  AOI22_X1 U23001 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20005), .B1(
        n20036), .B2(n20202), .ZN(n19999) );
  OAI211_X1 U23002 ( .C1(n20284), .C2(n20008), .A(n20000), .B(n19999), .ZN(
        P2_U3101) );
  AOI22_X1 U23003 ( .A1(n20004), .A2(n20350), .B1(n20003), .B2(n20349), .ZN(
        n20002) );
  AOI22_X1 U23004 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20005), .B1(
        n20036), .B2(n20205), .ZN(n20001) );
  OAI211_X1 U23005 ( .C1(n20289), .C2(n20008), .A(n20002), .B(n20001), .ZN(
        P2_U3102) );
  AOI22_X1 U23006 ( .A1(n20004), .A2(n20359), .B1(n20003), .B2(n20357), .ZN(
        n20007) );
  AOI22_X1 U23007 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20005), .B1(
        n20036), .B2(n20361), .ZN(n20006) );
  OAI211_X1 U23008 ( .C1(n20367), .C2(n20008), .A(n20007), .B(n20006), .ZN(
        P2_U3103) );
  INV_X1 U23009 ( .A(n20009), .ZN(n20016) );
  OAI21_X1 U23010 ( .B1(n20010), .B2(n20458), .A(n20016), .ZN(n20013) );
  AND2_X1 U23011 ( .A1(n20011), .A2(n20253), .ZN(n20012) );
  INV_X1 U23012 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n21514) );
  OAI21_X1 U23013 ( .B1(n20014), .B2(n9805), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20015) );
  AOI22_X1 U23014 ( .A1(n20035), .A2(n20307), .B1(n9805), .B2(n20306), .ZN(
        n20019) );
  INV_X1 U23015 ( .A(n20072), .ZN(n20026) );
  AOI22_X1 U23016 ( .A1(n20026), .A2(n20189), .B1(n20036), .B2(n20315), .ZN(
        n20018) );
  OAI211_X1 U23017 ( .C1(n20030), .C2(n21514), .A(n20019), .B(n20018), .ZN(
        P2_U3104) );
  AOI22_X1 U23018 ( .A1(n20035), .A2(n20320), .B1(n9805), .B2(n20319), .ZN(
        n20021) );
  AOI22_X1 U23019 ( .A1(n20026), .A2(n20321), .B1(n20036), .B2(n20226), .ZN(
        n20020) );
  OAI211_X1 U23020 ( .C1(n20030), .C2(n10798), .A(n20021), .B(n20020), .ZN(
        P2_U3105) );
  AOI22_X1 U23021 ( .A1(n20035), .A2(n20326), .B1(n9805), .B2(n20325), .ZN(
        n20023) );
  AOI22_X1 U23022 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20037), .B1(
        n20036), .B2(n20327), .ZN(n20022) );
  OAI211_X1 U23023 ( .C1(n20330), .C2(n20072), .A(n20023), .B(n20022), .ZN(
        P2_U3106) );
  AOI22_X1 U23024 ( .A1(n20035), .A2(n20332), .B1(n9805), .B2(n20331), .ZN(
        n20025) );
  AOI22_X1 U23025 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20037), .B1(
        n20036), .B2(n20231), .ZN(n20024) );
  OAI211_X1 U23026 ( .C1(n20274), .C2(n20072), .A(n20025), .B(n20024), .ZN(
        P2_U3107) );
  AOI22_X1 U23027 ( .A1(n20035), .A2(n20338), .B1(n9805), .B2(n20337), .ZN(
        n20028) );
  AOI22_X1 U23028 ( .A1(n20026), .A2(n20199), .B1(n20036), .B2(n20339), .ZN(
        n20027) );
  OAI211_X1 U23029 ( .C1(n20030), .C2(n20029), .A(n20028), .B(n20027), .ZN(
        P2_U3108) );
  AOI22_X1 U23030 ( .A1(n20035), .A2(n20344), .B1(n9805), .B2(n20343), .ZN(
        n20032) );
  AOI22_X1 U23031 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20037), .B1(
        n20036), .B2(n20345), .ZN(n20031) );
  OAI211_X1 U23032 ( .C1(n20348), .C2(n20072), .A(n20032), .B(n20031), .ZN(
        P2_U3109) );
  AOI22_X1 U23033 ( .A1(n20035), .A2(n20350), .B1(n9805), .B2(n20349), .ZN(
        n20034) );
  AOI22_X1 U23034 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20037), .B1(
        n20036), .B2(n20351), .ZN(n20033) );
  OAI211_X1 U23035 ( .C1(n20356), .C2(n20072), .A(n20034), .B(n20033), .ZN(
        P2_U3110) );
  AOI22_X1 U23036 ( .A1(n20035), .A2(n20359), .B1(n9805), .B2(n20357), .ZN(
        n20039) );
  AOI22_X1 U23037 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20037), .B1(
        n20036), .B2(n20241), .ZN(n20038) );
  OAI211_X1 U23038 ( .C1(n20295), .C2(n20072), .A(n20039), .B(n20038), .ZN(
        P2_U3111) );
  NOR2_X1 U23039 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20121), .ZN(
        n20086) );
  AND2_X1 U23040 ( .A1(n20086), .A2(n20248), .ZN(n20047) );
  INV_X1 U23041 ( .A(n20047), .ZN(n20071) );
  OAI22_X1 U23042 ( .A1(n20072), .A2(n20262), .B1(n20071), .B2(n20249), .ZN(
        n20040) );
  INV_X1 U23043 ( .A(n20040), .ZN(n20052) );
  NAND2_X1 U23044 ( .A1(n20111), .A2(n20072), .ZN(n20041) );
  AOI21_X1 U23045 ( .B1(n20041), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20252), 
        .ZN(n20046) );
  INV_X1 U23046 ( .A(n20042), .ZN(n20048) );
  OAI21_X1 U23047 ( .B1(n20048), .B2(n20463), .A(n20304), .ZN(n20043) );
  AOI21_X1 U23048 ( .B1(n20046), .B2(n20044), .A(n20043), .ZN(n20045) );
  OAI21_X2 U23049 ( .B1(n20045), .B2(n20047), .A(n20253), .ZN(n20075) );
  OAI21_X1 U23050 ( .B1(n9805), .B2(n20047), .A(n20046), .ZN(n20050) );
  OAI21_X1 U23051 ( .B1(n20048), .B2(n20047), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20049) );
  AOI22_X1 U23052 ( .A1(n20075), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n20307), .B2(n20074), .ZN(n20051) );
  OAI211_X1 U23053 ( .C1(n20318), .C2(n20111), .A(n20052), .B(n20051), .ZN(
        P2_U3112) );
  OAI22_X1 U23054 ( .A1(n20111), .A2(n20264), .B1(n20071), .B2(n20263), .ZN(
        n20053) );
  INV_X1 U23055 ( .A(n20053), .ZN(n20055) );
  AOI22_X1 U23056 ( .A1(n20075), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n20320), .B2(n20074), .ZN(n20054) );
  OAI211_X1 U23057 ( .C1(n20324), .C2(n20072), .A(n20055), .B(n20054), .ZN(
        P2_U3113) );
  OAI22_X1 U23058 ( .A1(n20072), .A2(n20272), .B1(n20071), .B2(n20268), .ZN(
        n20056) );
  INV_X1 U23059 ( .A(n20056), .ZN(n20058) );
  AOI22_X1 U23060 ( .A1(n20075), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n20326), .B2(n20074), .ZN(n20057) );
  OAI211_X1 U23061 ( .C1(n20330), .C2(n20111), .A(n20058), .B(n20057), .ZN(
        P2_U3114) );
  OAI22_X1 U23062 ( .A1(n20072), .A2(n20336), .B1(n20071), .B2(n20273), .ZN(
        n20059) );
  INV_X1 U23063 ( .A(n20059), .ZN(n20061) );
  AOI22_X1 U23064 ( .A1(n20075), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n20332), .B2(n20074), .ZN(n20060) );
  OAI211_X1 U23065 ( .C1(n20274), .C2(n20111), .A(n20061), .B(n20060), .ZN(
        P2_U3115) );
  OAI22_X1 U23066 ( .A1(n20111), .A2(n20342), .B1(n20071), .B2(n20278), .ZN(
        n20062) );
  INV_X1 U23067 ( .A(n20062), .ZN(n20064) );
  AOI22_X1 U23068 ( .A1(n20075), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n20338), .B2(n20074), .ZN(n20063) );
  OAI211_X1 U23069 ( .C1(n20282), .C2(n20072), .A(n20064), .B(n20063), .ZN(
        P2_U3116) );
  OAI22_X1 U23070 ( .A1(n20072), .A2(n20284), .B1(n20071), .B2(n20283), .ZN(
        n20065) );
  INV_X1 U23071 ( .A(n20065), .ZN(n20067) );
  AOI22_X1 U23072 ( .A1(n20075), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n20344), .B2(n20074), .ZN(n20066) );
  OAI211_X1 U23073 ( .C1(n20348), .C2(n20111), .A(n20067), .B(n20066), .ZN(
        P2_U3117) );
  OAI22_X1 U23074 ( .A1(n20072), .A2(n20289), .B1(n20071), .B2(n20288), .ZN(
        n20068) );
  INV_X1 U23075 ( .A(n20068), .ZN(n20070) );
  AOI22_X1 U23076 ( .A1(n20075), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n20350), .B2(n20074), .ZN(n20069) );
  OAI211_X1 U23077 ( .C1(n20356), .C2(n20111), .A(n20070), .B(n20069), .ZN(
        P2_U3118) );
  OAI22_X1 U23078 ( .A1(n20072), .A2(n20367), .B1(n20071), .B2(n20293), .ZN(
        n20073) );
  INV_X1 U23079 ( .A(n20073), .ZN(n20077) );
  AOI22_X1 U23080 ( .A1(n20075), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n20359), .B2(n20074), .ZN(n20076) );
  OAI211_X1 U23081 ( .C1(n20295), .C2(n20111), .A(n20077), .B(n20076), .ZN(
        P2_U3119) );
  NAND2_X1 U23082 ( .A1(n20312), .A2(n20078), .ZN(n20087) );
  INV_X1 U23083 ( .A(n20086), .ZN(n20079) );
  NAND2_X1 U23084 ( .A1(n20087), .A2(n20079), .ZN(n20084) );
  OR2_X1 U23085 ( .A1(n20088), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20082) );
  AND2_X1 U23086 ( .A1(n20080), .A2(n20117), .ZN(n20125) );
  NOR2_X1 U23087 ( .A1(n20125), .A2(n20463), .ZN(n20081) );
  AOI21_X1 U23088 ( .B1(n20082), .B2(n20081), .A(n20309), .ZN(n20083) );
  INV_X1 U23089 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n20094) );
  INV_X1 U23090 ( .A(n20125), .ZN(n20110) );
  OAI22_X1 U23091 ( .A1(n20111), .A2(n20262), .B1(n20249), .B2(n20110), .ZN(
        n20085) );
  INV_X1 U23092 ( .A(n20085), .ZN(n20093) );
  NAND3_X1 U23093 ( .A1(n20087), .A2(n20086), .A3(n20463), .ZN(n20090) );
  OAI21_X1 U23094 ( .B1(n10648), .B2(n20125), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20089) );
  AOI22_X1 U23095 ( .A1(n20307), .A2(n20113), .B1(n20147), .B2(n20189), .ZN(
        n20092) );
  OAI211_X1 U23096 ( .C1(n20095), .C2(n20094), .A(n20093), .B(n20092), .ZN(
        P2_U3120) );
  AOI22_X1 U23097 ( .A1(n20147), .A2(n20321), .B1(n20319), .B2(n20125), .ZN(
        n20097) );
  AOI22_X1 U23098 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20114), .B1(
        n20320), .B2(n20113), .ZN(n20096) );
  OAI211_X1 U23099 ( .C1(n20324), .C2(n20111), .A(n20097), .B(n20096), .ZN(
        P2_U3121) );
  OAI22_X1 U23100 ( .A1(n20111), .A2(n20272), .B1(n20110), .B2(n20268), .ZN(
        n20098) );
  INV_X1 U23101 ( .A(n20098), .ZN(n20100) );
  AOI22_X1 U23102 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20114), .B1(
        n20326), .B2(n20113), .ZN(n20099) );
  OAI211_X1 U23103 ( .C1(n20330), .C2(n20123), .A(n20100), .B(n20099), .ZN(
        P2_U3122) );
  OAI22_X1 U23104 ( .A1(n20111), .A2(n20336), .B1(n20110), .B2(n20273), .ZN(
        n20101) );
  INV_X1 U23105 ( .A(n20101), .ZN(n20103) );
  AOI22_X1 U23106 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20114), .B1(
        n20332), .B2(n20113), .ZN(n20102) );
  OAI211_X1 U23107 ( .C1(n20274), .C2(n20123), .A(n20103), .B(n20102), .ZN(
        P2_U3123) );
  AOI22_X1 U23108 ( .A1(n20147), .A2(n20199), .B1(n20337), .B2(n20125), .ZN(
        n20105) );
  AOI22_X1 U23109 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20114), .B1(
        n20338), .B2(n20113), .ZN(n20104) );
  OAI211_X1 U23110 ( .C1(n20282), .C2(n20111), .A(n20105), .B(n20104), .ZN(
        P2_U3124) );
  AOI22_X1 U23111 ( .A1(n20147), .A2(n20202), .B1(n20343), .B2(n20125), .ZN(
        n20107) );
  AOI22_X1 U23112 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20114), .B1(
        n20344), .B2(n20113), .ZN(n20106) );
  OAI211_X1 U23113 ( .C1(n20284), .C2(n20111), .A(n20107), .B(n20106), .ZN(
        P2_U3125) );
  AOI22_X1 U23114 ( .A1(n20147), .A2(n20205), .B1(n20349), .B2(n20125), .ZN(
        n20109) );
  AOI22_X1 U23115 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20114), .B1(
        n20350), .B2(n20113), .ZN(n20108) );
  OAI211_X1 U23116 ( .C1(n20289), .C2(n20111), .A(n20109), .B(n20108), .ZN(
        P2_U3126) );
  OAI22_X1 U23117 ( .A1(n20111), .A2(n20367), .B1(n20110), .B2(n20293), .ZN(
        n20112) );
  INV_X1 U23118 ( .A(n20112), .ZN(n20116) );
  AOI22_X1 U23119 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20114), .B1(
        n20359), .B2(n20113), .ZN(n20115) );
  OAI211_X1 U23120 ( .C1(n20295), .C2(n20123), .A(n20116), .B(n20115), .ZN(
        P2_U3127) );
  AND2_X1 U23121 ( .A1(n20118), .A2(n20117), .ZN(n20144) );
  OAI21_X1 U23122 ( .B1(n10789), .B2(n20144), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20119) );
  OAI21_X1 U23123 ( .B1(n20121), .B2(n20120), .A(n20119), .ZN(n20145) );
  AOI22_X1 U23124 ( .A1(n20145), .A2(n20307), .B1(n20306), .B2(n20144), .ZN(
        n20131) );
  AOI21_X1 U23125 ( .B1(n20123), .B2(n20175), .A(n20122), .ZN(n20124) );
  OAI21_X1 U23126 ( .B1(n20125), .B2(n20124), .A(n20304), .ZN(n20126) );
  AOI21_X1 U23127 ( .B1(n20127), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n20126), 
        .ZN(n20129) );
  OAI21_X1 U23128 ( .B1(n20129), .B2(n20144), .A(n20128), .ZN(n20146) );
  AOI22_X1 U23129 ( .A1(n20147), .A2(n20315), .B1(
        P2_INSTQUEUE_REG_10__0__SCAN_IN), .B2(n20146), .ZN(n20130) );
  OAI211_X1 U23130 ( .C1(n20318), .C2(n20175), .A(n20131), .B(n20130), .ZN(
        P2_U3128) );
  AOI22_X1 U23131 ( .A1(n20145), .A2(n20320), .B1(n20319), .B2(n20144), .ZN(
        n20133) );
  AOI22_X1 U23132 ( .A1(n20147), .A2(n20226), .B1(
        P2_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n20146), .ZN(n20132) );
  OAI211_X1 U23133 ( .C1(n20264), .C2(n20175), .A(n20133), .B(n20132), .ZN(
        P2_U3129) );
  AOI22_X1 U23134 ( .A1(n20145), .A2(n20326), .B1(n20325), .B2(n20144), .ZN(
        n20135) );
  AOI22_X1 U23135 ( .A1(n20147), .A2(n20327), .B1(
        P2_INSTQUEUE_REG_10__2__SCAN_IN), .B2(n20146), .ZN(n20134) );
  OAI211_X1 U23136 ( .C1(n20330), .C2(n20175), .A(n20135), .B(n20134), .ZN(
        P2_U3130) );
  AOI22_X1 U23137 ( .A1(n20145), .A2(n20332), .B1(n20331), .B2(n20144), .ZN(
        n20137) );
  AOI22_X1 U23138 ( .A1(n20147), .A2(n20231), .B1(
        P2_INSTQUEUE_REG_10__3__SCAN_IN), .B2(n20146), .ZN(n20136) );
  OAI211_X1 U23139 ( .C1(n20274), .C2(n20175), .A(n20137), .B(n20136), .ZN(
        P2_U3131) );
  AOI22_X1 U23140 ( .A1(n20145), .A2(n20338), .B1(n20337), .B2(n20144), .ZN(
        n20139) );
  AOI22_X1 U23141 ( .A1(n20147), .A2(n20339), .B1(
        P2_INSTQUEUE_REG_10__4__SCAN_IN), .B2(n20146), .ZN(n20138) );
  OAI211_X1 U23142 ( .C1(n20342), .C2(n20175), .A(n20139), .B(n20138), .ZN(
        P2_U3132) );
  AOI22_X1 U23143 ( .A1(n20145), .A2(n20344), .B1(n20343), .B2(n20144), .ZN(
        n20141) );
  AOI22_X1 U23144 ( .A1(n20147), .A2(n20345), .B1(
        P2_INSTQUEUE_REG_10__5__SCAN_IN), .B2(n20146), .ZN(n20140) );
  OAI211_X1 U23145 ( .C1(n20348), .C2(n20175), .A(n20141), .B(n20140), .ZN(
        P2_U3133) );
  AOI22_X1 U23146 ( .A1(n20145), .A2(n20350), .B1(n20349), .B2(n20144), .ZN(
        n20143) );
  AOI22_X1 U23147 ( .A1(n20147), .A2(n20351), .B1(
        P2_INSTQUEUE_REG_10__6__SCAN_IN), .B2(n20146), .ZN(n20142) );
  OAI211_X1 U23148 ( .C1(n20356), .C2(n20175), .A(n20143), .B(n20142), .ZN(
        P2_U3134) );
  AOI22_X1 U23149 ( .A1(n20145), .A2(n20359), .B1(n20357), .B2(n20144), .ZN(
        n20149) );
  AOI22_X1 U23150 ( .A1(n20147), .A2(n20241), .B1(
        P2_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n20146), .ZN(n20148) );
  OAI211_X1 U23151 ( .C1(n20295), .C2(n20175), .A(n20149), .B(n20148), .ZN(
        P2_U3135) );
  INV_X1 U23152 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n20153) );
  NOR2_X1 U23153 ( .A1(n20249), .A2(n20169), .ZN(n20150) );
  AOI21_X1 U23154 ( .B1(n20171), .B2(n20307), .A(n20150), .ZN(n20152) );
  AOI22_X1 U23155 ( .A1(n20166), .A2(n20315), .B1(n20184), .B2(n20189), .ZN(
        n20151) );
  OAI211_X1 U23156 ( .C1(n20154), .C2(n20153), .A(n20152), .B(n20151), .ZN(
        P2_U3136) );
  NOR2_X1 U23157 ( .A1(n20268), .A2(n20169), .ZN(n20155) );
  AOI21_X1 U23158 ( .B1(n20171), .B2(n20326), .A(n20155), .ZN(n20157) );
  AOI22_X1 U23159 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20172), .B1(
        n20166), .B2(n20327), .ZN(n20156) );
  OAI211_X1 U23160 ( .C1(n20330), .C2(n20213), .A(n20157), .B(n20156), .ZN(
        P2_U3138) );
  NOR2_X1 U23161 ( .A1(n20273), .A2(n20169), .ZN(n20158) );
  AOI21_X1 U23162 ( .B1(n20171), .B2(n20332), .A(n20158), .ZN(n20160) );
  AOI22_X1 U23163 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20172), .B1(
        n20184), .B2(n20333), .ZN(n20159) );
  OAI211_X1 U23164 ( .C1(n20336), .C2(n20175), .A(n20160), .B(n20159), .ZN(
        P2_U3139) );
  AOI22_X1 U23165 ( .A1(n20171), .A2(n20338), .B1(n20165), .B2(n20337), .ZN(
        n20162) );
  AOI22_X1 U23166 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20172), .B1(
        n20166), .B2(n20339), .ZN(n20161) );
  OAI211_X1 U23167 ( .C1(n20342), .C2(n20213), .A(n20162), .B(n20161), .ZN(
        P2_U3140) );
  AOI22_X1 U23168 ( .A1(n20171), .A2(n20344), .B1(n20165), .B2(n20343), .ZN(
        n20164) );
  AOI22_X1 U23169 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20172), .B1(
        n20166), .B2(n20345), .ZN(n20163) );
  OAI211_X1 U23170 ( .C1(n20348), .C2(n20213), .A(n20164), .B(n20163), .ZN(
        P2_U3141) );
  AOI22_X1 U23171 ( .A1(n20171), .A2(n20350), .B1(n20165), .B2(n20349), .ZN(
        n20168) );
  AOI22_X1 U23172 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20172), .B1(
        n20166), .B2(n20351), .ZN(n20167) );
  OAI211_X1 U23173 ( .C1(n20356), .C2(n20213), .A(n20168), .B(n20167), .ZN(
        P2_U3142) );
  NOR2_X1 U23174 ( .A1(n20293), .A2(n20169), .ZN(n20170) );
  AOI21_X1 U23175 ( .B1(n20171), .B2(n20359), .A(n20170), .ZN(n20174) );
  AOI22_X1 U23176 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20172), .B1(
        n20184), .B2(n20361), .ZN(n20173) );
  OAI211_X1 U23177 ( .C1(n20367), .C2(n20175), .A(n20174), .B(n20173), .ZN(
        P2_U3143) );
  INV_X1 U23178 ( .A(n20183), .ZN(n20177) );
  AND2_X1 U23179 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20247) );
  NAND2_X1 U23180 ( .A1(n20247), .A2(n20176), .ZN(n20218) );
  NOR2_X1 U23181 ( .A1(n20218), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20208) );
  OAI21_X1 U23182 ( .B1(n20177), .B2(n20208), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20182) );
  NAND3_X1 U23183 ( .A1(n20180), .A2(n20179), .A3(n20178), .ZN(n20181) );
  NAND2_X1 U23184 ( .A1(n20182), .A2(n20181), .ZN(n20209) );
  AOI22_X1 U23185 ( .A1(n20209), .A2(n20307), .B1(n20208), .B2(n20306), .ZN(
        n20191) );
  AOI21_X1 U23186 ( .B1(n20183), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20188) );
  OAI21_X1 U23187 ( .B1(n20184), .B2(n20242), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20185) );
  OAI21_X1 U23188 ( .B1(n20471), .B2(n20186), .A(n20185), .ZN(n20187) );
  AOI22_X1 U23189 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20210), .B1(
        n20242), .B2(n20189), .ZN(n20190) );
  OAI211_X1 U23190 ( .C1(n20262), .C2(n20213), .A(n20191), .B(n20190), .ZN(
        P2_U3144) );
  AOI22_X1 U23191 ( .A1(n20209), .A2(n20320), .B1(n20208), .B2(n20319), .ZN(
        n20193) );
  AOI22_X1 U23192 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20210), .B1(
        n20242), .B2(n20321), .ZN(n20192) );
  OAI211_X1 U23193 ( .C1(n20324), .C2(n20213), .A(n20193), .B(n20192), .ZN(
        P2_U3145) );
  AOI22_X1 U23194 ( .A1(n20209), .A2(n20326), .B1(n20208), .B2(n20325), .ZN(
        n20196) );
  AOI22_X1 U23195 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20210), .B1(
        n20242), .B2(n20194), .ZN(n20195) );
  OAI211_X1 U23196 ( .C1(n20272), .C2(n20213), .A(n20196), .B(n20195), .ZN(
        P2_U3146) );
  AOI22_X1 U23197 ( .A1(n20209), .A2(n20332), .B1(n20208), .B2(n20331), .ZN(
        n20198) );
  AOI22_X1 U23198 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20210), .B1(
        n20242), .B2(n20333), .ZN(n20197) );
  OAI211_X1 U23199 ( .C1(n20336), .C2(n20213), .A(n20198), .B(n20197), .ZN(
        P2_U3147) );
  AOI22_X1 U23200 ( .A1(n20209), .A2(n20338), .B1(n20208), .B2(n20337), .ZN(
        n20201) );
  AOI22_X1 U23201 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20210), .B1(
        n20242), .B2(n20199), .ZN(n20200) );
  OAI211_X1 U23202 ( .C1(n20282), .C2(n20213), .A(n20201), .B(n20200), .ZN(
        P2_U3148) );
  AOI22_X1 U23203 ( .A1(n20209), .A2(n20344), .B1(n20208), .B2(n20343), .ZN(
        n20204) );
  AOI22_X1 U23204 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20210), .B1(
        n20242), .B2(n20202), .ZN(n20203) );
  OAI211_X1 U23205 ( .C1(n20284), .C2(n20213), .A(n20204), .B(n20203), .ZN(
        P2_U3149) );
  AOI22_X1 U23206 ( .A1(n20209), .A2(n20350), .B1(n20208), .B2(n20349), .ZN(
        n20207) );
  AOI22_X1 U23207 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20210), .B1(
        n20242), .B2(n20205), .ZN(n20206) );
  OAI211_X1 U23208 ( .C1(n20289), .C2(n20213), .A(n20207), .B(n20206), .ZN(
        P2_U3150) );
  AOI22_X1 U23209 ( .A1(n20209), .A2(n20359), .B1(n20208), .B2(n20357), .ZN(
        n20212) );
  AOI22_X1 U23210 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20210), .B1(
        n20242), .B2(n20361), .ZN(n20211) );
  OAI211_X1 U23211 ( .C1(n20367), .C2(n20213), .A(n20212), .B(n20211), .ZN(
        P2_U3151) );
  OR2_X2 U23212 ( .A1(n20214), .A2(n20219), .ZN(n20301) );
  NOR2_X1 U23213 ( .A1(n20218), .A2(n20248), .ZN(n20255) );
  NOR2_X1 U23214 ( .A1(n20255), .A2(n20302), .ZN(n20215) );
  NAND2_X1 U23215 ( .A1(n20216), .A2(n20215), .ZN(n20222) );
  OAI21_X1 U23216 ( .B1(n20218), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20302), 
        .ZN(n20217) );
  AOI22_X1 U23217 ( .A1(n20240), .A2(n20307), .B1(n20255), .B2(n20306), .ZN(
        n20225) );
  INV_X1 U23218 ( .A(n20312), .ZN(n20220) );
  OAI21_X1 U23219 ( .B1(n20220), .B2(n20219), .A(n20218), .ZN(n20223) );
  OR2_X1 U23220 ( .A1(n20255), .A2(n20304), .ZN(n20221) );
  NAND4_X1 U23221 ( .A1(n20223), .A2(n20253), .A3(n20222), .A4(n20221), .ZN(
        n20243) );
  AOI22_X1 U23222 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20243), .B1(
        n20242), .B2(n20315), .ZN(n20224) );
  OAI211_X1 U23223 ( .C1(n20318), .C2(n20301), .A(n20225), .B(n20224), .ZN(
        P2_U3152) );
  AOI22_X1 U23224 ( .A1(n20240), .A2(n20320), .B1(n20319), .B2(n20255), .ZN(
        n20228) );
  AOI22_X1 U23225 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20243), .B1(
        n20242), .B2(n20226), .ZN(n20227) );
  OAI211_X1 U23226 ( .C1(n20264), .C2(n20301), .A(n20228), .B(n20227), .ZN(
        P2_U3153) );
  AOI22_X1 U23227 ( .A1(n20240), .A2(n20326), .B1(n20255), .B2(n20325), .ZN(
        n20230) );
  AOI22_X1 U23228 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20243), .B1(
        n20242), .B2(n20327), .ZN(n20229) );
  OAI211_X1 U23229 ( .C1(n20330), .C2(n20301), .A(n20230), .B(n20229), .ZN(
        P2_U3154) );
  AOI22_X1 U23230 ( .A1(n20240), .A2(n20332), .B1(n20255), .B2(n20331), .ZN(
        n20233) );
  AOI22_X1 U23231 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20243), .B1(
        n20242), .B2(n20231), .ZN(n20232) );
  OAI211_X1 U23232 ( .C1(n20274), .C2(n20301), .A(n20233), .B(n20232), .ZN(
        P2_U3155) );
  AOI22_X1 U23233 ( .A1(n20240), .A2(n20338), .B1(n20255), .B2(n20337), .ZN(
        n20235) );
  AOI22_X1 U23234 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20243), .B1(
        n20242), .B2(n20339), .ZN(n20234) );
  OAI211_X1 U23235 ( .C1(n20342), .C2(n20301), .A(n20235), .B(n20234), .ZN(
        P2_U3156) );
  AOI22_X1 U23236 ( .A1(n20240), .A2(n20344), .B1(n20255), .B2(n20343), .ZN(
        n20237) );
  AOI22_X1 U23237 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20243), .B1(
        n20242), .B2(n20345), .ZN(n20236) );
  OAI211_X1 U23238 ( .C1(n20348), .C2(n20301), .A(n20237), .B(n20236), .ZN(
        P2_U3157) );
  AOI22_X1 U23239 ( .A1(n20240), .A2(n20350), .B1(n20255), .B2(n20349), .ZN(
        n20239) );
  AOI22_X1 U23240 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20243), .B1(
        n20242), .B2(n20351), .ZN(n20238) );
  OAI211_X1 U23241 ( .C1(n20356), .C2(n20301), .A(n20239), .B(n20238), .ZN(
        P2_U3158) );
  AOI22_X1 U23242 ( .A1(n20240), .A2(n20359), .B1(n20255), .B2(n20357), .ZN(
        n20245) );
  AOI22_X1 U23243 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20243), .B1(
        n20242), .B2(n20241), .ZN(n20244) );
  OAI211_X1 U23244 ( .C1(n20295), .C2(n20301), .A(n20245), .B(n20244), .ZN(
        P2_U3159) );
  AND2_X1 U23245 ( .A1(n20247), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20314) );
  AND2_X1 U23246 ( .A1(n20314), .A2(n20248), .ZN(n20254) );
  INV_X1 U23247 ( .A(n20254), .ZN(n20294) );
  OAI22_X1 U23248 ( .A1(n20366), .A2(n20318), .B1(n20294), .B2(n20249), .ZN(
        n20250) );
  INV_X1 U23249 ( .A(n20250), .ZN(n20261) );
  INV_X1 U23250 ( .A(n20301), .ZN(n20251) );
  OAI21_X2 U23251 ( .B1(n9685), .B2(n20254), .A(n20253), .ZN(n20298) );
  INV_X1 U23252 ( .A(n20255), .ZN(n20258) );
  NOR2_X1 U23253 ( .A1(n20256), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20257) );
  AOI22_X1 U23254 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20298), .B1(
        n20307), .B2(n20297), .ZN(n20260) );
  OAI211_X1 U23255 ( .C1(n20262), .C2(n20301), .A(n20261), .B(n20260), .ZN(
        P2_U3160) );
  OAI22_X1 U23256 ( .A1(n20366), .A2(n20264), .B1(n20263), .B2(n20294), .ZN(
        n20265) );
  INV_X1 U23257 ( .A(n20265), .ZN(n20267) );
  AOI22_X1 U23258 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20298), .B1(
        n20320), .B2(n20297), .ZN(n20266) );
  OAI211_X1 U23259 ( .C1(n20324), .C2(n20301), .A(n20267), .B(n20266), .ZN(
        P2_U3161) );
  OAI22_X1 U23260 ( .A1(n20366), .A2(n20330), .B1(n20294), .B2(n20268), .ZN(
        n20269) );
  INV_X1 U23261 ( .A(n20269), .ZN(n20271) );
  AOI22_X1 U23262 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20298), .B1(
        n20326), .B2(n20297), .ZN(n20270) );
  OAI211_X1 U23263 ( .C1(n20272), .C2(n20301), .A(n20271), .B(n20270), .ZN(
        P2_U3162) );
  OAI22_X1 U23264 ( .A1(n20366), .A2(n20274), .B1(n20294), .B2(n20273), .ZN(
        n20275) );
  INV_X1 U23265 ( .A(n20275), .ZN(n20277) );
  AOI22_X1 U23266 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20298), .B1(
        n20332), .B2(n20297), .ZN(n20276) );
  OAI211_X1 U23267 ( .C1(n20336), .C2(n20301), .A(n20277), .B(n20276), .ZN(
        P2_U3163) );
  OAI22_X1 U23268 ( .A1(n20366), .A2(n20342), .B1(n20294), .B2(n20278), .ZN(
        n20279) );
  INV_X1 U23269 ( .A(n20279), .ZN(n20281) );
  AOI22_X1 U23270 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20298), .B1(
        n20338), .B2(n20297), .ZN(n20280) );
  OAI211_X1 U23271 ( .C1(n20282), .C2(n20301), .A(n20281), .B(n20280), .ZN(
        P2_U3164) );
  OAI22_X1 U23272 ( .A1(n20301), .A2(n20284), .B1(n20294), .B2(n20283), .ZN(
        n20285) );
  INV_X1 U23273 ( .A(n20285), .ZN(n20287) );
  AOI22_X1 U23274 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20298), .B1(
        n20344), .B2(n20297), .ZN(n20286) );
  OAI211_X1 U23275 ( .C1(n20348), .C2(n20366), .A(n20287), .B(n20286), .ZN(
        P2_U3165) );
  OAI22_X1 U23276 ( .A1(n20301), .A2(n20289), .B1(n20294), .B2(n20288), .ZN(
        n20290) );
  INV_X1 U23277 ( .A(n20290), .ZN(n20292) );
  AOI22_X1 U23278 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20298), .B1(
        n20350), .B2(n20297), .ZN(n20291) );
  OAI211_X1 U23279 ( .C1(n20356), .C2(n20366), .A(n20292), .B(n20291), .ZN(
        P2_U3166) );
  OAI22_X1 U23280 ( .A1(n20366), .A2(n20295), .B1(n20294), .B2(n20293), .ZN(
        n20296) );
  INV_X1 U23281 ( .A(n20296), .ZN(n20300) );
  AOI22_X1 U23282 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20298), .B1(
        n20359), .B2(n20297), .ZN(n20299) );
  OAI211_X1 U23283 ( .C1(n20367), .C2(n20301), .A(n20300), .B(n20299), .ZN(
        P2_U3167) );
  NOR3_X1 U23284 ( .A1(n20303), .A2(n20358), .A3(n20302), .ZN(n20308) );
  AOI21_X1 U23285 ( .B1(n20314), .B2(n20304), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20305) );
  AOI22_X1 U23286 ( .A1(n20360), .A2(n20307), .B1(n20358), .B2(n20306), .ZN(
        n20317) );
  AOI211_X1 U23287 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20310), .A(n20309), 
        .B(n20308), .ZN(n20311) );
  OAI221_X1 U23288 ( .B1(n20314), .B2(n20313), .C1(n20314), .C2(n20312), .A(
        n20311), .ZN(n20363) );
  AOI22_X1 U23289 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20363), .B1(
        n20352), .B2(n20315), .ZN(n20316) );
  OAI211_X1 U23290 ( .C1(n20318), .C2(n20355), .A(n20317), .B(n20316), .ZN(
        P2_U3168) );
  AOI22_X1 U23291 ( .A1(n20360), .A2(n20320), .B1(n20319), .B2(n20358), .ZN(
        n20323) );
  AOI22_X1 U23292 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20363), .B1(
        n20362), .B2(n20321), .ZN(n20322) );
  OAI211_X1 U23293 ( .C1(n20324), .C2(n20366), .A(n20323), .B(n20322), .ZN(
        P2_U3169) );
  AOI22_X1 U23294 ( .A1(n20360), .A2(n20326), .B1(n20358), .B2(n20325), .ZN(
        n20329) );
  AOI22_X1 U23295 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20363), .B1(
        n20352), .B2(n20327), .ZN(n20328) );
  OAI211_X1 U23296 ( .C1(n20330), .C2(n20355), .A(n20329), .B(n20328), .ZN(
        P2_U3170) );
  AOI22_X1 U23297 ( .A1(n20360), .A2(n20332), .B1(n20358), .B2(n20331), .ZN(
        n20335) );
  AOI22_X1 U23298 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20363), .B1(
        n20362), .B2(n20333), .ZN(n20334) );
  OAI211_X1 U23299 ( .C1(n20336), .C2(n20366), .A(n20335), .B(n20334), .ZN(
        P2_U3171) );
  AOI22_X1 U23300 ( .A1(n20360), .A2(n20338), .B1(n20358), .B2(n20337), .ZN(
        n20341) );
  AOI22_X1 U23301 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20363), .B1(
        n20352), .B2(n20339), .ZN(n20340) );
  OAI211_X1 U23302 ( .C1(n20342), .C2(n20355), .A(n20341), .B(n20340), .ZN(
        P2_U3172) );
  AOI22_X1 U23303 ( .A1(n20360), .A2(n20344), .B1(n20358), .B2(n20343), .ZN(
        n20347) );
  AOI22_X1 U23304 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20363), .B1(
        n20352), .B2(n20345), .ZN(n20346) );
  OAI211_X1 U23305 ( .C1(n20348), .C2(n20355), .A(n20347), .B(n20346), .ZN(
        P2_U3173) );
  AOI22_X1 U23306 ( .A1(n20360), .A2(n20350), .B1(n20358), .B2(n20349), .ZN(
        n20354) );
  AOI22_X1 U23307 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20363), .B1(
        n20352), .B2(n20351), .ZN(n20353) );
  OAI211_X1 U23308 ( .C1(n20356), .C2(n20355), .A(n20354), .B(n20353), .ZN(
        P2_U3174) );
  AOI22_X1 U23309 ( .A1(n20360), .A2(n20359), .B1(n20358), .B2(n20357), .ZN(
        n20365) );
  AOI22_X1 U23310 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20363), .B1(
        n20362), .B2(n20361), .ZN(n20364) );
  OAI211_X1 U23311 ( .C1(n20367), .C2(n20366), .A(n20365), .B(n20364), .ZN(
        P2_U3175) );
  INV_X1 U23312 ( .A(P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n21506) );
  NOR2_X1 U23313 ( .A1(n21506), .A2(n20456), .ZN(P2_U3179) );
  AND2_X1 U23314 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20368), .ZN(
        P2_U3180) );
  AND2_X1 U23315 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20368), .ZN(
        P2_U3181) );
  AND2_X1 U23316 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20368), .ZN(
        P2_U3182) );
  AND2_X1 U23317 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20368), .ZN(
        P2_U3183) );
  AND2_X1 U23318 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20368), .ZN(
        P2_U3184) );
  AND2_X1 U23319 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20368), .ZN(
        P2_U3185) );
  AND2_X1 U23320 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20368), .ZN(
        P2_U3186) );
  AND2_X1 U23321 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20368), .ZN(
        P2_U3187) );
  AND2_X1 U23322 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20368), .ZN(
        P2_U3188) );
  AND2_X1 U23323 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20368), .ZN(
        P2_U3189) );
  AND2_X1 U23324 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20368), .ZN(
        P2_U3190) );
  AND2_X1 U23325 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20368), .ZN(
        P2_U3191) );
  AND2_X1 U23326 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20368), .ZN(
        P2_U3192) );
  AND2_X1 U23327 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20368), .ZN(
        P2_U3193) );
  AND2_X1 U23328 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20368), .ZN(
        P2_U3194) );
  AND2_X1 U23329 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20368), .ZN(
        P2_U3195) );
  AND2_X1 U23330 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20368), .ZN(
        P2_U3196) );
  AND2_X1 U23331 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20368), .ZN(
        P2_U3197) );
  AND2_X1 U23332 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20368), .ZN(
        P2_U3198) );
  AND2_X1 U23333 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20368), .ZN(
        P2_U3199) );
  AND2_X1 U23334 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20368), .ZN(
        P2_U3200) );
  AND2_X1 U23335 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20368), .ZN(P2_U3201) );
  AND2_X1 U23336 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20368), .ZN(P2_U3202) );
  AND2_X1 U23337 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20368), .ZN(P2_U3203) );
  AND2_X1 U23338 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20368), .ZN(P2_U3204) );
  AND2_X1 U23339 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20368), .ZN(P2_U3205) );
  AND2_X1 U23340 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20368), .ZN(P2_U3206) );
  AND2_X1 U23341 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20368), .ZN(P2_U3207) );
  AND2_X1 U23342 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20368), .ZN(P2_U3208) );
  NOR2_X1 U23343 ( .A1(n20370), .A2(n20369), .ZN(n20382) );
  INV_X1 U23344 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20386) );
  OR3_X1 U23345 ( .A1(n20382), .A2(n20386), .A3(n20385), .ZN(n20372) );
  INV_X2 U23346 ( .A(n20483), .ZN(n20446) );
  AOI211_X1 U23347 ( .C1(n21300), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n20383), .B(n20446), .ZN(n20371) );
  INV_X1 U23348 ( .A(NA), .ZN(n21307) );
  NOR2_X1 U23349 ( .A1(n21307), .A2(n20374), .ZN(n20390) );
  AOI211_X1 U23350 ( .C1(n20391), .C2(n20372), .A(n20371), .B(n20390), .ZN(
        n20373) );
  INV_X1 U23351 ( .A(n20373), .ZN(P2_U3209) );
  AOI21_X1 U23352 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21300), .A(n20391), 
        .ZN(n20379) );
  NOR2_X1 U23353 ( .A1(n20386), .A2(n20379), .ZN(n20375) );
  AOI21_X1 U23354 ( .B1(n20375), .B2(n20374), .A(n20382), .ZN(n20377) );
  OAI211_X1 U23355 ( .C1(n21300), .C2(n20378), .A(n20377), .B(n20376), .ZN(
        P2_U3210) );
  AOI21_X1 U23356 ( .B1(n20381), .B2(n20380), .A(n20379), .ZN(n20389) );
  AOI22_X1 U23357 ( .A1(n20386), .A2(n20383), .B1(n21307), .B2(n20382), .ZN(
        n20384) );
  AOI211_X1 U23358 ( .C1(n20386), .C2(n21300), .A(n20385), .B(n20384), .ZN(
        n20387) );
  INV_X1 U23359 ( .A(n20387), .ZN(n20388) );
  OAI21_X1 U23360 ( .B1(n20390), .B2(n20389), .A(n20388), .ZN(P2_U3211) );
  INV_X1 U23361 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20394) );
  NAND2_X1 U23362 ( .A1(n20446), .A2(n20391), .ZN(n20449) );
  CLKBUF_X1 U23363 ( .A(n20449), .Z(n20443) );
  OAI222_X1 U23364 ( .A1(n20444), .A2(n10612), .B1(n20392), .B2(n20446), .C1(
        n20394), .C2(n20443), .ZN(P2_U3212) );
  OAI222_X1 U23365 ( .A1(n20444), .A2(n20394), .B1(n20393), .B2(n20446), .C1(
        n20396), .C2(n20443), .ZN(P2_U3213) );
  OAI222_X1 U23366 ( .A1(n20444), .A2(n20396), .B1(n20395), .B2(n20446), .C1(
        n16417), .C2(n20443), .ZN(P2_U3214) );
  INV_X1 U23367 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n20398) );
  OAI222_X1 U23368 ( .A1(n20443), .A2(n20398), .B1(n20397), .B2(n20446), .C1(
        n16417), .C2(n20444), .ZN(P2_U3215) );
  OAI222_X1 U23369 ( .A1(n20449), .A2(n20400), .B1(n20399), .B2(n20446), .C1(
        n20398), .C2(n20444), .ZN(P2_U3216) );
  OAI222_X1 U23370 ( .A1(n20449), .A2(n20402), .B1(n20401), .B2(n20446), .C1(
        n20400), .C2(n20444), .ZN(P2_U3217) );
  INV_X1 U23371 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20404) );
  OAI222_X1 U23372 ( .A1(n20449), .A2(n20404), .B1(n20403), .B2(n20446), .C1(
        n20402), .C2(n20444), .ZN(P2_U3218) );
  INV_X1 U23373 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20406) );
  OAI222_X1 U23374 ( .A1(n20449), .A2(n20406), .B1(n20405), .B2(n20446), .C1(
        n20404), .C2(n20444), .ZN(P2_U3219) );
  OAI222_X1 U23375 ( .A1(n20449), .A2(n12372), .B1(n20407), .B2(n20446), .C1(
        n20406), .C2(n20444), .ZN(P2_U3220) );
  OAI222_X1 U23376 ( .A1(n20449), .A2(n20409), .B1(n20408), .B2(n20446), .C1(
        n12372), .C2(n20444), .ZN(P2_U3221) );
  OAI222_X1 U23377 ( .A1(n20443), .A2(n20411), .B1(n20410), .B2(n20446), .C1(
        n20409), .C2(n20444), .ZN(P2_U3222) );
  OAI222_X1 U23378 ( .A1(n20443), .A2(n20413), .B1(n20412), .B2(n20446), .C1(
        n20411), .C2(n20444), .ZN(P2_U3223) );
  OAI222_X1 U23379 ( .A1(n20443), .A2(n12434), .B1(n20414), .B2(n20446), .C1(
        n20413), .C2(n20444), .ZN(P2_U3224) );
  OAI222_X1 U23380 ( .A1(n20443), .A2(n20416), .B1(n20415), .B2(n20446), .C1(
        n12434), .C2(n20444), .ZN(P2_U3225) );
  OAI222_X1 U23381 ( .A1(n20443), .A2(n20418), .B1(n20417), .B2(n20446), .C1(
        n20416), .C2(n20444), .ZN(P2_U3226) );
  OAI222_X1 U23382 ( .A1(n20443), .A2(n20420), .B1(n20419), .B2(n20446), .C1(
        n20418), .C2(n20444), .ZN(P2_U3227) );
  OAI222_X1 U23383 ( .A1(n20443), .A2(n15751), .B1(n20421), .B2(n20446), .C1(
        n20420), .C2(n20444), .ZN(P2_U3228) );
  OAI222_X1 U23384 ( .A1(n20449), .A2(n20423), .B1(n20422), .B2(n20446), .C1(
        n15751), .C2(n20444), .ZN(P2_U3229) );
  OAI222_X1 U23385 ( .A1(n20449), .A2(n16236), .B1(n20424), .B2(n20446), .C1(
        n20423), .C2(n20444), .ZN(P2_U3230) );
  OAI222_X1 U23386 ( .A1(n20449), .A2(n20426), .B1(n20425), .B2(n20446), .C1(
        n16236), .C2(n20444), .ZN(P2_U3231) );
  OAI222_X1 U23387 ( .A1(n20449), .A2(n16221), .B1(n20427), .B2(n20446), .C1(
        n20426), .C2(n20444), .ZN(P2_U3232) );
  OAI222_X1 U23388 ( .A1(n20443), .A2(n20429), .B1(n20428), .B2(n20446), .C1(
        n16221), .C2(n20444), .ZN(P2_U3233) );
  OAI222_X1 U23389 ( .A1(n20443), .A2(n20431), .B1(n20430), .B2(n20446), .C1(
        n20429), .C2(n20444), .ZN(P2_U3234) );
  OAI222_X1 U23390 ( .A1(n20443), .A2(n20433), .B1(n20432), .B2(n20446), .C1(
        n20431), .C2(n20444), .ZN(P2_U3235) );
  INV_X1 U23391 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20435) );
  OAI222_X1 U23392 ( .A1(n20443), .A2(n20435), .B1(n20434), .B2(n20446), .C1(
        n20433), .C2(n20444), .ZN(P2_U3236) );
  OAI222_X1 U23393 ( .A1(n20443), .A2(n20438), .B1(n20436), .B2(n20446), .C1(
        n20435), .C2(n20444), .ZN(P2_U3237) );
  OAI222_X1 U23394 ( .A1(n20444), .A2(n20438), .B1(n20437), .B2(n20446), .C1(
        n20439), .C2(n20443), .ZN(P2_U3238) );
  OAI222_X1 U23395 ( .A1(n20443), .A2(n20441), .B1(n20440), .B2(n20446), .C1(
        n20439), .C2(n20444), .ZN(P2_U3239) );
  OAI222_X1 U23396 ( .A1(n20443), .A2(n20445), .B1(n20442), .B2(n20446), .C1(
        n20441), .C2(n20444), .ZN(P2_U3240) );
  OAI222_X1 U23397 ( .A1(n20449), .A2(n20448), .B1(n20447), .B2(n20446), .C1(
        n20445), .C2(n20444), .ZN(P2_U3241) );
  OAI22_X1 U23398 ( .A1(n20483), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20446), .ZN(n20450) );
  INV_X1 U23399 ( .A(n20450), .ZN(P2_U3585) );
  MUX2_X1 U23400 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20483), .Z(P2_U3586) );
  OAI22_X1 U23401 ( .A1(n20483), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20446), .ZN(n20451) );
  INV_X1 U23402 ( .A(n20451), .ZN(P2_U3587) );
  OAI22_X1 U23403 ( .A1(n20483), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20446), .ZN(n20452) );
  INV_X1 U23404 ( .A(n20452), .ZN(P2_U3588) );
  OAI21_X1 U23405 ( .B1(n20456), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20454), 
        .ZN(n20453) );
  INV_X1 U23406 ( .A(n20453), .ZN(P2_U3591) );
  OAI21_X1 U23407 ( .B1(n20456), .B2(n20455), .A(n20454), .ZN(P2_U3592) );
  NOR2_X1 U23408 ( .A1(n20458), .A2(n20457), .ZN(n20467) );
  NAND2_X1 U23409 ( .A1(n20460), .A2(n20459), .ZN(n20474) );
  NAND2_X1 U23410 ( .A1(n20461), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20464) );
  AOI21_X1 U23411 ( .B1(n20464), .B2(n20463), .A(n20462), .ZN(n20473) );
  NAND2_X1 U23412 ( .A1(n20474), .A2(n20473), .ZN(n20466) );
  MUX2_X1 U23413 ( .A(n20467), .B(n20466), .S(n20465), .Z(n20468) );
  AOI21_X1 U23414 ( .B1(n20469), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20468), 
        .ZN(n20470) );
  AOI22_X1 U23415 ( .A1(n20481), .A2(n20471), .B1(n20470), .B2(n20478), .ZN(
        P2_U3602) );
  NOR2_X1 U23416 ( .A1(n20473), .A2(n20472), .ZN(n20476) );
  INV_X1 U23417 ( .A(n20474), .ZN(n20475) );
  AOI211_X1 U23418 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20477), .A(n20476), 
        .B(n20475), .ZN(n20479) );
  AOI22_X1 U23419 ( .A1(n20481), .A2(n20480), .B1(n20479), .B2(n20478), .ZN(
        P2_U3603) );
  INV_X1 U23420 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20482) );
  AOI22_X1 U23421 ( .A1(n20446), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20482), 
        .B2(n20483), .ZN(P2_U3608) );
  OAI22_X1 U23422 ( .A1(n20483), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20446), .ZN(n20484) );
  INV_X1 U23423 ( .A(n20484), .ZN(P2_U3611) );
  AOI21_X1 U23424 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21315), .A(n21312), 
        .ZN(n20487) );
  INV_X1 U23425 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20485) );
  AND2_X1 U23426 ( .A1(n21312), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21375) );
  AOI21_X1 U23427 ( .B1(n20487), .B2(n20485), .A(n21375), .ZN(P1_U2802) );
  INV_X1 U23428 ( .A(n21375), .ZN(n21373) );
  NOR2_X1 U23429 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20488) );
  INV_X1 U23430 ( .A(n21375), .ZN(n21389) );
  OAI21_X1 U23431 ( .B1(n20488), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21389), .ZN(
        n20486) );
  OAI21_X1 U23432 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21373), .A(n20486), 
        .ZN(P1_U2804) );
  NOR2_X1 U23433 ( .A1(n21375), .A2(n20487), .ZN(n21363) );
  OAI21_X1 U23434 ( .B1(BS16), .B2(n20488), .A(n21363), .ZN(n21361) );
  OAI21_X1 U23435 ( .B1(n21363), .B2(n21191), .A(n21361), .ZN(P1_U2805) );
  AOI21_X1 U23436 ( .B1(n20489), .B2(P1_FLUSH_REG_SCAN_IN), .A(n20650), .ZN(
        n20490) );
  INV_X1 U23437 ( .A(n20490), .ZN(P1_U2806) );
  NOR4_X1 U23438 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_11__SCAN_IN), .A3(P1_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20500) );
  NOR4_X1 U23439 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_6__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20499) );
  NOR2_X1 U23440 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n21401) );
  AOI211_X1 U23441 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_3__SCAN_IN), .B(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n20491) );
  NAND2_X1 U23442 ( .A1(n21401), .A2(n20491), .ZN(n20497) );
  NOR4_X1 U23443 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20495) );
  NOR4_X1 U23444 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_14__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_17__SCAN_IN), .ZN(n20494) );
  NOR4_X1 U23445 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_27__SCAN_IN), .A3(P1_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20493) );
  NOR4_X1 U23446 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20492) );
  NAND4_X1 U23447 ( .A1(n20495), .A2(n20494), .A3(n20493), .A4(n20492), .ZN(
        n20496) );
  NOR4_X1 U23448 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_2__SCAN_IN), .A3(n20497), .A4(n20496), .ZN(n20498) );
  NAND3_X1 U23449 ( .A1(n20500), .A2(n20499), .A3(n20498), .ZN(n21366) );
  NOR2_X1 U23450 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n21366), .ZN(n20502) );
  INV_X1 U23451 ( .A(n21366), .ZN(n21371) );
  NOR2_X1 U23452 ( .A1(n21371), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20501)
         );
  NOR2_X1 U23453 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(n21366), .ZN(n21364) );
  INV_X1 U23454 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21368) );
  INV_X1 U23455 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21362) );
  NAND3_X1 U23456 ( .A1(n21364), .A2(n21368), .A3(n21362), .ZN(n20503) );
  OAI21_X1 U23457 ( .B1(n20502), .B2(n20501), .A(n20503), .ZN(P1_U2807) );
  INV_X1 U23458 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20504) );
  NAND2_X1 U23459 ( .A1(n20502), .A2(n21362), .ZN(n21369) );
  OAI211_X1 U23460 ( .C1(n21371), .C2(n20504), .A(n20503), .B(n21369), .ZN(
        P1_U2808) );
  AOI22_X1 U23461 ( .A1(n20506), .A2(n20575), .B1(n20505), .B2(n20510), .ZN(
        n20516) );
  OAI22_X1 U23462 ( .A1(n20508), .A2(n20565), .B1(n20589), .B2(n20507), .ZN(
        n20509) );
  AOI211_X1 U23463 ( .C1(n20541), .C2(P1_EBX_REG_9__SCAN_IN), .A(n20683), .B(
        n20509), .ZN(n20515) );
  NOR2_X1 U23464 ( .A1(n20511), .A2(n20510), .ZN(n20512) );
  AOI21_X1 U23465 ( .B1(n20513), .B2(n20536), .A(n20512), .ZN(n20514) );
  NAND3_X1 U23466 ( .A1(n20516), .A2(n20515), .A3(n20514), .ZN(P1_U2831) );
  NAND2_X1 U23467 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20519) );
  OAI21_X1 U23468 ( .B1(n20519), .B2(n20518), .A(n20517), .ZN(n20539) );
  NOR2_X1 U23469 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20519), .ZN(n20520) );
  AOI22_X1 U23470 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(n20541), .B1(n20540), .B2(
        n20520), .ZN(n20530) );
  INV_X1 U23471 ( .A(n20521), .ZN(n20524) );
  INV_X1 U23472 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20522) );
  OAI21_X1 U23473 ( .B1(n20565), .B2(n20522), .A(n20667), .ZN(n20523) );
  AOI21_X1 U23474 ( .B1(n20524), .B2(n20575), .A(n20523), .ZN(n20525) );
  OAI21_X1 U23475 ( .B1(n20589), .B2(n20526), .A(n20525), .ZN(n20527) );
  AOI21_X1 U23476 ( .B1(n20528), .B2(n20536), .A(n20527), .ZN(n20529) );
  OAI211_X1 U23477 ( .C1(n21438), .C2(n20539), .A(n20530), .B(n20529), .ZN(
        P1_U2833) );
  INV_X1 U23478 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21320) );
  NOR2_X1 U23479 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n21320), .ZN(n20531) );
  AOI22_X1 U23480 ( .A1(n20532), .A2(n10449), .B1(n20540), .B2(n20531), .ZN(
        n20538) );
  AOI22_X1 U23481 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20579), .B1(
        P1_EBX_REG_6__SCAN_IN), .B2(n20574), .ZN(n20533) );
  OAI211_X1 U23482 ( .C1(n20560), .C2(n20534), .A(n20533), .B(n20667), .ZN(
        n20535) );
  AOI21_X1 U23483 ( .B1(n20591), .B2(n20536), .A(n20535), .ZN(n20537) );
  OAI211_X1 U23484 ( .C1(n17365), .C2(n20539), .A(n20538), .B(n20537), .ZN(
        P1_U2834) );
  AOI22_X1 U23485 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n20541), .B1(n20540), .B2(
        n21320), .ZN(n20549) );
  OAI22_X1 U23486 ( .A1(n20543), .A2(n20560), .B1(n20589), .B2(n20542), .ZN(
        n20544) );
  AOI211_X1 U23487 ( .C1(n20579), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n20683), .B(n20544), .ZN(n20548) );
  INV_X1 U23488 ( .A(n20545), .ZN(n20556) );
  AOI22_X1 U23489 ( .A1(n20546), .A2(n20585), .B1(n20556), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n20547) );
  NAND3_X1 U23490 ( .A1(n20549), .A2(n20548), .A3(n20547), .ZN(P1_U2835) );
  OR2_X1 U23491 ( .A1(n14072), .A2(n20550), .ZN(n20551) );
  NAND2_X1 U23492 ( .A1(n14194), .A2(n20551), .ZN(n20655) );
  OAI222_X1 U23493 ( .A1(n20598), .A2(n20553), .B1(n20578), .B2(n20552), .C1(
        n20589), .C2(n20655), .ZN(n20554) );
  AOI211_X1 U23494 ( .C1(n20579), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20683), .B(n20554), .ZN(n20559) );
  NAND2_X1 U23495 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n20564) );
  NAND2_X1 U23496 ( .A1(n20555), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20583) );
  INV_X1 U23497 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21317) );
  OAI21_X1 U23498 ( .B1(n20564), .B2(n20583), .A(n21317), .ZN(n20557) );
  AOI22_X1 U23499 ( .A1(n20557), .A2(n20556), .B1(n20648), .B2(n20585), .ZN(
        n20558) );
  OAI211_X1 U23500 ( .C1(n20653), .C2(n20560), .A(n20559), .B(n20558), .ZN(
        P1_U2836) );
  AOI22_X1 U23501 ( .A1(n20561), .A2(n20575), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n20574), .ZN(n20573) );
  NAND2_X1 U23502 ( .A1(n20563), .A2(n20562), .ZN(n20577) );
  OAI21_X1 U23503 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(P1_REIP_REG_2__SCAN_IN), 
        .A(n20564), .ZN(n20567) );
  OAI22_X1 U23504 ( .A1(n20583), .A2(n20567), .B1(n20566), .B2(n20565), .ZN(
        n20568) );
  AOI21_X1 U23505 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(n20577), .A(n20568), .ZN(
        n20569) );
  OAI21_X1 U23506 ( .B1(n20994), .B2(n20578), .A(n20569), .ZN(n20570) );
  AOI21_X1 U23507 ( .B1(n20571), .B2(n20585), .A(n20570), .ZN(n20572) );
  OAI211_X1 U23508 ( .C1(n20589), .C2(n20669), .A(n20573), .B(n20572), .ZN(
        P1_U2837) );
  AOI22_X1 U23509 ( .A1(n20576), .A2(n20575), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n20574), .ZN(n20588) );
  NAND2_X1 U23510 ( .A1(n20577), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20582) );
  INV_X1 U23511 ( .A(n20578), .ZN(n20580) );
  INV_X1 U23512 ( .A(n21127), .ZN(n20993) );
  AOI22_X1 U23513 ( .A1(n20580), .A2(n20993), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20579), .ZN(n20581) );
  OAI211_X1 U23514 ( .C1(P1_REIP_REG_2__SCAN_IN), .C2(n20583), .A(n20582), .B(
        n20581), .ZN(n20584) );
  AOI21_X1 U23515 ( .B1(n20586), .B2(n20585), .A(n20584), .ZN(n20587) );
  OAI211_X1 U23516 ( .C1(n20589), .C2(n20682), .A(n20588), .B(n20587), .ZN(
        P1_U2838) );
  INV_X1 U23517 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20593) );
  AOI22_X1 U23518 ( .A1(n20591), .A2(n20596), .B1(n20590), .B2(n10449), .ZN(
        n20592) );
  OAI21_X1 U23519 ( .B1(n20599), .B2(n20593), .A(n20592), .ZN(P1_U2866) );
  NOR2_X1 U23520 ( .A1(n20594), .A2(n20655), .ZN(n20595) );
  AOI21_X1 U23521 ( .B1(n20648), .B2(n20596), .A(n20595), .ZN(n20597) );
  OAI21_X1 U23522 ( .B1(n20599), .B2(n20598), .A(n20597), .ZN(P1_U2868) );
  AOI22_X1 U23523 ( .A1(n20624), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20601) );
  OAI21_X1 U23524 ( .B1(n20602), .B2(n20626), .A(n20601), .ZN(P1_U2921) );
  AOI22_X1 U23525 ( .A1(n20612), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20603) );
  OAI21_X1 U23526 ( .B1(n20604), .B2(n20626), .A(n20603), .ZN(P1_U2922) );
  INV_X1 U23527 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20640) );
  AOI22_X1 U23528 ( .A1(n20612), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20605) );
  OAI21_X1 U23529 ( .B1(n20640), .B2(n20626), .A(n20605), .ZN(P1_U2923) );
  AOI22_X1 U23530 ( .A1(n20612), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20606) );
  OAI21_X1 U23531 ( .B1(n20607), .B2(n20626), .A(n20606), .ZN(P1_U2924) );
  AOI22_X1 U23532 ( .A1(n20612), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20608) );
  OAI21_X1 U23533 ( .B1(n11687), .B2(n20626), .A(n20608), .ZN(P1_U2925) );
  AOI22_X1 U23534 ( .A1(n20612), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20609) );
  OAI21_X1 U23535 ( .B1(n20610), .B2(n20626), .A(n20609), .ZN(P1_U2926) );
  AOI22_X1 U23536 ( .A1(n20612), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20611) );
  OAI21_X1 U23537 ( .B1(n11653), .B2(n20626), .A(n20611), .ZN(P1_U2927) );
  AOI22_X1 U23538 ( .A1(n20612), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20613) );
  OAI21_X1 U23539 ( .B1(n11637), .B2(n20626), .A(n20613), .ZN(P1_U2928) );
  AOI22_X1 U23540 ( .A1(n20624), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20614) );
  OAI21_X1 U23541 ( .B1(n11619), .B2(n20626), .A(n20614), .ZN(P1_U2929) );
  AOI22_X1 U23542 ( .A1(n20624), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20616) );
  OAI21_X1 U23543 ( .B1(n11568), .B2(n20626), .A(n20616), .ZN(P1_U2930) );
  AOI22_X1 U23544 ( .A1(n20624), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20617) );
  OAI21_X1 U23545 ( .B1(n11552), .B2(n20626), .A(n20617), .ZN(P1_U2931) );
  AOI22_X1 U23546 ( .A1(n20624), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20618) );
  OAI21_X1 U23547 ( .B1(n20619), .B2(n20626), .A(n20618), .ZN(P1_U2932) );
  AOI22_X1 U23548 ( .A1(n20624), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20620) );
  OAI21_X1 U23549 ( .B1(n20621), .B2(n20626), .A(n20620), .ZN(P1_U2933) );
  AOI22_X1 U23550 ( .A1(n20624), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20622) );
  OAI21_X1 U23551 ( .B1(n21432), .B2(n20626), .A(n20622), .ZN(P1_U2934) );
  AOI22_X1 U23552 ( .A1(n20624), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20623) );
  OAI21_X1 U23553 ( .B1(n11580), .B2(n20626), .A(n20623), .ZN(P1_U2935) );
  AOI22_X1 U23554 ( .A1(n20624), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20615), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20625) );
  OAI21_X1 U23555 ( .B1(n20627), .B2(n20626), .A(n20625), .ZN(P1_U2936) );
  AOI21_X1 U23556 ( .B1(P1_UWORD_REG_0__SCAN_IN), .B2(n20637), .A(n20628), 
        .ZN(n20629) );
  OAI21_X1 U23557 ( .B1(n20630), .B2(n20639), .A(n20629), .ZN(P1_U2937) );
  INV_X1 U23558 ( .A(n20631), .ZN(n20632) );
  NOR2_X1 U23559 ( .A1(n20633), .A2(n20632), .ZN(n20636) );
  AOI21_X1 U23560 ( .B1(P1_UWORD_REG_13__SCAN_IN), .B2(n20637), .A(n20636), 
        .ZN(n20634) );
  OAI21_X1 U23561 ( .B1(n20635), .B2(n20639), .A(n20634), .ZN(P1_U2950) );
  AOI21_X1 U23562 ( .B1(P1_LWORD_REG_13__SCAN_IN), .B2(n20637), .A(n20636), 
        .ZN(n20638) );
  OAI21_X1 U23563 ( .B1(n20640), .B2(n20639), .A(n20638), .ZN(P1_U2965) );
  NOR2_X1 U23564 ( .A1(n20667), .A2(n21317), .ZN(n20656) );
  AOI21_X1 U23565 ( .B1(n20641), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20656), .ZN(n20652) );
  NAND2_X1 U23566 ( .A1(n20642), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n20643) );
  NAND2_X1 U23567 ( .A1(n20644), .A2(n20643), .ZN(n20647) );
  XNOR2_X1 U23568 ( .A(n20645), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20646) );
  XNOR2_X1 U23569 ( .A(n20647), .B(n20646), .ZN(n20659) );
  AOI22_X1 U23570 ( .A1(n20659), .A2(n20650), .B1(n20649), .B2(n20648), .ZN(
        n20651) );
  OAI211_X1 U23571 ( .C1(n20654), .C2(n20653), .A(n20652), .B(n20651), .ZN(
        P1_U2995) );
  INV_X1 U23572 ( .A(n20655), .ZN(n20657) );
  AOI21_X1 U23573 ( .B1(n20696), .B2(n20657), .A(n20656), .ZN(n20663) );
  AOI211_X1 U23574 ( .C1(n20664), .C2(n20673), .A(n20658), .B(n20674), .ZN(
        n20661) );
  AND2_X1 U23575 ( .A1(n20659), .A2(n20699), .ZN(n20660) );
  NOR2_X1 U23576 ( .A1(n20661), .A2(n20660), .ZN(n20662) );
  OAI211_X1 U23577 ( .C1(n20672), .C2(n20664), .A(n20663), .B(n20662), .ZN(
        P1_U3027) );
  OAI222_X1 U23578 ( .A1(n20669), .A2(n20668), .B1(n20667), .B2(n14230), .C1(
        n20666), .C2(n20665), .ZN(n20670) );
  INV_X1 U23579 ( .A(n20670), .ZN(n20671) );
  OAI221_X1 U23580 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20674), .C1(
        n20673), .C2(n20672), .A(n20671), .ZN(P1_U3028) );
  NAND2_X1 U23581 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20675), .ZN(
        n20691) );
  NOR3_X1 U23582 ( .A1(n13458), .A2(n20703), .A3(n20676), .ZN(n20678) );
  AOI211_X1 U23583 ( .C1(n20703), .C2(n20679), .A(n20678), .B(n20677), .ZN(
        n20689) );
  NAND3_X1 U23584 ( .A1(n20681), .A2(n20680), .A3(n20699), .ZN(n20687) );
  INV_X1 U23585 ( .A(n20682), .ZN(n20684) );
  AOI22_X1 U23586 ( .A1(n20696), .A2(n20684), .B1(n20683), .B2(
        P1_REIP_REG_2__SCAN_IN), .ZN(n20686) );
  AND3_X1 U23587 ( .A1(n20687), .A2(n20686), .A3(n20685), .ZN(n20688) );
  OAI221_X1 U23588 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20691), .C1(
        n20690), .C2(n20689), .A(n20688), .ZN(P1_U3029) );
  INV_X1 U23589 ( .A(n20692), .ZN(n20695) );
  INV_X1 U23590 ( .A(n20693), .ZN(n20694) );
  AOI21_X1 U23591 ( .B1(n20696), .B2(n20695), .A(n20694), .ZN(n20706) );
  NOR2_X1 U23592 ( .A1(n20697), .A2(n20703), .ZN(n20698) );
  AOI21_X1 U23593 ( .B1(n20700), .B2(n20699), .A(n20698), .ZN(n20705) );
  NAND3_X1 U23594 ( .A1(n20703), .A2(n20702), .A3(n20701), .ZN(n20704) );
  NAND3_X1 U23595 ( .A1(n20706), .A2(n20705), .A3(n20704), .ZN(P1_U3030) );
  NOR2_X1 U23596 ( .A1(n20708), .A2(n20707), .ZN(P1_U3032) );
  AOI22_X1 U23597 ( .A1(DATAI_16_), .A2(n20710), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20762), .ZN(n21251) );
  AOI22_X1 U23598 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20762), .B1(DATAI_24_), 
        .B2(n20710), .ZN(n21202) );
  NOR3_X1 U23599 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20777) );
  INV_X1 U23600 ( .A(n20777), .ZN(n20773) );
  NOR2_X1 U23601 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20773), .ZN(
        n20722) );
  INV_X1 U23602 ( .A(n20722), .ZN(n20765) );
  NOR2_X2 U23603 ( .A1(n20764), .A2(n20715), .ZN(n21240) );
  INV_X1 U23604 ( .A(n21240), .ZN(n21046) );
  OAI22_X1 U23605 ( .A1(n21297), .A2(n21202), .B1(n20765), .B2(n21046), .ZN(
        n20716) );
  INV_X1 U23606 ( .A(n20716), .ZN(n20732) );
  INV_X1 U23607 ( .A(n20797), .ZN(n20718) );
  INV_X1 U23608 ( .A(n21297), .ZN(n20717) );
  OAI21_X1 U23609 ( .B1(n20718), .B2(n20717), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20719) );
  NAND2_X1 U23610 ( .A1(n20719), .A2(n21163), .ZN(n20730) );
  OR2_X1 U23611 ( .A1(n20720), .A2(n20993), .ZN(n20802) );
  NOR2_X1 U23612 ( .A1(n20802), .A2(n21194), .ZN(n20726) );
  INV_X1 U23613 ( .A(n20874), .ZN(n20995) );
  NAND2_X1 U23614 ( .A1(n20995), .A2(n21184), .ZN(n20728) );
  INV_X1 U23615 ( .A(n20727), .ZN(n20721) );
  NOR2_X1 U23616 ( .A1(n20721), .A2(n21239), .ZN(n20873) );
  OAI21_X1 U23617 ( .B1(n20722), .B2(n21000), .A(n21050), .ZN(n20723) );
  AOI21_X1 U23618 ( .B1(n20728), .B2(P1_STATE2_REG_2__SCAN_IN), .A(n20723), 
        .ZN(n20724) );
  NOR2_X2 U23619 ( .A1(n20775), .A2(n20725), .ZN(n21241) );
  INV_X1 U23620 ( .A(n20726), .ZN(n20729) );
  OR2_X1 U23621 ( .A1(n20727), .A2(n21239), .ZN(n21054) );
  AOI22_X1 U23622 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20769), .B1(
        n21241), .B2(n20768), .ZN(n20731) );
  OAI211_X1 U23623 ( .C1(n21251), .C2(n20797), .A(n20732), .B(n20731), .ZN(
        P1_U3033) );
  AOI22_X1 U23624 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20762), .B1(DATAI_25_), 
        .B2(n20710), .ZN(n21206) );
  OR2_X1 U23625 ( .A1(n20764), .A2(n20733), .ZN(n21059) );
  OAI22_X1 U23626 ( .A1(n21297), .A2(n21206), .B1(n20765), .B2(n21059), .ZN(
        n20734) );
  INV_X1 U23627 ( .A(n20734), .ZN(n20737) );
  NOR2_X2 U23628 ( .A1(n20775), .A2(n20735), .ZN(n21253) );
  AOI22_X1 U23629 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20769), .B1(
        n21253), .B2(n20768), .ZN(n20736) );
  OAI211_X1 U23630 ( .C1(n21257), .C2(n20797), .A(n20737), .B(n20736), .ZN(
        P1_U3034) );
  AOI22_X1 U23631 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20762), .B1(DATAI_18_), 
        .B2(n20710), .ZN(n21263) );
  OAI22_X1 U23632 ( .A1(n21297), .A2(n21210), .B1(n20765), .B2(n21063), .ZN(
        n20738) );
  INV_X1 U23633 ( .A(n20738), .ZN(n20741) );
  NOR2_X2 U23634 ( .A1(n20775), .A2(n20739), .ZN(n21259) );
  AOI22_X1 U23635 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20769), .B1(
        n21259), .B2(n20768), .ZN(n20740) );
  OAI211_X1 U23636 ( .C1(n21263), .C2(n20797), .A(n20741), .B(n20740), .ZN(
        P1_U3035) );
  AOI22_X1 U23637 ( .A1(DATAI_19_), .A2(n20710), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20762), .ZN(n21269) );
  NOR2_X2 U23638 ( .A1(n20764), .A2(n20742), .ZN(n21264) );
  INV_X1 U23639 ( .A(n21264), .ZN(n21067) );
  OAI22_X1 U23640 ( .A1(n21297), .A2(n21214), .B1(n20765), .B2(n21067), .ZN(
        n20743) );
  INV_X1 U23641 ( .A(n20743), .ZN(n20746) );
  NOR2_X2 U23642 ( .A1(n20775), .A2(n20744), .ZN(n21265) );
  AOI22_X1 U23643 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20769), .B1(
        n21265), .B2(n20768), .ZN(n20745) );
  OAI211_X1 U23644 ( .C1(n21269), .C2(n20797), .A(n20746), .B(n20745), .ZN(
        P1_U3036) );
  AOI22_X1 U23645 ( .A1(DATAI_20_), .A2(n20710), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20762), .ZN(n21275) );
  NOR2_X2 U23646 ( .A1(n20764), .A2(n20747), .ZN(n21270) );
  INV_X1 U23647 ( .A(n21270), .ZN(n21071) );
  OAI22_X1 U23648 ( .A1(n21297), .A2(n21218), .B1(n20765), .B2(n21071), .ZN(
        n20748) );
  INV_X1 U23649 ( .A(n20748), .ZN(n20751) );
  NOR2_X2 U23650 ( .A1(n20775), .A2(n20749), .ZN(n21271) );
  AOI22_X1 U23651 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20769), .B1(
        n21271), .B2(n20768), .ZN(n20750) );
  OAI211_X1 U23652 ( .C1(n21275), .C2(n20797), .A(n20751), .B(n20750), .ZN(
        P1_U3037) );
  AOI22_X1 U23653 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20762), .B1(DATAI_29_), 
        .B2(n20710), .ZN(n21222) );
  OR2_X1 U23654 ( .A1(n20764), .A2(n20752), .ZN(n21075) );
  OAI22_X1 U23655 ( .A1(n21297), .A2(n21222), .B1(n20765), .B2(n21075), .ZN(
        n20753) );
  INV_X1 U23656 ( .A(n20753), .ZN(n20756) );
  NOR2_X2 U23657 ( .A1(n20775), .A2(n20754), .ZN(n21277) );
  AOI22_X1 U23658 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20769), .B1(
        n21277), .B2(n20768), .ZN(n20755) );
  OAI211_X1 U23659 ( .C1(n21281), .C2(n20797), .A(n20756), .B(n20755), .ZN(
        P1_U3038) );
  AOI22_X1 U23660 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20762), .B1(DATAI_22_), 
        .B2(n20710), .ZN(n21287) );
  OR2_X1 U23661 ( .A1(n20764), .A2(n20757), .ZN(n21079) );
  OAI22_X1 U23662 ( .A1(n21297), .A2(n21226), .B1(n20765), .B2(n21079), .ZN(
        n20758) );
  INV_X1 U23663 ( .A(n20758), .ZN(n20761) );
  NOR2_X2 U23664 ( .A1(n20775), .A2(n20759), .ZN(n21283) );
  AOI22_X1 U23665 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20769), .B1(
        n21283), .B2(n20768), .ZN(n20760) );
  OAI211_X1 U23666 ( .C1(n21287), .C2(n20797), .A(n20761), .B(n20760), .ZN(
        P1_U3039) );
  AOI22_X1 U23667 ( .A1(DATAI_23_), .A2(n20710), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n20762), .ZN(n21298) );
  NOR2_X2 U23668 ( .A1(n20764), .A2(n20763), .ZN(n21288) );
  INV_X1 U23669 ( .A(n21288), .ZN(n21083) );
  OAI22_X1 U23670 ( .A1(n21297), .A2(n21234), .B1(n20765), .B2(n21083), .ZN(
        n20766) );
  INV_X1 U23671 ( .A(n20766), .ZN(n20771) );
  NOR2_X2 U23672 ( .A1(n20775), .A2(n20767), .ZN(n21290) );
  AOI22_X1 U23673 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20769), .B1(
        n21290), .B2(n20768), .ZN(n20770) );
  OAI211_X1 U23674 ( .C1(n21298), .C2(n20797), .A(n20771), .B(n20770), .ZN(
        P1_U3040) );
  INV_X1 U23675 ( .A(n20802), .ZN(n20839) );
  INV_X1 U23676 ( .A(n20772), .ZN(n21158) );
  NOR2_X1 U23677 ( .A1(n21157), .A2(n20773), .ZN(n20792) );
  AOI21_X1 U23678 ( .B1(n20839), .B2(n21158), .A(n20792), .ZN(n20774) );
  OAI22_X1 U23679 ( .A1(n20774), .A2(n21376), .B1(n20773), .B2(n21239), .ZN(
        n20793) );
  AOI22_X1 U23680 ( .A1(n20793), .A2(n21241), .B1(n21240), .B2(n20792), .ZN(
        n20779) );
  INV_X1 U23681 ( .A(n20834), .ZN(n20837) );
  OAI211_X1 U23682 ( .C1(n20837), .C2(n21191), .A(n21163), .B(n20774), .ZN(
        n20776) );
  INV_X1 U23683 ( .A(n21251), .ZN(n21199) );
  AOI22_X1 U23684 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20794), .B1(
        n20799), .B2(n21199), .ZN(n20778) );
  OAI211_X1 U23685 ( .C1(n21202), .C2(n20797), .A(n20779), .B(n20778), .ZN(
        P1_U3041) );
  AOI22_X1 U23686 ( .A1(n20793), .A2(n21253), .B1(n21252), .B2(n20792), .ZN(
        n20781) );
  INV_X1 U23687 ( .A(n21257), .ZN(n21203) );
  AOI22_X1 U23688 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20794), .B1(
        n20799), .B2(n21203), .ZN(n20780) );
  OAI211_X1 U23689 ( .C1(n21206), .C2(n20797), .A(n20781), .B(n20780), .ZN(
        P1_U3042) );
  AOI22_X1 U23690 ( .A1(n20793), .A2(n21259), .B1(n21258), .B2(n20792), .ZN(
        n20783) );
  INV_X1 U23691 ( .A(n21263), .ZN(n21207) );
  AOI22_X1 U23692 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20794), .B1(
        n20799), .B2(n21207), .ZN(n20782) );
  OAI211_X1 U23693 ( .C1(n21210), .C2(n20797), .A(n20783), .B(n20782), .ZN(
        P1_U3043) );
  AOI22_X1 U23694 ( .A1(n20793), .A2(n21265), .B1(n21264), .B2(n20792), .ZN(
        n20785) );
  INV_X1 U23695 ( .A(n21269), .ZN(n21211) );
  AOI22_X1 U23696 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20794), .B1(
        n20799), .B2(n21211), .ZN(n20784) );
  OAI211_X1 U23697 ( .C1(n21214), .C2(n20797), .A(n20785), .B(n20784), .ZN(
        P1_U3044) );
  AOI22_X1 U23698 ( .A1(n20793), .A2(n21271), .B1(n21270), .B2(n20792), .ZN(
        n20787) );
  INV_X1 U23699 ( .A(n21275), .ZN(n21215) );
  AOI22_X1 U23700 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20794), .B1(
        n20799), .B2(n21215), .ZN(n20786) );
  OAI211_X1 U23701 ( .C1(n21218), .C2(n20797), .A(n20787), .B(n20786), .ZN(
        P1_U3045) );
  AOI22_X1 U23702 ( .A1(n20793), .A2(n21277), .B1(n21276), .B2(n20792), .ZN(
        n20789) );
  INV_X1 U23703 ( .A(n21281), .ZN(n21219) );
  AOI22_X1 U23704 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20794), .B1(
        n20799), .B2(n21219), .ZN(n20788) );
  OAI211_X1 U23705 ( .C1(n21222), .C2(n20797), .A(n20789), .B(n20788), .ZN(
        P1_U3046) );
  AOI22_X1 U23706 ( .A1(n20793), .A2(n21283), .B1(n21282), .B2(n20792), .ZN(
        n20791) );
  INV_X1 U23707 ( .A(n21287), .ZN(n21223) );
  AOI22_X1 U23708 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20794), .B1(
        n20799), .B2(n21223), .ZN(n20790) );
  OAI211_X1 U23709 ( .C1(n21226), .C2(n20797), .A(n20791), .B(n20790), .ZN(
        P1_U3047) );
  AOI22_X1 U23710 ( .A1(n20793), .A2(n21290), .B1(n21288), .B2(n20792), .ZN(
        n20796) );
  INV_X1 U23711 ( .A(n21298), .ZN(n21229) );
  AOI22_X1 U23712 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20794), .B1(
        n20799), .B2(n21229), .ZN(n20795) );
  OAI211_X1 U23713 ( .C1(n21234), .C2(n20797), .A(n20796), .B(n20795), .ZN(
        P1_U3048) );
  NAND3_X1 U23714 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21186), .A3(
        n21123), .ZN(n20843) );
  OR2_X1 U23715 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20843), .ZN(
        n20827) );
  OAI22_X1 U23716 ( .A1(n20871), .A2(n21251), .B1(n21046), .B2(n20827), .ZN(
        n20798) );
  INV_X1 U23717 ( .A(n20798), .ZN(n20808) );
  INV_X1 U23718 ( .A(n20871), .ZN(n20800) );
  OAI21_X1 U23719 ( .B1(n20800), .B2(n20799), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20801) );
  NAND2_X1 U23720 ( .A1(n20801), .A2(n21163), .ZN(n20806) );
  NOR2_X1 U23721 ( .A1(n20802), .A2(n21188), .ZN(n20804) );
  OR2_X1 U23722 ( .A1(n21184), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20932) );
  AND2_X1 U23723 ( .A1(n20932), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20928) );
  AOI21_X1 U23724 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20827), .A(n20928), 
        .ZN(n20803) );
  INV_X1 U23725 ( .A(n20804), .ZN(n20805) );
  AOI22_X1 U23726 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20830), .B1(
        n21241), .B2(n20829), .ZN(n20807) );
  OAI211_X1 U23727 ( .C1(n21202), .C2(n20833), .A(n20808), .B(n20807), .ZN(
        P1_U3049) );
  OAI22_X1 U23728 ( .A1(n20833), .A2(n21206), .B1(n20827), .B2(n21059), .ZN(
        n20809) );
  INV_X1 U23729 ( .A(n20809), .ZN(n20811) );
  AOI22_X1 U23730 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20830), .B1(
        n21253), .B2(n20829), .ZN(n20810) );
  OAI211_X1 U23731 ( .C1(n21257), .C2(n20871), .A(n20811), .B(n20810), .ZN(
        P1_U3050) );
  OAI22_X1 U23732 ( .A1(n20833), .A2(n21210), .B1(n20827), .B2(n21063), .ZN(
        n20812) );
  INV_X1 U23733 ( .A(n20812), .ZN(n20814) );
  AOI22_X1 U23734 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20830), .B1(
        n21259), .B2(n20829), .ZN(n20813) );
  OAI211_X1 U23735 ( .C1(n21263), .C2(n20871), .A(n20814), .B(n20813), .ZN(
        P1_U3051) );
  OAI22_X1 U23736 ( .A1(n20833), .A2(n21214), .B1(n21067), .B2(n20827), .ZN(
        n20815) );
  INV_X1 U23737 ( .A(n20815), .ZN(n20817) );
  AOI22_X1 U23738 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20830), .B1(
        n21265), .B2(n20829), .ZN(n20816) );
  OAI211_X1 U23739 ( .C1(n21269), .C2(n20871), .A(n20817), .B(n20816), .ZN(
        P1_U3052) );
  OAI22_X1 U23740 ( .A1(n20833), .A2(n21218), .B1(n21071), .B2(n20827), .ZN(
        n20818) );
  INV_X1 U23741 ( .A(n20818), .ZN(n20820) );
  AOI22_X1 U23742 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20830), .B1(
        n21271), .B2(n20829), .ZN(n20819) );
  OAI211_X1 U23743 ( .C1(n21275), .C2(n20871), .A(n20820), .B(n20819), .ZN(
        P1_U3053) );
  OAI22_X1 U23744 ( .A1(n20871), .A2(n21281), .B1(n20827), .B2(n21075), .ZN(
        n20821) );
  INV_X1 U23745 ( .A(n20821), .ZN(n20823) );
  AOI22_X1 U23746 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20830), .B1(
        n21277), .B2(n20829), .ZN(n20822) );
  OAI211_X1 U23747 ( .C1(n21222), .C2(n20833), .A(n20823), .B(n20822), .ZN(
        P1_U3054) );
  OAI22_X1 U23748 ( .A1(n20871), .A2(n21287), .B1(n20827), .B2(n21079), .ZN(
        n20824) );
  INV_X1 U23749 ( .A(n20824), .ZN(n20826) );
  AOI22_X1 U23750 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20830), .B1(
        n21283), .B2(n20829), .ZN(n20825) );
  OAI211_X1 U23751 ( .C1(n21226), .C2(n20833), .A(n20826), .B(n20825), .ZN(
        P1_U3055) );
  OAI22_X1 U23752 ( .A1(n20871), .A2(n21298), .B1(n21083), .B2(n20827), .ZN(
        n20828) );
  INV_X1 U23753 ( .A(n20828), .ZN(n20832) );
  AOI22_X1 U23754 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20830), .B1(
        n21290), .B2(n20829), .ZN(n20831) );
  OAI211_X1 U23755 ( .C1(n21234), .C2(n20833), .A(n20832), .B(n20831), .ZN(
        P1_U3056) );
  OR2_X1 U23756 ( .A1(n21093), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20861) );
  INV_X1 U23757 ( .A(n20861), .ZN(n20866) );
  AOI22_X1 U23758 ( .A1(n20896), .A2(n21199), .B1(n20866), .B2(n21240), .ZN(
        n20847) );
  INV_X1 U23759 ( .A(n20835), .ZN(n20836) );
  AOI21_X1 U23760 ( .B1(n20837), .B2(n21163), .A(n20836), .ZN(n20844) );
  AND2_X1 U23761 ( .A1(n20838), .A2(n11586), .ZN(n21236) );
  AOI21_X1 U23762 ( .B1(n20839), .B2(n21236), .A(n20866), .ZN(n20845) );
  INV_X1 U23763 ( .A(n20845), .ZN(n20842) );
  AOI21_X1 U23764 ( .B1(n20843), .B2(n21376), .A(n20840), .ZN(n20841) );
  AOI22_X1 U23765 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20868), .B1(
        n21241), .B2(n20867), .ZN(n20846) );
  OAI211_X1 U23766 ( .C1(n21202), .C2(n20871), .A(n20847), .B(n20846), .ZN(
        P1_U3057) );
  OAI22_X1 U23767 ( .A1(n20871), .A2(n21206), .B1(n20861), .B2(n21059), .ZN(
        n20848) );
  INV_X1 U23768 ( .A(n20848), .ZN(n20850) );
  AOI22_X1 U23769 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20868), .B1(
        n21253), .B2(n20867), .ZN(n20849) );
  OAI211_X1 U23770 ( .C1(n21257), .C2(n20865), .A(n20850), .B(n20849), .ZN(
        P1_U3058) );
  OAI22_X1 U23771 ( .A1(n20871), .A2(n21210), .B1(n20861), .B2(n21063), .ZN(
        n20851) );
  INV_X1 U23772 ( .A(n20851), .ZN(n20853) );
  AOI22_X1 U23773 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20868), .B1(
        n21259), .B2(n20867), .ZN(n20852) );
  OAI211_X1 U23774 ( .C1(n21263), .C2(n20865), .A(n20853), .B(n20852), .ZN(
        P1_U3059) );
  AOI22_X1 U23775 ( .A1(n20896), .A2(n21211), .B1(n20866), .B2(n21264), .ZN(
        n20855) );
  AOI22_X1 U23776 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20868), .B1(
        n21265), .B2(n20867), .ZN(n20854) );
  OAI211_X1 U23777 ( .C1(n21214), .C2(n20871), .A(n20855), .B(n20854), .ZN(
        P1_U3060) );
  AOI22_X1 U23778 ( .A1(n20896), .A2(n21215), .B1(n20866), .B2(n21270), .ZN(
        n20857) );
  AOI22_X1 U23779 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20868), .B1(
        n21271), .B2(n20867), .ZN(n20856) );
  OAI211_X1 U23780 ( .C1(n21218), .C2(n20871), .A(n20857), .B(n20856), .ZN(
        P1_U3061) );
  OAI22_X1 U23781 ( .A1(n20871), .A2(n21222), .B1(n20861), .B2(n21075), .ZN(
        n20858) );
  INV_X1 U23782 ( .A(n20858), .ZN(n20860) );
  AOI22_X1 U23783 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20868), .B1(
        n21277), .B2(n20867), .ZN(n20859) );
  OAI211_X1 U23784 ( .C1(n21281), .C2(n20865), .A(n20860), .B(n20859), .ZN(
        P1_U3062) );
  OAI22_X1 U23785 ( .A1(n20871), .A2(n21226), .B1(n20861), .B2(n21079), .ZN(
        n20862) );
  INV_X1 U23786 ( .A(n20862), .ZN(n20864) );
  AOI22_X1 U23787 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20868), .B1(
        n21283), .B2(n20867), .ZN(n20863) );
  OAI211_X1 U23788 ( .C1(n21287), .C2(n20865), .A(n20864), .B(n20863), .ZN(
        P1_U3063) );
  AOI22_X1 U23789 ( .A1(n20896), .A2(n21229), .B1(n20866), .B2(n21288), .ZN(
        n20870) );
  AOI22_X1 U23790 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20868), .B1(
        n21290), .B2(n20867), .ZN(n20869) );
  OAI211_X1 U23791 ( .C1(n21234), .C2(n20871), .A(n20870), .B(n20869), .ZN(
        P1_U3064) );
  NOR2_X1 U23792 ( .A1(n21127), .A2(n20872), .ZN(n20964) );
  INV_X1 U23793 ( .A(n20964), .ZN(n20877) );
  INV_X1 U23794 ( .A(n20873), .ZN(n21185) );
  INV_X1 U23795 ( .A(n21184), .ZN(n21052) );
  OAI33_X1 U23796 ( .A1(n21376), .A2(n21194), .A3(n20877), .B1(n21185), .B2(
        n20874), .B3(n21052), .ZN(n20895) );
  NOR3_X1 U23797 ( .A1(n21123), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20904) );
  INV_X1 U23798 ( .A(n20904), .ZN(n20900) );
  NOR2_X1 U23799 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20900), .ZN(
        n20894) );
  AOI22_X1 U23800 ( .A1(n9779), .A2(n21241), .B1(n21240), .B2(n20894), .ZN(
        n20881) );
  INV_X1 U23801 ( .A(n20925), .ZN(n20875) );
  OAI21_X1 U23802 ( .B1(n20896), .B2(n20875), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20876) );
  OAI21_X1 U23803 ( .B1(n21194), .B2(n20877), .A(n20876), .ZN(n20879) );
  INV_X1 U23804 ( .A(n21202), .ZN(n21248) );
  AOI22_X1 U23805 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20897), .B1(
        n20896), .B2(n21248), .ZN(n20880) );
  OAI211_X1 U23806 ( .C1(n21251), .C2(n20925), .A(n20881), .B(n20880), .ZN(
        P1_U3065) );
  AOI22_X1 U23807 ( .A1(n9779), .A2(n21253), .B1(n21252), .B2(n20894), .ZN(
        n20883) );
  INV_X1 U23808 ( .A(n21206), .ZN(n21254) );
  AOI22_X1 U23809 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20897), .B1(
        n20896), .B2(n21254), .ZN(n20882) );
  OAI211_X1 U23810 ( .C1(n21257), .C2(n20925), .A(n20883), .B(n20882), .ZN(
        P1_U3066) );
  AOI22_X1 U23811 ( .A1(n9779), .A2(n21259), .B1(n21258), .B2(n20894), .ZN(
        n20885) );
  INV_X1 U23812 ( .A(n21210), .ZN(n21260) );
  AOI22_X1 U23813 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20897), .B1(
        n20896), .B2(n21260), .ZN(n20884) );
  OAI211_X1 U23814 ( .C1(n21263), .C2(n20925), .A(n20885), .B(n20884), .ZN(
        P1_U3067) );
  AOI22_X1 U23815 ( .A1(n9779), .A2(n21265), .B1(n21264), .B2(n20894), .ZN(
        n20887) );
  INV_X1 U23816 ( .A(n21214), .ZN(n21266) );
  AOI22_X1 U23817 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20897), .B1(
        n20896), .B2(n21266), .ZN(n20886) );
  OAI211_X1 U23818 ( .C1(n21269), .C2(n20925), .A(n20887), .B(n20886), .ZN(
        P1_U3068) );
  AOI22_X1 U23819 ( .A1(n9779), .A2(n21271), .B1(n21270), .B2(n20894), .ZN(
        n20889) );
  INV_X1 U23820 ( .A(n21218), .ZN(n21272) );
  AOI22_X1 U23821 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20897), .B1(
        n20896), .B2(n21272), .ZN(n20888) );
  OAI211_X1 U23822 ( .C1(n21275), .C2(n20925), .A(n20889), .B(n20888), .ZN(
        P1_U3069) );
  AOI22_X1 U23823 ( .A1(n9779), .A2(n21277), .B1(n21276), .B2(n20894), .ZN(
        n20891) );
  INV_X1 U23824 ( .A(n21222), .ZN(n21278) );
  AOI22_X1 U23825 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20897), .B1(
        n20896), .B2(n21278), .ZN(n20890) );
  OAI211_X1 U23826 ( .C1(n21281), .C2(n20925), .A(n20891), .B(n20890), .ZN(
        P1_U3070) );
  AOI22_X1 U23827 ( .A1(n9779), .A2(n21283), .B1(n21282), .B2(n20894), .ZN(
        n20893) );
  INV_X1 U23828 ( .A(n21226), .ZN(n21284) );
  AOI22_X1 U23829 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20897), .B1(
        n20896), .B2(n21284), .ZN(n20892) );
  OAI211_X1 U23830 ( .C1(n21287), .C2(n20925), .A(n20893), .B(n20892), .ZN(
        P1_U3071) );
  AOI22_X1 U23831 ( .A1(n9779), .A2(n21290), .B1(n21288), .B2(n20894), .ZN(
        n20899) );
  INV_X1 U23832 ( .A(n21234), .ZN(n21292) );
  AOI22_X1 U23833 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20897), .B1(
        n20896), .B2(n21292), .ZN(n20898) );
  OAI211_X1 U23834 ( .C1(n21298), .C2(n20925), .A(n20899), .B(n20898), .ZN(
        P1_U3072) );
  NOR2_X1 U23835 ( .A1(n21157), .A2(n20900), .ZN(n20919) );
  AOI21_X1 U23836 ( .B1(n20964), .B2(n21158), .A(n20919), .ZN(n20901) );
  OAI22_X1 U23837 ( .A1(n20901), .A2(n21376), .B1(n20900), .B2(n21239), .ZN(
        n20920) );
  AOI22_X1 U23838 ( .A1(n20920), .A2(n21241), .B1(n21240), .B2(n20919), .ZN(
        n20906) );
  OAI211_X1 U23839 ( .C1(n20902), .C2(n21191), .A(n21163), .B(n20901), .ZN(
        n20903) );
  OAI211_X1 U23840 ( .C1(n21163), .C2(n20904), .A(n20903), .B(n21245), .ZN(
        n20922) );
  AOI22_X1 U23841 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20922), .B1(
        n20921), .B2(n21199), .ZN(n20905) );
  OAI211_X1 U23842 ( .C1(n21202), .C2(n20925), .A(n20906), .B(n20905), .ZN(
        P1_U3073) );
  AOI22_X1 U23843 ( .A1(n20920), .A2(n21253), .B1(n21252), .B2(n20919), .ZN(
        n20908) );
  AOI22_X1 U23844 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20922), .B1(
        n20921), .B2(n21203), .ZN(n20907) );
  OAI211_X1 U23845 ( .C1(n21206), .C2(n20925), .A(n20908), .B(n20907), .ZN(
        P1_U3074) );
  AOI22_X1 U23846 ( .A1(n20920), .A2(n21259), .B1(n21258), .B2(n20919), .ZN(
        n20910) );
  AOI22_X1 U23847 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20922), .B1(
        n20921), .B2(n21207), .ZN(n20909) );
  OAI211_X1 U23848 ( .C1(n21210), .C2(n20925), .A(n20910), .B(n20909), .ZN(
        P1_U3075) );
  AOI22_X1 U23849 ( .A1(n20920), .A2(n21265), .B1(n21264), .B2(n20919), .ZN(
        n20912) );
  AOI22_X1 U23850 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20922), .B1(
        n20921), .B2(n21211), .ZN(n20911) );
  OAI211_X1 U23851 ( .C1(n21214), .C2(n20925), .A(n20912), .B(n20911), .ZN(
        P1_U3076) );
  AOI22_X1 U23852 ( .A1(n20920), .A2(n21271), .B1(n21270), .B2(n20919), .ZN(
        n20914) );
  AOI22_X1 U23853 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20922), .B1(
        n20921), .B2(n21215), .ZN(n20913) );
  OAI211_X1 U23854 ( .C1(n21218), .C2(n20925), .A(n20914), .B(n20913), .ZN(
        P1_U3077) );
  AOI22_X1 U23855 ( .A1(n20920), .A2(n21277), .B1(n21276), .B2(n20919), .ZN(
        n20916) );
  AOI22_X1 U23856 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20922), .B1(
        n20921), .B2(n21219), .ZN(n20915) );
  OAI211_X1 U23857 ( .C1(n21222), .C2(n20925), .A(n20916), .B(n20915), .ZN(
        P1_U3078) );
  AOI22_X1 U23858 ( .A1(n20920), .A2(n21283), .B1(n21282), .B2(n20919), .ZN(
        n20918) );
  AOI22_X1 U23859 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20922), .B1(
        n20921), .B2(n21223), .ZN(n20917) );
  OAI211_X1 U23860 ( .C1(n21226), .C2(n20925), .A(n20918), .B(n20917), .ZN(
        P1_U3079) );
  AOI22_X1 U23861 ( .A1(n20920), .A2(n21290), .B1(n21288), .B2(n20919), .ZN(
        n20924) );
  AOI22_X1 U23862 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20922), .B1(
        n20921), .B2(n21229), .ZN(n20923) );
  OAI211_X1 U23863 ( .C1(n21234), .C2(n20925), .A(n20924), .B(n20923), .ZN(
        P1_U3080) );
  NOR2_X1 U23864 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20965), .ZN(
        n20930) );
  INV_X1 U23865 ( .A(n20930), .ZN(n20955) );
  OAI22_X1 U23866 ( .A1(n20956), .A2(n21202), .B1(n21046), .B2(n20955), .ZN(
        n20926) );
  INV_X1 U23867 ( .A(n20926), .ZN(n20936) );
  NAND2_X1 U23868 ( .A1(n20991), .A2(n20956), .ZN(n20927) );
  AOI21_X1 U23869 ( .B1(n20927), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21376), 
        .ZN(n20931) );
  NAND2_X1 U23870 ( .A1(n20964), .A2(n21194), .ZN(n20933) );
  AOI21_X1 U23871 ( .B1(n20931), .B2(n20933), .A(n20928), .ZN(n20929) );
  INV_X1 U23872 ( .A(n20931), .ZN(n20934) );
  AOI22_X1 U23873 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20959), .B1(
        n21241), .B2(n20958), .ZN(n20935) );
  OAI211_X1 U23874 ( .C1(n21251), .C2(n20991), .A(n20936), .B(n20935), .ZN(
        P1_U3081) );
  OAI22_X1 U23875 ( .A1(n20991), .A2(n21257), .B1(n21059), .B2(n20955), .ZN(
        n20937) );
  INV_X1 U23876 ( .A(n20937), .ZN(n20939) );
  AOI22_X1 U23877 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20959), .B1(
        n21253), .B2(n20958), .ZN(n20938) );
  OAI211_X1 U23878 ( .C1(n21206), .C2(n20956), .A(n20939), .B(n20938), .ZN(
        P1_U3082) );
  OAI22_X1 U23879 ( .A1(n20956), .A2(n21210), .B1(n21063), .B2(n20955), .ZN(
        n20940) );
  INV_X1 U23880 ( .A(n20940), .ZN(n20942) );
  AOI22_X1 U23881 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20959), .B1(
        n21259), .B2(n20958), .ZN(n20941) );
  OAI211_X1 U23882 ( .C1(n21263), .C2(n20991), .A(n20942), .B(n20941), .ZN(
        P1_U3083) );
  OAI22_X1 U23883 ( .A1(n20956), .A2(n21214), .B1(n21067), .B2(n20955), .ZN(
        n20943) );
  INV_X1 U23884 ( .A(n20943), .ZN(n20945) );
  AOI22_X1 U23885 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20959), .B1(
        n21265), .B2(n20958), .ZN(n20944) );
  OAI211_X1 U23886 ( .C1(n21269), .C2(n20991), .A(n20945), .B(n20944), .ZN(
        P1_U3084) );
  OAI22_X1 U23887 ( .A1(n20991), .A2(n21275), .B1(n21071), .B2(n20955), .ZN(
        n20946) );
  INV_X1 U23888 ( .A(n20946), .ZN(n20948) );
  AOI22_X1 U23889 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20959), .B1(
        n21271), .B2(n20958), .ZN(n20947) );
  OAI211_X1 U23890 ( .C1(n21218), .C2(n20956), .A(n20948), .B(n20947), .ZN(
        P1_U3085) );
  OAI22_X1 U23891 ( .A1(n20991), .A2(n21281), .B1(n21075), .B2(n20955), .ZN(
        n20949) );
  INV_X1 U23892 ( .A(n20949), .ZN(n20951) );
  AOI22_X1 U23893 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20959), .B1(
        n21277), .B2(n20958), .ZN(n20950) );
  OAI211_X1 U23894 ( .C1(n21222), .C2(n20956), .A(n20951), .B(n20950), .ZN(
        P1_U3086) );
  OAI22_X1 U23895 ( .A1(n20956), .A2(n21226), .B1(n21079), .B2(n20955), .ZN(
        n20952) );
  INV_X1 U23896 ( .A(n20952), .ZN(n20954) );
  AOI22_X1 U23897 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20959), .B1(
        n21283), .B2(n20958), .ZN(n20953) );
  OAI211_X1 U23898 ( .C1(n21287), .C2(n20991), .A(n20954), .B(n20953), .ZN(
        P1_U3087) );
  OAI22_X1 U23899 ( .A1(n20956), .A2(n21234), .B1(n21083), .B2(n20955), .ZN(
        n20957) );
  INV_X1 U23900 ( .A(n20957), .ZN(n20961) );
  AOI22_X1 U23901 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20959), .B1(
        n21290), .B2(n20958), .ZN(n20960) );
  OAI211_X1 U23902 ( .C1(n21298), .C2(n20991), .A(n20961), .B(n20960), .ZN(
        P1_U3088) );
  INV_X1 U23903 ( .A(n20963), .ZN(n20986) );
  AOI21_X1 U23904 ( .B1(n20964), .B2(n21236), .A(n20986), .ZN(n20967) );
  OAI22_X1 U23905 ( .A1(n20967), .A2(n21376), .B1(n20965), .B2(n21239), .ZN(
        n20987) );
  AOI22_X1 U23906 ( .A1(n20987), .A2(n21241), .B1(n20986), .B2(n21240), .ZN(
        n20971) );
  INV_X1 U23907 ( .A(n20966), .ZN(n20968) );
  NAND3_X1 U23908 ( .A1(n20968), .A2(n21163), .A3(n20967), .ZN(n20969) );
  INV_X1 U23909 ( .A(n20991), .ZN(n20980) );
  AOI22_X1 U23910 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20988), .B1(
        n20980), .B2(n21248), .ZN(n20970) );
  OAI211_X1 U23911 ( .C1(n21251), .C2(n20983), .A(n20971), .B(n20970), .ZN(
        P1_U3089) );
  AOI22_X1 U23912 ( .A1(n20987), .A2(n21253), .B1(n20986), .B2(n21252), .ZN(
        n20973) );
  AOI22_X1 U23913 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20988), .B1(
        n20980), .B2(n21254), .ZN(n20972) );
  OAI211_X1 U23914 ( .C1(n21257), .C2(n20983), .A(n20973), .B(n20972), .ZN(
        P1_U3090) );
  AOI22_X1 U23915 ( .A1(n20987), .A2(n21259), .B1(n20986), .B2(n21258), .ZN(
        n20975) );
  AOI22_X1 U23916 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20988), .B1(
        n21017), .B2(n21207), .ZN(n20974) );
  OAI211_X1 U23917 ( .C1(n21210), .C2(n20991), .A(n20975), .B(n20974), .ZN(
        P1_U3091) );
  AOI22_X1 U23918 ( .A1(n20987), .A2(n21265), .B1(n20986), .B2(n21264), .ZN(
        n20977) );
  AOI22_X1 U23919 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20988), .B1(
        n21017), .B2(n21211), .ZN(n20976) );
  OAI211_X1 U23920 ( .C1(n21214), .C2(n20991), .A(n20977), .B(n20976), .ZN(
        P1_U3092) );
  AOI22_X1 U23921 ( .A1(n20987), .A2(n21271), .B1(n20986), .B2(n21270), .ZN(
        n20979) );
  AOI22_X1 U23922 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20988), .B1(
        n21017), .B2(n21215), .ZN(n20978) );
  OAI211_X1 U23923 ( .C1(n21218), .C2(n20991), .A(n20979), .B(n20978), .ZN(
        P1_U3093) );
  AOI22_X1 U23924 ( .A1(n20987), .A2(n21277), .B1(n20986), .B2(n21276), .ZN(
        n20982) );
  AOI22_X1 U23925 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20988), .B1(
        n20980), .B2(n21278), .ZN(n20981) );
  OAI211_X1 U23926 ( .C1(n21281), .C2(n20983), .A(n20982), .B(n20981), .ZN(
        P1_U3094) );
  AOI22_X1 U23927 ( .A1(n20987), .A2(n21283), .B1(n20986), .B2(n21282), .ZN(
        n20985) );
  AOI22_X1 U23928 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20988), .B1(
        n21017), .B2(n21223), .ZN(n20984) );
  OAI211_X1 U23929 ( .C1(n21226), .C2(n20991), .A(n20985), .B(n20984), .ZN(
        P1_U3095) );
  AOI22_X1 U23930 ( .A1(n20987), .A2(n21290), .B1(n20986), .B2(n21288), .ZN(
        n20990) );
  AOI22_X1 U23931 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20988), .B1(
        n21017), .B2(n21229), .ZN(n20989) );
  OAI211_X1 U23932 ( .C1(n21234), .C2(n20991), .A(n20990), .B(n20989), .ZN(
        P1_U3096) );
  NOR3_X1 U23933 ( .A1(n21186), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21024) );
  INV_X1 U23934 ( .A(n21024), .ZN(n21021) );
  NOR2_X1 U23935 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21021), .ZN(
        n21015) );
  AOI21_X1 U23936 ( .B1(n21094), .B2(n21188), .A(n21015), .ZN(n20997) );
  NOR2_X1 U23937 ( .A1(n20995), .A2(n21052), .ZN(n21130) );
  INV_X1 U23938 ( .A(n21130), .ZN(n21132) );
  OAI22_X1 U23939 ( .A1(n20997), .A2(n21376), .B1(n21054), .B2(n21132), .ZN(
        n21016) );
  AOI22_X1 U23940 ( .A1(n21016), .A2(n21241), .B1(n21240), .B2(n21015), .ZN(
        n21002) );
  INV_X1 U23941 ( .A(n21045), .ZN(n20996) );
  OAI21_X1 U23942 ( .B1(n20996), .B2(n21017), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20998) );
  NAND2_X1 U23943 ( .A1(n20998), .A2(n20997), .ZN(n20999) );
  AOI22_X1 U23944 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n21018), .B1(
        n21017), .B2(n21248), .ZN(n21001) );
  OAI211_X1 U23945 ( .C1(n21251), .C2(n21045), .A(n21002), .B(n21001), .ZN(
        P1_U3097) );
  AOI22_X1 U23946 ( .A1(n21016), .A2(n21253), .B1(n21252), .B2(n21015), .ZN(
        n21004) );
  AOI22_X1 U23947 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n21018), .B1(
        n21017), .B2(n21254), .ZN(n21003) );
  OAI211_X1 U23948 ( .C1(n21257), .C2(n21045), .A(n21004), .B(n21003), .ZN(
        P1_U3098) );
  AOI22_X1 U23949 ( .A1(n21016), .A2(n21259), .B1(n21258), .B2(n21015), .ZN(
        n21006) );
  AOI22_X1 U23950 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n21018), .B1(
        n21017), .B2(n21260), .ZN(n21005) );
  OAI211_X1 U23951 ( .C1(n21263), .C2(n21045), .A(n21006), .B(n21005), .ZN(
        P1_U3099) );
  AOI22_X1 U23952 ( .A1(n21016), .A2(n21265), .B1(n21264), .B2(n21015), .ZN(
        n21008) );
  AOI22_X1 U23953 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n21018), .B1(
        n21017), .B2(n21266), .ZN(n21007) );
  OAI211_X1 U23954 ( .C1(n21269), .C2(n21045), .A(n21008), .B(n21007), .ZN(
        P1_U3100) );
  AOI22_X1 U23955 ( .A1(n21016), .A2(n21271), .B1(n21270), .B2(n21015), .ZN(
        n21010) );
  AOI22_X1 U23956 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n21018), .B1(
        n21017), .B2(n21272), .ZN(n21009) );
  OAI211_X1 U23957 ( .C1(n21275), .C2(n21045), .A(n21010), .B(n21009), .ZN(
        P1_U3101) );
  AOI22_X1 U23958 ( .A1(n21016), .A2(n21277), .B1(n21276), .B2(n21015), .ZN(
        n21012) );
  AOI22_X1 U23959 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n21018), .B1(
        n21017), .B2(n21278), .ZN(n21011) );
  OAI211_X1 U23960 ( .C1(n21281), .C2(n21045), .A(n21012), .B(n21011), .ZN(
        P1_U3102) );
  AOI22_X1 U23961 ( .A1(n21016), .A2(n21283), .B1(n21282), .B2(n21015), .ZN(
        n21014) );
  AOI22_X1 U23962 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n21018), .B1(
        n21017), .B2(n21284), .ZN(n21013) );
  OAI211_X1 U23963 ( .C1(n21287), .C2(n21045), .A(n21014), .B(n21013), .ZN(
        P1_U3103) );
  AOI22_X1 U23964 ( .A1(n21016), .A2(n21290), .B1(n21288), .B2(n21015), .ZN(
        n21020) );
  AOI22_X1 U23965 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n21018), .B1(
        n21017), .B2(n21292), .ZN(n21019) );
  OAI211_X1 U23966 ( .C1(n21298), .C2(n21045), .A(n21020), .B(n21019), .ZN(
        P1_U3104) );
  NOR2_X1 U23967 ( .A1(n21157), .A2(n21021), .ZN(n21039) );
  AOI21_X1 U23968 ( .B1(n21094), .B2(n21158), .A(n21039), .ZN(n21022) );
  OAI22_X1 U23969 ( .A1(n21022), .A2(n21376), .B1(n21021), .B2(n21239), .ZN(
        n21040) );
  AOI22_X1 U23970 ( .A1(n21040), .A2(n21241), .B1(n21240), .B2(n21039), .ZN(
        n21026) );
  OAI211_X1 U23971 ( .C1(n21097), .C2(n21191), .A(n21163), .B(n21022), .ZN(
        n21023) );
  AOI22_X1 U23972 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n21042), .B1(
        n21041), .B2(n21199), .ZN(n21025) );
  OAI211_X1 U23973 ( .C1(n21202), .C2(n21045), .A(n21026), .B(n21025), .ZN(
        P1_U3105) );
  AOI22_X1 U23974 ( .A1(n21040), .A2(n21253), .B1(n21252), .B2(n21039), .ZN(
        n21028) );
  AOI22_X1 U23975 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n21042), .B1(
        n21041), .B2(n21203), .ZN(n21027) );
  OAI211_X1 U23976 ( .C1(n21206), .C2(n21045), .A(n21028), .B(n21027), .ZN(
        P1_U3106) );
  AOI22_X1 U23977 ( .A1(n21040), .A2(n21259), .B1(n21258), .B2(n21039), .ZN(
        n21030) );
  AOI22_X1 U23978 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n21042), .B1(
        n21041), .B2(n21207), .ZN(n21029) );
  OAI211_X1 U23979 ( .C1(n21210), .C2(n21045), .A(n21030), .B(n21029), .ZN(
        P1_U3107) );
  AOI22_X1 U23980 ( .A1(n21040), .A2(n21265), .B1(n21264), .B2(n21039), .ZN(
        n21032) );
  AOI22_X1 U23981 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n21042), .B1(
        n21041), .B2(n21211), .ZN(n21031) );
  OAI211_X1 U23982 ( .C1(n21214), .C2(n21045), .A(n21032), .B(n21031), .ZN(
        P1_U3108) );
  AOI22_X1 U23983 ( .A1(n21040), .A2(n21271), .B1(n21270), .B2(n21039), .ZN(
        n21034) );
  AOI22_X1 U23984 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n21042), .B1(
        n21041), .B2(n21215), .ZN(n21033) );
  OAI211_X1 U23985 ( .C1(n21218), .C2(n21045), .A(n21034), .B(n21033), .ZN(
        P1_U3109) );
  AOI22_X1 U23986 ( .A1(n21040), .A2(n21277), .B1(n21276), .B2(n21039), .ZN(
        n21036) );
  AOI22_X1 U23987 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n21042), .B1(
        n21041), .B2(n21219), .ZN(n21035) );
  OAI211_X1 U23988 ( .C1(n21222), .C2(n21045), .A(n21036), .B(n21035), .ZN(
        P1_U3110) );
  AOI22_X1 U23989 ( .A1(n21040), .A2(n21283), .B1(n21282), .B2(n21039), .ZN(
        n21038) );
  AOI22_X1 U23990 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n21042), .B1(
        n21041), .B2(n21223), .ZN(n21037) );
  OAI211_X1 U23991 ( .C1(n21226), .C2(n21045), .A(n21038), .B(n21037), .ZN(
        P1_U3111) );
  AOI22_X1 U23992 ( .A1(n21040), .A2(n21290), .B1(n21288), .B2(n21039), .ZN(
        n21044) );
  AOI22_X1 U23993 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n21042), .B1(
        n21041), .B2(n21229), .ZN(n21043) );
  OAI211_X1 U23994 ( .C1(n21234), .C2(n21045), .A(n21044), .B(n21043), .ZN(
        P1_U3112) );
  NOR3_X1 U23995 ( .A1(n21186), .A2(n13998), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21099) );
  NAND2_X1 U23996 ( .A1(n21157), .A2(n21099), .ZN(n21084) );
  OAI22_X1 U23997 ( .A1(n21115), .A2(n21251), .B1(n21084), .B2(n21046), .ZN(
        n21047) );
  INV_X1 U23998 ( .A(n21047), .ZN(n21058) );
  NAND2_X1 U23999 ( .A1(n21115), .A2(n21085), .ZN(n21048) );
  AOI21_X1 U24000 ( .B1(n21048), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21376), 
        .ZN(n21051) );
  NAND2_X1 U24001 ( .A1(n21094), .A2(n21194), .ZN(n21055) );
  AOI22_X1 U24002 ( .A1(n21051), .A2(n21055), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21084), .ZN(n21049) );
  OAI21_X1 U24003 ( .B1(n21186), .B2(n21184), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n21196) );
  NAND3_X1 U24004 ( .A1(n21050), .A2(n21049), .A3(n21196), .ZN(n21088) );
  INV_X1 U24005 ( .A(n21051), .ZN(n21056) );
  NAND2_X1 U24006 ( .A1(n21052), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21053) );
  AOI22_X1 U24007 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n21088), .B1(
        n21241), .B2(n21087), .ZN(n21057) );
  OAI211_X1 U24008 ( .C1(n21202), .C2(n21085), .A(n21058), .B(n21057), .ZN(
        P1_U3113) );
  OAI22_X1 U24009 ( .A1(n21115), .A2(n21257), .B1(n21084), .B2(n21059), .ZN(
        n21060) );
  INV_X1 U24010 ( .A(n21060), .ZN(n21062) );
  AOI22_X1 U24011 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n21088), .B1(
        n21253), .B2(n21087), .ZN(n21061) );
  OAI211_X1 U24012 ( .C1(n21206), .C2(n21085), .A(n21062), .B(n21061), .ZN(
        P1_U3114) );
  OAI22_X1 U24013 ( .A1(n21085), .A2(n21210), .B1(n21084), .B2(n21063), .ZN(
        n21064) );
  INV_X1 U24014 ( .A(n21064), .ZN(n21066) );
  AOI22_X1 U24015 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n21088), .B1(
        n21259), .B2(n21087), .ZN(n21065) );
  OAI211_X1 U24016 ( .C1(n21263), .C2(n21115), .A(n21066), .B(n21065), .ZN(
        P1_U3115) );
  OAI22_X1 U24017 ( .A1(n21115), .A2(n21269), .B1(n21084), .B2(n21067), .ZN(
        n21068) );
  INV_X1 U24018 ( .A(n21068), .ZN(n21070) );
  AOI22_X1 U24019 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n21088), .B1(
        n21265), .B2(n21087), .ZN(n21069) );
  OAI211_X1 U24020 ( .C1(n21214), .C2(n21085), .A(n21070), .B(n21069), .ZN(
        P1_U3116) );
  OAI22_X1 U24021 ( .A1(n21085), .A2(n21218), .B1(n21084), .B2(n21071), .ZN(
        n21072) );
  INV_X1 U24022 ( .A(n21072), .ZN(n21074) );
  AOI22_X1 U24023 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n21088), .B1(
        n21271), .B2(n21087), .ZN(n21073) );
  OAI211_X1 U24024 ( .C1(n21275), .C2(n21115), .A(n21074), .B(n21073), .ZN(
        P1_U3117) );
  OAI22_X1 U24025 ( .A1(n21115), .A2(n21281), .B1(n21084), .B2(n21075), .ZN(
        n21076) );
  INV_X1 U24026 ( .A(n21076), .ZN(n21078) );
  AOI22_X1 U24027 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n21088), .B1(
        n21277), .B2(n21087), .ZN(n21077) );
  OAI211_X1 U24028 ( .C1(n21222), .C2(n21085), .A(n21078), .B(n21077), .ZN(
        P1_U3118) );
  OAI22_X1 U24029 ( .A1(n21085), .A2(n21226), .B1(n21084), .B2(n21079), .ZN(
        n21080) );
  INV_X1 U24030 ( .A(n21080), .ZN(n21082) );
  AOI22_X1 U24031 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n21088), .B1(
        n21283), .B2(n21087), .ZN(n21081) );
  OAI211_X1 U24032 ( .C1(n21287), .C2(n21115), .A(n21082), .B(n21081), .ZN(
        P1_U3119) );
  OAI22_X1 U24033 ( .A1(n21085), .A2(n21234), .B1(n21084), .B2(n21083), .ZN(
        n21086) );
  INV_X1 U24034 ( .A(n21086), .ZN(n21090) );
  AOI22_X1 U24035 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n21088), .B1(
        n21290), .B2(n21087), .ZN(n21089) );
  OAI211_X1 U24036 ( .C1(n21298), .C2(n21115), .A(n21090), .B(n21089), .ZN(
        P1_U3120) );
  NOR2_X1 U24037 ( .A1(n21093), .A2(n21186), .ZN(n21116) );
  AOI21_X1 U24038 ( .B1(n21094), .B2(n21236), .A(n21116), .ZN(n21096) );
  INV_X1 U24039 ( .A(n21099), .ZN(n21095) );
  OAI22_X1 U24040 ( .A1(n21096), .A2(n21376), .B1(n21095), .B2(n21239), .ZN(
        n21117) );
  AOI22_X1 U24041 ( .A1(n21117), .A2(n21241), .B1(n21240), .B2(n21116), .ZN(
        n21101) );
  OAI211_X1 U24042 ( .C1(n21097), .C2(n21243), .A(n21163), .B(n21096), .ZN(
        n21098) );
  AOI22_X1 U24043 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n21119), .B1(
        n21118), .B2(n21248), .ZN(n21100) );
  OAI211_X1 U24044 ( .C1(n21251), .C2(n21154), .A(n21101), .B(n21100), .ZN(
        P1_U3121) );
  AOI22_X1 U24045 ( .A1(n21117), .A2(n21253), .B1(n21252), .B2(n21116), .ZN(
        n21103) );
  AOI22_X1 U24046 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n21119), .B1(
        n21118), .B2(n21254), .ZN(n21102) );
  OAI211_X1 U24047 ( .C1(n21257), .C2(n21154), .A(n21103), .B(n21102), .ZN(
        P1_U3122) );
  AOI22_X1 U24048 ( .A1(n21117), .A2(n21259), .B1(n21258), .B2(n21116), .ZN(
        n21105) );
  INV_X1 U24049 ( .A(n21154), .ZN(n21112) );
  AOI22_X1 U24050 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n21119), .B1(
        n21112), .B2(n21207), .ZN(n21104) );
  OAI211_X1 U24051 ( .C1(n21210), .C2(n21115), .A(n21105), .B(n21104), .ZN(
        P1_U3123) );
  AOI22_X1 U24052 ( .A1(n21117), .A2(n21265), .B1(n21264), .B2(n21116), .ZN(
        n21107) );
  AOI22_X1 U24053 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n21119), .B1(
        n21112), .B2(n21211), .ZN(n21106) );
  OAI211_X1 U24054 ( .C1(n21214), .C2(n21115), .A(n21107), .B(n21106), .ZN(
        P1_U3124) );
  AOI22_X1 U24055 ( .A1(n21117), .A2(n21271), .B1(n21270), .B2(n21116), .ZN(
        n21109) );
  AOI22_X1 U24056 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n21119), .B1(
        n21118), .B2(n21272), .ZN(n21108) );
  OAI211_X1 U24057 ( .C1(n21275), .C2(n21154), .A(n21109), .B(n21108), .ZN(
        P1_U3125) );
  AOI22_X1 U24058 ( .A1(n21117), .A2(n21277), .B1(n21276), .B2(n21116), .ZN(
        n21111) );
  AOI22_X1 U24059 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n21119), .B1(
        n21118), .B2(n21278), .ZN(n21110) );
  OAI211_X1 U24060 ( .C1(n21281), .C2(n21154), .A(n21111), .B(n21110), .ZN(
        P1_U3126) );
  AOI22_X1 U24061 ( .A1(n21117), .A2(n21283), .B1(n21282), .B2(n21116), .ZN(
        n21114) );
  AOI22_X1 U24062 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n21119), .B1(
        n21112), .B2(n21223), .ZN(n21113) );
  OAI211_X1 U24063 ( .C1(n21226), .C2(n21115), .A(n21114), .B(n21113), .ZN(
        P1_U3127) );
  AOI22_X1 U24064 ( .A1(n21117), .A2(n21290), .B1(n21288), .B2(n21116), .ZN(
        n21121) );
  AOI22_X1 U24065 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n21119), .B1(
        n21118), .B2(n21292), .ZN(n21120) );
  OAI211_X1 U24066 ( .C1(n21298), .C2(n21154), .A(n21121), .B(n21120), .ZN(
        P1_U3128) );
  NOR3_X1 U24067 ( .A1(n21123), .A2(n21186), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21162) );
  NAND2_X1 U24068 ( .A1(n21157), .A2(n21162), .ZN(n21128) );
  INV_X1 U24069 ( .A(n21128), .ZN(n21149) );
  AOI22_X1 U24070 ( .A1(n21180), .A2(n21199), .B1(n21149), .B2(n21240), .ZN(
        n21136) );
  INV_X1 U24071 ( .A(n21180), .ZN(n21124) );
  NAND2_X1 U24072 ( .A1(n21124), .A2(n21154), .ZN(n21125) );
  AOI21_X1 U24073 ( .B1(n21125), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21376), 
        .ZN(n21131) );
  NAND2_X1 U24074 ( .A1(n21237), .A2(n21188), .ZN(n21133) );
  AOI22_X1 U24075 ( .A1(n21131), .A2(n21133), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21128), .ZN(n21129) );
  INV_X1 U24076 ( .A(n21131), .ZN(n21134) );
  AOI22_X1 U24077 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n21151), .B1(
        n21241), .B2(n21150), .ZN(n21135) );
  OAI211_X1 U24078 ( .C1(n21202), .C2(n21154), .A(n21136), .B(n21135), .ZN(
        P1_U3129) );
  AOI22_X1 U24079 ( .A1(n21180), .A2(n21203), .B1(n21149), .B2(n21252), .ZN(
        n21138) );
  AOI22_X1 U24080 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n21151), .B1(
        n21253), .B2(n21150), .ZN(n21137) );
  OAI211_X1 U24081 ( .C1(n21206), .C2(n21154), .A(n21138), .B(n21137), .ZN(
        P1_U3130) );
  AOI22_X1 U24082 ( .A1(n21180), .A2(n21207), .B1(n21149), .B2(n21258), .ZN(
        n21140) );
  AOI22_X1 U24083 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n21151), .B1(
        n21259), .B2(n21150), .ZN(n21139) );
  OAI211_X1 U24084 ( .C1(n21210), .C2(n21154), .A(n21140), .B(n21139), .ZN(
        P1_U3131) );
  AOI22_X1 U24085 ( .A1(n21180), .A2(n21211), .B1(n21149), .B2(n21264), .ZN(
        n21142) );
  AOI22_X1 U24086 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n21151), .B1(
        n21265), .B2(n21150), .ZN(n21141) );
  OAI211_X1 U24087 ( .C1(n21214), .C2(n21154), .A(n21142), .B(n21141), .ZN(
        P1_U3132) );
  AOI22_X1 U24088 ( .A1(n21180), .A2(n21215), .B1(n21149), .B2(n21270), .ZN(
        n21144) );
  AOI22_X1 U24089 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n21151), .B1(
        n21271), .B2(n21150), .ZN(n21143) );
  OAI211_X1 U24090 ( .C1(n21218), .C2(n21154), .A(n21144), .B(n21143), .ZN(
        P1_U3133) );
  AOI22_X1 U24091 ( .A1(n21180), .A2(n21219), .B1(n21149), .B2(n21276), .ZN(
        n21146) );
  AOI22_X1 U24092 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n21151), .B1(
        n21277), .B2(n21150), .ZN(n21145) );
  OAI211_X1 U24093 ( .C1(n21222), .C2(n21154), .A(n21146), .B(n21145), .ZN(
        P1_U3134) );
  AOI22_X1 U24094 ( .A1(n21180), .A2(n21223), .B1(n21149), .B2(n21282), .ZN(
        n21148) );
  AOI22_X1 U24095 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n21151), .B1(
        n21283), .B2(n21150), .ZN(n21147) );
  OAI211_X1 U24096 ( .C1(n21226), .C2(n21154), .A(n21148), .B(n21147), .ZN(
        P1_U3135) );
  AOI22_X1 U24097 ( .A1(n21180), .A2(n21229), .B1(n21149), .B2(n21288), .ZN(
        n21153) );
  AOI22_X1 U24098 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n21151), .B1(
        n21290), .B2(n21150), .ZN(n21152) );
  OAI211_X1 U24099 ( .C1(n21234), .C2(n21154), .A(n21153), .B(n21152), .ZN(
        P1_U3136) );
  INV_X1 U24100 ( .A(n21162), .ZN(n21159) );
  NOR2_X1 U24101 ( .A1(n21157), .A2(n21159), .ZN(n21178) );
  AOI21_X1 U24102 ( .B1(n21237), .B2(n21158), .A(n21178), .ZN(n21160) );
  OAI22_X1 U24103 ( .A1(n21160), .A2(n21376), .B1(n21159), .B2(n21239), .ZN(
        n21179) );
  AOI22_X1 U24104 ( .A1(n21179), .A2(n21241), .B1(n21240), .B2(n21178), .ZN(
        n21165) );
  OAI211_X1 U24105 ( .C1(n21244), .C2(n21191), .A(n21163), .B(n21160), .ZN(
        n21161) );
  AOI22_X1 U24106 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n21181), .B1(
        n21180), .B2(n21248), .ZN(n21164) );
  OAI211_X1 U24107 ( .C1(n21251), .C2(n21233), .A(n21165), .B(n21164), .ZN(
        P1_U3137) );
  AOI22_X1 U24108 ( .A1(n21179), .A2(n21253), .B1(n21252), .B2(n21178), .ZN(
        n21167) );
  AOI22_X1 U24109 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n21181), .B1(
        n21180), .B2(n21254), .ZN(n21166) );
  OAI211_X1 U24110 ( .C1(n21257), .C2(n21233), .A(n21167), .B(n21166), .ZN(
        P1_U3138) );
  AOI22_X1 U24111 ( .A1(n21179), .A2(n21259), .B1(n21258), .B2(n21178), .ZN(
        n21169) );
  AOI22_X1 U24112 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n21181), .B1(
        n21180), .B2(n21260), .ZN(n21168) );
  OAI211_X1 U24113 ( .C1(n21263), .C2(n21233), .A(n21169), .B(n21168), .ZN(
        P1_U3139) );
  AOI22_X1 U24114 ( .A1(n21179), .A2(n21265), .B1(n21264), .B2(n21178), .ZN(
        n21171) );
  AOI22_X1 U24115 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21181), .B1(
        n21180), .B2(n21266), .ZN(n21170) );
  OAI211_X1 U24116 ( .C1(n21269), .C2(n21233), .A(n21171), .B(n21170), .ZN(
        P1_U3140) );
  AOI22_X1 U24117 ( .A1(n21179), .A2(n21271), .B1(n21270), .B2(n21178), .ZN(
        n21173) );
  AOI22_X1 U24118 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n21181), .B1(
        n21180), .B2(n21272), .ZN(n21172) );
  OAI211_X1 U24119 ( .C1(n21275), .C2(n21233), .A(n21173), .B(n21172), .ZN(
        P1_U3141) );
  AOI22_X1 U24120 ( .A1(n21179), .A2(n21277), .B1(n21276), .B2(n21178), .ZN(
        n21175) );
  AOI22_X1 U24121 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n21181), .B1(
        n21180), .B2(n21278), .ZN(n21174) );
  OAI211_X1 U24122 ( .C1(n21281), .C2(n21233), .A(n21175), .B(n21174), .ZN(
        P1_U3142) );
  AOI22_X1 U24123 ( .A1(n21179), .A2(n21283), .B1(n21282), .B2(n21178), .ZN(
        n21177) );
  AOI22_X1 U24124 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n21181), .B1(
        n21180), .B2(n21284), .ZN(n21176) );
  OAI211_X1 U24125 ( .C1(n21287), .C2(n21233), .A(n21177), .B(n21176), .ZN(
        P1_U3143) );
  AOI22_X1 U24126 ( .A1(n21179), .A2(n21290), .B1(n21288), .B2(n21178), .ZN(
        n21183) );
  AOI22_X1 U24127 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n21181), .B1(
        n21180), .B2(n21292), .ZN(n21182) );
  OAI211_X1 U24128 ( .C1(n21298), .C2(n21233), .A(n21183), .B(n21182), .ZN(
        P1_U3144) );
  INV_X1 U24129 ( .A(n21237), .ZN(n21187) );
  OAI33_X1 U24130 ( .A1(n21188), .A2(n21187), .A3(n21376), .B1(n21186), .B2(
        n21185), .B3(n21184), .ZN(n21228) );
  INV_X1 U24131 ( .A(n21247), .ZN(n21238) );
  NOR2_X1 U24132 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21238), .ZN(
        n21227) );
  AOI22_X1 U24133 ( .A1(n9778), .A2(n21241), .B1(n21240), .B2(n21227), .ZN(
        n21201) );
  INV_X1 U24134 ( .A(n21189), .ZN(n21190) );
  INV_X1 U24135 ( .A(n21293), .ZN(n21192) );
  AOI21_X1 U24136 ( .B1(n21192), .B2(n21233), .A(n21191), .ZN(n21193) );
  AOI21_X1 U24137 ( .B1(n21237), .B2(n21194), .A(n21193), .ZN(n21195) );
  NOR2_X1 U24138 ( .A1(n21195), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21198) );
  AOI22_X1 U24139 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n21230), .B1(
        n21293), .B2(n21199), .ZN(n21200) );
  OAI211_X1 U24140 ( .C1(n21202), .C2(n21233), .A(n21201), .B(n21200), .ZN(
        P1_U3145) );
  AOI22_X1 U24141 ( .A1(n9778), .A2(n21253), .B1(n21252), .B2(n21227), .ZN(
        n21205) );
  AOI22_X1 U24142 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21230), .B1(
        n21293), .B2(n21203), .ZN(n21204) );
  OAI211_X1 U24143 ( .C1(n21206), .C2(n21233), .A(n21205), .B(n21204), .ZN(
        P1_U3146) );
  AOI22_X1 U24144 ( .A1(n9778), .A2(n21259), .B1(n21258), .B2(n21227), .ZN(
        n21209) );
  AOI22_X1 U24145 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n21230), .B1(
        n21293), .B2(n21207), .ZN(n21208) );
  OAI211_X1 U24146 ( .C1(n21210), .C2(n21233), .A(n21209), .B(n21208), .ZN(
        P1_U3147) );
  AOI22_X1 U24147 ( .A1(n9778), .A2(n21265), .B1(n21264), .B2(n21227), .ZN(
        n21213) );
  AOI22_X1 U24148 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n21230), .B1(
        n21293), .B2(n21211), .ZN(n21212) );
  OAI211_X1 U24149 ( .C1(n21214), .C2(n21233), .A(n21213), .B(n21212), .ZN(
        P1_U3148) );
  AOI22_X1 U24150 ( .A1(n9778), .A2(n21271), .B1(n21270), .B2(n21227), .ZN(
        n21217) );
  AOI22_X1 U24151 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n21230), .B1(
        n21293), .B2(n21215), .ZN(n21216) );
  OAI211_X1 U24152 ( .C1(n21218), .C2(n21233), .A(n21217), .B(n21216), .ZN(
        P1_U3149) );
  AOI22_X1 U24153 ( .A1(n9778), .A2(n21277), .B1(n21276), .B2(n21227), .ZN(
        n21221) );
  AOI22_X1 U24154 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n21230), .B1(
        n21293), .B2(n21219), .ZN(n21220) );
  OAI211_X1 U24155 ( .C1(n21222), .C2(n21233), .A(n21221), .B(n21220), .ZN(
        P1_U3150) );
  AOI22_X1 U24156 ( .A1(n9778), .A2(n21283), .B1(n21282), .B2(n21227), .ZN(
        n21225) );
  AOI22_X1 U24157 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n21230), .B1(
        n21293), .B2(n21223), .ZN(n21224) );
  OAI211_X1 U24158 ( .C1(n21226), .C2(n21233), .A(n21225), .B(n21224), .ZN(
        P1_U3151) );
  AOI22_X1 U24159 ( .A1(n9778), .A2(n21290), .B1(n21288), .B2(n21227), .ZN(
        n21232) );
  AOI22_X1 U24160 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n21230), .B1(
        n21293), .B2(n21229), .ZN(n21231) );
  OAI211_X1 U24161 ( .C1(n21234), .C2(n21233), .A(n21232), .B(n21231), .ZN(
        P1_U3152) );
  INV_X1 U24162 ( .A(n21235), .ZN(n21289) );
  AOI21_X1 U24163 ( .B1(n21237), .B2(n21236), .A(n21289), .ZN(n21242) );
  OAI22_X1 U24164 ( .A1(n21242), .A2(n21376), .B1(n21239), .B2(n21238), .ZN(
        n21291) );
  AOI22_X1 U24165 ( .A1(n21291), .A2(n21241), .B1(n21289), .B2(n21240), .ZN(
        n21250) );
  OAI211_X1 U24166 ( .C1(n21244), .C2(n21243), .A(n21163), .B(n21242), .ZN(
        n21246) );
  AOI22_X1 U24167 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21294), .B1(
        n21293), .B2(n21248), .ZN(n21249) );
  OAI211_X1 U24168 ( .C1(n21251), .C2(n21297), .A(n21250), .B(n21249), .ZN(
        P1_U3153) );
  AOI22_X1 U24169 ( .A1(n21291), .A2(n21253), .B1(n21289), .B2(n21252), .ZN(
        n21256) );
  AOI22_X1 U24170 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21294), .B1(
        n21293), .B2(n21254), .ZN(n21255) );
  OAI211_X1 U24171 ( .C1(n21257), .C2(n21297), .A(n21256), .B(n21255), .ZN(
        P1_U3154) );
  AOI22_X1 U24172 ( .A1(n21291), .A2(n21259), .B1(n21289), .B2(n21258), .ZN(
        n21262) );
  AOI22_X1 U24173 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21294), .B1(
        n21293), .B2(n21260), .ZN(n21261) );
  OAI211_X1 U24174 ( .C1(n21263), .C2(n21297), .A(n21262), .B(n21261), .ZN(
        P1_U3155) );
  AOI22_X1 U24175 ( .A1(n21291), .A2(n21265), .B1(n21289), .B2(n21264), .ZN(
        n21268) );
  AOI22_X1 U24176 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21294), .B1(
        n21293), .B2(n21266), .ZN(n21267) );
  OAI211_X1 U24177 ( .C1(n21269), .C2(n21297), .A(n21268), .B(n21267), .ZN(
        P1_U3156) );
  AOI22_X1 U24178 ( .A1(n21291), .A2(n21271), .B1(n21289), .B2(n21270), .ZN(
        n21274) );
  AOI22_X1 U24179 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21294), .B1(
        n21293), .B2(n21272), .ZN(n21273) );
  OAI211_X1 U24180 ( .C1(n21275), .C2(n21297), .A(n21274), .B(n21273), .ZN(
        P1_U3157) );
  AOI22_X1 U24181 ( .A1(n21291), .A2(n21277), .B1(n21289), .B2(n21276), .ZN(
        n21280) );
  AOI22_X1 U24182 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21294), .B1(
        n21293), .B2(n21278), .ZN(n21279) );
  OAI211_X1 U24183 ( .C1(n21281), .C2(n21297), .A(n21280), .B(n21279), .ZN(
        P1_U3158) );
  AOI22_X1 U24184 ( .A1(n21291), .A2(n21283), .B1(n21289), .B2(n21282), .ZN(
        n21286) );
  AOI22_X1 U24185 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21294), .B1(
        n21293), .B2(n21284), .ZN(n21285) );
  OAI211_X1 U24186 ( .C1(n21287), .C2(n21297), .A(n21286), .B(n21285), .ZN(
        P1_U3159) );
  AOI22_X1 U24187 ( .A1(n21291), .A2(n21290), .B1(n21289), .B2(n21288), .ZN(
        n21296) );
  AOI22_X1 U24188 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21294), .B1(
        n21293), .B2(n21292), .ZN(n21295) );
  OAI211_X1 U24189 ( .C1(n21298), .C2(n21297), .A(n21296), .B(n21295), .ZN(
        P1_U3160) );
  AND2_X1 U24190 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21299), .ZN(
        P1_U3164) );
  AND2_X1 U24191 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21299), .ZN(
        P1_U3165) );
  AND2_X1 U24192 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21299), .ZN(
        P1_U3166) );
  INV_X1 U24193 ( .A(P1_DATAWIDTH_REG_28__SCAN_IN), .ZN(n21431) );
  NOR2_X1 U24194 ( .A1(n21363), .A2(n21431), .ZN(P1_U3167) );
  AND2_X1 U24195 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21299), .ZN(
        P1_U3168) );
  AND2_X1 U24196 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21299), .ZN(
        P1_U3169) );
  AND2_X1 U24197 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21299), .ZN(
        P1_U3170) );
  AND2_X1 U24198 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21299), .ZN(
        P1_U3171) );
  AND2_X1 U24199 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21299), .ZN(
        P1_U3172) );
  AND2_X1 U24200 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21299), .ZN(
        P1_U3173) );
  AND2_X1 U24201 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21299), .ZN(
        P1_U3174) );
  AND2_X1 U24202 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21299), .ZN(
        P1_U3175) );
  INV_X1 U24203 ( .A(P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n21482) );
  NOR2_X1 U24204 ( .A1(n21363), .A2(n21482), .ZN(P1_U3176) );
  AND2_X1 U24205 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21299), .ZN(
        P1_U3177) );
  AND2_X1 U24206 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21299), .ZN(
        P1_U3178) );
  AND2_X1 U24207 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21299), .ZN(
        P1_U3179) );
  AND2_X1 U24208 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21299), .ZN(
        P1_U3180) );
  AND2_X1 U24209 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21299), .ZN(
        P1_U3181) );
  AND2_X1 U24210 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21299), .ZN(
        P1_U3182) );
  AND2_X1 U24211 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21299), .ZN(
        P1_U3183) );
  AND2_X1 U24212 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21299), .ZN(
        P1_U3184) );
  AND2_X1 U24213 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21299), .ZN(
        P1_U3185) );
  AND2_X1 U24214 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21299), .ZN(P1_U3186) );
  INV_X1 U24215 ( .A(P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n21527) );
  NOR2_X1 U24216 ( .A1(n21363), .A2(n21527), .ZN(P1_U3187) );
  AND2_X1 U24217 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21299), .ZN(P1_U3188) );
  AND2_X1 U24218 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21299), .ZN(P1_U3189) );
  AND2_X1 U24219 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21299), .ZN(P1_U3190) );
  AND2_X1 U24220 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21299), .ZN(P1_U3191) );
  AND2_X1 U24221 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21299), .ZN(P1_U3192) );
  AND2_X1 U24222 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21299), .ZN(P1_U3193) );
  AOI21_X1 U24223 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21379), .A(n21312), 
        .ZN(n21314) );
  OAI22_X1 U24224 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21307), .B1(n21315), 
        .B2(n21300), .ZN(n21301) );
  NOR3_X1 U24225 ( .A1(n21302), .A2(n21310), .A3(n21301), .ZN(n21303) );
  OAI22_X1 U24226 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21314), .B1(n21375), 
        .B2(n21303), .ZN(P1_U3194) );
  NOR2_X1 U24227 ( .A1(n21304), .A2(n21315), .ZN(n21305) );
  AOI221_X1 U24228 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n21307), .C1(n21306), 
        .C2(n21307), .A(n21305), .ZN(n21313) );
  OAI211_X1 U24229 ( .C1(NA), .C2(n21308), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n21315), .ZN(n21309) );
  OAI211_X1 U24230 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21310), .A(HOLD), .B(
        n21309), .ZN(n21311) );
  OAI22_X1 U24231 ( .A1(n21314), .A2(n21313), .B1(n21312), .B2(n21311), .ZN(
        P1_U3196) );
  NOR2_X1 U24232 ( .A1(n21389), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21342) );
  INV_X1 U24233 ( .A(n21342), .ZN(n21357) );
  INV_X1 U24234 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n21497) );
  INV_X1 U24235 ( .A(n21355), .ZN(n21353) );
  OAI222_X1 U24236 ( .A1(n21357), .A2(n13835), .B1(n21497), .B2(n21375), .C1(
        n15005), .C2(n21353), .ZN(P1_U3197) );
  AOI222_X1 U24237 ( .A1(n21355), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n21342), .ZN(n21316) );
  INV_X1 U24238 ( .A(n21316), .ZN(P1_U3198) );
  INV_X1 U24239 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21498) );
  OAI222_X1 U24240 ( .A1(n21353), .A2(n14230), .B1(n21498), .B2(n21375), .C1(
        n21317), .C2(n21357), .ZN(P1_U3199) );
  AOI222_X1 U24241 ( .A1(n21351), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n21355), .ZN(n21318) );
  INV_X1 U24242 ( .A(n21318), .ZN(P1_U3200) );
  OAI222_X1 U24243 ( .A1(n21353), .A2(n21320), .B1(n21319), .B2(n21375), .C1(
        n17365), .C2(n21357), .ZN(P1_U3201) );
  AOI222_X1 U24244 ( .A1(n21355), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n21342), .ZN(n21321) );
  INV_X1 U24245 ( .A(n21321), .ZN(P1_U3202) );
  AOI222_X1 U24246 ( .A1(n21355), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n21351), .ZN(n21322) );
  INV_X1 U24247 ( .A(n21322), .ZN(P1_U3203) );
  AOI222_X1 U24248 ( .A1(n21351), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n21355), .ZN(n21323) );
  INV_X1 U24249 ( .A(n21323), .ZN(P1_U3204) );
  AOI222_X1 U24250 ( .A1(n21355), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n21351), .ZN(n21324) );
  INV_X1 U24251 ( .A(n21324), .ZN(P1_U3205) );
  AOI222_X1 U24252 ( .A1(n21342), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n21355), .ZN(n21325) );
  INV_X1 U24253 ( .A(n21325), .ZN(P1_U3206) );
  AOI222_X1 U24254 ( .A1(n21355), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n21351), .ZN(n21326) );
  INV_X1 U24255 ( .A(n21326), .ZN(P1_U3207) );
  AOI22_X1 U24256 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n21389), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(n21342), .ZN(n21327) );
  OAI21_X1 U24257 ( .B1(n21328), .B2(n21353), .A(n21327), .ZN(P1_U3208) );
  AOI22_X1 U24258 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n21389), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(n21355), .ZN(n21329) );
  OAI21_X1 U24259 ( .B1(n21330), .B2(n21357), .A(n21329), .ZN(P1_U3209) );
  AOI222_X1 U24260 ( .A1(n21342), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n21355), .ZN(n21331) );
  INV_X1 U24261 ( .A(n21331), .ZN(P1_U3210) );
  AOI222_X1 U24262 ( .A1(n21355), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n21351), .ZN(n21332) );
  INV_X1 U24263 ( .A(n21332), .ZN(P1_U3211) );
  AOI222_X1 U24264 ( .A1(n21355), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n21351), .ZN(n21333) );
  INV_X1 U24265 ( .A(n21333), .ZN(P1_U3212) );
  AOI222_X1 U24266 ( .A1(n21351), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n21355), .ZN(n21334) );
  INV_X1 U24267 ( .A(n21334), .ZN(P1_U3213) );
  AOI222_X1 U24268 ( .A1(n21355), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n21351), .ZN(n21335) );
  INV_X1 U24269 ( .A(n21335), .ZN(P1_U3214) );
  AOI222_X1 U24270 ( .A1(n21355), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n21351), .ZN(n21336) );
  INV_X1 U24271 ( .A(n21336), .ZN(P1_U3215) );
  AOI222_X1 U24272 ( .A1(n21355), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n21351), .ZN(n21337) );
  INV_X1 U24273 ( .A(n21337), .ZN(P1_U3216) );
  AOI222_X1 U24274 ( .A1(n21351), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n21355), .ZN(n21338) );
  INV_X1 U24275 ( .A(n21338), .ZN(P1_U3217) );
  AOI22_X1 U24276 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n21389), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21342), .ZN(n21339) );
  OAI21_X1 U24277 ( .B1(n21340), .B2(n21353), .A(n21339), .ZN(P1_U3218) );
  AOI22_X1 U24278 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n21389), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21355), .ZN(n21341) );
  OAI21_X1 U24279 ( .B1(n21344), .B2(n21357), .A(n21341), .ZN(P1_U3219) );
  AOI22_X1 U24280 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n21342), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n21373), .ZN(n21343) );
  OAI21_X1 U24281 ( .B1(n21344), .B2(n21353), .A(n21343), .ZN(P1_U3220) );
  INV_X1 U24282 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21347) );
  AOI22_X1 U24283 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n21355), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21373), .ZN(n21345) );
  OAI21_X1 U24284 ( .B1(n21347), .B2(n21357), .A(n21345), .ZN(P1_U3221) );
  AOI22_X1 U24285 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n21351), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21373), .ZN(n21346) );
  OAI21_X1 U24286 ( .B1(n21347), .B2(n21353), .A(n21346), .ZN(P1_U3222) );
  AOI22_X1 U24287 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n21355), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21373), .ZN(n21348) );
  OAI21_X1 U24288 ( .B1(n21349), .B2(n21357), .A(n21348), .ZN(P1_U3223) );
  AOI222_X1 U24289 ( .A1(n21355), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21373), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21351), .ZN(n21350) );
  INV_X1 U24290 ( .A(n21350), .ZN(P1_U3224) );
  AOI22_X1 U24291 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n21351), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21373), .ZN(n21352) );
  OAI21_X1 U24292 ( .B1(n21354), .B2(n21353), .A(n21352), .ZN(P1_U3225) );
  AOI22_X1 U24293 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n21355), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21389), .ZN(n21356) );
  OAI21_X1 U24294 ( .B1(n21358), .B2(n21357), .A(n21356), .ZN(P1_U3226) );
  OAI22_X1 U24295 ( .A1(n21389), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21375), .ZN(n21359) );
  INV_X1 U24296 ( .A(n21359), .ZN(P1_U3458) );
  MUX2_X1 U24297 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .B(P1_BE_N_REG_2__SCAN_IN), .S(n21389), .Z(P1_U3459) );
  MUX2_X1 U24298 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .B(P1_BE_N_REG_1__SCAN_IN), .S(n21389), .Z(P1_U3460) );
  MUX2_X1 U24299 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .B(P1_BE_N_REG_0__SCAN_IN), .S(n21389), .Z(P1_U3461) );
  OAI21_X1 U24300 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21363), .A(n21361), 
        .ZN(n21360) );
  INV_X1 U24301 ( .A(n21360), .ZN(P1_U3464) );
  OAI21_X1 U24302 ( .B1(n21363), .B2(n21362), .A(n21361), .ZN(P1_U3465) );
  NAND2_X1 U24303 ( .A1(n21364), .A2(n15005), .ZN(n21370) );
  AND2_X1 U24304 ( .A1(n21371), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n21365) );
  AOI22_X1 U24305 ( .A1(P1_BYTEENABLE_REG_2__SCAN_IN), .A2(n21366), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(n21365), .ZN(n21367) );
  OAI221_X1 U24306 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21369), .C1(n21368), .C2(n21370), .A(n21367), .ZN(P1_U3481) );
  OAI21_X1 U24307 ( .B1(n21371), .B2(P1_BYTEENABLE_REG_0__SCAN_IN), .A(n21370), 
        .ZN(n21372) );
  INV_X1 U24308 ( .A(n21372), .ZN(P1_U3482) );
  AOI22_X1 U24309 ( .A1(n21375), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21374), 
        .B2(n21373), .ZN(P1_U3483) );
  OAI211_X1 U24310 ( .C1(n21379), .C2(n21378), .A(n21377), .B(n21376), .ZN(
        n21380) );
  INV_X1 U24311 ( .A(n21380), .ZN(n21381) );
  AND2_X1 U24312 ( .A1(n21382), .A2(n21381), .ZN(n21388) );
  OAI211_X1 U24313 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n12108), .A(n21383), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21385) );
  AOI21_X1 U24314 ( .B1(n21385), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n21384), 
        .ZN(n21387) );
  NAND2_X1 U24315 ( .A1(n21388), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21386) );
  OAI21_X1 U24316 ( .B1(n21388), .B2(n21387), .A(n21386), .ZN(P1_U3485) );
  MUX2_X1 U24317 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n21389), .Z(P1_U3486) );
  NAND4_X1 U24318 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_19__SCAN_IN), .A3(n21479), .A4(n21476), .ZN(n21394)
         );
  NAND4_X1 U24319 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(DATAI_15_), .A3(
        P3_EBX_REG_18__SCAN_IN), .A4(P2_DATAO_REG_14__SCAN_IN), .ZN(n21393) );
  NAND4_X1 U24320 ( .A1(P2_EBX_REG_5__SCAN_IN), .A2(P1_UWORD_REG_8__SCAN_IN), 
        .A3(n10798), .A4(n21464), .ZN(n21390) );
  NOR2_X1 U24321 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n21390), .ZN(
        n21391) );
  NAND4_X1 U24322 ( .A1(n21391), .A2(P1_ADDRESS_REG_2__SCAN_IN), .A3(
        P1_ADDRESS_REG_0__SCAN_IN), .A4(n21496), .ZN(n21392) );
  NOR3_X1 U24323 ( .A1(n21394), .A2(n21393), .A3(n21392), .ZN(n21543) );
  NAND4_X1 U24324 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P2_DATAO_REG_8__SCAN_IN), 
        .A3(n21428), .A4(n21429), .ZN(n21399) );
  NAND2_X1 U24325 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21509), .ZN(
        n21395) );
  NOR2_X1 U24326 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n21395), .ZN(n21397) );
  INV_X1 U24327 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n21414) );
  AND2_X1 U24328 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21396) );
  NAND4_X1 U24329 ( .A1(n21397), .A2(n13557), .A3(n21414), .A4(n21396), .ZN(
        n21398) );
  NOR3_X1 U24330 ( .A1(n21399), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A3(
        n21398), .ZN(n21400) );
  NAND4_X1 U24331 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21401), .A3(
        n21400), .A4(n13258), .ZN(n21412) );
  INV_X1 U24332 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21450) );
  NAND4_X1 U24333 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(
        P2_DATAO_REG_16__SCAN_IN), .A3(n11619), .A4(n21450), .ZN(n21411) );
  NOR4_X1 U24334 ( .A1(P1_EAX_REG_2__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .A3(n21438), .A4(n21435), .ZN(n21404) );
  NOR3_X1 U24335 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(
        BUF2_REG_2__SCAN_IN), .A3(P3_LWORD_REG_1__SCAN_IN), .ZN(n21403) );
  INV_X1 U24336 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n21458) );
  NOR4_X1 U24337 ( .A1(P1_EAX_REG_17__SCAN_IN), .A2(P3_MORE_REG_SCAN_IN), .A3(
        P1_UWORD_REG_13__SCAN_IN), .A4(n21458), .ZN(n21402) );
  NAND4_X1 U24338 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n21404), .A3(n21403), 
        .A4(n21402), .ZN(n21410) );
  NOR4_X1 U24339 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A4(n21475), .ZN(n21408) );
  NOR4_X1 U24340 ( .A1(P1_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(n21521), .A4(n21522), .ZN(n21407) );
  NOR4_X1 U24341 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_DATAO_REG_23__SCAN_IN), .A3(P2_DATAWIDTH_REG_31__SCAN_IN), .A4(
        n21507), .ZN(n21406) );
  NOR4_X1 U24342 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(
        P1_EAX_REG_6__SCAN_IN), .A3(P3_EAX_REG_0__SCAN_IN), .A4(
        P2_LWORD_REG_11__SCAN_IN), .ZN(n21405) );
  NAND4_X1 U24343 ( .A1(n21408), .A2(n21407), .A3(n21406), .A4(n21405), .ZN(
        n21409) );
  NOR4_X1 U24344 ( .A1(n21412), .A2(n21411), .A3(n21410), .A4(n21409), .ZN(
        n21542) );
  AOI22_X1 U24345 ( .A1(n21415), .A2(keyinput29), .B1(n21414), .B2(keyinput57), 
        .ZN(n21413) );
  OAI221_X1 U24346 ( .B1(n21415), .B2(keyinput29), .C1(n21414), .C2(keyinput57), .A(n21413), .ZN(n21426) );
  INV_X1 U24347 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n21417) );
  AOI22_X1 U24348 ( .A1(n21417), .A2(keyinput9), .B1(n13258), .B2(keyinput27), 
        .ZN(n21416) );
  OAI221_X1 U24349 ( .B1(n21417), .B2(keyinput9), .C1(n13258), .C2(keyinput27), 
        .A(n21416), .ZN(n21425) );
  INV_X1 U24350 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n21419) );
  AOI22_X1 U24351 ( .A1(n21420), .A2(keyinput5), .B1(n21419), .B2(keyinput60), 
        .ZN(n21418) );
  OAI221_X1 U24352 ( .B1(n21420), .B2(keyinput5), .C1(n21419), .C2(keyinput60), 
        .A(n21418), .ZN(n21424) );
  XOR2_X1 U24353 ( .A(n13557), .B(keyinput11), .Z(n21422) );
  XNOR2_X1 U24354 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B(keyinput0), .ZN(
        n21421) );
  NAND2_X1 U24355 ( .A1(n21422), .A2(n21421), .ZN(n21423) );
  NOR4_X1 U24356 ( .A1(n21426), .A2(n21425), .A3(n21424), .A4(n21423), .ZN(
        n21473) );
  AOI22_X1 U24357 ( .A1(n21429), .A2(keyinput36), .B1(n21428), .B2(keyinput53), 
        .ZN(n21427) );
  OAI221_X1 U24358 ( .B1(n21429), .B2(keyinput36), .C1(n21428), .C2(keyinput53), .A(n21427), .ZN(n21442) );
  AOI22_X1 U24359 ( .A1(n21432), .A2(keyinput10), .B1(keyinput63), .B2(n21431), 
        .ZN(n21430) );
  OAI221_X1 U24360 ( .B1(n21432), .B2(keyinput10), .C1(n21431), .C2(keyinput63), .A(n21430), .ZN(n21441) );
  AOI22_X1 U24361 ( .A1(n21435), .A2(keyinput30), .B1(n21434), .B2(keyinput62), 
        .ZN(n21433) );
  OAI221_X1 U24362 ( .B1(n21435), .B2(keyinput30), .C1(n21434), .C2(keyinput62), .A(n21433), .ZN(n21440) );
  AOI22_X1 U24363 ( .A1(n21438), .A2(keyinput19), .B1(n21437), .B2(keyinput31), 
        .ZN(n21436) );
  OAI221_X1 U24364 ( .B1(n21438), .B2(keyinput19), .C1(n21437), .C2(keyinput31), .A(n21436), .ZN(n21439) );
  NOR4_X1 U24365 ( .A1(n21442), .A2(n21441), .A3(n21440), .A4(n21439), .ZN(
        n21472) );
  INV_X1 U24366 ( .A(P3_LWORD_REG_1__SCAN_IN), .ZN(n21445) );
  AOI22_X1 U24367 ( .A1(n21445), .A2(keyinput12), .B1(n21444), .B2(keyinput40), 
        .ZN(n21443) );
  OAI221_X1 U24368 ( .B1(n21445), .B2(keyinput12), .C1(n21444), .C2(keyinput40), .A(n21443), .ZN(n21456) );
  INV_X1 U24369 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n21448) );
  INV_X1 U24370 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n21447) );
  AOI22_X1 U24371 ( .A1(n21448), .A2(keyinput7), .B1(keyinput15), .B2(n21447), 
        .ZN(n21446) );
  OAI221_X1 U24372 ( .B1(n21448), .B2(keyinput7), .C1(n21447), .C2(keyinput15), 
        .A(n21446), .ZN(n21455) );
  AOI22_X1 U24373 ( .A1(n21450), .A2(keyinput20), .B1(n10742), .B2(keyinput24), 
        .ZN(n21449) );
  OAI221_X1 U24374 ( .B1(n21450), .B2(keyinput20), .C1(n10742), .C2(keyinput24), .A(n21449), .ZN(n21454) );
  AOI22_X1 U24375 ( .A1(n11619), .A2(keyinput55), .B1(keyinput16), .B2(n21452), 
        .ZN(n21451) );
  OAI221_X1 U24376 ( .B1(n11619), .B2(keyinput55), .C1(n21452), .C2(keyinput16), .A(n21451), .ZN(n21453) );
  NOR4_X1 U24377 ( .A1(n21456), .A2(n21455), .A3(n21454), .A4(n21453), .ZN(
        n21471) );
  AOI22_X1 U24378 ( .A1(n15126), .A2(keyinput17), .B1(keyinput50), .B2(n21458), 
        .ZN(n21457) );
  OAI221_X1 U24379 ( .B1(n15126), .B2(keyinput17), .C1(n21458), .C2(keyinput50), .A(n21457), .ZN(n21469) );
  INV_X1 U24380 ( .A(P1_UWORD_REG_13__SCAN_IN), .ZN(n21461) );
  AOI22_X1 U24381 ( .A1(n21461), .A2(keyinput43), .B1(n21460), .B2(keyinput61), 
        .ZN(n21459) );
  OAI221_X1 U24382 ( .B1(n21461), .B2(keyinput43), .C1(n21460), .C2(keyinput61), .A(n21459), .ZN(n21468) );
  INV_X1 U24383 ( .A(P1_UWORD_REG_8__SCAN_IN), .ZN(n21463) );
  AOI22_X1 U24384 ( .A1(n21464), .A2(keyinput44), .B1(keyinput59), .B2(n21463), 
        .ZN(n21462) );
  OAI221_X1 U24385 ( .B1(n21464), .B2(keyinput44), .C1(n21463), .C2(keyinput59), .A(n21462), .ZN(n21467) );
  AOI22_X1 U24386 ( .A1(n11071), .A2(keyinput4), .B1(n10798), .B2(keyinput37), 
        .ZN(n21465) );
  OAI221_X1 U24387 ( .B1(n11071), .B2(keyinput4), .C1(n10798), .C2(keyinput37), 
        .A(n21465), .ZN(n21466) );
  NOR4_X1 U24388 ( .A1(n21469), .A2(n21468), .A3(n21467), .A4(n21466), .ZN(
        n21470) );
  NAND4_X1 U24389 ( .A1(n21473), .A2(n21472), .A3(n21471), .A4(n21470), .ZN(
        n21541) );
  AOI22_X1 U24390 ( .A1(n21476), .A2(keyinput6), .B1(n21475), .B2(keyinput49), 
        .ZN(n21474) );
  OAI221_X1 U24391 ( .B1(n21476), .B2(keyinput6), .C1(n21475), .C2(keyinput49), 
        .A(n21474), .ZN(n21489) );
  AOI22_X1 U24392 ( .A1(n21479), .A2(keyinput13), .B1(n21478), .B2(keyinput33), 
        .ZN(n21477) );
  OAI221_X1 U24393 ( .B1(n21479), .B2(keyinput13), .C1(n21478), .C2(keyinput33), .A(n21477), .ZN(n21488) );
  AOI22_X1 U24394 ( .A1(n21482), .A2(keyinput28), .B1(n21481), .B2(keyinput26), 
        .ZN(n21480) );
  OAI221_X1 U24395 ( .B1(n21482), .B2(keyinput28), .C1(n21481), .C2(keyinput26), .A(n21480), .ZN(n21487) );
  XOR2_X1 U24396 ( .A(n21483), .B(keyinput41), .Z(n21485) );
  XNOR2_X1 U24397 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B(keyinput58), .ZN(
        n21484) );
  NAND2_X1 U24398 ( .A1(n21485), .A2(n21484), .ZN(n21486) );
  NOR4_X1 U24399 ( .A1(n21489), .A2(n21488), .A3(n21487), .A4(n21486), .ZN(
        n21539) );
  AOI22_X1 U24400 ( .A1(n12981), .A2(keyinput1), .B1(keyinput51), .B2(n21491), 
        .ZN(n21490) );
  OAI221_X1 U24401 ( .B1(n12981), .B2(keyinput1), .C1(n21491), .C2(keyinput51), 
        .A(n21490), .ZN(n21504) );
  INV_X1 U24402 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n21494) );
  AOI22_X1 U24403 ( .A1(n21494), .A2(keyinput46), .B1(keyinput2), .B2(n21493), 
        .ZN(n21492) );
  OAI221_X1 U24404 ( .B1(n21494), .B2(keyinput46), .C1(n21493), .C2(keyinput2), 
        .A(n21492), .ZN(n21503) );
  AOI22_X1 U24405 ( .A1(n21497), .A2(keyinput38), .B1(n21496), .B2(keyinput54), 
        .ZN(n21495) );
  OAI221_X1 U24406 ( .B1(n21497), .B2(keyinput38), .C1(n21496), .C2(keyinput54), .A(n21495), .ZN(n21502) );
  XOR2_X1 U24407 ( .A(n21498), .B(keyinput39), .Z(n21500) );
  XNOR2_X1 U24408 ( .A(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B(keyinput14), .ZN(
        n21499) );
  NAND2_X1 U24409 ( .A1(n21500), .A2(n21499), .ZN(n21501) );
  NOR4_X1 U24410 ( .A1(n21504), .A2(n21503), .A3(n21502), .A4(n21501), .ZN(
        n21538) );
  AOI22_X1 U24411 ( .A1(n21507), .A2(keyinput34), .B1(keyinput3), .B2(n21506), 
        .ZN(n21505) );
  OAI221_X1 U24412 ( .B1(n21507), .B2(keyinput34), .C1(n21506), .C2(keyinput3), 
        .A(n21505), .ZN(n21519) );
  AOI22_X1 U24413 ( .A1(n21510), .A2(keyinput56), .B1(n21509), .B2(keyinput35), 
        .ZN(n21508) );
  OAI221_X1 U24414 ( .B1(n21510), .B2(keyinput56), .C1(n21509), .C2(keyinput35), .A(n21508), .ZN(n21518) );
  AOI22_X1 U24415 ( .A1(n21512), .A2(keyinput48), .B1(n11568), .B2(keyinput42), 
        .ZN(n21511) );
  OAI221_X1 U24416 ( .B1(n21512), .B2(keyinput48), .C1(n11568), .C2(keyinput42), .A(n21511), .ZN(n21517) );
  INV_X1 U24417 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n21515) );
  AOI22_X1 U24418 ( .A1(n21515), .A2(keyinput45), .B1(n21514), .B2(keyinput18), 
        .ZN(n21513) );
  OAI221_X1 U24419 ( .B1(n21515), .B2(keyinput45), .C1(n21514), .C2(keyinput18), .A(n21513), .ZN(n21516) );
  NOR4_X1 U24420 ( .A1(n21519), .A2(n21518), .A3(n21517), .A4(n21516), .ZN(
        n21537) );
  AOI22_X1 U24421 ( .A1(n21522), .A2(keyinput52), .B1(keyinput23), .B2(n21521), 
        .ZN(n21520) );
  OAI221_X1 U24422 ( .B1(n21522), .B2(keyinput52), .C1(n21521), .C2(keyinput23), .A(n21520), .ZN(n21535) );
  AOI22_X1 U24423 ( .A1(n21525), .A2(keyinput22), .B1(keyinput21), .B2(n21524), 
        .ZN(n21523) );
  OAI221_X1 U24424 ( .B1(n21525), .B2(keyinput22), .C1(n21524), .C2(keyinput21), .A(n21523), .ZN(n21534) );
  INV_X1 U24425 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n21528) );
  AOI22_X1 U24426 ( .A1(n21528), .A2(keyinput47), .B1(keyinput25), .B2(n21527), 
        .ZN(n21526) );
  OAI221_X1 U24427 ( .B1(n21528), .B2(keyinput47), .C1(n21527), .C2(keyinput25), .A(n21526), .ZN(n21533) );
  AOI22_X1 U24428 ( .A1(n21531), .A2(keyinput32), .B1(keyinput8), .B2(n21530), 
        .ZN(n21529) );
  OAI221_X1 U24429 ( .B1(n21531), .B2(keyinput32), .C1(n21530), .C2(keyinput8), 
        .A(n21529), .ZN(n21532) );
  NOR4_X1 U24430 ( .A1(n21535), .A2(n21534), .A3(n21533), .A4(n21532), .ZN(
        n21536) );
  NAND4_X1 U24431 ( .A1(n21539), .A2(n21538), .A3(n21537), .A4(n21536), .ZN(
        n21540) );
  AOI211_X1 U24432 ( .C1(n21543), .C2(n21542), .A(n21541), .B(n21540), .ZN(
        n21557) );
  AOI22_X1 U24433 ( .A1(n21547), .A2(n21546), .B1(n21545), .B2(n21544), .ZN(
        n21548) );
  INV_X1 U24434 ( .A(n21548), .ZN(n21554) );
  OAI22_X1 U24435 ( .A1(n21552), .A2(n21551), .B1(n21550), .B2(n21549), .ZN(
        n21553) );
  AOI211_X1 U24436 ( .C1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .C2(n21555), .A(
        n21554), .B(n21553), .ZN(n21556) );
  XNOR2_X1 U24437 ( .A(n21557), .B(n21556), .ZN(P3_U2915) );
  AND2_X1 U13216 ( .A1(n10186), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10691) );
  INV_X1 U11031 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20304) );
  BUF_X1 U11160 ( .A(n14474), .Z(n9590) );
  CLKBUF_X3 U11021 ( .A(n12477), .Z(n9594) );
  NAND2_X1 U11147 ( .A1(n12012), .A2(n11995), .ZN(n13240) );
  AND2_X2 U11114 ( .A1(n14625), .A2(n10551), .ZN(n14473) );
  AND4_X1 U11020 ( .A1(n10581), .A2(n10589), .A3(n12512), .A4(n10585), .ZN(
        n10582) );
  CLKBUF_X1 U11026 ( .A(n14481), .Z(n9584) );
  CLKBUF_X1 U11053 ( .A(n10594), .Z(n11022) );
  CLKBUF_X1 U11064 ( .A(n14474), .Z(n9589) );
  CLKBUF_X1 U11069 ( .A(n11068), .Z(n11144) );
  CLKBUF_X1 U11149 ( .A(n17497), .Z(n17509) );
  AND4_X1 U11350 ( .A1(n10787), .A2(n10792), .A3(n9674), .A4(n10009), .ZN(
        n21558) );
  INV_X1 U12583 ( .A(n11995), .ZN(n12782) );
endmodule

