

module b21_C_AntiSAT_k_256_2 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, 
        keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, 
        keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, 
        keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, 
        keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, 
        keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, 
        keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, 
        keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, 
        keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, 
        keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, 
        keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, 
        keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, 
        keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, 
        keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, 
        keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, 
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, 
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, 
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, 
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, 
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, 
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, 
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, 
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, 
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, 
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249, 
        keyinput250, keyinput251, keyinput252, keyinput253, keyinput254, 
        keyinput255, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, 
        ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, 
        ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, 
        ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, 
        ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, 
        P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, 
        P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, 
        P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, 
        P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, 
        P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, 
        P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, 
        P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, 
        P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, 
        P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, 
        P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, 
        P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, 
        P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, 
        P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, 
        P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, 
        P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, 
        P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, 
        P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, 
        P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, 
        P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, 
        P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430;

  OAI211_X1 U4984 ( .C1(n5015), .C2(n4896), .A(n5012), .B(n5009), .ZN(n9753)
         );
  AND2_X1 U4985 ( .A1(n9309), .A2(n9308), .ZN(n9319) );
  AND4_X1 U4986 ( .A1(n6234), .A2(n6233), .A3(n6232), .A4(n6231), .ZN(n9618)
         );
  BUF_X2 U4987 ( .A(n6255), .Z(n4490) );
  INV_X1 U4988 ( .A(n4486), .ZN(n6216) );
  INV_X1 U4989 ( .A(n8559), .ZN(n6245) );
  CLKBUF_X2 U4990 ( .A(n6301), .Z(n6527) );
  BUF_X2 U4991 ( .A(n6294), .Z(n4481) );
  INV_X2 U4992 ( .A(n10296), .ZN(n10272) );
  INV_X1 U4993 ( .A(n8465), .ZN(n8478) );
  INV_X4 U4994 ( .A(n6329), .ZN(n6422) );
  NAND2_X1 U4995 ( .A1(n5357), .A2(n7493), .ZN(n8360) );
  NAND2_X1 U4996 ( .A1(n7497), .A2(n6368), .ZN(n7646) );
  NAND2_X1 U4997 ( .A1(n5644), .A2(n8349), .ZN(n8488) );
  AND2_X1 U4998 ( .A1(n4489), .A2(n4483), .ZN(n9214) );
  INV_X1 U4999 ( .A(n5764), .ZN(n5765) );
  INV_X1 U5000 ( .A(n6252), .ZN(n7574) );
  NAND2_X1 U5001 ( .A1(n4481), .A2(n9987), .ZN(n6545) );
  INV_X1 U5002 ( .A(n5326), .ZN(n8318) );
  NAND2_X1 U5003 ( .A1(n5413), .A2(n5412), .ZN(n10321) );
  NAND2_X1 U5004 ( .A1(n5090), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5092) );
  NAND2_X1 U5005 ( .A1(n4481), .A2(n9987), .ZN(n4489) );
  XNOR2_X1 U5006 ( .A(n5018), .B(P1_IR_REG_28__SCAN_IN), .ZN(n6294) );
  INV_X1 U5007 ( .A(n8271), .ZN(n10315) );
  INV_X2 U5008 ( .A(n9728), .ZN(n9703) );
  XNOR2_X1 U5009 ( .A(n5734), .B(n5733), .ZN(n9987) );
  NOR2_X4 U5010 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5824) );
  MUX2_X2 U5011 ( .A(n8788), .B(n8787), .S(n8856), .Z(n8790) );
  AND4_X2 U5012 ( .A1(n5079), .A2(n5259), .A3(n5471), .A4(n5398), .ZN(n5080)
         );
  AND4_X2 U5013 ( .A1(n5243), .A2(n5078), .A3(n5077), .A4(n5076), .ZN(n5081)
         );
  OAI21_X2 U5014 ( .B1(n7646), .B2(n4602), .A(n4603), .ZN(n6376) );
  AOI21_X2 U5015 ( .B1(n4926), .B2(n4605), .A(n4604), .ZN(n4603) );
  AND2_X2 U5016 ( .A1(n10248), .A2(n10261), .ZN(n10250) );
  INV_X1 U5017 ( .A(n7240), .ZN(n6328) );
  OAI21_X2 U5018 ( .B1(n7126), .B2(n4579), .A(n4570), .ZN(n7240) );
  OAI21_X2 U5020 ( .B1(n7612), .B2(n4973), .A(n4972), .ZN(n4975) );
  OR2_X2 U5021 ( .A1(n7999), .A2(n9972), .ZN(n8167) );
  NAND2_X2 U5022 ( .A1(n6027), .A2(n6026), .ZN(n9972) );
  OAI21_X2 U5023 ( .B1(n5484), .B2(n5167), .A(n5172), .ZN(n5219) );
  CLKBUF_X1 U5024 ( .A(n6338), .Z(n4479) );
  CLKBUF_X1 U5025 ( .A(n6338), .Z(n4480) );
  AOI21_X2 U5026 ( .B1(n7136), .B2(P2_REG2_REG_4__SCAN_IN), .A(n7135), .ZN(
        n7157) );
  AND2_X2 U5027 ( .A1(n5770), .A2(n6543), .ZN(n4486) );
  AND2_X2 U5028 ( .A1(n5770), .A2(n6543), .ZN(n4487) );
  OAI21_X2 U5029 ( .B1(n9177), .B2(n9179), .A(n9178), .ZN(n9084) );
  NAND2_X2 U5030 ( .A1(n6136), .A2(n6135), .ZN(n9178) );
  OAI22_X2 U5031 ( .A1(n9724), .A2(n8534), .B1(n9182), .B2(n9730), .ZN(n9707)
         );
  NOR2_X2 U5032 ( .A1(n8533), .A2(n8532), .ZN(n9724) );
  AOI211_X2 U5033 ( .C1(n9733), .C2(n9592), .A(n9562), .B(n9561), .ZN(n9757)
         );
  AOI21_X2 U5034 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n8767), .A(n8766), .ZN(
        n8775) );
  OAI21_X1 U5035 ( .B1(n8880), .B2(n4988), .A(n4985), .ZN(n8858) );
  NAND2_X1 U5036 ( .A1(n8902), .A2(n8901), .ZN(n8989) );
  NAND2_X1 U5037 ( .A1(n7978), .A2(n8482), .ZN(n8068) );
  INV_X1 U5038 ( .A(n9607), .ZN(n9102) );
  NAND2_X1 U5039 ( .A1(n7211), .A2(n8487), .ZN(n7210) );
  NAND2_X1 U5041 ( .A1(n10315), .A2(n8679), .ZN(n5644) );
  INV_X1 U5042 ( .A(n6236), .ZN(n6255) );
  NAND2_X2 U5043 ( .A1(n8348), .A2(n8372), .ZN(n8487) );
  NAND2_X2 U5044 ( .A1(n8360), .A2(n8363), .ZN(n8484) );
  NAND3_X1 U5045 ( .A1(n4659), .A2(n4660), .A3(n5795), .ZN(n9492) );
  INV_X1 U5046 ( .A(n4479), .ZN(n6638) );
  NAND2_X1 U5047 ( .A1(n7279), .A2(n8681), .ZN(n8363) );
  BUF_X1 U5049 ( .A(n6360), .Z(n6398) );
  INV_X1 U5051 ( .A(n7493), .ZN(n7279) );
  INV_X2 U5053 ( .A(n6642), .ZN(n6672) );
  NAND2_X2 U5054 ( .A1(n6283), .A2(n5775), .ZN(n5770) );
  BUF_X2 U5055 ( .A(n5334), .Z(n5377) );
  NOR2_X1 U5056 ( .A1(n5018), .A2(n5756), .ZN(n5758) );
  NOR2_X1 U5057 ( .A1(n8963), .A2(n4909), .ZN(n8966) );
  OR2_X1 U5058 ( .A1(n9074), .A2(n4834), .ZN(n4833) );
  AND2_X1 U5059 ( .A1(n4991), .A2(n4990), .ZN(n8864) );
  AND2_X1 U5060 ( .A1(n4991), .A2(n4576), .ZN(n8983) );
  OR2_X1 U5061 ( .A1(n5014), .A2(n10233), .ZN(n5007) );
  AOI21_X1 U5062 ( .B1(n4895), .B2(n9738), .A(n4892), .ZN(n9752) );
  XNOR2_X1 U5063 ( .A(n4897), .B(n4896), .ZN(n4895) );
  NOR2_X1 U5064 ( .A1(n9558), .A2(n8554), .ZN(n4897) );
  OR2_X1 U5065 ( .A1(n8776), .A2(n8777), .ZN(n4692) );
  NOR2_X1 U5066 ( .A1(n8770), .A2(n5496), .ZN(n8776) );
  AND2_X1 U5067 ( .A1(n9197), .A2(n9196), .ZN(n9201) );
  NAND2_X1 U5068 ( .A1(n5016), .A2(n4555), .ZN(n9659) );
  AOI21_X1 U5069 ( .B1(n4985), .B2(n4988), .A(n4984), .ZN(n4983) );
  NAND2_X1 U5070 ( .A1(n9416), .A2(n9411), .ZN(n9575) );
  NAND2_X1 U5071 ( .A1(n6513), .A2(n6512), .ZN(n9755) );
  NAND2_X1 U5072 ( .A1(n4937), .A2(n4934), .ZN(n8594) );
  OR2_X1 U5073 ( .A1(n9769), .A2(n9618), .ZN(n9293) );
  NAND2_X1 U5074 ( .A1(n7555), .A2(n5959), .ZN(n5963) );
  NAND2_X1 U5075 ( .A1(n8176), .A2(n4696), .ZN(n8734) );
  NAND2_X1 U5076 ( .A1(n5020), .A2(n5019), .ZN(n8206) );
  AND2_X1 U5077 ( .A1(n8012), .A2(n9333), .ZN(n8216) );
  AND4_X1 U5078 ( .A1(n6306), .A2(n6305), .A3(n6304), .A4(n6303), .ZN(n8541)
         );
  AOI21_X1 U5079 ( .B1(n4852), .B2(n4854), .A(n4538), .ZN(n4851) );
  OAI21_X1 U5080 ( .B1(n4878), .B2(n7910), .A(n4877), .ZN(n8162) );
  NAND2_X1 U5081 ( .A1(n7376), .A2(n4965), .ZN(n7413) );
  NAND4_X1 U5082 ( .A1(n6249), .A2(n6248), .A3(n6247), .A4(n6246), .ZN(n9607)
         );
  NAND2_X1 U5083 ( .A1(n7716), .A2(n7715), .ZN(n7877) );
  AND2_X1 U5084 ( .A1(n7660), .A2(n9443), .ZN(n7718) );
  OR2_X1 U5085 ( .A1(n7845), .A2(n7655), .ZN(n7660) );
  AND2_X2 U5086 ( .A1(n7455), .A2(n8903), .ZN(n10296) );
  AND2_X1 U5087 ( .A1(n6009), .A2(n6008), .ZN(n9952) );
  NAND2_X1 U5088 ( .A1(n6044), .A2(n6043), .ZN(n9825) );
  OAI21_X1 U5089 ( .B1(n5257), .B2(n5154), .A(n5153), .ZN(n5470) );
  NAND2_X1 U5090 ( .A1(n5266), .A2(n5265), .ZN(n5468) );
  NAND2_X2 U5091 ( .A1(n7569), .A2(n9669), .ZN(n9728) );
  NAND2_X1 U5092 ( .A1(n5311), .A2(n5310), .ZN(n7389) );
  OAI211_X1 U5093 ( .C1(n6545), .C2(n6613), .A(n5970), .B(n5969), .ZN(n7881)
         );
  XNOR2_X1 U5094 ( .A(n5263), .B(n5053), .ZN(n6661) );
  AND3_X1 U5095 ( .A1(n5879), .A2(n5878), .A3(n5877), .ZN(n7602) );
  AND2_X2 U5096 ( .A1(n4486), .A2(n7627), .ZN(n5923) );
  AND3_X1 U5097 ( .A1(n5861), .A2(n5860), .A3(n5859), .ZN(n10172) );
  AND2_X2 U5098 ( .A1(n6580), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  INV_X1 U5099 ( .A(n9209), .ZN(n6282) );
  NAND2_X1 U5100 ( .A1(n5389), .A2(n4508), .ZN(n8679) );
  AND3_X1 U5101 ( .A1(n5843), .A2(n5842), .A3(n5841), .ZN(n10167) );
  CLKBUF_X1 U5102 ( .A(n5917), .Z(n6627) );
  NAND3_X4 U5103 ( .A1(n6271), .A2(n6266), .A3(n6275), .ZN(n6543) );
  NAND2_X1 U5104 ( .A1(n5773), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5774) );
  INV_X2 U5105 ( .A(n5917), .ZN(n8555) );
  AND2_X1 U5106 ( .A1(n5755), .A2(n4506), .ZN(n6271) );
  AND2_X1 U5107 ( .A1(n5749), .A2(n5748), .ZN(n6266) );
  XNOR2_X1 U5108 ( .A(n5772), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6283) );
  INV_X1 U5109 ( .A(n9855), .ZN(n5763) );
  NAND2_X1 U5110 ( .A1(n5741), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5772) );
  XNOR2_X1 U5111 ( .A(n5758), .B(n5757), .ZN(n5764) );
  BUF_X2 U5112 ( .A(n5328), .Z(n4485) );
  OR2_X1 U5113 ( .A1(n6278), .A2(n5750), .ZN(n5753) );
  XNOR2_X1 U5114 ( .A(n5636), .B(n5635), .ZN(n8330) );
  AND2_X1 U5115 ( .A1(n4675), .A2(n4674), .ZN(n5018) );
  NAND2_X1 U5116 ( .A1(n4679), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5734) );
  XNOR2_X1 U5117 ( .A(n4869), .B(SI_3_), .ZN(n5369) );
  XNOR2_X1 U5118 ( .A(n5120), .B(SI_6_), .ZN(n5408) );
  INV_X2 U5119 ( .A(n4568), .ZN(n8311) );
  AND2_X1 U5120 ( .A1(n5992), .A2(n4866), .ZN(n5776) );
  INV_X2 U5121 ( .A(n4567), .ZN(n9857) );
  NAND2_X1 U5122 ( .A1(n5201), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5205) );
  CLKBUF_X1 U5123 ( .A(n5991), .Z(n5992) );
  NOR2_X1 U5124 ( .A1(n5730), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n5038) );
  NOR2_X2 U5125 ( .A1(n5875), .A2(n5721), .ZN(n5967) );
  BUF_X8 U5126 ( .A(n5112), .Z(n4483) );
  AND3_X1 U5127 ( .A1(n5040), .A2(n5050), .A3(n4544), .ZN(n4866) );
  AND4_X1 U5128 ( .A1(n5742), .A2(n5739), .A3(n5738), .A4(n5740), .ZN(n5726)
         );
  NAND3_X1 U5129 ( .A1(n5101), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4819) );
  AND2_X1 U5130 ( .A1(n4769), .A2(n4768), .ZN(n5083) );
  AND2_X1 U5131 ( .A1(n5351), .A2(n5075), .ZN(n5378) );
  AND2_X1 U5132 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4579), .ZN(n4535) );
  INV_X1 U5133 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5740) );
  NOR2_X1 U5134 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5720) );
  INV_X1 U5135 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5742) );
  INV_X1 U5136 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5757) );
  AND2_X1 U5137 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n5756) );
  INV_X1 U5138 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5950) );
  INV_X1 U5139 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5718) );
  INV_X1 U5140 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5738) );
  INV_X1 U5141 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5398) );
  NOR2_X1 U5142 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n4768) );
  NOR2_X1 U5143 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4769) );
  INV_X1 U5144 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9537) );
  NOR2_X1 U5145 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5040) );
  INV_X4 U5146 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  BUF_X4 U5147 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n4579) );
  INV_X4 U5148 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U5149 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5078) );
  NOR2_X1 U5150 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5077) );
  NOR2_X1 U5151 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5076) );
  NOR2_X1 U5152 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5079) );
  INV_X2 U5153 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5101) );
  INV_X1 U5154 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5471) );
  INV_X1 U5155 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5259) );
  XNOR2_X2 U5156 ( .A(n5564), .B(n5559), .ZN(n7824) );
  AOI21_X1 U5157 ( .B1(n4929), .B2(n4931), .A(n4539), .ZN(n4928) );
  AOI21_X2 U5158 ( .B1(n7834), .B2(n7830), .A(n7831), .ZN(n7924) );
  INV_X4 U5159 ( .A(n4485), .ZN(n5663) );
  OAI22_X2 U5160 ( .A1(n7934), .A2(n8414), .B1(n8060), .B2(n8670), .ZN(n7981)
         );
  NAND3_X2 U5161 ( .A1(n5824), .A2(n5042), .A3(n5718), .ZN(n5875) );
  NAND2_X1 U5162 ( .A1(n9166), .A2(n5839), .ZN(n7296) );
  AND2_X1 U5163 ( .A1(n4486), .A2(n7627), .ZN(n4484) );
  NOR2_X2 U5164 ( .A1(n6069), .A2(n6068), .ZN(n6083) );
  OR2_X2 U5165 ( .A1(n6046), .A2(n6045), .ZN(n6069) );
  NOR2_X2 U5166 ( .A1(n9560), .A2(n9559), .ZN(n9558) );
  OAI21_X2 U5167 ( .B1(n9110), .B2(n4863), .A(n4861), .ZN(n4864) );
  XNOR2_X1 U5168 ( .A(n10167), .B(n7846), .ZN(n7803) );
  NAND4_X2 U5169 ( .A1(n5847), .A2(n5846), .A3(n5845), .A4(n5844), .ZN(n7846)
         );
  OR2_X1 U5170 ( .A1(n4839), .A2(n9075), .ZN(n9127) );
  NAND2_X1 U5171 ( .A1(n4481), .A2(n9987), .ZN(n4488) );
  OAI222_X1 U5172 ( .A1(n9857), .A2(n8232), .B1(P1_U3084), .B2(n5764), .C1(
        n8543), .C2(n8257), .ZN(P1_U3324) );
  AND2_X1 U5173 ( .A1(n5763), .A2(n5764), .ZN(n5880) );
  NOR2_X2 U5174 ( .A1(n6104), .A2(n6877), .ZN(n6127) );
  OR2_X2 U5175 ( .A1(n6102), .A2(n9111), .ZN(n6104) );
  NOR3_X2 U5176 ( .A1(n9619), .A2(n9755), .A3(n4765), .ZN(n4763) );
  OR2_X2 U5177 ( .A1(n9627), .A2(n9776), .ZN(n9619) );
  CLKBUF_X1 U5178 ( .A(n9987), .Z(n4491) );
  NOR2_X2 U5179 ( .A1(n9084), .A2(n9085), .ZN(n9149) );
  NOR2_X2 U5180 ( .A1(n5972), .A2(n5971), .ZN(n5996) );
  OR2_X2 U5181 ( .A1(n5943), .A2(n7004), .ZN(n5972) );
  NOR2_X1 U5182 ( .A1(n8007), .A2(n5026), .ZN(n5025) );
  INV_X1 U5183 ( .A(n5028), .ZN(n5026) );
  OR2_X1 U5184 ( .A1(n9348), .A2(n5056), .ZN(n8007) );
  NAND2_X1 U5185 ( .A1(n8194), .A2(n8193), .ZN(n8281) );
  NAND2_X1 U5186 ( .A1(n8189), .A2(n8188), .ZN(n8194) );
  INV_X1 U5187 ( .A(n4789), .ZN(n4788) );
  OAI21_X1 U5188 ( .B1(n5655), .B2(n4502), .A(n8430), .ZN(n4789) );
  BUF_X1 U5189 ( .A(n5337), .Z(n5429) );
  NAND2_X1 U5190 ( .A1(n4540), .A2(n4631), .ZN(n4630) );
  NAND2_X1 U5191 ( .A1(n4496), .A2(n4632), .ZN(n4631) );
  NAND2_X1 U5192 ( .A1(n5141), .A2(n5140), .ZN(n5144) );
  NOR2_X1 U5193 ( .A1(n7734), .A2(n4930), .ZN(n4929) );
  NOR2_X1 U5194 ( .A1(n4931), .A2(n7644), .ZN(n4930) );
  INV_X1 U5195 ( .A(n8231), .ZN(n5094) );
  INV_X1 U5196 ( .A(n5093), .ZN(n5095) );
  OR2_X1 U5197 ( .A1(n7458), .A2(n5445), .ZN(n8386) );
  AND2_X1 U5198 ( .A1(n9540), .A2(n9539), .ZN(n9422) );
  OAI21_X1 U5199 ( .B1(n9417), .B2(n4890), .A(n9413), .ZN(n4889) );
  OR2_X1 U5200 ( .A1(n9764), .A2(n9607), .ZN(n9325) );
  AND2_X1 U5201 ( .A1(n9764), .A2(n9607), .ZN(n9326) );
  NOR2_X1 U5202 ( .A1(n9779), .A2(n9477), .ZN(n8552) );
  OR2_X1 U5203 ( .A1(n9816), .A2(n9193), .ZN(n9388) );
  XNOR2_X1 U5204 ( .A(n8284), .B(n8282), .ZN(n8296) );
  OAI21_X1 U5205 ( .B1(n5581), .B2(n5580), .A(n5579), .ZN(n5601) );
  NAND2_X1 U5206 ( .A1(n5312), .A2(n5128), .ZN(n4624) );
  NOR2_X2 U5207 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5042) );
  NAND3_X1 U5208 ( .A1(n4958), .A2(n4957), .A3(n4956), .ZN(n6436) );
  INV_X1 U5209 ( .A(n6440), .ZN(n4956) );
  XNOR2_X1 U5210 ( .A(n6329), .B(n7511), .ZN(n6325) );
  INV_X1 U5211 ( .A(n6376), .ZN(n6379) );
  NOR2_X1 U5212 ( .A1(n9035), .A2(n8658), .ZN(n8474) );
  CLKBUF_X1 U5213 ( .A(n5553), .Z(n5578) );
  OR2_X1 U5214 ( .A1(n8177), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4696) );
  NAND2_X1 U5215 ( .A1(n8437), .A2(n4907), .ZN(n4905) );
  OAI21_X1 U5216 ( .B1(n8935), .B2(n4908), .A(n8437), .ZN(n4904) );
  INV_X1 U5217 ( .A(n8336), .ZN(n4790) );
  NAND2_X1 U5218 ( .A1(n8071), .A2(n4978), .ZN(n8119) );
  OR2_X1 U5219 ( .A1(n8203), .A2(n8668), .ZN(n4978) );
  NAND2_X1 U5220 ( .A1(n8291), .A2(n8290), .ZN(n8323) );
  NAND2_X1 U5221 ( .A1(n9853), .A2(n8297), .ZN(n8291) );
  XNOR2_X1 U5222 ( .A(n5631), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8327) );
  AND2_X1 U5223 ( .A1(n4846), .A2(n9092), .ZN(n4845) );
  OR2_X1 U5224 ( .A1(n4847), .A2(n9147), .ZN(n4846) );
  NAND2_X1 U5225 ( .A1(n9074), .A2(n9077), .ZN(n4840) );
  INV_X1 U5226 ( .A(n4482), .ZN(n6296) );
  XNOR2_X1 U5227 ( .A(n9510), .B(n9509), .ZN(n10077) );
  NAND2_X1 U5228 ( .A1(n9675), .A2(n5017), .ZN(n5016) );
  OR2_X1 U5229 ( .A1(n9796), .A2(n9701), .ZN(n5017) );
  AOI21_X1 U5230 ( .B1(n4494), .B2(n5024), .A(n4533), .ZN(n5019) );
  AND2_X1 U5231 ( .A1(n9220), .A2(n9228), .ZN(n9340) );
  NAND2_X1 U5232 ( .A1(n8545), .A2(n8544), .ZN(n9749) );
  NAND2_X1 U5233 ( .A1(n9755), .A2(n9476), .ZN(n5015) );
  AND2_X1 U5234 ( .A1(n7570), .A2(n6285), .ZN(n9964) );
  XNOR2_X1 U5235 ( .A(n5117), .B(SI_5_), .ZN(n5395) );
  NAND2_X1 U5236 ( .A1(n7365), .A2(n4925), .ZN(n4921) );
  NAND2_X1 U5237 ( .A1(n6646), .A2(n6645), .ZN(n4592) );
  NAND2_X1 U5238 ( .A1(n4894), .A2(n4893), .ZN(n4892) );
  NAND2_X1 U5239 ( .A1(n9538), .A2(n9474), .ZN(n4893) );
  NAND2_X1 U5240 ( .A1(n8340), .A2(n7500), .ZN(n4648) );
  NAND2_X1 U5241 ( .A1(n8406), .A2(n8478), .ZN(n4641) );
  AOI21_X1 U5242 ( .B1(n8407), .B2(n8465), .A(n8410), .ZN(n4642) );
  NAND2_X1 U5243 ( .A1(n9919), .A2(n8409), .ZN(n4640) );
  NOR2_X1 U5244 ( .A1(n4630), .A2(n4528), .ZN(n4629) );
  NAND2_X1 U5245 ( .A1(n8437), .A2(n8439), .ZN(n4633) );
  NAND2_X1 U5246 ( .A1(n4628), .A2(n8438), .ZN(n4627) );
  INV_X1 U5247 ( .A(n4630), .ZN(n4628) );
  AND2_X1 U5248 ( .A1(n4830), .A2(n4828), .ZN(n8434) );
  NOR2_X1 U5249 ( .A1(n8633), .A2(n4829), .ZN(n4828) );
  INV_X1 U5250 ( .A(n5515), .ZN(n4829) );
  NAND2_X1 U5251 ( .A1(n9277), .A2(n4689), .ZN(n4688) );
  NOR2_X1 U5252 ( .A1(n9328), .A2(n9318), .ZN(n4689) );
  NAND2_X1 U5253 ( .A1(n4671), .A2(n9279), .ZN(n9276) );
  NAND2_X1 U5254 ( .A1(n9283), .A2(n4521), .ZN(n4687) );
  AND2_X1 U5255 ( .A1(n4824), .A2(n4547), .ZN(n8448) );
  NAND2_X1 U5256 ( .A1(n4818), .A2(n8478), .ZN(n4817) );
  INV_X1 U5257 ( .A(n9317), .ZN(n4657) );
  INV_X1 U5258 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5722) );
  AOI22_X1 U5259 ( .A1(n8594), .A2(n8593), .B1(n6401), .B2(n6400), .ZN(n6404)
         );
  INV_X1 U5260 ( .A(n6375), .ZN(n4604) );
  OR2_X1 U5261 ( .A1(n8323), .A2(n8322), .ZN(n8477) );
  NAND2_X1 U5262 ( .A1(n8398), .A2(n4776), .ZN(n4775) );
  INV_X1 U5263 ( .A(n8341), .ZN(n4776) );
  OR2_X1 U5264 ( .A1(n5468), .A2(n7856), .ZN(n8408) );
  OR2_X1 U5265 ( .A1(n5461), .A2(n8712), .ZN(n5289) );
  NAND2_X1 U5266 ( .A1(n5064), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5460) );
  OR2_X1 U5267 ( .A1(n7389), .A2(n8583), .ZN(n8340) );
  OR2_X1 U5268 ( .A1(n8588), .A2(n7379), .ZN(n8390) );
  NAND2_X1 U5269 ( .A1(n9575), .A2(n4998), .ZN(n4997) );
  INV_X1 U5270 ( .A(n5002), .ZN(n4998) );
  NAND2_X1 U5271 ( .A1(n4999), .A2(n4995), .ZN(n4994) );
  INV_X1 U5272 ( .A(n5006), .ZN(n4995) );
  OR2_X1 U5273 ( .A1(n6527), .A2(n9553), .ZN(n6503) );
  INV_X1 U5274 ( .A(n9326), .ZN(n5005) );
  NAND2_X1 U5275 ( .A1(n8539), .A2(n9638), .ZN(n5006) );
  AOI21_X1 U5276 ( .B1(n9646), .B2(n9400), .A(n9328), .ZN(n9634) );
  OR2_X1 U5277 ( .A1(n9786), .A2(n9665), .ZN(n9400) );
  OR2_X1 U5278 ( .A1(n9791), .A2(n9682), .ZN(n9396) );
  NOR2_X1 U5279 ( .A1(n4758), .A2(n9809), .ZN(n4757) );
  INV_X1 U5280 ( .A(n4759), .ZN(n4758) );
  NOR2_X1 U5281 ( .A1(n9816), .A2(n9204), .ZN(n4759) );
  NAND2_X1 U5282 ( .A1(n10202), .A2(n9485), .ZN(n9233) );
  NAND2_X1 U5283 ( .A1(n5035), .A2(n7587), .ZN(n5034) );
  INV_X1 U5284 ( .A(n9340), .ZN(n5035) );
  OAI21_X1 U5285 ( .B1(n8281), .B2(n8280), .A(n8279), .ZN(n8284) );
  NAND2_X1 U5286 ( .A1(n5603), .A2(n5602), .ZN(n5617) );
  NAND2_X1 U5287 ( .A1(n5601), .A2(n5600), .ZN(n5603) );
  OAI21_X1 U5288 ( .B1(n5564), .B2(n5563), .A(n5562), .ZN(n5581) );
  OAI21_X1 U5289 ( .B1(n5219), .B2(n5218), .A(n5177), .ZN(n5502) );
  AND2_X1 U5290 ( .A1(n5181), .A2(n5180), .ZN(n5501) );
  AND2_X1 U5291 ( .A1(n5165), .A2(n5164), .ZN(n5238) );
  INV_X1 U5292 ( .A(n5256), .ZN(n5154) );
  NAND2_X1 U5293 ( .A1(n5159), .A2(n5158), .ZN(n5469) );
  NOR2_X1 U5294 ( .A1(n5047), .A2(n4509), .ZN(n4806) );
  NAND2_X1 U5295 ( .A1(n5144), .A2(n5143), .ZN(n5282) );
  XNOR2_X1 U5296 ( .A(n5138), .B(SI_11_), .ZN(n5296) );
  AND2_X1 U5297 ( .A1(n5447), .A2(n5450), .ZN(n5294) );
  NAND2_X1 U5298 ( .A1(n4618), .A2(n4623), .ZN(n5448) );
  NAND2_X1 U5299 ( .A1(n5111), .A2(n5110), .ZN(n4869) );
  OR2_X1 U5300 ( .A1(n4483), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5111) );
  AOI21_X1 U5301 ( .B1(n6421), .B2(n6420), .A(n6430), .ZN(n6467) );
  AND2_X1 U5302 ( .A1(n4928), .A2(n4932), .ZN(n4926) );
  INV_X1 U5303 ( .A(n7855), .ZN(n4932) );
  NOR2_X1 U5304 ( .A1(n4939), .A2(n8621), .ZN(n4938) );
  INV_X1 U5305 ( .A(n4940), .ZN(n4939) );
  NOR2_X1 U5306 ( .A1(n8621), .A2(n4943), .ZN(n4936) );
  NAND2_X1 U5307 ( .A1(n5073), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5552) );
  AOI21_X1 U5308 ( .B1(n8564), .B2(n8565), .A(n6409), .ZN(n6412) );
  INV_X1 U5309 ( .A(n6339), .ZN(n4593) );
  INV_X1 U5310 ( .A(n6340), .ZN(n4594) );
  NAND2_X1 U5311 ( .A1(n8581), .A2(n8580), .ZN(n4923) );
  AOI21_X1 U5312 ( .B1(n4943), .B2(n4941), .A(n6394), .ZN(n4940) );
  INV_X1 U5313 ( .A(n8233), .ZN(n4941) );
  XNOR2_X1 U5314 ( .A(n6404), .B(n6402), .ZN(n8630) );
  INV_X1 U5315 ( .A(n8680), .ZN(n6688) );
  XNOR2_X1 U5316 ( .A(n7493), .B(n6422), .ZN(n6336) );
  INV_X1 U5317 ( .A(n4954), .ZN(n4950) );
  NAND2_X1 U5318 ( .A1(n6415), .A2(n8602), .ZN(n4958) );
  NAND2_X1 U5319 ( .A1(n6417), .A2(n6416), .ZN(n4957) );
  NAND2_X1 U5320 ( .A1(n5326), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5332) );
  AND4_X1 U5321 ( .A1(n5345), .A2(n5344), .A3(n5343), .A4(n5342), .ZN(n6327)
         );
  OR2_X1 U5322 ( .A1(n4485), .A2(n5341), .ZN(n5343) );
  INV_X1 U5323 ( .A(n8739), .ZN(n4703) );
  NAND2_X1 U5324 ( .A1(n8294), .A2(n8293), .ZN(n8965) );
  NOR2_X1 U5325 ( .A1(n8929), .A2(n8920), .ZN(n8898) );
  NAND2_X1 U5326 ( .A1(n8898), .A2(n8445), .ZN(n8899) );
  NAND2_X1 U5327 ( .A1(n8916), .A2(n8915), .ZN(n8914) );
  NAND2_X1 U5328 ( .A1(n5045), .A2(n4963), .ZN(n4959) );
  NAND2_X1 U5329 ( .A1(n4906), .A2(n4907), .ZN(n8945) );
  AOI21_X1 U5330 ( .B1(n4788), .B2(n4502), .A(n4787), .ZN(n4786) );
  INV_X1 U5331 ( .A(n8506), .ZN(n4787) );
  AND2_X1 U5332 ( .A1(n9025), .A2(n8669), .ZN(n4979) );
  OR2_X1 U5333 ( .A1(n7983), .A2(n9025), .ZN(n8073) );
  AND2_X1 U5334 ( .A1(n8419), .A2(n8418), .ZN(n8482) );
  INV_X1 U5335 ( .A(n4974), .ZN(n4973) );
  AOI21_X1 U5336 ( .B1(n4974), .B2(n8500), .A(n4499), .ZN(n4972) );
  NOR2_X1 U5337 ( .A1(n9919), .A2(n4977), .ZN(n4974) );
  AND2_X1 U5338 ( .A1(n8412), .A2(n8411), .ZN(n9919) );
  AOI21_X1 U5339 ( .B1(n7736), .B2(n10363), .A(n7473), .ZN(n7612) );
  NAND2_X1 U5340 ( .A1(n7612), .A2(n8410), .ZN(n7611) );
  OR2_X1 U5341 ( .A1(n7389), .A2(n10257), .ZN(n4965) );
  OR2_X1 U5342 ( .A1(n10252), .A2(n7389), .ZN(n7421) );
  AOI21_X1 U5343 ( .B1(n8380), .B2(n4782), .A(n4781), .ZN(n4780) );
  INV_X1 U5344 ( .A(n8389), .ZN(n4781) );
  NOR2_X1 U5345 ( .A1(n10289), .A2(n7458), .ZN(n10253) );
  OR2_X1 U5346 ( .A1(n5424), .A2(n5423), .ZN(n5425) );
  NAND2_X1 U5347 ( .A1(n5383), .A2(n5382), .ZN(n8271) );
  OR2_X1 U5348 ( .A1(n5856), .A2(n5429), .ZN(n5383) );
  AND2_X1 U5349 ( .A1(n5381), .A2(n5054), .ZN(n5382) );
  NOR2_X1 U5350 ( .A1(n7271), .A2(n4726), .ZN(n8270) );
  NAND2_X1 U5351 ( .A1(n6638), .A2(n10315), .ZN(n4726) );
  NAND2_X1 U5352 ( .A1(n7126), .A2(n9072), .ZN(n4570) );
  OR2_X1 U5353 ( .A1(n5710), .A2(n10309), .ZN(n6426) );
  INV_X1 U5354 ( .A(n8964), .ZN(n4911) );
  NAND2_X1 U5355 ( .A1(n8965), .A2(n9026), .ZN(n4910) );
  NAND2_X1 U5356 ( .A1(n5222), .A2(n5221), .ZN(n8248) );
  INV_X1 U5357 ( .A(n5084), .ZN(n4981) );
  NAND2_X1 U5358 ( .A1(n4504), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5681) );
  NOR2_X1 U5359 ( .A1(n4530), .A2(n4947), .ZN(n4946) );
  INV_X1 U5360 ( .A(n6023), .ZN(n4858) );
  NAND2_X1 U5361 ( .A1(n5941), .A2(n5940), .ZN(n7555) );
  NAND2_X1 U5362 ( .A1(n4848), .A2(n6169), .ZN(n4847) );
  NAND2_X1 U5363 ( .A1(n9147), .A2(n9148), .ZN(n4848) );
  NAND2_X1 U5364 ( .A1(n4840), .A2(n9128), .ZN(n4839) );
  AOI21_X1 U5365 ( .B1(n5802), .B2(n7600), .A(n4511), .ZN(n5800) );
  NAND2_X1 U5366 ( .A1(n4835), .A2(n4837), .ZN(n6289) );
  NAND2_X1 U5367 ( .A1(n4833), .A2(n4831), .ZN(n4837) );
  INV_X1 U5368 ( .A(n9099), .ZN(n4836) );
  NAND2_X1 U5369 ( .A1(n4684), .A2(n4683), .ZN(n4682) );
  NAND2_X1 U5370 ( .A1(n9428), .A2(n9532), .ZN(n4683) );
  AND4_X1 U5371 ( .A1(n5922), .A2(n5921), .A3(n5920), .A4(n5919), .ZN(n7714)
         );
  OR2_X1 U5372 ( .A1(n6729), .A2(n6728), .ZN(n4710) );
  NAND2_X1 U5373 ( .A1(n10052), .A2(n10051), .ZN(n4723) );
  AOI21_X1 U5374 ( .B1(n4721), .B2(n4720), .A(n4725), .ZN(n4719) );
  INV_X1 U5375 ( .A(n10051), .ZN(n4720) );
  AND2_X1 U5376 ( .A1(n6741), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4725) );
  NOR2_X1 U5377 ( .A1(n9507), .A2(n9508), .ZN(n9510) );
  INV_X1 U5378 ( .A(n4714), .ZN(n9506) );
  OR2_X1 U5379 ( .A1(n10077), .A2(n8140), .ZN(n4705) );
  NAND2_X1 U5380 ( .A1(n4883), .A2(n9416), .ZN(n4882) );
  INV_X1 U5381 ( .A(n4886), .ZN(n4883) );
  NAND2_X1 U5382 ( .A1(n9614), .A2(n4891), .ZN(n4887) );
  NOR2_X1 U5383 ( .A1(n4889), .A2(n9575), .ZN(n4886) );
  NAND2_X1 U5384 ( .A1(n4887), .A2(n4888), .ZN(n9574) );
  INV_X1 U5385 ( .A(n4889), .ZN(n4888) );
  NAND2_X1 U5386 ( .A1(n5005), .A2(n5003), .ZN(n5002) );
  NAND2_X1 U5387 ( .A1(n9325), .A2(n5004), .ZN(n5003) );
  NAND2_X1 U5388 ( .A1(n9602), .A2(n9618), .ZN(n5004) );
  OR2_X1 U5389 ( .A1(n9327), .A2(n9326), .ZN(n9589) );
  NOR2_X1 U5390 ( .A1(n9619), .A2(n9769), .ZN(n9598) );
  NAND2_X1 U5391 ( .A1(n9293), .A2(n9298), .ZN(n9605) );
  OAI21_X1 U5392 ( .B1(n9677), .B2(n9330), .A(n9331), .ZN(n9662) );
  AOI21_X1 U5393 ( .B1(n9691), .B2(n8537), .A(n8536), .ZN(n9675) );
  NOR2_X1 U5394 ( .A1(n9800), .A2(n9718), .ZN(n8536) );
  OAI21_X1 U5395 ( .B1(n8551), .B2(n8550), .A(n9388), .ZN(n9731) );
  AND2_X1 U5396 ( .A1(n9816), .A2(n9734), .ZN(n8532) );
  AOI21_X1 U5397 ( .B1(n8162), .B2(n8161), .A(n8011), .ZN(n8012) );
  AOI21_X1 U5398 ( .B1(n5025), .B2(n5023), .A(n4531), .ZN(n5022) );
  INV_X1 U5399 ( .A(n5029), .ZN(n5023) );
  INV_X1 U5400 ( .A(n5025), .ZN(n5024) );
  AND2_X1 U5401 ( .A1(n9255), .A2(n9253), .ZN(n9333) );
  NAND2_X1 U5402 ( .A1(n4881), .A2(n9226), .ZN(n4880) );
  INV_X1 U5403 ( .A(n5822), .ZN(n6137) );
  NAND2_X1 U5404 ( .A1(n7678), .A2(n7592), .ZN(n7801) );
  NAND2_X1 U5405 ( .A1(n7622), .A2(n7581), .ZN(n7677) );
  OR2_X1 U5406 ( .A1(n9368), .A2(n9998), .ZN(n9683) );
  NAND2_X1 U5407 ( .A1(n7590), .A2(n9430), .ZN(n9336) );
  AND2_X1 U5408 ( .A1(n7598), .A2(n9998), .ZN(n9733) );
  INV_X1 U5409 ( .A(n9683), .ZN(n9735) );
  NAND2_X1 U5410 ( .A1(n9216), .A2(n9215), .ZN(n9746) );
  NAND2_X1 U5411 ( .A1(n9212), .A2(n9211), .ZN(n9310) );
  NAND2_X1 U5412 ( .A1(n5731), .A2(n5732), .ZN(n4674) );
  INV_X1 U5413 ( .A(n5041), .ZN(n4676) );
  NAND2_X1 U5414 ( .A1(n4678), .A2(n5991), .ZN(n4679) );
  NOR2_X1 U5415 ( .A1(n5039), .A2(n5041), .ZN(n4678) );
  XNOR2_X1 U5416 ( .A(n5617), .B(n5616), .ZN(n8064) );
  XNOR2_X1 U5417 ( .A(n5601), .B(n5600), .ZN(n7972) );
  XNOR2_X1 U5418 ( .A(n5581), .B(n5580), .ZN(n7950) );
  OR2_X1 U5419 ( .A1(n5745), .A2(n5724), .ZN(n5749) );
  NOR2_X1 U5420 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5746) );
  OR2_X1 U5421 ( .A1(n5193), .A2(n5192), .ZN(n5543) );
  XNOR2_X1 U5422 ( .A(n5532), .B(n5531), .ZN(n7799) );
  CLKBUF_X1 U5423 ( .A(n6283), .Z(n6284) );
  NAND2_X1 U5424 ( .A1(n5779), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5743) );
  OAI22_X1 U5425 ( .A1(n4617), .A2(n4616), .B1(n4619), .B2(n5451), .ZN(n4615)
         );
  NAND2_X1 U5426 ( .A1(n4622), .A2(n5128), .ZN(n5308) );
  AOI22_X2 U5427 ( .A1(n4809), .A2(n4807), .B1(n4810), .B2(n4505), .ZN(n5314)
         );
  NOR2_X1 U5428 ( .A1(n4808), .A2(n4872), .ZN(n4807) );
  OAI21_X1 U5429 ( .B1(n4872), .B2(n5408), .A(n5427), .ZN(n4810) );
  INV_X1 U5430 ( .A(n5122), .ZN(n4872) );
  XNOR2_X1 U5431 ( .A(n5123), .B(n7018), .ZN(n5427) );
  NAND2_X1 U5432 ( .A1(n4809), .A2(n5119), .ZN(n5409) );
  NAND2_X1 U5433 ( .A1(n5374), .A2(n4637), .ZN(n4636) );
  AND2_X1 U5434 ( .A1(n5373), .A2(n5113), .ZN(n4637) );
  AND2_X1 U5435 ( .A1(n5899), .A2(n5898), .ZN(n6563) );
  XNOR2_X1 U5436 ( .A(n5115), .B(n5114), .ZN(n5375) );
  NAND2_X1 U5437 ( .A1(n8581), .A2(n4922), .ZN(n4919) );
  INV_X1 U5438 ( .A(n4918), .ZN(n4922) );
  AND2_X1 U5439 ( .A1(n4917), .A2(n7407), .ZN(n4916) );
  NAND2_X1 U5440 ( .A1(n4918), .A2(n4920), .ZN(n4917) );
  NAND2_X1 U5441 ( .A1(n4596), .A2(n4599), .ZN(n8197) );
  AND2_X1 U5442 ( .A1(n4597), .A2(n6385), .ZN(n4596) );
  NAND2_X1 U5443 ( .A1(n5232), .A2(n5231), .ZN(n8203) );
  OR2_X1 U5444 ( .A1(n6685), .A2(n6684), .ZN(n4955) );
  AND2_X1 U5445 ( .A1(n6456), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8639) );
  NOR2_X1 U5446 ( .A1(n6665), .A2(n6333), .ZN(n6645) );
  XNOR2_X1 U5447 ( .A(n6336), .B(n6334), .ZN(n6646) );
  XNOR2_X1 U5448 ( .A(n4793), .B(n8327), .ZN(n4792) );
  INV_X1 U5449 ( .A(n8474), .ZN(n4794) );
  NAND2_X1 U5450 ( .A1(n4651), .A2(n8521), .ZN(n4580) );
  OR2_X1 U5451 ( .A1(n8520), .A2(n4569), .ZN(n4651) );
  OR2_X1 U5452 ( .A1(n5385), .A2(n5384), .ZN(n5387) );
  NAND2_X1 U5453 ( .A1(n4695), .A2(n9065), .ZN(n4694) );
  NAND2_X1 U5454 ( .A1(n4535), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n4693) );
  XNOR2_X1 U5455 ( .A(n8734), .B(n8726), .ZN(n8178) );
  NAND2_X1 U5456 ( .A1(n4512), .A2(n9922), .ZN(n8794) );
  AOI21_X1 U5457 ( .B1(n4969), .B2(n4971), .A(n4523), .ZN(n4967) );
  NAND2_X1 U5458 ( .A1(n4912), .A2(n8816), .ZN(n8963) );
  OR2_X1 U5459 ( .A1(n4913), .A2(n9910), .ZN(n4912) );
  XNOR2_X1 U5460 ( .A(n8812), .B(n8811), .ZN(n4913) );
  NAND2_X1 U5461 ( .A1(n8880), .A2(n8881), .ZN(n4576) );
  NAND2_X1 U5462 ( .A1(n5548), .A2(n5547), .ZN(n8991) );
  OR2_X1 U5463 ( .A1(n7112), .A2(n6452), .ZN(n8903) );
  NAND2_X1 U5464 ( .A1(n5401), .A2(n5400), .ZN(n7302) );
  NAND2_X1 U5465 ( .A1(n8794), .A2(n8958), .ZN(n9032) );
  XNOR2_X1 U5466 ( .A(n5634), .B(n5633), .ZN(n8479) );
  INV_X1 U5467 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U5468 ( .A1(n5631), .A2(n5630), .ZN(n5632) );
  NAND2_X1 U5469 ( .A1(n5736), .A2(n5735), .ZN(n9779) );
  INV_X1 U5470 ( .A(n9655), .ZN(n9786) );
  NAND2_X1 U5471 ( .A1(n9543), .A2(n4749), .ZN(n9962) );
  OR2_X1 U5472 ( .A1(n9544), .A2(n9545), .ZN(n4749) );
  NAND2_X1 U5473 ( .A1(n10180), .A2(n7587), .ZN(n7666) );
  AND2_X1 U5474 ( .A1(n9751), .A2(n9752), .ZN(n5014) );
  OR2_X1 U5475 ( .A1(n9551), .A2(n4896), .ZN(n5012) );
  NOR2_X1 U5476 ( .A1(n9364), .A2(n5011), .ZN(n5010) );
  NAND2_X1 U5477 ( .A1(n4672), .A2(n9340), .ZN(n9229) );
  XNOR2_X1 U5478 ( .A(n9218), .B(n4673), .ZN(n4672) );
  NOR2_X1 U5479 ( .A1(n8339), .A2(n4649), .ZN(n8395) );
  NAND2_X1 U5480 ( .A1(n8337), .A2(n8465), .ZN(n4650) );
  INV_X1 U5481 ( .A(n4527), .ZN(n4632) );
  NAND2_X1 U5482 ( .A1(n9274), .A2(n9318), .ZN(n4670) );
  NAND2_X1 U5483 ( .A1(n9271), .A2(n4673), .ZN(n4669) );
  OAI21_X1 U5484 ( .B1(n4639), .B2(n4638), .A(n4532), .ZN(n8422) );
  NAND2_X1 U5485 ( .A1(n8414), .A2(n8413), .ZN(n4638) );
  AOI21_X1 U5486 ( .B1(n4642), .B2(n4641), .A(n4640), .ZN(n4639) );
  OAI21_X1 U5487 ( .B1(n9274), .B2(n4495), .A(n4667), .ZN(n4666) );
  OR2_X1 U5488 ( .A1(n9271), .A2(n4668), .ZN(n4667) );
  NAND2_X1 U5489 ( .A1(n4498), .A2(n4673), .ZN(n4668) );
  NAND2_X1 U5490 ( .A1(n4664), .A2(n4662), .ZN(n4671) );
  NOR2_X1 U5491 ( .A1(n4666), .A2(n4663), .ZN(n4662) );
  INV_X1 U5492 ( .A(n9331), .ZN(n4663) );
  NAND2_X1 U5493 ( .A1(n4664), .A2(n4665), .ZN(n9278) );
  INV_X1 U5494 ( .A(n4666), .ZN(n4665) );
  AOI21_X1 U5495 ( .B1(n4534), .B2(n8438), .A(n8478), .ZN(n4625) );
  NAND2_X1 U5496 ( .A1(n8442), .A2(n8441), .ZN(n4825) );
  NOR2_X1 U5497 ( .A1(n8901), .A2(n4827), .ZN(n4826) );
  AND2_X1 U5498 ( .A1(n8440), .A2(n8478), .ZN(n4827) );
  AND2_X1 U5499 ( .A1(n8444), .A2(n8465), .ZN(n4823) );
  NAND2_X1 U5500 ( .A1(n9292), .A2(n4686), .ZN(n9303) );
  INV_X1 U5501 ( .A(n8459), .ZN(n4812) );
  AOI21_X1 U5502 ( .B1(n8450), .B2(n4645), .A(n4644), .ZN(n4643) );
  AND2_X1 U5503 ( .A1(n8875), .A2(n8449), .ZN(n4645) );
  NAND2_X1 U5504 ( .A1(n4817), .A2(n8451), .ZN(n4644) );
  NAND2_X1 U5505 ( .A1(n8453), .A2(n8465), .ZN(n4816) );
  NOR2_X1 U5506 ( .A1(n8451), .A2(n8478), .ZN(n4814) );
  INV_X1 U5507 ( .A(n4929), .ZN(n4605) );
  AOI21_X1 U5508 ( .B1(n4815), .B2(n4813), .A(n4811), .ZN(n8464) );
  NOR2_X1 U5509 ( .A1(n8510), .A2(n4814), .ZN(n4813) );
  OAI21_X1 U5510 ( .B1(n4643), .B2(n5657), .A(n4816), .ZN(n4815) );
  NAND2_X1 U5511 ( .A1(n4812), .A2(n8312), .ZN(n4811) );
  NOR2_X2 U5512 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5243) );
  INV_X1 U5513 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5739) );
  INV_X1 U5514 ( .A(n5053), .ZN(n4798) );
  NOR2_X1 U5515 ( .A1(n4804), .A2(n5282), .ZN(n4803) );
  NAND2_X1 U5516 ( .A1(n4583), .A2(n4582), .ZN(n5138) );
  NAND2_X1 U5517 ( .A1(n4483), .A2(n6878), .ZN(n4582) );
  OR2_X1 U5518 ( .A1(n4483), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n4583) );
  NAND2_X1 U5519 ( .A1(n5130), .A2(n5129), .ZN(n5447) );
  OR2_X1 U5520 ( .A1(n8965), .A2(n8314), .ZN(n8466) );
  NOR2_X1 U5521 ( .A1(n8827), .A2(n5671), .ZN(n8295) );
  INV_X1 U5522 ( .A(n8857), .ZN(n4984) );
  AND2_X1 U5523 ( .A1(n8898), .A2(n4546), .ZN(n8837) );
  NOR2_X1 U5524 ( .A1(n8872), .A2(n8863), .ZN(n8848) );
  NOR2_X1 U5525 ( .A1(n8980), .A2(n4733), .ZN(n4731) );
  NOR2_X1 U5526 ( .A1(n8333), .A2(n8901), .ZN(n4903) );
  NAND2_X1 U5527 ( .A1(n5045), .A2(n4962), .ZN(n4961) );
  INV_X1 U5528 ( .A(n4964), .ZN(n4962) );
  NOR2_X1 U5529 ( .A1(n9020), .A2(n8248), .ZN(n4740) );
  NOR2_X1 U5530 ( .A1(n9921), .A2(n9917), .ZN(n7935) );
  OR2_X1 U5531 ( .A1(n7528), .A2(n4745), .ZN(n4744) );
  NAND2_X1 U5532 ( .A1(n10363), .A2(n10348), .ZN(n4745) );
  NAND2_X1 U5533 ( .A1(n5066), .A2(n5065), .ZN(n5461) );
  INV_X1 U5534 ( .A(n8386), .ZN(n4783) );
  NAND2_X1 U5535 ( .A1(n5220), .A2(n4948), .ZN(n4947) );
  INV_X1 U5536 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4948) );
  NAND3_X1 U5537 ( .A1(n4822), .A2(n9537), .A3(n4821), .ZN(n4820) );
  INV_X1 U5538 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4821) );
  INV_X1 U5539 ( .A(n6543), .ZN(n5799) );
  NAND2_X1 U5540 ( .A1(n9492), .A2(n5802), .ZN(n5805) );
  AND2_X1 U5541 ( .A1(n5803), .A2(n5058), .ZN(n5804) );
  NAND2_X1 U5542 ( .A1(n4843), .A2(n6185), .ZN(n4842) );
  OR2_X1 U5543 ( .A1(n6184), .A2(n6183), .ZN(n6185) );
  NAND2_X1 U5544 ( .A1(n4845), .A2(n4847), .ZN(n4843) );
  INV_X1 U5545 ( .A(n9128), .ZN(n4834) );
  AOI21_X1 U5546 ( .B1(n9128), .B2(n4832), .A(n6222), .ZN(n4831) );
  INV_X1 U5547 ( .A(n9077), .ZN(n4832) );
  NOR2_X1 U5548 ( .A1(n4857), .A2(n6094), .ZN(n4852) );
  NOR2_X1 U5549 ( .A1(n9310), .A2(n9365), .ZN(n9454) );
  OAI21_X1 U5550 ( .B1(n9467), .B2(n9368), .A(n9367), .ZN(n4685) );
  AOI22_X1 U5551 ( .A1(n4658), .A2(n4520), .B1(n9319), .B2(n9320), .ZN(n9322)
         );
  OR2_X1 U5552 ( .A1(n9319), .A2(n4542), .ZN(n4658) );
  OR2_X1 U5553 ( .A1(n9865), .A2(n9866), .ZN(n4711) );
  OR2_X1 U5554 ( .A1(n10061), .A2(n4715), .ZN(n4714) );
  AND2_X1 U5555 ( .A1(n10066), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4715) );
  NOR2_X1 U5556 ( .A1(n9414), .A2(n9417), .ZN(n4885) );
  OR2_X1 U5557 ( .A1(n9755), .A2(n9572), .ZN(n9419) );
  NAND2_X1 U5558 ( .A1(n9571), .A2(n4766), .ZN(n4765) );
  INV_X1 U5559 ( .A(n4767), .ZN(n4766) );
  NAND2_X1 U5560 ( .A1(n9586), .A2(n9602), .ZN(n4767) );
  OR2_X1 U5561 ( .A1(n9776), .A2(n9638), .ZN(n9407) );
  AND2_X1 U5562 ( .A1(n9252), .A2(n9241), .ZN(n8161) );
  NAND2_X1 U5563 ( .A1(n9952), .A2(n8049), .ZN(n5028) );
  NAND2_X1 U5564 ( .A1(n7912), .A2(n5030), .ZN(n5029) );
  NOR2_X1 U5565 ( .A1(n5891), .A2(n5881), .ZN(n5915) );
  NAND2_X1 U5566 ( .A1(n7678), .A2(n4654), .ZN(n4652) );
  NOR2_X1 U5567 ( .A1(n4656), .A2(n7593), .ZN(n4654) );
  OR2_X1 U5568 ( .A1(n9749), .A2(n9557), .ZN(n9418) );
  NAND2_X1 U5569 ( .A1(n4754), .A2(n4753), .ZN(n9666) );
  INV_X1 U5570 ( .A(n5753), .ZN(n5747) );
  OR2_X1 U5571 ( .A1(n5483), .A2(n5487), .ZN(n5167) );
  AND2_X1 U5572 ( .A1(n5171), .A2(n5170), .ZN(n5172) );
  INV_X1 U5573 ( .A(n4803), .ZN(n4802) );
  AOI21_X1 U5574 ( .B1(n4803), .B2(n4801), .A(n4800), .ZN(n4799) );
  INV_X1 U5575 ( .A(n5144), .ZN(n4800) );
  INV_X1 U5576 ( .A(n5137), .ZN(n4801) );
  NAND2_X1 U5577 ( .A1(n5135), .A2(SI_10_), .ZN(n5449) );
  INV_X1 U5578 ( .A(n4619), .ZN(n4617) );
  NOR2_X1 U5579 ( .A1(n4623), .A2(n5451), .ZN(n4616) );
  AOI21_X1 U5580 ( .B1(n4623), .B2(n4621), .A(n4620), .ZN(n4619) );
  INV_X1 U5581 ( .A(n5447), .ZN(n4620) );
  INV_X1 U5582 ( .A(n5128), .ZN(n4621) );
  INV_X1 U5583 ( .A(n5451), .ZN(n4614) );
  INV_X1 U5584 ( .A(n5314), .ZN(n4612) );
  INV_X1 U5585 ( .A(n6372), .ZN(n4933) );
  NAND2_X1 U5586 ( .A1(n7646), .A2(n4929), .ZN(n4927) );
  NAND2_X1 U5587 ( .A1(n4924), .A2(n8580), .ZN(n4918) );
  NOR2_X1 U5588 ( .A1(n7309), .A2(n6349), .ZN(n6350) );
  NAND2_X1 U5589 ( .A1(n4610), .A2(n6354), .ZN(n8581) );
  XNOR2_X1 U5590 ( .A(n9002), .B(n6422), .ZN(n6400) );
  AND2_X1 U5591 ( .A1(n8148), .A2(n4600), .ZN(n4598) );
  NAND2_X1 U5592 ( .A1(n8149), .A2(n8148), .ZN(n4599) );
  OR2_X1 U5593 ( .A1(n5535), .A2(n8636), .ZN(n5550) );
  AND2_X1 U5594 ( .A1(n6694), .A2(n6343), .ZN(n4953) );
  NAND2_X1 U5595 ( .A1(n6345), .A2(n6346), .ZN(n4954) );
  NAND2_X1 U5596 ( .A1(n4958), .A2(n4957), .ZN(n8644) );
  NAND2_X1 U5597 ( .A1(n8480), .A2(n8479), .ZN(n8520) );
  NAND2_X1 U5598 ( .A1(n5440), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U5599 ( .A1(n5440), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U5600 ( .A1(n5440), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5096) );
  AND2_X1 U5601 ( .A1(n5558), .A2(n5557), .ZN(n8634) );
  INV_X1 U5602 ( .A(n5440), .ZN(n5666) );
  NAND2_X1 U5603 ( .A1(n5440), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5364) );
  INV_X1 U5604 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4695) );
  XNOR2_X1 U5605 ( .A(n9879), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n9876) );
  OR2_X1 U5606 ( .A1(n7155), .A2(n4560), .ZN(n4700) );
  NAND2_X1 U5607 ( .A1(n4700), .A2(n7139), .ZN(n4699) );
  AOI21_X1 U5608 ( .B1(n7330), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7322), .ZN(
        n8688) );
  NOR2_X1 U5609 ( .A1(n7757), .A2(n4691), .ZN(n8715) );
  AND2_X1 U5610 ( .A1(n7758), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4691) );
  NAND2_X1 U5611 ( .A1(n8715), .A2(n8716), .ZN(n8714) );
  AOI21_X1 U5612 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7866), .A(n7865), .ZN(
        n7869) );
  NAND2_X1 U5613 ( .A1(n7961), .A2(n4697), .ZN(n7963) );
  OR2_X1 U5614 ( .A1(n7962), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4697) );
  NAND2_X1 U5615 ( .A1(n7963), .A2(n7964), .ZN(n8176) );
  AND2_X1 U5616 ( .A1(n8800), .A2(n4970), .ZN(n4969) );
  NAND2_X1 U5617 ( .A1(n8833), .A2(n5615), .ZN(n4970) );
  INV_X1 U5618 ( .A(n5615), .ZN(n4971) );
  NOR2_X1 U5619 ( .A1(n8313), .A2(n8460), .ZN(n8812) );
  AND2_X1 U5620 ( .A1(n8295), .A2(n8806), .ZN(n8804) );
  OR3_X1 U5621 ( .A1(n5623), .A2(n6471), .A3(n5622), .ZN(n8808) );
  NAND2_X1 U5622 ( .A1(n8312), .A2(n8456), .ZN(n8800) );
  AND2_X1 U5623 ( .A1(n4986), .A2(n4559), .ZN(n4985) );
  NAND2_X1 U5624 ( .A1(n8863), .A2(n4987), .ZN(n4986) );
  INV_X1 U5625 ( .A(n4990), .ZN(n4987) );
  NAND2_X1 U5626 ( .A1(n8863), .A2(n4989), .ZN(n4988) );
  INV_X1 U5627 ( .A(n8881), .ZN(n4989) );
  NAND2_X1 U5628 ( .A1(n8451), .A2(n8454), .ZN(n8857) );
  OR2_X1 U5629 ( .A1(n5571), .A2(n8607), .ZN(n5589) );
  NAND2_X1 U5630 ( .A1(n4772), .A2(n4770), .ZN(n8872) );
  NAND2_X1 U5631 ( .A1(n4771), .A2(n5656), .ZN(n4770) );
  NAND2_X1 U5632 ( .A1(n8914), .A2(n4524), .ZN(n4772) );
  INV_X1 U5633 ( .A(n4899), .ZN(n4771) );
  NAND2_X1 U5634 ( .A1(n8898), .A2(n4731), .ZN(n8865) );
  AND2_X1 U5635 ( .A1(n5656), .A2(n8332), .ZN(n8881) );
  NOR2_X1 U5636 ( .A1(n4898), .A2(n8444), .ZN(n8882) );
  INV_X1 U5637 ( .A(n4901), .ZN(n4898) );
  AND2_X1 U5638 ( .A1(n8881), .A2(n4900), .ZN(n4899) );
  INV_X1 U5639 ( .A(n8444), .ZN(n4900) );
  NAND2_X1 U5640 ( .A1(n8914), .A2(n4903), .ZN(n4901) );
  OR2_X1 U5641 ( .A1(n9002), .A2(n8664), .ZN(n5525) );
  OR2_X1 U5642 ( .A1(n8934), .A2(n8633), .ZN(n5046) );
  NAND2_X1 U5643 ( .A1(n8123), .A2(n4736), .ZN(n8929) );
  NOR2_X1 U5644 ( .A1(n9002), .A2(n4738), .ZN(n4736) );
  NAND2_X1 U5645 ( .A1(n5071), .A2(n5070), .ZN(n5505) );
  NAND2_X1 U5646 ( .A1(n8123), .A2(n8128), .ZN(n8247) );
  NAND2_X1 U5647 ( .A1(n8123), .A2(n4740), .ZN(n8949) );
  OR2_X1 U5648 ( .A1(n5235), .A2(n8748), .ZN(n5493) );
  NOR2_X1 U5649 ( .A1(n8203), .A2(n8073), .ZN(n8123) );
  NAND2_X1 U5650 ( .A1(n5069), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5235) );
  INV_X1 U5651 ( .A(n5479), .ZN(n5069) );
  NAND2_X1 U5652 ( .A1(n5067), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5269) );
  INV_X1 U5653 ( .A(n5277), .ZN(n5067) );
  NAND2_X1 U5654 ( .A1(n5068), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5477) );
  INV_X1 U5655 ( .A(n5269), .ZN(n5068) );
  NAND2_X1 U5656 ( .A1(n7515), .A2(n8398), .ZN(n7606) );
  NAND2_X1 U5657 ( .A1(n5648), .A2(n8398), .ZN(n4773) );
  AND2_X1 U5658 ( .A1(n5650), .A2(n4775), .ZN(n4774) );
  NAND2_X1 U5659 ( .A1(n4743), .A2(n4742), .ZN(n9921) );
  NOR2_X1 U5660 ( .A1(n4744), .A2(n5468), .ZN(n4742) );
  INV_X1 U5661 ( .A(n7421), .ZN(n4743) );
  AND2_X1 U5662 ( .A1(n8399), .A2(n8402), .ZN(n8499) );
  NOR3_X1 U5663 ( .A1(n7421), .A2(n7528), .A3(n7425), .ZN(n7523) );
  NAND2_X1 U5664 ( .A1(n7415), .A2(n8341), .ZN(n7515) );
  NOR2_X1 U5665 ( .A1(n7421), .A2(n7425), .ZN(n7522) );
  NAND2_X1 U5666 ( .A1(n7377), .A2(n8495), .ZN(n7376) );
  NAND2_X1 U5667 ( .A1(n8340), .A2(n8392), .ZN(n8495) );
  NAND2_X1 U5668 ( .A1(n8390), .A2(n8389), .ZN(n10261) );
  NAND2_X1 U5669 ( .A1(n7450), .A2(n8386), .ZN(n10262) );
  NAND2_X1 U5670 ( .A1(n4784), .A2(n8492), .ZN(n7450) );
  INV_X1 U5671 ( .A(n7448), .ZN(n4784) );
  NOR2_X1 U5672 ( .A1(n5392), .A2(n8488), .ZN(n5393) );
  INV_X1 U5673 ( .A(n8649), .ZN(n10258) );
  NAND2_X1 U5674 ( .A1(n8299), .A2(n8298), .ZN(n8795) );
  NAND2_X1 U5675 ( .A1(n9210), .A2(n8297), .ZN(n8299) );
  NAND2_X1 U5676 ( .A1(n5609), .A2(n5608), .ZN(n8970) );
  NAND2_X1 U5677 ( .A1(n5534), .A2(n5533), .ZN(n8920) );
  NAND2_X1 U5678 ( .A1(n5249), .A2(n5248), .ZN(n9025) );
  NAND2_X1 U5679 ( .A1(n10266), .A2(n10335), .ZN(n10368) );
  NOR2_X1 U5680 ( .A1(n5227), .A2(n4778), .ZN(n4777) );
  NAND2_X1 U5681 ( .A1(n5089), .A2(n5687), .ZN(n4778) );
  CLKBUF_X1 U5682 ( .A(n5660), .Z(n5661) );
  NAND2_X1 U5683 ( .A1(n4601), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U5684 ( .A1(n4980), .A2(n4945), .ZN(n4601) );
  INV_X1 U5685 ( .A(n4947), .ZN(n4945) );
  INV_X1 U5686 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5630) );
  AOI21_X1 U5687 ( .B1(n4857), .B2(n4855), .A(n4529), .ZN(n4854) );
  INV_X1 U5688 ( .A(n7923), .ZN(n4855) );
  AND2_X1 U5689 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5892) );
  AND2_X1 U5690 ( .A1(n5988), .A2(n5962), .ZN(n4859) );
  OR2_X1 U5691 ( .A1(n8559), .A2(n6566), .ZN(n7579) );
  AOI21_X1 U5692 ( .B1(n4862), .B2(n9120), .A(n6135), .ZN(n4861) );
  AOI21_X1 U5693 ( .B1(n9110), .B2(n4860), .A(n4863), .ZN(n6136) );
  INV_X1 U5694 ( .A(n9120), .ZN(n4860) );
  NAND2_X1 U5695 ( .A1(n9136), .A2(n5874), .ZN(n7534) );
  NAND2_X1 U5696 ( .A1(n5829), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4660) );
  INV_X1 U5697 ( .A(n4718), .ZN(n4717) );
  AOI21_X1 U5698 ( .B1(n4719), .B2(n4722), .A(n6757), .ZN(n4718) );
  NOR2_X1 U5699 ( .A1(n7790), .A2(n4716), .ZN(n10063) );
  AND2_X1 U5700 ( .A1(n7791), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4716) );
  NOR2_X1 U5701 ( .A1(n10063), .A2(n10062), .ZN(n10061) );
  XNOR2_X1 U5702 ( .A(n4714), .B(n7796), .ZN(n7793) );
  NOR2_X1 U5703 ( .A1(n10100), .A2(n4565), .ZN(n9514) );
  NOR2_X1 U5704 ( .A1(n9514), .A2(n9515), .ZN(n9520) );
  NOR2_X1 U5705 ( .A1(n9552), .A2(n9749), .ZN(n9544) );
  NAND2_X1 U5706 ( .A1(n9476), .A2(n9733), .ZN(n4894) );
  NAND2_X1 U5707 ( .A1(n9419), .A2(n9412), .ZN(n9559) );
  NAND2_X1 U5708 ( .A1(n4541), .A2(n4994), .ZN(n4993) );
  NOR3_X1 U5709 ( .A1(n9613), .A2(n8540), .A3(n5000), .ZN(n4992) );
  NOR2_X1 U5710 ( .A1(n9619), .A2(n4767), .ZN(n9582) );
  NOR2_X1 U5711 ( .A1(n9666), .A2(n9786), .ZN(n9650) );
  NAND2_X1 U5712 ( .A1(n9650), .A2(n9633), .ZN(n9627) );
  NAND2_X1 U5713 ( .A1(n6173), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U5714 ( .A1(n9396), .A2(n9279), .ZN(n9658) );
  AND2_X1 U5715 ( .A1(n6155), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6173) );
  AND2_X1 U5716 ( .A1(n9273), .A2(n9369), .ZN(n9700) );
  AND2_X1 U5717 ( .A1(n9804), .A2(n9736), .ZN(n8535) );
  AND2_X1 U5718 ( .A1(n8141), .A2(n4755), .ZN(n9708) );
  NOR2_X1 U5719 ( .A1(n9804), .A2(n4756), .ZN(n4755) );
  INV_X1 U5720 ( .A(n4757), .ZN(n4756) );
  NAND2_X1 U5721 ( .A1(n8141), .A2(n4759), .ZN(n9725) );
  NAND2_X1 U5722 ( .A1(n8141), .A2(n9820), .ZN(n8211) );
  NOR2_X1 U5723 ( .A1(n8208), .A2(n9355), .ZN(n8533) );
  AND2_X1 U5724 ( .A1(n9388), .A2(n9385), .ZN(n9355) );
  AND2_X1 U5725 ( .A1(n8166), .A2(n9966), .ZN(n8141) );
  NOR2_X1 U5726 ( .A1(n8167), .A2(n9825), .ZN(n8166) );
  NAND2_X1 U5727 ( .A1(n9245), .A2(n9226), .ZN(n4878) );
  NAND2_X1 U5728 ( .A1(n4874), .A2(n9244), .ZN(n4873) );
  NAND2_X1 U5729 ( .A1(n6011), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U5730 ( .A1(n5027), .A2(n5028), .ZN(n8008) );
  NAND2_X1 U5731 ( .A1(n7989), .A2(n5029), .ZN(n5027) );
  NAND2_X1 U5732 ( .A1(n4880), .A2(n4879), .ZN(n8010) );
  NOR2_X1 U5733 ( .A1(n4876), .A2(n7992), .ZN(n4879) );
  AND2_X1 U5734 ( .A1(n7893), .A2(n9901), .ZN(n7902) );
  AND2_X1 U5735 ( .A1(n5996), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6011) );
  OAI21_X1 U5736 ( .B1(n7877), .B2(n4536), .A(n5060), .ZN(n7885) );
  NOR2_X1 U5737 ( .A1(n7751), .A2(n7881), .ZN(n7893) );
  INV_X1 U5738 ( .A(n9343), .ZN(n7878) );
  OR2_X1 U5739 ( .A1(n7727), .A2(n7741), .ZN(n7751) );
  NAND2_X1 U5740 ( .A1(n9230), .A2(n9233), .ZN(n9343) );
  AND4_X1 U5741 ( .A1(n5948), .A2(n5947), .A3(n5946), .A4(n5945), .ZN(n7745)
         );
  NAND2_X1 U5742 ( .A1(n5032), .A2(n5033), .ZN(n5031) );
  AND2_X1 U5743 ( .A1(n4492), .A2(n4761), .ZN(n7669) );
  NOR2_X1 U5744 ( .A1(n7842), .A2(n7665), .ZN(n4761) );
  NAND2_X1 U5745 ( .A1(n4762), .A2(n4492), .ZN(n7700) );
  NAND2_X1 U5746 ( .A1(n7801), .A2(n9338), .ZN(n4655) );
  NAND2_X1 U5747 ( .A1(n4762), .A2(n10172), .ZN(n7843) );
  NOR2_X1 U5748 ( .A1(n7684), .A2(n9172), .ZN(n7807) );
  INV_X1 U5749 ( .A(n5015), .ZN(n5011) );
  NAND2_X1 U5750 ( .A1(n6101), .A2(n6100), .ZN(n9816) );
  AND2_X1 U5751 ( .A1(n7570), .A2(n5775), .ZN(n10187) );
  AND2_X1 U5752 ( .A1(n6282), .A2(n9423), .ZN(n7570) );
  AND3_X1 U5753 ( .A1(n6275), .A2(n6268), .A3(n6267), .ZN(n10118) );
  XNOR2_X1 U5754 ( .A(n8296), .B(n4584), .ZN(n9210) );
  INV_X1 U5755 ( .A(SI_30_), .ZN(n4584) );
  XNOR2_X1 U5756 ( .A(n8281), .B(n8195), .ZN(n8542) );
  NAND2_X1 U5757 ( .A1(n5619), .A2(n5618), .ZN(n8189) );
  NAND2_X1 U5758 ( .A1(n5617), .A2(n5616), .ZN(n5619) );
  XNOR2_X1 U5759 ( .A(n5514), .B(n5527), .ZN(n7620) );
  XNOR2_X1 U5760 ( .A(n5488), .B(n5487), .ZN(n7318) );
  OR2_X1 U5761 ( .A1(n5484), .A2(n5483), .ZN(n5486) );
  NAND2_X1 U5762 ( .A1(n5991), .A2(n4865), .ZN(n6098) );
  NOR2_X1 U5763 ( .A1(n5039), .A2(n4867), .ZN(n4865) );
  NAND2_X1 U5764 ( .A1(n4805), .A2(n4806), .ZN(n5283) );
  NAND2_X1 U5765 ( .A1(n5448), .A2(n5137), .ZN(n4805) );
  INV_X1 U5766 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5719) );
  OR2_X1 U5767 ( .A1(n5949), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5952) );
  OR2_X1 U5768 ( .A1(n5952), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5964) );
  INV_X1 U5769 ( .A(n4869), .ZN(n4868) );
  NAND2_X1 U5770 ( .A1(n4870), .A2(n5109), .ZN(n5370) );
  INV_X1 U5771 ( .A(n6436), .ZN(n6463) );
  NAND2_X1 U5772 ( .A1(n8645), .A2(n6468), .ZN(n6469) );
  NAND2_X1 U5773 ( .A1(n4928), .A2(n4927), .ZN(n7854) );
  NAND2_X1 U5774 ( .A1(n4944), .A2(n4943), .ZN(n8570) );
  AND2_X1 U5775 ( .A1(n4944), .A2(n4519), .ZN(n8572) );
  NAND2_X1 U5776 ( .A1(n8234), .A2(n8233), .ZN(n4944) );
  NOR2_X1 U5777 ( .A1(n6434), .A2(n6433), .ZN(n6435) );
  NAND2_X1 U5778 ( .A1(n5318), .A2(n5317), .ZN(n8588) );
  OR2_X1 U5779 ( .A1(n6607), .A2(n5429), .ZN(n5318) );
  NAND2_X1 U5780 ( .A1(n6332), .A2(n4606), .ZN(n6666) );
  NAND2_X1 U5781 ( .A1(n4608), .A2(n4607), .ZN(n4606) );
  INV_X1 U5782 ( .A(n6325), .ZN(n4608) );
  INV_X1 U5783 ( .A(n6326), .ZN(n4607) );
  NAND2_X1 U5784 ( .A1(n6329), .A2(n7240), .ZN(n6330) );
  AOI21_X1 U5785 ( .B1(n4936), .B2(n4940), .A(n4935), .ZN(n4934) );
  NOR2_X1 U5786 ( .A1(n6397), .A2(n6396), .ZN(n4935) );
  OR2_X1 U5787 ( .A1(n6412), .A2(n6411), .ZN(n6413) );
  XNOR2_X1 U5788 ( .A(n6412), .B(n6410), .ZN(n8612) );
  NAND2_X1 U5789 ( .A1(n4591), .A2(n6337), .ZN(n4589) );
  AND2_X1 U5790 ( .A1(n4923), .A2(n4925), .ZN(n7369) );
  OAI21_X1 U5791 ( .B1(n8234), .B2(n4942), .A(n4940), .ZN(n8622) );
  AOI21_X1 U5792 ( .B1(n7646), .B2(n7644), .A(n4931), .ZN(n7733) );
  NAND2_X1 U5793 ( .A1(n7406), .A2(n6364), .ZN(n7499) );
  OAI21_X1 U5794 ( .B1(n6685), .B2(n4951), .A(n4949), .ZN(n7228) );
  NAND2_X1 U5795 ( .A1(n4952), .A2(n4954), .ZN(n4951) );
  OR2_X1 U5796 ( .A1(n4953), .A2(n4950), .ZN(n4949) );
  INV_X1 U5797 ( .A(n6684), .ZN(n4952) );
  NAND2_X1 U5798 ( .A1(n7228), .A2(n7229), .ZN(n7308) );
  AND2_X1 U5799 ( .A1(n6450), .A2(n6449), .ZN(n8654) );
  NAND2_X1 U5800 ( .A1(n5440), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8317) );
  NAND2_X1 U5801 ( .A1(n5440), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U5802 ( .A1(n5440), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U5803 ( .A1(n5440), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U5804 ( .A1(n5440), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U5805 ( .A1(n5440), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5418) );
  NAND4_X1 U5806 ( .A1(n5407), .A2(n5406), .A3(n5405), .A4(n5404), .ZN(n8678)
         );
  NAND2_X1 U5807 ( .A1(n5440), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5404) );
  AOI21_X1 U5808 ( .B1(n9892), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9888), .ZN(
        n7183) );
  INV_X1 U5809 ( .A(n4699), .ZN(n7167) );
  INV_X1 U5810 ( .A(n4700), .ZN(n7141) );
  NOR2_X1 U5811 ( .A1(n7171), .A2(n7170), .ZN(n7322) );
  AND2_X1 U5812 ( .A1(n4699), .A2(n4698), .ZN(n7171) );
  NAND2_X1 U5813 ( .A1(n7168), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4698) );
  OR2_X1 U5814 ( .A1(n8689), .A2(n8688), .ZN(n8691) );
  AOI21_X1 U5815 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n8706), .A(n7326), .ZN(
        n7329) );
  NOR2_X1 U5816 ( .A1(n7329), .A2(n7328), .ZN(n7757) );
  NAND2_X1 U5817 ( .A1(n8714), .A2(n4690), .ZN(n7762) );
  OR2_X1 U5818 ( .A1(n8711), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4690) );
  NAND2_X1 U5819 ( .A1(n8736), .A2(n8737), .ZN(n8740) );
  INV_X1 U5820 ( .A(n4702), .ZN(n8745) );
  NAND2_X1 U5821 ( .A1(n4515), .A2(n8736), .ZN(n4702) );
  XNOR2_X1 U5822 ( .A(n4692), .B(n8778), .ZN(n8786) );
  AND2_X1 U5823 ( .A1(n7119), .A2(n7116), .ZN(n10238) );
  NOR2_X1 U5824 ( .A1(n4902), .A2(n8333), .ZN(n8895) );
  INV_X1 U5825 ( .A(n8914), .ZN(n4902) );
  NAND2_X1 U5826 ( .A1(n8945), .A2(n8436), .ZN(n8936) );
  CLKBUF_X1 U5827 ( .A(n8927), .Z(n8928) );
  NAND2_X1 U5828 ( .A1(n4960), .A2(n5045), .ZN(n8942) );
  NAND2_X1 U5829 ( .A1(n8245), .A2(n4964), .ZN(n4960) );
  OAI21_X1 U5830 ( .B1(n8068), .B2(n4502), .A(n4788), .ZN(n8242) );
  NAND2_X1 U5831 ( .A1(n4791), .A2(n8336), .ZN(n8120) );
  NAND2_X1 U5832 ( .A1(n8068), .A2(n5655), .ZN(n4791) );
  NAND2_X1 U5833 ( .A1(n7611), .A2(n4976), .ZN(n9918) );
  NAND2_X1 U5834 ( .A1(n5435), .A2(n5434), .ZN(n7458) );
  OR2_X1 U5835 ( .A1(n8261), .A2(n5429), .ZN(n5413) );
  NOR2_X1 U5836 ( .A1(n4729), .A2(n10315), .ZN(n4728) );
  NAND2_X1 U5837 ( .A1(n10272), .A2(n7353), .ZN(n10270) );
  NAND2_X1 U5838 ( .A1(n4727), .A2(n7218), .ZN(n7360) );
  INV_X1 U5839 ( .A(n4729), .ZN(n4727) );
  INV_X1 U5840 ( .A(n8956), .ZN(n10293) );
  OR2_X1 U5841 ( .A1(n5337), .A2(n6589), .ZN(n5356) );
  INV_X1 U5842 ( .A(n8795), .ZN(n8300) );
  NAND2_X1 U5843 ( .A1(n4911), .A2(n4910), .ZN(n4909) );
  AOI211_X1 U5844 ( .C1(n8986), .C2(n10368), .A(n8985), .B(n8984), .ZN(n9046)
         );
  NAND2_X1 U5845 ( .A1(n5476), .A2(n5475), .ZN(n8060) );
  INV_X1 U5846 ( .A(n7302), .ZN(n7465) );
  AND3_X2 U5847 ( .A1(n5338), .A2(n5339), .A3(n4574), .ZN(n7263) );
  NAND2_X1 U5848 ( .A1(n4575), .A2(n9879), .ZN(n4574) );
  AND2_X1 U5849 ( .A1(n6603), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10313) );
  NAND2_X1 U5850 ( .A1(n9066), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5088) );
  INV_X1 U5851 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5635) );
  INV_X1 U5852 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6992) );
  NAND2_X1 U5853 ( .A1(n6482), .A2(n6481), .ZN(n9759) );
  NAND2_X1 U5854 ( .A1(n8064), .A2(n9214), .ZN(n6482) );
  NAND2_X1 U5855 ( .A1(n6067), .A2(n6066), .ZN(n8131) );
  AND4_X1 U5856 ( .A1(n6196), .A2(n6195), .A3(n6194), .A4(n6193), .ZN(n9665)
         );
  NAND2_X1 U5857 ( .A1(n6536), .A2(n6535), .ZN(n6537) );
  NAND2_X1 U5858 ( .A1(n6495), .A2(n6494), .ZN(n6522) );
  INV_X1 U5859 ( .A(n7741), .ZN(n10202) );
  INV_X1 U5860 ( .A(n4844), .ZN(n9091) );
  AOI21_X1 U5861 ( .B1(n9149), .B2(n9147), .A(n4847), .ZN(n4844) );
  NAND2_X1 U5862 ( .A1(n7922), .A2(n6023), .ZN(n8044) );
  NAND2_X1 U5863 ( .A1(n9127), .A2(n6223), .ZN(n9098) );
  NAND2_X1 U5864 ( .A1(n7950), .A2(n9214), .ZN(n6225) );
  AND4_X1 U5865 ( .A1(n6089), .A2(n6088), .A3(n6087), .A4(n6086), .ZN(n9113)
         );
  NOR2_X1 U5866 ( .A1(n9110), .A2(n6119), .ZN(n9121) );
  NOR2_X1 U5867 ( .A1(n9121), .A2(n9120), .ZN(n9119) );
  NAND2_X1 U5868 ( .A1(n5785), .A2(n5784), .ZN(n9809) );
  AND2_X1 U5869 ( .A1(n4838), .A2(n4840), .ZN(n9129) );
  INV_X1 U5870 ( .A(n9075), .ZN(n4838) );
  AND4_X2 U5871 ( .A1(n7577), .A2(n7578), .A3(n7579), .A4(n7576), .ZN(n7679)
         );
  NAND2_X1 U5872 ( .A1(n6154), .A2(n6153), .ZN(n9796) );
  OR2_X1 U5873 ( .A1(n6315), .A2(n6314), .ZN(n9189) );
  OAI21_X1 U5874 ( .B1(n9149), .B2(n9148), .A(n9147), .ZN(n9146) );
  AND4_X1 U5875 ( .A1(n6178), .A2(n6177), .A3(n6176), .A4(n6175), .ZN(n9682)
         );
  INV_X1 U5876 ( .A(n9189), .ZN(n9181) );
  NAND2_X1 U5877 ( .A1(n6243), .A2(n6242), .ZN(n9764) );
  AND4_X1 U5878 ( .A1(n6108), .A2(n6107), .A3(n6106), .A4(n6105), .ZN(n9193)
         );
  INV_X1 U5879 ( .A(n9170), .ZN(n9194) );
  NAND2_X1 U5880 ( .A1(n9463), .A2(n5775), .ZN(n4680) );
  AND4_X1 U5881 ( .A1(n9467), .A2(n9466), .A3(n6282), .A4(n9465), .ZN(n9469)
         );
  NAND2_X1 U5882 ( .A1(n5829), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5830) );
  XNOR2_X1 U5883 ( .A(n5825), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10014) );
  OR2_X1 U5884 ( .A1(n9864), .A2(n6552), .ZN(n10021) );
  NAND2_X1 U5885 ( .A1(n10037), .A2(n4558), .ZN(n6729) );
  INV_X1 U5886 ( .A(n4710), .ZN(n6727) );
  NAND2_X1 U5887 ( .A1(n6701), .A2(n6702), .ZN(n6700) );
  AND2_X1 U5888 ( .A1(n4710), .A2(n4709), .ZN(n6701) );
  NAND2_X1 U5889 ( .A1(n6732), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4709) );
  AND2_X1 U5890 ( .A1(n4723), .A2(n4513), .ZN(n6560) );
  AND2_X1 U5891 ( .A1(n4723), .A2(n4721), .ZN(n6740) );
  AND2_X1 U5892 ( .A1(n6751), .A2(n6737), .ZN(n6739) );
  INV_X1 U5893 ( .A(n4705), .ZN(n10076) );
  AND2_X1 U5894 ( .A1(n4705), .A2(n4543), .ZN(n10089) );
  OR3_X1 U5895 ( .A1(n9988), .A2(n4481), .A3(n9995), .ZN(n10070) );
  NOR2_X1 U5896 ( .A1(n9523), .A2(n4571), .ZN(n9526) );
  NOR2_X1 U5897 ( .A1(n9521), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n4571) );
  XNOR2_X1 U5898 ( .A(n4707), .B(n4706), .ZN(n9531) );
  INV_X1 U5899 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n4706) );
  OR2_X1 U5900 ( .A1(n9520), .A2(n4708), .ZN(n4707) );
  AND2_X1 U5901 ( .A1(n9521), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4708) );
  INV_X1 U5902 ( .A(n9310), .ZN(n9545) );
  AND2_X1 U5903 ( .A1(n4887), .A2(n4886), .ZN(n9573) );
  NAND2_X1 U5904 ( .A1(n4996), .A2(n5002), .ZN(n9566) );
  NAND2_X1 U5905 ( .A1(n9597), .A2(n4507), .ZN(n4996) );
  NOR2_X1 U5906 ( .A1(n9614), .A2(n9409), .ZN(n9588) );
  INV_X1 U5907 ( .A(n9764), .ZN(n9586) );
  AOI21_X1 U5908 ( .B1(n9597), .B2(n9605), .A(n5001), .ZN(n9581) );
  INV_X1 U5909 ( .A(n5004), .ZN(n5001) );
  AND2_X1 U5910 ( .A1(n6187), .A2(n6186), .ZN(n9655) );
  NAND2_X1 U5911 ( .A1(n5021), .A2(n5022), .ZN(n8132) );
  OR2_X1 U5912 ( .A1(n7989), .A2(n5024), .ZN(n5021) );
  NAND2_X1 U5913 ( .A1(n4880), .A2(n9370), .ZN(n7993) );
  NAND2_X1 U5914 ( .A1(n5995), .A2(n5994), .ZN(n7908) );
  INV_X1 U5915 ( .A(n9218), .ZN(n9219) );
  NAND2_X1 U5916 ( .A1(n7586), .A2(n5036), .ZN(n10180) );
  NAND2_X1 U5917 ( .A1(n7586), .A2(n7585), .ZN(n7706) );
  NAND2_X1 U5918 ( .A1(n6545), .A2(n4751), .ZN(n4750) );
  OAI21_X1 U5919 ( .B1(n6593), .B2(n4635), .A(n4752), .ZN(n4751) );
  INV_X1 U5920 ( .A(n9951), .ZN(n9660) );
  AND2_X1 U5921 ( .A1(n4748), .A2(n4747), .ZN(n9979) );
  AOI21_X1 U5922 ( .B1(n9310), .B2(n9964), .A(n9963), .ZN(n4747) );
  OR2_X1 U5923 ( .A1(n9962), .A2(n10210), .ZN(n4748) );
  INV_X1 U5924 ( .A(n4679), .ZN(n5759) );
  XNOR2_X1 U5925 ( .A(n8289), .B(n8288), .ZN(n9853) );
  NAND2_X1 U5926 ( .A1(n8286), .A2(n8285), .ZN(n8289) );
  XNOR2_X1 U5927 ( .A(n8189), .B(n8188), .ZN(n8220) );
  INV_X1 U5928 ( .A(n6266), .ZN(n7829) );
  XNOR2_X1 U5929 ( .A(n5546), .B(n5545), .ZN(n7779) );
  XNOR2_X1 U5930 ( .A(n5428), .B(n5427), .ZN(n6599) );
  NAND2_X1 U5931 ( .A1(n4871), .A2(n5122), .ZN(n5428) );
  NAND2_X1 U5932 ( .A1(n5409), .A2(n5408), .ZN(n4871) );
  AND2_X1 U5933 ( .A1(n4526), .A2(n4636), .ZN(n5396) );
  NAND2_X1 U5934 ( .A1(n4634), .A2(n5796), .ZN(n5798) );
  NOR2_X1 U5935 ( .A1(n8107), .A2(n10420), .ZN(n10409) );
  NAND2_X1 U5936 ( .A1(n4919), .A2(n4920), .ZN(n7408) );
  AND2_X1 U5937 ( .A1(n4592), .A2(n4595), .ZN(n6634) );
  AOI21_X1 U5938 ( .B1(n4792), .B2(n8522), .A(n4580), .ZN(n8531) );
  OAI21_X1 U5939 ( .B1(n9032), .B2(n10380), .A(n4730), .ZN(n8308) );
  AND2_X1 U5940 ( .A1(n5713), .A2(n4586), .ZN(n4585) );
  NAND2_X1 U5941 ( .A1(n10380), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n4586) );
  NAND2_X1 U5942 ( .A1(n8859), .A2(n5712), .ZN(n4578) );
  AND2_X1 U5943 ( .A1(n5717), .A2(n4588), .ZN(n4587) );
  NAND2_X1 U5944 ( .A1(n10370), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n4588) );
  NAND2_X1 U5945 ( .A1(n8859), .A2(n5716), .ZN(n4577) );
  OAI211_X1 U5946 ( .C1(n9753), .C2(n5008), .A(n5013), .B(n5007), .ZN(P1_U3552) );
  NAND2_X1 U5947 ( .A1(n10236), .A2(n10199), .ZN(n5008) );
  AND2_X1 U5948 ( .A1(n7701), .A2(n10172), .ZN(n4492) );
  NAND2_X1 U5949 ( .A1(n8408), .A2(n9909), .ZN(n8410) );
  NAND2_X1 U5950 ( .A1(n5262), .A2(n5261), .ZN(n9917) );
  AND2_X1 U5951 ( .A1(n5880), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4493) );
  INV_X1 U5952 ( .A(n4722), .ZN(n4721) );
  NAND2_X1 U5953 ( .A1(n6559), .A2(n4513), .ZN(n4722) );
  AND2_X1 U5954 ( .A1(n5022), .A2(n4525), .ZN(n4494) );
  OR2_X1 U5955 ( .A1(n9275), .A2(n4673), .ZN(n4495) );
  INV_X1 U5956 ( .A(n9244), .ZN(n4875) );
  AND2_X1 U5957 ( .A1(n8433), .A2(n8432), .ZN(n4496) );
  NAND2_X1 U5958 ( .A1(n5570), .A2(n5569), .ZN(n8980) );
  AND2_X1 U5959 ( .A1(n4514), .A2(n5726), .ZN(n4497) );
  OR2_X1 U5960 ( .A1(n8980), .A2(n8648), .ZN(n8849) );
  INV_X1 U5961 ( .A(n8849), .ZN(n4818) );
  NAND2_X1 U5962 ( .A1(n9273), .A2(n9269), .ZN(n4498) );
  NOR2_X1 U5963 ( .A1(n9917), .A2(n8671), .ZN(n4499) );
  AND2_X1 U5964 ( .A1(n8944), .A2(n4961), .ZN(n4500) );
  INV_X1 U5965 ( .A(n5648), .ZN(n5649) );
  NAND2_X1 U5966 ( .A1(n8331), .A2(n5672), .ZN(n8465) );
  INV_X2 U5967 ( .A(n8539), .ZN(n9776) );
  AND2_X1 U5968 ( .A1(n6207), .A2(n6206), .ZN(n8539) );
  INV_X1 U5969 ( .A(n8944), .ZN(n4907) );
  AND4_X1 U5970 ( .A1(n6505), .A2(n6504), .A3(n6503), .A4(n6502), .ZN(n9572)
         );
  NAND2_X1 U5971 ( .A1(n5963), .A2(n5962), .ZN(n7814) );
  OR2_X1 U5972 ( .A1(n8738), .A2(n8747), .ZN(n4501) );
  BUF_X1 U5973 ( .A(n5340), .Z(n7126) );
  INV_X2 U5974 ( .A(n5340), .ZN(n4575) );
  OR2_X1 U5975 ( .A1(n8425), .A2(n4790), .ZN(n4502) );
  NAND2_X2 U5976 ( .A1(n4488), .A2(n4635), .ZN(n5822) );
  NOR2_X1 U5977 ( .A1(n8118), .A2(n8425), .ZN(n4503) );
  OR2_X1 U5978 ( .A1(n5637), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n4504) );
  NAND4_X1 U5979 ( .A1(n5361), .A2(n5360), .A3(n5359), .A4(n5358), .ZN(n8681)
         );
  NAND2_X1 U5980 ( .A1(n5123), .A2(SI_7_), .ZN(n4505) );
  NAND2_X2 U5981 ( .A1(n5095), .A2(n5094), .ZN(n5553) );
  OR2_X1 U5982 ( .A1(n6278), .A2(n5751), .ZN(n4506) );
  AND2_X1 U5983 ( .A1(n5005), .A2(n9605), .ZN(n4507) );
  AND3_X1 U5984 ( .A1(n5388), .A2(n5387), .A3(n5386), .ZN(n4508) );
  INV_X4 U5985 ( .A(n5385), .ZN(n5326) );
  NAND2_X1 U5986 ( .A1(n4489), .A2(n4483), .ZN(n5823) );
  AND2_X1 U5987 ( .A1(n5139), .A2(SI_11_), .ZN(n4509) );
  NOR2_X1 U5988 ( .A1(n8559), .A2(n10220), .ZN(n4510) );
  INV_X1 U5989 ( .A(n4863), .ZN(n4862) );
  OAI21_X1 U5990 ( .B1(n9120), .B2(n6118), .A(n4537), .ZN(n4863) );
  AND2_X1 U5991 ( .A1(n5799), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n4511) );
  XOR2_X1 U5992 ( .A(n8323), .B(n8796), .Z(n4512) );
  NAND2_X1 U5993 ( .A1(n5492), .A2(n5491), .ZN(n9020) );
  INV_X1 U5994 ( .A(n5770), .ZN(n7625) );
  AND2_X1 U5995 ( .A1(n8849), .A2(n8452), .ZN(n8875) );
  INV_X1 U5996 ( .A(n8875), .ZN(n8863) );
  NAND2_X1 U5997 ( .A1(n10049), .A2(n7726), .ZN(n4513) );
  AND2_X1 U5998 ( .A1(n4624), .A2(n5052), .ZN(n4623) );
  NAND2_X1 U5999 ( .A1(n5457), .A2(n5456), .ZN(n7425) );
  AND3_X1 U6000 ( .A1(n5728), .A2(n5727), .A3(n5729), .ZN(n4514) );
  AND2_X1 U6001 ( .A1(n8737), .A2(n4703), .ZN(n4515) );
  NAND2_X1 U6002 ( .A1(n9418), .A2(n9455), .ZN(n9364) );
  INV_X1 U6003 ( .A(n9364), .ZN(n4896) );
  INV_X1 U6004 ( .A(n9409), .ZN(n4890) );
  INV_X1 U6005 ( .A(n9417), .ZN(n4891) );
  OR2_X1 U6006 ( .A1(n8920), .A2(n8596), .ZN(n8438) );
  OR3_X1 U6007 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n4516) );
  OR3_X1 U6008 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        n4579), .ZN(n4517) );
  OR2_X1 U6009 ( .A1(n7665), .A2(n9487), .ZN(n4518) );
  NAND2_X1 U6010 ( .A1(n6390), .A2(n6391), .ZN(n4519) );
  AND2_X1 U6011 ( .A1(n9425), .A2(n4657), .ZN(n4520) );
  AND2_X1 U6012 ( .A1(n9400), .A2(n9318), .ZN(n4521) );
  INV_X1 U6013 ( .A(n4483), .ZN(n4635) );
  OR2_X1 U6014 ( .A1(n9759), .A2(n9592), .ZN(n4522) );
  OR2_X1 U6015 ( .A1(n8950), .A2(n8595), .ZN(n8436) );
  INV_X1 U6016 ( .A(n8436), .ZN(n4908) );
  NAND2_X1 U6017 ( .A1(n5992), .A2(n5723), .ZN(n6024) );
  NAND2_X1 U6018 ( .A1(n5042), .A2(n5824), .ZN(n5857) );
  AND2_X1 U6019 ( .A1(n8802), .A2(n8461), .ZN(n4523) );
  AND2_X1 U6020 ( .A1(n4903), .A2(n5656), .ZN(n4524) );
  NAND2_X1 U6021 ( .A1(n6126), .A2(n6125), .ZN(n9804) );
  AND2_X1 U6022 ( .A1(n6082), .A2(n6081), .ZN(n9820) );
  INV_X1 U6023 ( .A(n9820), .ZN(n9204) );
  OR2_X1 U6024 ( .A1(n9759), .A2(n8541), .ZN(n9416) );
  OR2_X1 U6025 ( .A1(n8887), .A2(n8605), .ZN(n5656) );
  NAND2_X1 U6026 ( .A1(n8131), .A2(n9481), .ZN(n4525) );
  INV_X1 U6027 ( .A(n9879), .ZN(n7122) );
  AND3_X1 U6028 ( .A1(n5333), .A2(n4694), .A3(n4693), .ZN(n9879) );
  INV_X1 U6029 ( .A(n4857), .ZN(n4856) );
  NOR2_X1 U6030 ( .A1(n6061), .A2(n4858), .ZN(n4857) );
  OR2_X1 U6031 ( .A1(n5116), .A2(n5375), .ZN(n4526) );
  INV_X1 U6032 ( .A(n4977), .ZN(n4976) );
  OR2_X1 U6033 ( .A1(n8827), .A2(n8461), .ZN(n8312) );
  AND2_X1 U6034 ( .A1(n8427), .A2(n8426), .ZN(n4527) );
  INV_X1 U6035 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9065) );
  AND2_X1 U6036 ( .A1(n4496), .A2(n8430), .ZN(n4528) );
  AND2_X1 U6037 ( .A1(n9786), .A2(n9665), .ZN(n9328) );
  NOR2_X1 U6038 ( .A1(n5051), .A2(n6060), .ZN(n4529) );
  INV_X1 U6039 ( .A(n4764), .ZN(n9567) );
  NOR2_X1 U6040 ( .A1(n9619), .A2(n4765), .ZN(n4764) );
  INV_X1 U6041 ( .A(n5227), .ZN(n4980) );
  AOI21_X1 U6042 ( .B1(n9149), .B2(n4845), .A(n4842), .ZN(n4841) );
  INV_X1 U6043 ( .A(n6337), .ZN(n4595) );
  AND2_X1 U6044 ( .A1(n6336), .A2(n6335), .ZN(n6337) );
  INV_X1 U6045 ( .A(n4943), .ZN(n4942) );
  AND2_X1 U6046 ( .A1(n4519), .A2(n8571), .ZN(n4943) );
  INV_X1 U6047 ( .A(n5000), .ZN(n4999) );
  NAND2_X1 U6048 ( .A1(n9575), .A2(n4507), .ZN(n5000) );
  OR2_X1 U6049 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n4530) );
  NOR2_X1 U6050 ( .A1(n5056), .A2(n8006), .ZN(n4531) );
  AND2_X1 U6051 ( .A1(n8417), .A2(n8482), .ZN(n4532) );
  INV_X1 U6052 ( .A(n7992), .ZN(n4874) );
  NOR2_X1 U6053 ( .A1(n8131), .A2(n9481), .ZN(n4533) );
  NAND2_X1 U6054 ( .A1(n8386), .A2(n8385), .ZN(n8380) );
  INV_X1 U6055 ( .A(n4733), .ZN(n4732) );
  NAND2_X1 U6056 ( .A1(n8445), .A2(n4734), .ZN(n4733) );
  INV_X1 U6057 ( .A(n4738), .ZN(n4737) );
  NAND2_X1 U6058 ( .A1(n4740), .A2(n4739), .ZN(n4738) );
  OR2_X1 U6059 ( .A1(n4633), .A2(n4629), .ZN(n4534) );
  OR2_X1 U6060 ( .A1(n7878), .A2(n7880), .ZN(n4536) );
  NAND2_X1 U6061 ( .A1(n6121), .A2(n6122), .ZN(n4537) );
  NAND2_X1 U6062 ( .A1(n6097), .A2(n6093), .ZN(n4538) );
  AND2_X1 U6063 ( .A1(n6371), .A2(n4933), .ZN(n4539) );
  AND2_X1 U6064 ( .A1(n8435), .A2(n8436), .ZN(n4540) );
  AND2_X1 U6065 ( .A1(n4997), .A2(n4522), .ZN(n4541) );
  INV_X1 U6066 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5731) );
  OR2_X1 U6067 ( .A1(n9749), .A2(n9475), .ZN(n4542) );
  OR2_X1 U6068 ( .A1(n9510), .A2(n9509), .ZN(n4543) );
  AND3_X1 U6069 ( .A1(n5739), .A2(n5781), .A3(n6940), .ZN(n4544) );
  AND3_X1 U6070 ( .A1(n4670), .A2(n9267), .A3(n4669), .ZN(n4545) );
  INV_X1 U6071 ( .A(n6094), .ZN(n4853) );
  AND2_X1 U6072 ( .A1(n4731), .A2(n9044), .ZN(n4546) );
  NOR2_X1 U6073 ( .A1(n4823), .A2(n8443), .ZN(n4547) );
  AND2_X1 U6074 ( .A1(n8588), .A2(n8676), .ZN(n4548) );
  INV_X1 U6075 ( .A(n9439), .ZN(n4656) );
  AND2_X1 U6076 ( .A1(n8415), .A2(n8416), .ZN(n8414) );
  NOR2_X1 U6077 ( .A1(n10261), .A2(n4783), .ZN(n4782) );
  AND2_X1 U6078 ( .A1(n10018), .A2(n4713), .ZN(n4549) );
  NAND2_X1 U6079 ( .A1(n4921), .A2(n4924), .ZN(n4920) );
  NAND2_X1 U6080 ( .A1(n4626), .A2(n4625), .ZN(n4550) );
  AND2_X1 U6081 ( .A1(n5732), .A2(n5722), .ZN(n4551) );
  NAND2_X1 U6082 ( .A1(n4594), .A2(n4593), .ZN(n4552) );
  AND2_X1 U6083 ( .A1(n4901), .A2(n4899), .ZN(n4553) );
  NAND2_X1 U6084 ( .A1(n5209), .A2(n5208), .ZN(n8887) );
  INV_X1 U6085 ( .A(n8887), .ZN(n4734) );
  NAND2_X1 U6086 ( .A1(n6282), .A2(n9670), .ZN(n9318) );
  INV_X1 U6087 ( .A(n9318), .ZN(n4673) );
  NAND2_X1 U6088 ( .A1(n5621), .A2(n5620), .ZN(n8827) );
  INV_X1 U6089 ( .A(n5040), .ZN(n5039) );
  NAND2_X1 U6090 ( .A1(n6139), .A2(n6138), .ZN(n9800) );
  NAND2_X1 U6091 ( .A1(n4980), .A2(n5220), .ZN(n5229) );
  XNOR2_X1 U6092 ( .A(n8970), .B(n8650), .ZN(n8510) );
  AND4_X1 U6093 ( .A1(n6016), .A2(n6015), .A3(n6014), .A4(n6013), .ZN(n8049)
         );
  INV_X1 U6094 ( .A(n8049), .ZN(n5030) );
  AND3_X1 U6095 ( .A1(n6380), .A2(n6381), .A3(n4600), .ZN(n4554) );
  NAND2_X1 U6096 ( .A1(n7924), .A2(n7923), .ZN(n7922) );
  NAND2_X1 U6097 ( .A1(n6225), .A2(n6224), .ZN(n9769) );
  INV_X1 U6098 ( .A(n9769), .ZN(n9602) );
  OR2_X1 U6099 ( .A1(n9688), .A2(n9664), .ZN(n4555) );
  INV_X1 U6100 ( .A(n4754), .ZN(n9684) );
  NOR2_X1 U6101 ( .A1(n9692), .A2(n9796), .ZN(n4754) );
  NAND2_X1 U6102 ( .A1(n8898), .A2(n4732), .ZN(n4735) );
  NAND2_X1 U6103 ( .A1(n8123), .A2(n4737), .ZN(n4741) );
  AND2_X1 U6104 ( .A1(n4702), .A2(n8738), .ZN(n4556) );
  NAND2_X1 U6105 ( .A1(n8141), .A2(n4757), .ZN(n4760) );
  NAND2_X1 U6106 ( .A1(n4599), .A2(n4597), .ZN(n4557) );
  OR2_X1 U6107 ( .A1(n6563), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4558) );
  INV_X1 U6108 ( .A(n9370), .ZN(n4876) );
  NAND2_X1 U6109 ( .A1(n8241), .A2(n8432), .ZN(n8943) );
  INV_X1 U6110 ( .A(n8943), .ZN(n4906) );
  OR2_X1 U6111 ( .A1(n8980), .A2(n8661), .ZN(n4559) );
  AND2_X1 U6112 ( .A1(n7143), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4560) );
  AND2_X1 U6113 ( .A1(n7611), .A2(n4974), .ZN(n4561) );
  INV_X1 U6114 ( .A(n5513), .ZN(n4963) );
  NAND2_X1 U6115 ( .A1(n5504), .A2(n5503), .ZN(n8950) );
  INV_X1 U6116 ( .A(n8950), .ZN(n4739) );
  NAND2_X1 U6117 ( .A1(n7308), .A2(n7307), .ZN(n4562) );
  NAND2_X1 U6118 ( .A1(n6171), .A2(n6170), .ZN(n9791) );
  INV_X1 U6119 ( .A(n9791), .ZN(n4753) );
  NAND2_X1 U6120 ( .A1(n5963), .A2(n4859), .ZN(n7815) );
  AND2_X1 U6121 ( .A1(n4927), .A2(n4926), .ZN(n4563) );
  NAND2_X1 U6122 ( .A1(n7744), .A2(n9233), .ZN(n7910) );
  INV_X1 U6123 ( .A(n7910), .ZN(n4881) );
  INV_X1 U6124 ( .A(n4746), .ZN(n7615) );
  NOR2_X1 U6125 ( .A1(n7421), .A2(n4744), .ZN(n4746) );
  INV_X1 U6126 ( .A(n8859), .ZN(n9044) );
  NAND2_X1 U6127 ( .A1(n5587), .A2(n5586), .ZN(n8859) );
  AND2_X2 U6128 ( .A1(n5711), .A2(n8479), .ZN(n9922) );
  INV_X1 U6129 ( .A(n6322), .ZN(n5711) );
  NOR2_X1 U6130 ( .A1(n7271), .A2(n4480), .ZN(n4729) );
  AND2_X1 U6131 ( .A1(n7998), .A2(n10155), .ZN(n10192) );
  AND2_X1 U6132 ( .A1(n5801), .A2(n5800), .ZN(n7203) );
  OR2_X1 U6133 ( .A1(n6370), .A2(n6369), .ZN(n4564) );
  INV_X1 U6134 ( .A(n7842), .ZN(n4762) );
  AND2_X1 U6135 ( .A1(n5821), .A2(n7394), .ZN(n9165) );
  INV_X1 U6136 ( .A(n8747), .ZN(n4704) );
  AND2_X1 U6137 ( .A1(n9513), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4565) );
  AND2_X1 U6138 ( .A1(n4955), .A2(n6343), .ZN(n4566) );
  AND2_X1 U6139 ( .A1(n4483), .A2(P1_U3084), .ZN(n4567) );
  AND2_X1 U6140 ( .A1(n4483), .A2(P2_U3152), .ZN(n4568) );
  INV_X1 U6141 ( .A(n9532), .ZN(n9670) );
  INV_X1 U6142 ( .A(n10018), .ZN(n4712) );
  OR2_X1 U6143 ( .A1(n8481), .A2(n5711), .ZN(n4569) );
  INV_X1 U6144 ( .A(n6552), .ZN(n4713) );
  NAND2_X1 U6145 ( .A1(n7520), .A2(n8497), .ZN(n7519) );
  AOI21_X1 U6146 ( .B1(n7210), .B2(n5394), .A(n5393), .ZN(n7282) );
  NAND2_X1 U6147 ( .A1(n7238), .A2(n5350), .ZN(n7269) );
  OAI22_X1 U6148 ( .A1(n8245), .A2(n4959), .B1(n4500), .B2(n5513), .ZN(n8927)
         );
  NOR2_X1 U6149 ( .A1(n7980), .A2(n4979), .ZN(n8072) );
  AOI21_X2 U6150 ( .B1(n7459), .B2(n8380), .A(n5446), .ZN(n10248) );
  NAND2_X2 U6151 ( .A1(n8989), .A2(n5048), .ZN(n8880) );
  OAI21_X1 U6152 ( .B1(n9497), .B2(n9496), .A(n10094), .ZN(n10112) );
  NAND2_X1 U6153 ( .A1(n4572), .A2(n6570), .ZN(n9870) );
  NAND2_X1 U6154 ( .A1(n10006), .A2(n6569), .ZN(n4572) );
  NOR2_X1 U6155 ( .A1(n10022), .A2(n6571), .ZN(n10043) );
  NOR2_X1 U6156 ( .A1(n6574), .A2(n6703), .ZN(n10056) );
  NAND2_X1 U6157 ( .A1(n10081), .A2(n9495), .ZN(n10096) );
  NOR2_X1 U6158 ( .A1(n6735), .A2(n6734), .ZN(n6754) );
  NAND2_X1 U6159 ( .A1(n4981), .A2(n4777), .ZN(n5090) );
  AOI21_X1 U6160 ( .B1(n8259), .B2(n10227), .A(n6722), .ZN(n6705) );
  AOI21_X1 U6161 ( .B1(n9505), .B2(n9970), .A(n9493), .ZN(n9494) );
  AOI21_X1 U6162 ( .B1(n6010), .B2(n7248), .A(n7247), .ZN(n7250) );
  AOI21_X1 U6163 ( .B1(n6028), .B2(n7784), .A(n7783), .ZN(n10069) );
  AOI21_X1 U6164 ( .B1(n7786), .B2(n7785), .A(n10067), .ZN(n7788) );
  NAND2_X1 U6165 ( .A1(n4573), .A2(n6459), .ZN(P2_U3222) );
  NAND3_X1 U6166 ( .A1(n6446), .A2(n6447), .A3(n6445), .ZN(n4573) );
  NAND2_X1 U6167 ( .A1(n6414), .A2(n6413), .ZN(n8601) );
  INV_X1 U6168 ( .A(n8644), .ZN(n6443) );
  OR2_X1 U6169 ( .A1(n8880), .A2(n8881), .ZN(n4991) );
  NAND2_X1 U6170 ( .A1(n9043), .A2(n4577), .ZN(P2_U3514) );
  NAND2_X1 U6171 ( .A1(n8977), .A2(n4578), .ZN(P2_U3546) );
  NOR2_X2 U6172 ( .A1(n7474), .A2(n8499), .ZN(n7473) );
  NAND2_X1 U6173 ( .A1(n8072), .A2(n8504), .ZN(n8071) );
  NAND2_X1 U6174 ( .A1(n4796), .A2(n4797), .ZN(n5150) );
  NAND2_X1 U6175 ( .A1(n4795), .A2(n4794), .ZN(n4793) );
  NOR2_X1 U6176 ( .A1(n8850), .A2(n5657), .ZN(n8834) );
  NAND3_X2 U6177 ( .A1(n4581), .A2(n5831), .A3(n5830), .ZN(n9490) );
  NOR2_X2 U6178 ( .A1(n4493), .A2(n4510), .ZN(n4581) );
  INV_X2 U6179 ( .A(n6301), .ZN(n5829) );
  NAND2_X2 U6180 ( .A1(n5763), .A2(n5765), .ZN(n6301) );
  NAND2_X1 U6181 ( .A1(n4884), .A2(n4882), .ZN(n9560) );
  INV_X1 U6182 ( .A(n6522), .ZN(n6539) );
  OR2_X2 U6183 ( .A1(n7924), .A2(n4856), .ZN(n4850) );
  AOI21_X2 U6184 ( .B1(n8025), .B2(n6097), .A(n6096), .ZN(n9195) );
  NAND2_X1 U6185 ( .A1(n5744), .A2(n4497), .ZN(n6278) );
  INV_X1 U6186 ( .A(n4841), .ZN(n6201) );
  NAND2_X1 U6187 ( .A1(n5528), .A2(n5184), .ZN(n5544) );
  AOI21_X1 U6188 ( .B1(n4799), .B2(n4802), .A(n4798), .ZN(n4797) );
  NAND2_X1 U6189 ( .A1(n5200), .A2(n5199), .ZN(n5564) );
  OAI21_X1 U6190 ( .B1(n5470), .B2(n5469), .A(n5159), .ZN(n5239) );
  NAND2_X1 U6191 ( .A1(n4685), .A2(n9670), .ZN(n4684) );
  NAND2_X1 U6192 ( .A1(n4682), .A2(n7588), .ZN(n4681) );
  NAND2_X1 U6193 ( .A1(n4681), .A2(n4680), .ZN(n9470) );
  INV_X1 U6194 ( .A(n4806), .ZN(n4804) );
  OAI21_X1 U6195 ( .B1(n5715), .B2(n10380), .A(n4585), .ZN(P2_U3548) );
  OAI21_X1 U6196 ( .B1(n5715), .B2(n10370), .A(n4587), .ZN(P2_U3516) );
  NAND2_X1 U6197 ( .A1(n4968), .A2(n5615), .ZN(n8801) );
  NAND2_X1 U6198 ( .A1(n4779), .A2(n4780), .ZN(n7378) );
  NAND2_X1 U6199 ( .A1(n8326), .A2(n8513), .ZN(n4795) );
  NAND2_X1 U6200 ( .A1(n7608), .A2(n5652), .ZN(n9908) );
  INV_X1 U6201 ( .A(n6633), .ZN(n4591) );
  NAND3_X1 U6202 ( .A1(n4590), .A2(n4589), .A3(n4552), .ZN(n6685) );
  NAND3_X1 U6203 ( .A1(n4591), .A2(n6645), .A3(n6646), .ZN(n4590) );
  NAND3_X1 U6204 ( .A1(n6380), .A2(n6381), .A3(n4598), .ZN(n4597) );
  NAND2_X1 U6205 ( .A1(n6380), .A2(n6381), .ZN(n8054) );
  INV_X1 U6206 ( .A(n8055), .ZN(n4600) );
  INV_X1 U6207 ( .A(n4926), .ZN(n4602) );
  AND2_X2 U6208 ( .A1(n8524), .A2(n6324), .ZN(n6329) );
  NAND3_X1 U6209 ( .A1(n4958), .A2(n4957), .A3(n6464), .ZN(n8645) );
  NAND2_X1 U6210 ( .A1(n7308), .A2(n6350), .ZN(n4610) );
  NAND2_X1 U6211 ( .A1(n4916), .A2(n4609), .ZN(n7406) );
  NAND3_X1 U6212 ( .A1(n4920), .A2(n6354), .A3(n4610), .ZN(n4609) );
  NAND3_X1 U6213 ( .A1(n4619), .A2(n4614), .A3(n5314), .ZN(n4613) );
  NAND2_X1 U6214 ( .A1(n5314), .A2(n5128), .ZN(n4618) );
  OR2_X1 U6215 ( .A1(n5314), .A2(n5312), .ZN(n4622) );
  NAND3_X1 U6216 ( .A1(n4615), .A2(n4613), .A3(n4611), .ZN(n6614) );
  NAND3_X1 U6217 ( .A1(n4612), .A2(n4623), .A3(n5451), .ZN(n4611) );
  OR2_X1 U6218 ( .A1(n8431), .A2(n4627), .ZN(n4626) );
  NAND2_X2 U6219 ( .A1(n4820), .A2(n4819), .ZN(n5112) );
  NAND3_X1 U6220 ( .A1(n4819), .A2(n4820), .A3(n5103), .ZN(n5348) );
  NAND2_X1 U6221 ( .A1(n4635), .A2(SI_0_), .ZN(n5347) );
  NAND2_X1 U6222 ( .A1(n4635), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4752) );
  NAND2_X1 U6223 ( .A1(n4483), .A2(SI_0_), .ZN(n4634) );
  MUX2_X1 U6224 ( .A(n9071), .B(n9858), .S(n4483), .Z(n8282) );
  MUX2_X1 U6225 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4483), .Z(n8287) );
  AND2_X1 U6226 ( .A1(P2_U3152), .A2(n4635), .ZN(n8114) );
  NAND2_X1 U6227 ( .A1(P1_U3084), .A2(n4635), .ZN(n8257) );
  NAND2_X1 U6228 ( .A1(n5340), .A2(n4635), .ZN(n5337) );
  NAND2_X1 U6229 ( .A1(n5370), .A2(n5369), .ZN(n5374) );
  NAND3_X1 U6230 ( .A1(n4526), .A2(n5395), .A3(n4636), .ZN(n4809) );
  NAND2_X1 U6231 ( .A1(n4868), .A2(SI_3_), .ZN(n5373) );
  AOI21_X1 U6232 ( .B1(n7425), .B2(n8340), .A(n8465), .ZN(n4647) );
  NAND2_X1 U6233 ( .A1(n4646), .A2(n4650), .ZN(n4649) );
  NAND2_X1 U6234 ( .A1(n4647), .A2(n4648), .ZN(n4646) );
  OR2_X1 U6235 ( .A1(n7425), .A2(n7500), .ZN(n8341) );
  NAND2_X1 U6236 ( .A1(n4653), .A2(n4652), .ZN(n7595) );
  AOI21_X1 U6237 ( .B1(n7803), .B2(n9439), .A(n7659), .ZN(n4653) );
  NAND2_X1 U6238 ( .A1(n4655), .A2(n9439), .ZN(n7845) );
  NAND4_X1 U6239 ( .A1(n4659), .A2(n4660), .A3(n7600), .A4(n5795), .ZN(n7630)
         );
  AND2_X1 U6240 ( .A1(n4661), .A2(n5794), .ZN(n4659) );
  OR2_X1 U6241 ( .A1(n8559), .A2(n9991), .ZN(n4661) );
  NAND2_X1 U6242 ( .A1(n9268), .A2(n4545), .ZN(n4664) );
  AND2_X1 U6243 ( .A1(n5967), .A2(n4551), .ZN(n4677) );
  AND2_X2 U6244 ( .A1(n5967), .A2(n5722), .ZN(n5991) );
  NAND3_X1 U6245 ( .A1(n4677), .A2(n5040), .A3(n4676), .ZN(n4675) );
  OR2_X2 U6246 ( .A1(n9324), .A2(n9323), .ZN(n9467) );
  NAND3_X1 U6247 ( .A1(n4688), .A2(n9286), .A3(n4687), .ZN(n4686) );
  XNOR2_X2 U6248 ( .A(n8768), .B(n8769), .ZN(n8770) );
  NAND2_X1 U6249 ( .A1(n4701), .A2(n4501), .ZN(n8766) );
  NAND3_X1 U6250 ( .A1(n4515), .A2(n8736), .A3(n4704), .ZN(n4701) );
  NAND2_X1 U6251 ( .A1(n4711), .A2(n4549), .ZN(n10019) );
  INV_X1 U6252 ( .A(n4711), .ZN(n9864) );
  AOI21_X1 U6253 ( .B1(n10052), .B2(n4719), .A(n4717), .ZN(n6756) );
  OAI21_X1 U6254 ( .B1(n10052), .B2(n4722), .A(n4719), .ZN(n4724) );
  INV_X1 U6255 ( .A(n4724), .ZN(n6758) );
  OAI211_X2 U6256 ( .C1(n7126), .C2(n6585), .A(n5355), .B(n5356), .ZN(n7493)
         );
  NOR2_X1 U6257 ( .A1(n8270), .A2(n4728), .ZN(n10314) );
  NAND2_X1 U6258 ( .A1(n10380), .A2(n8307), .ZN(n4730) );
  INV_X1 U6259 ( .A(n4735), .ZN(n8886) );
  INV_X1 U6260 ( .A(n4741), .ZN(n8948) );
  NAND2_X1 U6261 ( .A1(n9544), .A2(n9545), .ZN(n9543) );
  OAI21_X2 U6262 ( .B1(n6545), .B2(n6721), .A(n4750), .ZN(n7641) );
  INV_X1 U6263 ( .A(n4760), .ZN(n9727) );
  NAND2_X1 U6264 ( .A1(n7669), .A2(n7713), .ZN(n7727) );
  INV_X1 U6265 ( .A(n4763), .ZN(n9552) );
  OAI22_X1 U6266 ( .A1(n7415), .A2(n4773), .B1(n5649), .B2(n4774), .ZN(n7608)
         );
  NAND2_X1 U6267 ( .A1(n7378), .A2(n8340), .ZN(n7414) );
  NAND2_X1 U6268 ( .A1(n4782), .A2(n7448), .ZN(n4779) );
  NAND2_X1 U6269 ( .A1(n8068), .A2(n4788), .ZN(n4785) );
  NAND2_X1 U6270 ( .A1(n4785), .A2(n4786), .ZN(n8241) );
  NAND2_X1 U6271 ( .A1(n5448), .A2(n4799), .ZN(n4796) );
  OAI21_X1 U6272 ( .B1(n5448), .B2(n4802), .A(n4799), .ZN(n5263) );
  NAND2_X1 U6273 ( .A1(n4505), .A2(n5119), .ZN(n4808) );
  INV_X1 U6274 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4822) );
  NAND3_X1 U6275 ( .A1(n4550), .A2(n4826), .A3(n4825), .ZN(n4824) );
  NAND2_X1 U6276 ( .A1(n7620), .A2(n8297), .ZN(n4830) );
  NAND2_X1 U6277 ( .A1(n4830), .A2(n5515), .ZN(n9002) );
  NAND2_X1 U6278 ( .A1(n5166), .A2(n5165), .ZN(n5484) );
  INV_X1 U6279 ( .A(n5528), .ZN(n5514) );
  NAND2_X1 U6280 ( .A1(n8837), .A2(n8842), .ZN(n5671) );
  NAND2_X1 U6281 ( .A1(n5150), .A2(n5149), .ZN(n5257) );
  OAI21_X1 U6282 ( .B1(n9753), .B2(n10192), .A(n5014), .ZN(n9832) );
  AOI21_X1 U6283 ( .B1(n9075), .B2(n6223), .A(n4836), .ZN(n4835) );
  OAI21_X1 U6284 ( .B1(n9149), .B2(n4847), .A(n4845), .ZN(n9090) );
  NAND2_X1 U6285 ( .A1(n4851), .A2(n4849), .ZN(n9197) );
  NAND3_X1 U6286 ( .A1(n7924), .A2(n4853), .A3(n4854), .ZN(n4849) );
  NAND2_X2 U6287 ( .A1(n4850), .A2(n4854), .ZN(n8025) );
  NAND2_X1 U6288 ( .A1(n7815), .A2(n5989), .ZN(n7834) );
  INV_X1 U6289 ( .A(n4864), .ZN(n9177) );
  NAND2_X1 U6290 ( .A1(n5991), .A2(n5040), .ZN(n6041) );
  INV_X1 U6291 ( .A(n5050), .ZN(n4867) );
  NAND2_X1 U6292 ( .A1(n5353), .A2(n5354), .ZN(n4870) );
  NAND2_X1 U6293 ( .A1(n5112), .A2(n5102), .ZN(n5797) );
  OAI22_X1 U6294 ( .A1(n9245), .A2(n4875), .B1(n4873), .B2(n4876), .ZN(n4877)
         );
  NAND2_X1 U6295 ( .A1(n9614), .A2(n4885), .ZN(n4884) );
  OAI21_X1 U6296 ( .B1(n4905), .B2(n8943), .A(n4904), .ZN(n8916) );
  INV_X1 U6297 ( .A(n9909), .ZN(n4914) );
  NOR2_X1 U6298 ( .A1(n8402), .A2(n4914), .ZN(n4915) );
  NAND2_X1 U6299 ( .A1(n4915), .A2(n8408), .ZN(n5648) );
  INV_X1 U6300 ( .A(n7367), .ZN(n4924) );
  NAND2_X1 U6301 ( .A1(n6356), .A2(n6357), .ZN(n4925) );
  INV_X1 U6302 ( .A(n4564), .ZN(n4931) );
  NAND2_X1 U6303 ( .A1(n8234), .A2(n4938), .ZN(n4937) );
  NAND2_X1 U6304 ( .A1(n4980), .A2(n4946), .ZN(n5637) );
  INV_X1 U6305 ( .A(n4955), .ZN(n6683) );
  NAND2_X1 U6306 ( .A1(n8927), .A2(n5046), .ZN(n5526) );
  OR2_X1 U6307 ( .A1(n8248), .A2(n8666), .ZN(n4964) );
  OAI22_X2 U6308 ( .A1(n7413), .A2(n7416), .B1(n7500), .B2(n10348), .ZN(n7520)
         );
  NOR2_X1 U6309 ( .A1(n10250), .A2(n4548), .ZN(n7377) );
  NAND2_X1 U6310 ( .A1(n8831), .A2(n4969), .ZN(n4966) );
  NAND2_X1 U6311 ( .A1(n4966), .A2(n4967), .ZN(n8803) );
  NAND2_X1 U6312 ( .A1(n8831), .A2(n8510), .ZN(n4968) );
  INV_X1 U6313 ( .A(n4975), .ZN(n7934) );
  NOR2_X1 U6314 ( .A1(n9936), .A2(n7856), .ZN(n4977) );
  NOR2_X2 U6315 ( .A1(n7981), .A2(n8482), .ZN(n7980) );
  NAND4_X1 U6316 ( .A1(n4980), .A2(n4981), .A3(n5687), .A4(n5086), .ZN(n9066)
         );
  NOR2_X2 U6317 ( .A1(n5227), .A2(n5084), .ZN(n5678) );
  NAND2_X1 U6318 ( .A1(n4982), .A2(n4983), .ZN(n5599) );
  NAND2_X1 U6319 ( .A1(n8880), .A2(n4985), .ZN(n4982) );
  NAND2_X1 U6320 ( .A1(n4734), .A2(n8605), .ZN(n4990) );
  OAI21_X1 U6321 ( .B1(n9613), .B2(n8540), .A(n5006), .ZN(n9597) );
  NOR2_X1 U6322 ( .A1(n4992), .A2(n4993), .ZN(n9550) );
  NAND2_X1 U6323 ( .A1(n9551), .A2(n5010), .ZN(n5009) );
  OR2_X1 U6324 ( .A1(n10236), .A2(n6526), .ZN(n5013) );
  AOI21_X2 U6325 ( .B1(n9707), .B2(n9717), .A(n8535), .ZN(n9691) );
  NAND2_X1 U6326 ( .A1(n9336), .A2(n7623), .ZN(n7622) );
  NAND2_X1 U6327 ( .A1(n7675), .A2(n7582), .ZN(n7802) );
  OR2_X1 U6328 ( .A1(n7677), .A2(n7591), .ZN(n7675) );
  NAND2_X1 U6329 ( .A1(n7989), .A2(n4494), .ZN(n5020) );
  OAI211_X2 U6330 ( .C1(n7586), .C2(n5034), .A(n4518), .B(n5031), .ZN(n7712)
         );
  INV_X1 U6331 ( .A(n5034), .ZN(n5032) );
  INV_X1 U6332 ( .A(n5033), .ZN(n5036) );
  NAND2_X1 U6333 ( .A1(n5037), .A2(n7585), .ZN(n5033) );
  INV_X1 U6334 ( .A(n9339), .ZN(n5037) );
  NAND3_X1 U6335 ( .A1(n4514), .A2(n5726), .A3(n5038), .ZN(n5041) );
  NAND2_X1 U6336 ( .A1(n8520), .A2(n8519), .ZN(n8521) );
  NAND2_X1 U6337 ( .A1(n5239), .A2(n5238), .ZN(n5166) );
  AOI211_X1 U6338 ( .C1(n4491), .C2(n9991), .A(n9986), .B(n9985), .ZN(n9990)
         );
  OAI222_X1 U6339 ( .A1(P1_U3084), .A2(n4491), .B1(n9857), .B2(n8066), .C1(
        n8065), .C2(n8257), .ZN(P1_U3326) );
  AOI21_X1 U6340 ( .B1(n6443), .B2(n5049), .A(n5055), .ZN(n6446) );
  NAND2_X1 U6341 ( .A1(n6672), .A2(n6360), .ZN(n6326) );
  NAND2_X1 U6342 ( .A1(n6379), .A2(n6378), .ZN(n6380) );
  CLKBUF_X1 U6343 ( .A(n7237), .Z(n8483) );
  NAND2_X1 U6344 ( .A1(n7302), .A2(n6687), .ZN(n8352) );
  OR2_X1 U6345 ( .A1(n5328), .A2(n5327), .ZN(n5329) );
  NAND2_X1 U6346 ( .A1(n7511), .A2(n6642), .ZN(n8361) );
  INV_X1 U6347 ( .A(n5422), .ZN(n5423) );
  NOR2_X1 U6348 ( .A1(n6666), .A2(n6667), .ZN(n6665) );
  NAND2_X1 U6349 ( .A1(n5093), .A2(n8231), .ZN(n5328) );
  OAI22_X2 U6350 ( .A1(n8119), .A2(n5500), .B1(n8128), .B2(n8243), .ZN(n8245)
         );
  OAI22_X2 U6351 ( .A1(n8197), .A2(n8196), .B1(n6388), .B2(n6387), .ZN(n8234)
         );
  INV_X1 U6352 ( .A(n7817), .ZN(n5988) );
  AND2_X1 U6353 ( .A1(n6451), .A2(n8654), .ZN(n5043) );
  INV_X1 U6354 ( .A(n8642), .ZN(n8631) );
  NOR2_X1 U6355 ( .A1(n5909), .A2(n5907), .ZN(n5044) );
  OR2_X1 U6356 ( .A1(n9062), .A2(n8237), .ZN(n5045) );
  NOR2_X1 U6357 ( .A1(n5136), .A2(n5449), .ZN(n5047) );
  OR2_X1 U6358 ( .A1(n8445), .A2(n8634), .ZN(n5048) );
  NOR2_X1 U6359 ( .A1(n6440), .A2(n6442), .ZN(n5049) );
  AND3_X1 U6360 ( .A1(n7039), .A2(n5738), .A3(n5737), .ZN(n5050) );
  AND2_X1 U6361 ( .A1(n6057), .A2(n6056), .ZN(n5051) );
  AND2_X1 U6362 ( .A1(n5447), .A2(n5132), .ZN(n5052) );
  AND2_X1 U6363 ( .A1(n5149), .A2(n5148), .ZN(n5053) );
  OR2_X1 U6364 ( .A1(n7126), .A2(n7146), .ZN(n5054) );
  NOR2_X1 U6365 ( .A1(n6442), .A2(n6441), .ZN(n5055) );
  NOR2_X1 U6366 ( .A1(n9825), .A2(n9482), .ZN(n5056) );
  NAND2_X1 U6367 ( .A1(n8034), .A2(n8033), .ZN(n5057) );
  INV_X1 U6368 ( .A(n9017), .ZN(n5712) );
  INV_X1 U6369 ( .A(n9061), .ZN(n5716) );
  INV_X1 U6370 ( .A(n9199), .ZN(n9168) );
  OR2_X1 U6371 ( .A1(n6543), .A2(n9991), .ZN(n5058) );
  OR2_X1 U6372 ( .A1(n6278), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n5059) );
  AND2_X1 U6373 ( .A1(n7883), .A2(n7882), .ZN(n5060) );
  AND2_X1 U6374 ( .A1(n6320), .A2(n6319), .ZN(n5061) );
  OAI21_X1 U6375 ( .B1(n8677), .B2(n10321), .A(n10284), .ZN(n5422) );
  INV_X1 U6376 ( .A(n8827), .ZN(n8802) );
  INV_X1 U6377 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U6378 ( .A1(n9217), .A2(n9746), .ZN(n9425) );
  INV_X1 U6379 ( .A(n5550), .ZN(n5073) );
  INV_X1 U6380 ( .A(n6352), .ZN(n6353) );
  INV_X1 U6381 ( .A(n5517), .ZN(n5072) );
  INV_X1 U6382 ( .A(n5589), .ZN(n5588) );
  INV_X1 U6383 ( .A(n5493), .ZN(n5071) );
  INV_X1 U6384 ( .A(n5460), .ZN(n5066) );
  NAND2_X1 U6385 ( .A1(n5658), .A2(n8327), .ZN(n6323) );
  INV_X1 U6386 ( .A(n8679), .ZN(n5391) );
  INV_X1 U6387 ( .A(n6128), .ZN(n6140) );
  INV_X1 U6388 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5881) );
  INV_X1 U6389 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7004) );
  AND2_X1 U6390 ( .A1(n5543), .A2(n5545), .ZN(n5198) );
  NAND2_X1 U6391 ( .A1(n5502), .A2(n5501), .ZN(n5182) );
  OR2_X1 U6392 ( .A1(n5487), .A2(n5485), .ZN(n5171) );
  AND2_X1 U6393 ( .A1(n5294), .A2(n5296), .ZN(n5137) );
  INV_X1 U6394 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5924) );
  INV_X1 U6395 ( .A(n6465), .ZN(n6466) );
  INV_X1 U6396 ( .A(n6441), .ZN(n6433) );
  INV_X1 U6397 ( .A(n6377), .ZN(n6378) );
  OR2_X1 U6398 ( .A1(n5552), .A2(n8615), .ZN(n5571) );
  NAND2_X1 U6399 ( .A1(n5072), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U6400 ( .A1(n5672), .A2(n8330), .ZN(n6322) );
  NAND2_X1 U6401 ( .A1(n5588), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5623) );
  AND2_X1 U6402 ( .A1(n8950), .A2(n8665), .ZN(n5513) );
  OR2_X1 U6403 ( .A1(n5477), .A2(n8056), .ZN(n5479) );
  OR2_X1 U6404 ( .A1(n5289), .A2(n5275), .ZN(n5277) );
  INV_X1 U6405 ( .A(n8898), .ZN(n8919) );
  NOR2_X1 U6406 ( .A1(n6189), .A2(n9160), .ZN(n6190) );
  NOR2_X1 U6407 ( .A1(n6227), .A2(n9101), .ZN(n6244) );
  AND2_X1 U6408 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(n6140), .ZN(n6155) );
  OR2_X1 U6409 ( .A1(n6209), .A2(n9131), .ZN(n6227) );
  OR2_X1 U6410 ( .A1(n6030), .A2(n6029), .ZN(n6046) );
  NAND2_X1 U6411 ( .A1(n5892), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U6412 ( .A1(n5544), .A2(n5198), .ZN(n5200) );
  NAND2_X1 U6413 ( .A1(n5156), .A2(n5155), .ZN(n5159) );
  NAND2_X1 U6414 ( .A1(n5125), .A2(n5124), .ZN(n5128) );
  NAND2_X1 U6415 ( .A1(n4483), .A2(n8253), .ZN(n5110) );
  NOR2_X1 U6416 ( .A1(n6467), .A2(n6466), .ZN(n6468) );
  NAND2_X1 U6417 ( .A1(n6325), .A2(n6326), .ZN(n6332) );
  OR2_X1 U6418 ( .A1(n6384), .A2(n6383), .ZN(n6385) );
  OR2_X1 U6419 ( .A1(n5505), .A2(n8623), .ZN(n5517) );
  INV_X1 U6420 ( .A(n8329), .ZN(n6673) );
  AND2_X1 U6421 ( .A1(n5624), .A2(n8808), .ZN(n8821) );
  INV_X1 U6422 ( .A(n8659), .ZN(n8650) );
  INV_X1 U6423 ( .A(n8837), .ZN(n8845) );
  AND2_X1 U6424 ( .A1(n8426), .A2(n8432), .ZN(n8506) );
  INV_X1 U6425 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5087) );
  NOR2_X1 U6426 ( .A1(n6489), .A2(n6488), .ZN(n6523) );
  AND2_X1 U6427 ( .A1(n6318), .A2(n6317), .ZN(n6319) );
  INV_X1 U6428 ( .A(n6545), .ZN(n9986) );
  OR2_X1 U6429 ( .A1(n6754), .A2(n6753), .ZN(n6751) );
  INV_X1 U6430 ( .A(n9800), .ZN(n9697) );
  AND2_X1 U6431 ( .A1(n9242), .A2(n9244), .ZN(n9348) );
  OR2_X1 U6432 ( .A1(n9703), .A2(n7568), .ZN(n9951) );
  NAND2_X1 U6433 ( .A1(n5530), .A2(n5529), .ZN(n5532) );
  NAND2_X1 U6434 ( .A1(n5486), .A2(n5485), .ZN(n5488) );
  XNOR2_X1 U6435 ( .A(n5151), .B(SI_14_), .ZN(n5256) );
  NAND2_X1 U6436 ( .A1(n5128), .A2(n5127), .ZN(n5312) );
  OAI21_X1 U6437 ( .B1(n8842), .B2(n8657), .A(n6473), .ZN(n6474) );
  INV_X1 U6438 ( .A(n6457), .ZN(n6458) );
  INV_X1 U6439 ( .A(n8657), .ZN(n8618) );
  INV_X1 U6440 ( .A(n10238), .ZN(n9887) );
  NAND2_X1 U6441 ( .A1(n8804), .A2(n8300), .ZN(n8796) );
  INV_X1 U6442 ( .A(n8510), .ZN(n8833) );
  AND2_X1 U6443 ( .A1(n8341), .A2(n8338), .ZN(n7416) );
  INV_X1 U6444 ( .A(n10270), .ZN(n10283) );
  INV_X1 U6445 ( .A(n6426), .ZN(n7344) );
  AND2_X1 U6446 ( .A1(n5690), .A2(n5689), .ZN(n10297) );
  INV_X1 U6447 ( .A(n5678), .ZN(n5686) );
  AND2_X1 U6448 ( .A1(n5410), .A2(n5399), .ZN(n7143) );
  AND2_X1 U6449 ( .A1(n7544), .A2(n9964), .ZN(n9205) );
  AND4_X1 U6450 ( .A1(n6532), .A2(n6531), .A3(n6530), .A4(n6529), .ZN(n9557)
         );
  AND4_X1 U6451 ( .A1(n6133), .A2(n6132), .A3(n6131), .A4(n6130), .ZN(n9123)
         );
  AND4_X1 U6452 ( .A1(n6036), .A2(n6035), .A3(n6034), .A4(n6033), .ZN(n7990)
         );
  AND2_X1 U6453 ( .A1(n9713), .A2(n9715), .ZN(n9732) );
  OR2_X1 U6454 ( .A1(n7564), .A2(n10155), .ZN(n9669) );
  INV_X1 U6455 ( .A(n10187), .ZN(n10210) );
  OR2_X1 U6456 ( .A1(n9318), .A2(n7588), .ZN(n10155) );
  AND2_X1 U6457 ( .A1(n6653), .A2(n6652), .ZN(n7919) );
  NOR2_X1 U6458 ( .A1(n5747), .A2(n5746), .ZN(n5748) );
  NOR2_X1 U6459 ( .A1(n8104), .A2(n10423), .ZN(n8106) );
  INV_X1 U6460 ( .A(n6474), .ZN(n6475) );
  NOR2_X1 U6461 ( .A1(n5043), .A2(n6458), .ZN(n6459) );
  INV_X1 U6462 ( .A(n8639), .ZN(n8652) );
  AND2_X1 U6463 ( .A1(n6428), .A2(n8903), .ZN(n8657) );
  AND2_X1 U6464 ( .A1(n5100), .A2(n5099), .ZN(n8605) );
  NAND2_X1 U6465 ( .A1(n8827), .A2(n5712), .ZN(n5713) );
  OR2_X1 U6466 ( .A1(n5714), .A2(n6426), .ZN(n10380) );
  INV_X1 U6467 ( .A(n8323), .ZN(n9035) );
  OR2_X1 U6468 ( .A1(n5714), .A2(n7344), .ZN(n10370) );
  INV_X1 U6469 ( .A(n10307), .ZN(n10310) );
  AND2_X1 U6470 ( .A1(n6508), .A2(n6507), .ZN(n6509) );
  OR2_X1 U6471 ( .A1(n6293), .A2(n6308), .ZN(n9199) );
  INV_X1 U6472 ( .A(n8541), .ZN(n9592) );
  INV_X1 U6473 ( .A(n9682), .ZN(n9479) );
  INV_X1 U6474 ( .A(n7745), .ZN(n9485) );
  OR2_X1 U6475 ( .A1(P1_U3083), .A2(n6580), .ZN(n10116) );
  OR2_X1 U6476 ( .A1(n9703), .A2(n7575), .ZN(n9745) );
  OR2_X1 U6477 ( .A1(n9703), .A2(n7624), .ZN(n9953) );
  INV_X1 U6478 ( .A(n10236), .ZN(n10233) );
  OR3_X1 U6479 ( .A1(n9824), .A2(n9823), .A3(n9822), .ZN(n9846) );
  INV_X1 U6480 ( .A(n10218), .ZN(n10216) );
  CLKBUF_X1 U6481 ( .A(n10144), .Z(n10151) );
  INV_X1 U6482 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6878) );
  NOR2_X1 U6483 ( .A1(n10422), .A2(n10421), .ZN(n10420) );
  NOR2_X1 U6484 ( .A1(n10409), .A2(n10408), .ZN(n10407) );
  NAND3_X1 U6485 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5414) );
  INV_X1 U6486 ( .A(n5414), .ZN(n5062) );
  NAND2_X1 U6487 ( .A1(n5062), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5437) );
  INV_X1 U6488 ( .A(n5437), .ZN(n5063) );
  NAND2_X1 U6489 ( .A1(n5063), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5439) );
  INV_X1 U6490 ( .A(n5439), .ZN(n5064) );
  AND2_X1 U6491 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5065) );
  INV_X1 U6492 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8712) );
  INV_X1 U6493 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5275) );
  INV_X1 U6494 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8056) );
  INV_X1 U6495 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8748) );
  AND2_X1 U6496 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n5070) );
  INV_X1 U6497 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8623) );
  INV_X1 U6498 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8636) );
  INV_X1 U6499 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U6500 ( .A1(n5552), .A2(n8615), .ZN(n5074) );
  NAND2_X1 U6501 ( .A1(n5571), .A2(n5074), .ZN(n8888) );
  NOR2_X2 U6502 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5351) );
  NOR2_X1 U6503 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5075) );
  NAND3_X2 U6504 ( .A1(n5378), .A2(n5081), .A3(n5080), .ZN(n5227) );
  NOR2_X1 U6505 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5082) );
  NOR2_X1 U6506 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5674) );
  INV_X1 U6507 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5676) );
  NAND4_X1 U6508 ( .A1(n5083), .A2(n5082), .A3(n5674), .A4(n5676), .ZN(n5084)
         );
  INV_X1 U6509 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5687) );
  NOR2_X1 U6510 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n5089) );
  INV_X1 U6511 ( .A(n5089), .ZN(n5085) );
  NOR2_X1 U6512 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(n5085), .ZN(n5086) );
  XNOR2_X2 U6513 ( .A(n5088), .B(n5087), .ZN(n5093) );
  INV_X1 U6514 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5091) );
  OR2_X1 U6515 ( .A1(n8888), .A2(n5578), .ZN(n5100) );
  INV_X1 U6516 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9047) );
  NAND2_X2 U6517 ( .A1(n5093), .A2(n5094), .ZN(n5385) );
  NAND2_X1 U6518 ( .A1(n5326), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5097) );
  AND2_X2 U6519 ( .A1(n5095), .A2(n8231), .ZN(n5440) );
  OAI211_X1 U6520 ( .C1(n9047), .C2(n4485), .A(n5097), .B(n5096), .ZN(n5098)
         );
  INV_X1 U6521 ( .A(n5098), .ZN(n5099) );
  AND2_X1 U6522 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5102) );
  AND2_X1 U6523 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6524 ( .A1(n5797), .A2(n5348), .ZN(n5104) );
  XNOR2_X1 U6525 ( .A(n5104), .B(n6907), .ZN(n5336) );
  MUX2_X1 U6526 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5112), .Z(n5335) );
  NAND2_X1 U6527 ( .A1(n5336), .A2(n5335), .ZN(n5106) );
  NAND2_X1 U6528 ( .A1(n5104), .A2(SI_1_), .ZN(n5105) );
  NAND2_X1 U6529 ( .A1(n5106), .A2(n5105), .ZN(n5353) );
  INV_X1 U6530 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6586) );
  INV_X1 U6531 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6590) );
  MUX2_X1 U6532 ( .A(n6586), .B(n6590), .S(n5112), .Z(n5107) );
  XNOR2_X1 U6533 ( .A(n5107), .B(SI_2_), .ZN(n5354) );
  INV_X1 U6534 ( .A(n5107), .ZN(n5108) );
  NAND2_X1 U6535 ( .A1(n5108), .A2(SI_2_), .ZN(n5109) );
  INV_X1 U6536 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8256) );
  INV_X1 U6537 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n8253) );
  MUX2_X1 U6538 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5112), .Z(n5115) );
  NAND2_X1 U6539 ( .A1(n5115), .A2(SI_4_), .ZN(n5113) );
  INV_X1 U6540 ( .A(n5113), .ZN(n5116) );
  INV_X1 U6541 ( .A(SI_4_), .ZN(n5114) );
  INV_X1 U6542 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6592) );
  MUX2_X1 U6543 ( .A(n6992), .B(n6592), .S(n4483), .Z(n5117) );
  INV_X1 U6544 ( .A(n5117), .ZN(n5118) );
  NAND2_X1 U6545 ( .A1(n5118), .A2(SI_5_), .ZN(n5119) );
  INV_X1 U6546 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n8262) );
  INV_X1 U6547 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n8258) );
  MUX2_X1 U6548 ( .A(n8262), .B(n8258), .S(n4483), .Z(n5120) );
  INV_X1 U6549 ( .A(n5120), .ZN(n5121) );
  NAND2_X1 U6550 ( .A1(n5121), .A2(SI_6_), .ZN(n5122) );
  MUX2_X1 U6551 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4483), .Z(n5123) );
  INV_X1 U6552 ( .A(SI_7_), .ZN(n7018) );
  INV_X1 U6553 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6608) );
  INV_X1 U6554 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6606) );
  MUX2_X1 U6555 ( .A(n6608), .B(n6606), .S(n4483), .Z(n5125) );
  INV_X1 U6556 ( .A(SI_8_), .ZN(n5124) );
  INV_X1 U6557 ( .A(n5125), .ZN(n5126) );
  NAND2_X1 U6558 ( .A1(n5126), .A2(SI_8_), .ZN(n5127) );
  INV_X1 U6559 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6610) );
  INV_X1 U6560 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6611) );
  MUX2_X1 U6561 ( .A(n6610), .B(n6611), .S(n4483), .Z(n5130) );
  INV_X1 U6562 ( .A(SI_9_), .ZN(n5129) );
  INV_X1 U6563 ( .A(n5130), .ZN(n5131) );
  NAND2_X1 U6564 ( .A1(n5131), .A2(SI_9_), .ZN(n5132) );
  INV_X1 U6565 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6615) );
  INV_X1 U6566 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6616) );
  MUX2_X1 U6567 ( .A(n6615), .B(n6616), .S(n4483), .Z(n5134) );
  INV_X1 U6568 ( .A(SI_10_), .ZN(n5133) );
  NAND2_X1 U6569 ( .A1(n5134), .A2(n5133), .ZN(n5450) );
  INV_X1 U6570 ( .A(n5296), .ZN(n5136) );
  INV_X1 U6571 ( .A(n5134), .ZN(n5135) );
  INV_X1 U6572 ( .A(n5138), .ZN(n5139) );
  INV_X1 U6573 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6622) );
  INV_X1 U6574 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6623) );
  MUX2_X1 U6575 ( .A(n6622), .B(n6623), .S(n4483), .Z(n5141) );
  INV_X1 U6576 ( .A(SI_12_), .ZN(n5140) );
  INV_X1 U6577 ( .A(n5141), .ZN(n5142) );
  NAND2_X1 U6578 ( .A1(n5142), .A2(SI_12_), .ZN(n5143) );
  INV_X1 U6579 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6971) );
  INV_X1 U6580 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6662) );
  MUX2_X1 U6581 ( .A(n6971), .B(n6662), .S(n4483), .Z(n5146) );
  INV_X1 U6582 ( .A(SI_13_), .ZN(n5145) );
  NAND2_X1 U6583 ( .A1(n5146), .A2(n5145), .ZN(n5149) );
  INV_X1 U6584 ( .A(n5146), .ZN(n5147) );
  NAND2_X1 U6585 ( .A1(n5147), .A2(SI_13_), .ZN(n5148) );
  INV_X1 U6586 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6682) );
  INV_X1 U6587 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6680) );
  MUX2_X1 U6588 ( .A(n6682), .B(n6680), .S(n4483), .Z(n5151) );
  INV_X1 U6589 ( .A(n5151), .ZN(n5152) );
  NAND2_X1 U6590 ( .A1(n5152), .A2(SI_14_), .ZN(n5153) );
  INV_X1 U6591 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7193) );
  INV_X1 U6592 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7194) );
  MUX2_X1 U6593 ( .A(n7193), .B(n7194), .S(n4483), .Z(n5156) );
  INV_X1 U6594 ( .A(SI_15_), .ZN(n5155) );
  INV_X1 U6595 ( .A(n5156), .ZN(n5157) );
  NAND2_X1 U6596 ( .A1(n5157), .A2(SI_15_), .ZN(n5158) );
  INV_X1 U6597 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7227) );
  INV_X1 U6598 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5160) );
  MUX2_X1 U6599 ( .A(n7227), .B(n5160), .S(n4483), .Z(n5162) );
  INV_X1 U6600 ( .A(SI_16_), .ZN(n5161) );
  NAND2_X1 U6601 ( .A1(n5162), .A2(n5161), .ZN(n5165) );
  INV_X1 U6602 ( .A(n5162), .ZN(n5163) );
  NAND2_X1 U6603 ( .A1(n5163), .A2(SI_16_), .ZN(n5164) );
  MUX2_X1 U6604 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n4483), .Z(n5168) );
  INV_X1 U6605 ( .A(SI_17_), .ZN(n7051) );
  XNOR2_X1 U6606 ( .A(n5168), .B(n7051), .ZN(n5226) );
  INV_X1 U6607 ( .A(n5226), .ZN(n5483) );
  MUX2_X1 U6608 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4483), .Z(n5169) );
  XNOR2_X1 U6609 ( .A(n5169), .B(SI_18_), .ZN(n5487) );
  NAND2_X1 U6610 ( .A1(n5168), .A2(SI_17_), .ZN(n5485) );
  NAND2_X1 U6611 ( .A1(n5169), .A2(SI_18_), .ZN(n5170) );
  INV_X1 U6612 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7405) );
  INV_X1 U6613 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7403) );
  MUX2_X1 U6614 ( .A(n7405), .B(n7403), .S(n4483), .Z(n5174) );
  INV_X1 U6615 ( .A(SI_19_), .ZN(n5173) );
  NAND2_X1 U6616 ( .A1(n5174), .A2(n5173), .ZN(n5177) );
  INV_X1 U6617 ( .A(n5174), .ZN(n5175) );
  NAND2_X1 U6618 ( .A1(n5175), .A2(SI_19_), .ZN(n5176) );
  NAND2_X1 U6619 ( .A1(n5177), .A2(n5176), .ZN(n5218) );
  INV_X1 U6620 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7551) );
  INV_X1 U6621 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7549) );
  MUX2_X1 U6622 ( .A(n7551), .B(n7549), .S(n4483), .Z(n5178) );
  INV_X1 U6623 ( .A(SI_20_), .ZN(n6991) );
  NAND2_X1 U6624 ( .A1(n5178), .A2(n6991), .ZN(n5181) );
  INV_X1 U6625 ( .A(n5178), .ZN(n5179) );
  NAND2_X1 U6626 ( .A1(n5179), .A2(SI_20_), .ZN(n5180) );
  AND2_X2 U6627 ( .A1(n5182), .A2(n5181), .ZN(n5528) );
  INV_X1 U6628 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7711) );
  INV_X1 U6629 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7621) );
  MUX2_X1 U6630 ( .A(n7711), .B(n7621), .S(n4483), .Z(n5189) );
  XNOR2_X1 U6631 ( .A(n5189), .B(SI_21_), .ZN(n5527) );
  INV_X1 U6632 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8310) );
  INV_X1 U6633 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7800) );
  MUX2_X1 U6634 ( .A(n8310), .B(n7800), .S(n4483), .Z(n5185) );
  INV_X1 U6635 ( .A(SI_22_), .ZN(n5183) );
  NAND2_X1 U6636 ( .A1(n5185), .A2(n5183), .ZN(n5188) );
  AND2_X1 U6637 ( .A1(n5527), .A2(n5188), .ZN(n5184) );
  INV_X1 U6638 ( .A(n5188), .ZN(n5193) );
  INV_X1 U6639 ( .A(n5185), .ZN(n5186) );
  NAND2_X1 U6640 ( .A1(n5186), .A2(SI_22_), .ZN(n5187) );
  NAND2_X1 U6641 ( .A1(n5188), .A2(n5187), .ZN(n5531) );
  INV_X1 U6642 ( .A(n5531), .ZN(n5191) );
  INV_X1 U6643 ( .A(n5189), .ZN(n5190) );
  NAND2_X1 U6644 ( .A1(n5190), .A2(SI_21_), .ZN(n5529) );
  AND2_X1 U6645 ( .A1(n5191), .A2(n5529), .ZN(n5192) );
  INV_X1 U6646 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7778) );
  INV_X1 U6647 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7782) );
  MUX2_X1 U6648 ( .A(n7778), .B(n7782), .S(n4483), .Z(n5195) );
  INV_X1 U6649 ( .A(SI_23_), .ZN(n5194) );
  NAND2_X1 U6650 ( .A1(n5195), .A2(n5194), .ZN(n5199) );
  INV_X1 U6651 ( .A(n5195), .ZN(n5196) );
  NAND2_X1 U6652 ( .A1(n5196), .A2(SI_23_), .ZN(n5197) );
  AND2_X1 U6653 ( .A1(n5199), .A2(n5197), .ZN(n5545) );
  INV_X1 U6654 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7825) );
  INV_X1 U6655 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7827) );
  MUX2_X1 U6656 ( .A(n7825), .B(n7827), .S(n4483), .Z(n5560) );
  XNOR2_X1 U6657 ( .A(n5560), .B(SI_24_), .ZN(n5559) );
  NAND2_X1 U6658 ( .A1(n5678), .A2(n5687), .ZN(n5201) );
  INV_X1 U6659 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5204) );
  OR2_X1 U6660 ( .A1(n9065), .A2(n5204), .ZN(n5202) );
  NAND2_X1 U6661 ( .A1(n5205), .A2(n5202), .ZN(n5203) );
  XNOR2_X2 U6662 ( .A(n5203), .B(P2_IR_REG_28__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U6663 ( .A1(n5205), .A2(n5204), .ZN(n5207) );
  OR2_X1 U6664 ( .A1(n5205), .A2(n5204), .ZN(n5206) );
  NAND2_X1 U6665 ( .A1(n5207), .A2(n5206), .ZN(n8301) );
  NAND2_X2 U6666 ( .A1(n5660), .A2(n8301), .ZN(n5340) );
  INV_X2 U6667 ( .A(n5429), .ZN(n8297) );
  NAND2_X1 U6668 ( .A1(n7824), .A2(n8297), .ZN(n5209) );
  NAND2_X1 U6669 ( .A1(n5340), .A2(n4483), .ZN(n5334) );
  OR2_X1 U6670 ( .A1(n5377), .A2(n7825), .ZN(n5208) );
  INV_X1 U6671 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5211) );
  INV_X1 U6672 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5210) );
  OAI21_X1 U6673 ( .B1(n5493), .B2(n5211), .A(n5210), .ZN(n5212) );
  NAND2_X1 U6674 ( .A1(n5212), .A2(n5505), .ZN(n8574) );
  OR2_X1 U6675 ( .A1(n8574), .A2(n5578), .ZN(n5217) );
  INV_X1 U6676 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U6677 ( .A1(n5326), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6678 ( .A1(n5663), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5213) );
  OAI211_X1 U6679 ( .C1(n8778), .C2(n5666), .A(n5214), .B(n5213), .ZN(n5215)
         );
  INV_X1 U6680 ( .A(n5215), .ZN(n5216) );
  NAND2_X1 U6681 ( .A1(n5217), .A2(n5216), .ZN(n8666) );
  XNOR2_X1 U6682 ( .A(n5219), .B(n5218), .ZN(n7402) );
  NAND2_X1 U6683 ( .A1(n7402), .A2(n8297), .ZN(n5222) );
  INV_X2 U6684 ( .A(n5377), .ZN(n5490) );
  AOI22_X1 U6685 ( .A1(n5490), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8327), .B2(
        n4575), .ZN(n5221) );
  NAND2_X1 U6686 ( .A1(n5235), .A2(n8748), .ZN(n5223) );
  NAND2_X1 U6687 ( .A1(n5493), .A2(n5223), .ZN(n8198) );
  AOI22_X1 U6688 ( .A1(n5326), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n5663), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n5225) );
  INV_X1 U6689 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8074) );
  OR2_X1 U6690 ( .A1(n5666), .A2(n8074), .ZN(n5224) );
  OAI211_X1 U6691 ( .C1(n8198), .C2(n5553), .A(n5225), .B(n5224), .ZN(n8668)
         );
  XNOR2_X1 U6692 ( .A(n5484), .B(n5226), .ZN(n7264) );
  NAND2_X1 U6693 ( .A1(n7264), .A2(n8297), .ZN(n5232) );
  NAND2_X1 U6694 ( .A1(n5227), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5228) );
  MUX2_X1 U6695 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5228), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5230) );
  AND2_X1 U6696 ( .A1(n5230), .A2(n5229), .ZN(n8767) );
  AOI22_X1 U6697 ( .A1(n5490), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n4575), .B2(
        n8767), .ZN(n5231) );
  INV_X1 U6698 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7984) );
  INV_X1 U6699 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U6700 ( .A1(n5479), .A2(n5233), .ZN(n5234) );
  NAND2_X1 U6701 ( .A1(n5235), .A2(n5234), .ZN(n8151) );
  OR2_X1 U6702 ( .A1(n8151), .A2(n5553), .ZN(n5237) );
  AOI22_X1 U6703 ( .A1(n5326), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n5663), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n5236) );
  OAI211_X1 U6704 ( .C1(n5666), .C2(n7984), .A(n5237), .B(n5236), .ZN(n8669)
         );
  XNOR2_X1 U6705 ( .A(n5239), .B(n5238), .ZN(n7200) );
  NAND2_X1 U6706 ( .A1(n7200), .A2(n8297), .ZN(n5249) );
  INV_X1 U6707 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6708 ( .A1(n5378), .A2(n5379), .ZN(n5397) );
  INV_X1 U6709 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5240) );
  INV_X1 U6710 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5432) );
  NAND3_X1 U6711 ( .A1(n5240), .A2(n5398), .A3(n5432), .ZN(n5241) );
  NOR2_X1 U6712 ( .A1(n5397), .A2(n5241), .ZN(n5315) );
  INV_X1 U6713 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5242) );
  NAND2_X1 U6714 ( .A1(n5315), .A2(n5242), .ZN(n5298) );
  INV_X1 U6715 ( .A(n5243), .ZN(n5244) );
  OR3_X1 U6716 ( .A1(n5298), .A2(P2_IR_REG_10__SCAN_IN), .A3(n5244), .ZN(n5284) );
  OR2_X1 U6717 ( .A1(n5284), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5258) );
  INV_X1 U6718 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5245) );
  NAND3_X1 U6719 ( .A1(n5471), .A2(n5259), .A3(n5245), .ZN(n5246) );
  OAI21_X1 U6720 ( .B1(n5258), .B2(n5246), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5247) );
  XNOR2_X1 U6721 ( .A(n5247), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8746) );
  AOI22_X1 U6722 ( .A1(n5490), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n4575), .B2(
        n8746), .ZN(n5248) );
  NAND2_X1 U6723 ( .A1(n5326), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5255) );
  NAND2_X1 U6724 ( .A1(n5663), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5254) );
  INV_X1 U6725 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U6726 ( .A1(n5269), .A2(n5250), .ZN(n5251) );
  NAND2_X1 U6727 ( .A1(n5477), .A2(n5251), .ZN(n9915) );
  OR2_X1 U6728 ( .A1(n5578), .A2(n9915), .ZN(n5253) );
  NAND4_X1 U6729 ( .A1(n5255), .A2(n5254), .A3(n5253), .A4(n5252), .ZN(n8671)
         );
  INV_X1 U6730 ( .A(n8671), .ZN(n8058) );
  XNOR2_X1 U6731 ( .A(n5257), .B(n5256), .ZN(n6679) );
  NAND2_X1 U6732 ( .A1(n6679), .A2(n8297), .ZN(n5262) );
  NAND2_X1 U6733 ( .A1(n5258), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5264) );
  NAND2_X1 U6734 ( .A1(n5264), .A2(n5259), .ZN(n5260) );
  NAND2_X1 U6735 ( .A1(n5260), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5472) );
  XNOR2_X1 U6736 ( .A(n5472), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8177) );
  AOI22_X1 U6737 ( .A1(n5490), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8177), .B2(
        n4575), .ZN(n5261) );
  INV_X1 U6738 ( .A(n9917), .ZN(n9930) );
  NAND2_X1 U6739 ( .A1(n6661), .A2(n8297), .ZN(n5266) );
  XNOR2_X1 U6740 ( .A(n5264), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7962) );
  AOI22_X1 U6741 ( .A1(n5490), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n4575), .B2(
        n7962), .ZN(n5265) );
  INV_X1 U6742 ( .A(n5468), .ZN(n9936) );
  NAND2_X1 U6743 ( .A1(n5326), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5273) );
  INV_X1 U6744 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U6745 ( .A1(n5277), .A2(n5267), .ZN(n5268) );
  NAND2_X1 U6746 ( .A1(n5269), .A2(n5268), .ZN(n7735) );
  OR2_X1 U6747 ( .A1(n5553), .A2(n7735), .ZN(n5272) );
  INV_X1 U6748 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7614) );
  OR2_X1 U6749 ( .A1(n5666), .A2(n7614), .ZN(n5271) );
  NAND2_X1 U6750 ( .A1(n5663), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5270) );
  NAND4_X1 U6751 ( .A1(n5273), .A2(n5272), .A3(n5271), .A4(n5270), .ZN(n8672)
         );
  INV_X1 U6752 ( .A(n8672), .ZN(n7856) );
  INV_X1 U6753 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5274) );
  OR2_X1 U6754 ( .A1(n4485), .A2(n5274), .ZN(n5281) );
  INV_X1 U6755 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7767) );
  OR2_X1 U6756 ( .A1(n8318), .A2(n7767), .ZN(n5280) );
  NAND2_X1 U6757 ( .A1(n5289), .A2(n5275), .ZN(n5276) );
  NAND2_X1 U6758 ( .A1(n5277), .A2(n5276), .ZN(n7649) );
  OR2_X1 U6759 ( .A1(n5578), .A2(n7649), .ZN(n5279) );
  INV_X1 U6760 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7475) );
  OR2_X1 U6761 ( .A1(n5666), .A2(n7475), .ZN(n5278) );
  NAND4_X1 U6762 ( .A1(n5281), .A2(n5280), .A3(n5279), .A4(n5278), .ZN(n8673)
         );
  INV_X1 U6763 ( .A(n8673), .ZN(n7736) );
  XNOR2_X1 U6764 ( .A(n5283), .B(n5282), .ZN(n6621) );
  NAND2_X1 U6765 ( .A1(n6621), .A2(n8297), .ZN(n5287) );
  NAND2_X1 U6766 ( .A1(n5284), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5285) );
  XNOR2_X1 U6767 ( .A(n5285), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7866) );
  AOI22_X1 U6768 ( .A1(n5490), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n4575), .B2(
        n7866), .ZN(n5286) );
  NAND2_X1 U6769 ( .A1(n5287), .A2(n5286), .ZN(n7479) );
  INV_X1 U6770 ( .A(n7479), .ZN(n10363) );
  NAND2_X1 U6771 ( .A1(n5663), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6772 ( .A1(n5461), .A2(n8712), .ZN(n5288) );
  NAND2_X1 U6773 ( .A1(n5289), .A2(n5288), .ZN(n7525) );
  OR2_X1 U6774 ( .A1(n5553), .A2(n7525), .ZN(n5292) );
  INV_X1 U6775 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7526) );
  OR2_X1 U6776 ( .A1(n5666), .A2(n7526), .ZN(n5291) );
  NAND2_X1 U6777 ( .A1(n5326), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5290) );
  NAND4_X1 U6778 ( .A1(n5293), .A2(n5292), .A3(n5291), .A4(n5290), .ZN(n8674)
         );
  INV_X1 U6779 ( .A(n8674), .ZN(n5467) );
  NAND2_X1 U6780 ( .A1(n5448), .A2(n5294), .ZN(n5295) );
  AND2_X1 U6781 ( .A1(n5295), .A2(n5449), .ZN(n5297) );
  XNOR2_X1 U6782 ( .A(n5297), .B(n5296), .ZN(n6618) );
  NAND2_X1 U6783 ( .A1(n6618), .A2(n8297), .ZN(n5303) );
  NAND2_X1 U6784 ( .A1(n5298), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5309) );
  INV_X1 U6785 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6786 ( .A1(n5309), .A2(n5299), .ZN(n5300) );
  NAND2_X1 U6787 ( .A1(n5300), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5453) );
  INV_X1 U6788 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U6789 ( .A1(n5453), .A2(n5452), .ZN(n5455) );
  NAND2_X1 U6790 ( .A1(n5455), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5301) );
  XNOR2_X1 U6791 ( .A(n5301), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8711) );
  AOI22_X1 U6792 ( .A1(n5490), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n4575), .B2(
        n8711), .ZN(n5302) );
  NAND2_X1 U6793 ( .A1(n5303), .A2(n5302), .ZN(n7528) );
  INV_X1 U6794 ( .A(n7528), .ZN(n10356) );
  NAND2_X1 U6795 ( .A1(n5663), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U6796 ( .A1(n5326), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5306) );
  INV_X1 U6797 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5459) );
  XNOR2_X1 U6798 ( .A(n5460), .B(n5459), .ZN(n7384) );
  OR2_X1 U6799 ( .A1(n5553), .A2(n7384), .ZN(n5305) );
  NAND4_X1 U6800 ( .A1(n5307), .A2(n5306), .A3(n5305), .A4(n5304), .ZN(n10257)
         );
  XNOR2_X1 U6801 ( .A(n5308), .B(n5052), .ZN(n6609) );
  NAND2_X1 U6802 ( .A1(n6609), .A2(n8297), .ZN(n5311) );
  XNOR2_X1 U6803 ( .A(n5309), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8706) );
  AOI22_X1 U6804 ( .A1(n5490), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n4575), .B2(
        n8706), .ZN(n5310) );
  INV_X1 U6805 ( .A(n5312), .ZN(n5313) );
  XNOR2_X1 U6806 ( .A(n5314), .B(n5313), .ZN(n6607) );
  OR2_X1 U6807 ( .A1(n5315), .A2(n9065), .ZN(n5316) );
  XNOR2_X1 U6808 ( .A(n5316), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7333) );
  AOI22_X1 U6809 ( .A1(n5490), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n4575), .B2(
        n7333), .ZN(n5317) );
  NAND2_X1 U6810 ( .A1(n5326), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5325) );
  INV_X1 U6811 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U6812 ( .A1(n5439), .A2(n5319), .ZN(n5320) );
  NAND2_X1 U6813 ( .A1(n5460), .A2(n5320), .ZN(n8586) );
  OR2_X1 U6814 ( .A1(n5578), .A2(n8586), .ZN(n5324) );
  INV_X1 U6815 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5321) );
  OR2_X1 U6816 ( .A1(n4485), .A2(n5321), .ZN(n5323) );
  NAND4_X1 U6817 ( .A1(n5325), .A2(n5324), .A3(n5323), .A4(n5322), .ZN(n8676)
         );
  INV_X1 U6818 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7506) );
  OR2_X1 U6819 ( .A1(n5553), .A2(n7506), .ZN(n5331) );
  NAND2_X1 U6820 ( .A1(n5440), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5330) );
  INV_X1 U6821 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5327) );
  AND4_X2 U6822 ( .A1(n5332), .A2(n5331), .A3(n5330), .A4(n5329), .ZN(n6642)
         );
  INV_X1 U6823 ( .A(n5351), .ZN(n5333) );
  INV_X1 U6824 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6584) );
  OR2_X1 U6825 ( .A1(n5334), .A2(n6584), .ZN(n5339) );
  XNOR2_X1 U6826 ( .A(n5336), .B(n5335), .ZN(n6593) );
  OR2_X1 U6827 ( .A1(n5337), .A2(n6593), .ZN(n5338) );
  NAND2_X1 U6828 ( .A1(n8358), .A2(n8361), .ZN(n7237) );
  NAND2_X1 U6829 ( .A1(n5440), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5345) );
  INV_X1 U6830 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9880) );
  OR2_X1 U6831 ( .A1(n5385), .A2(n9880), .ZN(n5344) );
  INV_X1 U6832 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5341) );
  INV_X1 U6833 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7349) );
  OR2_X1 U6834 ( .A1(n5553), .A2(n7349), .ZN(n5342) );
  INV_X1 U6835 ( .A(n6327), .ZN(n8683) );
  INV_X1 U6836 ( .A(n4579), .ZN(n10246) );
  INV_X1 U6837 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6838 ( .A1(n5347), .A2(n5346), .ZN(n5349) );
  NAND2_X1 U6839 ( .A1(n5349), .A2(n5348), .ZN(n9072) );
  NAND2_X1 U6840 ( .A1(n8683), .A2(n6328), .ZN(n7239) );
  NAND2_X1 U6841 ( .A1(n7237), .A2(n7239), .ZN(n7238) );
  NAND2_X1 U6842 ( .A1(n7263), .A2(n6642), .ZN(n5350) );
  INV_X1 U6843 ( .A(n5553), .ZN(n5668) );
  NAND2_X1 U6844 ( .A1(n5668), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5361) );
  INV_X1 U6845 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7121) );
  OR2_X1 U6846 ( .A1(n5385), .A2(n7121), .ZN(n5360) );
  NAND2_X1 U6847 ( .A1(n5440), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U6848 ( .A1(n5663), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5358) );
  AND4_X1 U6849 ( .A1(n5361), .A2(n5360), .A3(n5359), .A4(n5358), .ZN(n5357)
         );
  OR2_X1 U6850 ( .A1(n5351), .A2(n9065), .ZN(n5352) );
  XNOR2_X1 U6851 ( .A(n5352), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9892) );
  INV_X1 U6852 ( .A(n9892), .ZN(n6585) );
  XNOR2_X1 U6853 ( .A(n5353), .B(n5354), .ZN(n6589) );
  OR2_X1 U6854 ( .A1(n5334), .A2(n6586), .ZN(n5355) );
  NAND2_X1 U6855 ( .A1(n7269), .A2(n8484), .ZN(n7268) );
  NAND2_X1 U6856 ( .A1(n7279), .A2(n5357), .ZN(n5362) );
  NAND2_X1 U6857 ( .A1(n7268), .A2(n5362), .ZN(n7211) );
  NAND2_X1 U6858 ( .A1(n5326), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5367) );
  INV_X1 U6859 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5363) );
  OR2_X1 U6860 ( .A1(n4485), .A2(n5363), .ZN(n5366) );
  OR2_X1 U6861 ( .A1(n5553), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5365) );
  NAND4_X1 U6862 ( .A1(n5367), .A2(n5366), .A3(n5365), .A4(n5364), .ZN(n8680)
         );
  INV_X1 U6863 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6910) );
  NAND2_X1 U6864 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4517), .ZN(n5368) );
  XNOR2_X1 U6865 ( .A(n6910), .B(n5368), .ZN(n8254) );
  XNOR2_X1 U6866 ( .A(n5370), .B(n5369), .ZN(n8255) );
  OR2_X1 U6867 ( .A1(n8255), .A2(n5429), .ZN(n5372) );
  OR2_X1 U6868 ( .A1(n5377), .A2(n8256), .ZN(n5371) );
  OAI211_X1 U6869 ( .C1(n7126), .C2(n8254), .A(n5372), .B(n5371), .ZN(n6338)
         );
  NAND2_X1 U6870 ( .A1(n6688), .A2(n4480), .ZN(n8348) );
  NAND2_X1 U6871 ( .A1(n6638), .A2(n8680), .ZN(n8372) );
  NAND2_X1 U6872 ( .A1(n6638), .A2(n6688), .ZN(n8263) );
  NAND2_X1 U6873 ( .A1(n5374), .A2(n5373), .ZN(n5376) );
  XNOR2_X1 U6874 ( .A(n5376), .B(n5375), .ZN(n5856) );
  INV_X1 U6875 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6587) );
  OR2_X1 U6876 ( .A1(n5377), .A2(n6587), .ZN(n5381) );
  OR2_X1 U6877 ( .A1(n5378), .A2(n9065), .ZN(n5380) );
  XNOR2_X1 U6878 ( .A(n5380), .B(n5379), .ZN(n7146) );
  XNOR2_X1 U6879 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8272) );
  OR2_X1 U6880 ( .A1(n5578), .A2(n8272), .ZN(n5389) );
  NAND2_X1 U6881 ( .A1(n5663), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5388) );
  INV_X1 U6882 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6883 ( .A1(n5440), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U6884 ( .A1(n10315), .A2(n5391), .ZN(n5390) );
  AND2_X1 U6885 ( .A1(n8263), .A2(n5390), .ZN(n5394) );
  INV_X1 U6886 ( .A(n5390), .ZN(n5392) );
  NAND2_X1 U6887 ( .A1(n5391), .A2(n8271), .ZN(n8349) );
  XNOR2_X1 U6888 ( .A(n5396), .B(n5395), .ZN(n6591) );
  OR2_X1 U6889 ( .A1(n6591), .A2(n5429), .ZN(n5401) );
  NAND2_X1 U6890 ( .A1(n5397), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6891 ( .A1(n5431), .A2(n5398), .ZN(n5410) );
  OR2_X1 U6892 ( .A1(n5431), .A2(n5398), .ZN(n5399) );
  AOI22_X1 U6893 ( .A1(n5490), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n4575), .B2(
        n7143), .ZN(n5400) );
  NAND2_X1 U6894 ( .A1(n5663), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5407) );
  INV_X1 U6895 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7144) );
  OR2_X1 U6896 ( .A1(n8318), .A2(n7144), .ZN(n5406) );
  INV_X1 U6897 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6695) );
  NAND2_X1 U6898 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5402) );
  NAND2_X1 U6899 ( .A1(n6695), .A2(n5402), .ZN(n5403) );
  NAND2_X1 U6900 ( .A1(n5414), .A2(n5403), .ZN(n7463) );
  OR2_X1 U6901 ( .A1(n5553), .A2(n7463), .ZN(n5405) );
  NAND2_X1 U6902 ( .A1(n7465), .A2(n8678), .ZN(n8371) );
  INV_X1 U6903 ( .A(n8678), .ZN(n6687) );
  NAND2_X1 U6904 ( .A1(n8371), .A2(n8352), .ZN(n8489) );
  XNOR2_X1 U6905 ( .A(n5409), .B(n5408), .ZN(n8261) );
  NAND2_X1 U6906 ( .A1(n5410), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5411) );
  XNOR2_X1 U6907 ( .A(n5411), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7168) );
  AOI22_X1 U6908 ( .A1(n5490), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n4575), .B2(
        n7168), .ZN(n5412) );
  INV_X1 U6909 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7148) );
  OR2_X1 U6910 ( .A1(n8318), .A2(n7148), .ZN(n5419) );
  INV_X1 U6911 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7233) );
  NAND2_X1 U6912 ( .A1(n5414), .A2(n7233), .ZN(n5415) );
  NAND2_X1 U6913 ( .A1(n5437), .A2(n5415), .ZN(n10280) );
  OR2_X1 U6914 ( .A1(n5578), .A2(n10280), .ZN(n5417) );
  NAND2_X1 U6915 ( .A1(n5663), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5416) );
  NAND4_X1 U6916 ( .A1(n5419), .A2(n5418), .A3(n5417), .A4(n5416), .ZN(n8677)
         );
  NAND2_X1 U6917 ( .A1(n10321), .A2(n8677), .ZN(n5421) );
  AND2_X1 U6918 ( .A1(n8489), .A2(n5421), .ZN(n5420) );
  NAND2_X1 U6919 ( .A1(n7282), .A2(n5420), .ZN(n5426) );
  INV_X1 U6920 ( .A(n5421), .ZN(n5424) );
  NAND2_X1 U6921 ( .A1(n7465), .A2(n6687), .ZN(n10284) );
  NAND2_X1 U6922 ( .A1(n5426), .A2(n5425), .ZN(n7459) );
  OR2_X1 U6923 ( .A1(n6599), .A2(n5429), .ZN(n5435) );
  OAI21_X1 U6924 ( .B1(P2_IR_REG_6__SCAN_IN), .B2(P2_IR_REG_5__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U6925 ( .A1(n5431), .A2(n5430), .ZN(n5433) );
  XNOR2_X1 U6926 ( .A(n5433), .B(n5432), .ZN(n7330) );
  AOI22_X1 U6927 ( .A1(n5490), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n4575), .B2(
        n7330), .ZN(n5434) );
  NAND2_X1 U6928 ( .A1(n5663), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5444) );
  INV_X1 U6929 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7173) );
  OR2_X1 U6930 ( .A1(n8318), .A2(n7173), .ZN(n5443) );
  INV_X1 U6931 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6932 ( .A1(n5437), .A2(n5436), .ZN(n5438) );
  NAND2_X1 U6933 ( .A1(n5439), .A2(n5438), .ZN(n7452) );
  OR2_X1 U6934 ( .A1(n5553), .A2(n7452), .ZN(n5442) );
  NAND2_X1 U6935 ( .A1(n5440), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5441) );
  NAND4_X1 U6936 ( .A1(n5444), .A2(n5443), .A3(n5442), .A4(n5441), .ZN(n10259)
         );
  INV_X1 U6937 ( .A(n10259), .ZN(n5445) );
  NAND2_X1 U6938 ( .A1(n7458), .A2(n5445), .ZN(n8385) );
  NOR2_X1 U6939 ( .A1(n7458), .A2(n10259), .ZN(n5446) );
  INV_X1 U6940 ( .A(n8676), .ZN(n7379) );
  NAND2_X1 U6941 ( .A1(n8588), .A2(n7379), .ZN(n8389) );
  INV_X1 U6942 ( .A(n10257), .ZN(n8583) );
  NAND2_X1 U6943 ( .A1(n7389), .A2(n8583), .ZN(n8392) );
  AND2_X1 U6944 ( .A1(n5450), .A2(n5449), .ZN(n5451) );
  NAND2_X1 U6945 ( .A1(n6614), .A2(n8297), .ZN(n5457) );
  OR2_X1 U6946 ( .A1(n5453), .A2(n5452), .ZN(n5454) );
  AND2_X1 U6947 ( .A1(n5455), .A2(n5454), .ZN(n7758) );
  AOI22_X1 U6948 ( .A1(n5490), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n4575), .B2(
        n7758), .ZN(n5456) );
  NAND2_X1 U6949 ( .A1(n5663), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U6950 ( .A1(n5326), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5465) );
  INV_X1 U6951 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5458) );
  OAI21_X1 U6952 ( .B1(n5460), .B2(n5459), .A(n5458), .ZN(n5462) );
  NAND2_X1 U6953 ( .A1(n5462), .A2(n5461), .ZN(n7420) );
  OR2_X1 U6954 ( .A1(n5578), .A2(n7420), .ZN(n5464) );
  NAND4_X1 U6955 ( .A1(n5466), .A2(n5465), .A3(n5464), .A4(n5463), .ZN(n8675)
         );
  INV_X1 U6956 ( .A(n8675), .ZN(n7500) );
  NAND2_X1 U6957 ( .A1(n7425), .A2(n7500), .ZN(n8338) );
  INV_X1 U6958 ( .A(n7425), .ZN(n10348) );
  OR2_X1 U6959 ( .A1(n7528), .A2(n5467), .ZN(n8342) );
  NAND2_X1 U6960 ( .A1(n7528), .A2(n5467), .ZN(n8398) );
  NAND2_X1 U6961 ( .A1(n8342), .A2(n8398), .ZN(n8497) );
  OAI21_X1 U6962 ( .B1(n5467), .B2(n10356), .A(n7519), .ZN(n7474) );
  OR2_X1 U6963 ( .A1(n7479), .A2(n7736), .ZN(n8399) );
  NAND2_X1 U6964 ( .A1(n7479), .A2(n7736), .ZN(n8402) );
  NAND2_X1 U6965 ( .A1(n5468), .A2(n7856), .ZN(n9909) );
  OR2_X1 U6966 ( .A1(n9917), .A2(n8058), .ZN(n8412) );
  NAND2_X1 U6967 ( .A1(n9917), .A2(n8058), .ZN(n8411) );
  XNOR2_X1 U6968 ( .A(n5470), .B(n5469), .ZN(n7192) );
  NAND2_X1 U6969 ( .A1(n7192), .A2(n8297), .ZN(n5476) );
  NAND2_X1 U6970 ( .A1(n5472), .A2(n5471), .ZN(n5473) );
  NAND2_X1 U6971 ( .A1(n5473), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5474) );
  XNOR2_X1 U6972 ( .A(n5474), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8726) );
  AOI22_X1 U6973 ( .A1(n8726), .A2(n4575), .B1(n5490), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U6974 ( .A1(n5477), .A2(n8056), .ZN(n5478) );
  NAND2_X1 U6975 ( .A1(n5479), .A2(n5478), .ZN(n8057) );
  INV_X1 U6976 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5480) );
  OAI22_X1 U6977 ( .A1(n8057), .A2(n5578), .B1(n8318), .B2(n5480), .ZN(n5482)
         );
  INV_X1 U6978 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7938) );
  INV_X1 U6979 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n6988) );
  OAI22_X1 U6980 ( .A1(n5666), .A2(n7938), .B1(n4485), .B2(n6988), .ZN(n5481)
         );
  OR2_X1 U6981 ( .A1(n5482), .A2(n5481), .ZN(n8670) );
  INV_X1 U6982 ( .A(n8670), .ZN(n8152) );
  OR2_X1 U6983 ( .A1(n8060), .A2(n8152), .ZN(n8415) );
  NAND2_X1 U6984 ( .A1(n8060), .A2(n8152), .ZN(n8416) );
  INV_X1 U6985 ( .A(n8669), .ZN(n8199) );
  OR2_X1 U6986 ( .A1(n9025), .A2(n8199), .ZN(n8419) );
  NAND2_X1 U6987 ( .A1(n9025), .A2(n8199), .ZN(n8418) );
  INV_X1 U6988 ( .A(n8668), .ZN(n8122) );
  OR2_X1 U6989 ( .A1(n8203), .A2(n8122), .ZN(n8336) );
  NAND2_X1 U6990 ( .A1(n8203), .A2(n8122), .ZN(n8334) );
  NAND2_X1 U6991 ( .A1(n8336), .A2(n8334), .ZN(n8504) );
  NAND2_X1 U6992 ( .A1(n7318), .A2(n8297), .ZN(n5492) );
  NAND2_X1 U6993 ( .A1(n5229), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5489) );
  XNOR2_X1 U6994 ( .A(n5489), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8769) );
  AOI22_X1 U6995 ( .A1(n5490), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n4575), .B2(
        n8769), .ZN(n5491) );
  XNOR2_X1 U6996 ( .A(n5493), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8235) );
  NAND2_X1 U6997 ( .A1(n8235), .A2(n5668), .ZN(n5499) );
  INV_X1 U6998 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U6999 ( .A1(n5663), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5495) );
  INV_X1 U7000 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8780) );
  OR2_X1 U7001 ( .A1(n8318), .A2(n8780), .ZN(n5494) );
  OAI211_X1 U7002 ( .C1(n5666), .C2(n5496), .A(n5495), .B(n5494), .ZN(n5497)
         );
  INV_X1 U7003 ( .A(n5497), .ZN(n5498) );
  NAND2_X1 U7004 ( .A1(n5499), .A2(n5498), .ZN(n8667) );
  NOR2_X1 U7005 ( .A1(n9020), .A2(n8667), .ZN(n5500) );
  INV_X1 U7006 ( .A(n9020), .ZN(n8128) );
  INV_X1 U7007 ( .A(n8667), .ZN(n8243) );
  INV_X1 U7008 ( .A(n8248), .ZN(n9062) );
  INV_X1 U7009 ( .A(n8666), .ZN(n8237) );
  XNOR2_X1 U7010 ( .A(n5502), .B(n5501), .ZN(n7548) );
  NAND2_X1 U7011 ( .A1(n7548), .A2(n8297), .ZN(n5504) );
  OR2_X1 U7012 ( .A1(n5377), .A2(n7551), .ZN(n5503) );
  NAND2_X1 U7013 ( .A1(n5505), .A2(n8623), .ZN(n5506) );
  AND2_X1 U7014 ( .A1(n5517), .A2(n5506), .ZN(n8951) );
  NAND2_X1 U7015 ( .A1(n8951), .A2(n5668), .ZN(n5512) );
  INV_X1 U7016 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U7017 ( .A1(n5663), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U7018 ( .A1(n5326), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5507) );
  OAI211_X1 U7019 ( .C1(n5509), .C2(n5666), .A(n5508), .B(n5507), .ZN(n5510)
         );
  INV_X1 U7020 ( .A(n5510), .ZN(n5511) );
  NAND2_X1 U7021 ( .A1(n5512), .A2(n5511), .ZN(n8665) );
  INV_X1 U7022 ( .A(n8665), .ZN(n8595) );
  NAND2_X1 U7023 ( .A1(n8950), .A2(n8595), .ZN(n8433) );
  NAND2_X1 U7024 ( .A1(n8436), .A2(n8433), .ZN(n8944) );
  OR2_X1 U7025 ( .A1(n5377), .A2(n7711), .ZN(n5515) );
  INV_X1 U7026 ( .A(n9002), .ZN(n8934) );
  INV_X1 U7027 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7028 ( .A1(n5517), .A2(n5516), .ZN(n5518) );
  NAND2_X1 U7029 ( .A1(n5535), .A2(n5518), .ZN(n8931) );
  OR2_X1 U7030 ( .A1(n8931), .A2(n5578), .ZN(n5524) );
  INV_X1 U7031 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7032 ( .A1(n5326), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5520) );
  INV_X1 U7033 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n6875) );
  OR2_X1 U7034 ( .A1(n4485), .A2(n6875), .ZN(n5519) );
  OAI211_X1 U7035 ( .C1(n5666), .C2(n5521), .A(n5520), .B(n5519), .ZN(n5522)
         );
  INV_X1 U7036 ( .A(n5522), .ZN(n5523) );
  NAND2_X1 U7037 ( .A1(n5524), .A2(n5523), .ZN(n8664) );
  INV_X1 U7038 ( .A(n8664), .ZN(n8633) );
  NAND2_X1 U7039 ( .A1(n5526), .A2(n5525), .ZN(n8913) );
  NAND2_X1 U7040 ( .A1(n5528), .A2(n5527), .ZN(n5530) );
  NAND2_X1 U7041 ( .A1(n7799), .A2(n8297), .ZN(n5534) );
  OR2_X1 U7042 ( .A1(n5377), .A2(n8310), .ZN(n5533) );
  NAND2_X1 U7043 ( .A1(n5535), .A2(n8636), .ZN(n5536) );
  AND2_X1 U7044 ( .A1(n5550), .A2(n5536), .ZN(n8921) );
  NAND2_X1 U7045 ( .A1(n8921), .A2(n5668), .ZN(n5542) );
  INV_X1 U7046 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U7047 ( .A1(n5326), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7048 ( .A1(n5663), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5537) );
  OAI211_X1 U7049 ( .C1(n5666), .C2(n5539), .A(n5538), .B(n5537), .ZN(n5540)
         );
  INV_X1 U7050 ( .A(n5540), .ZN(n5541) );
  NAND2_X1 U7051 ( .A1(n5542), .A2(n5541), .ZN(n8663) );
  INV_X1 U7052 ( .A(n8663), .ZN(n8596) );
  NAND2_X1 U7053 ( .A1(n8920), .A2(n8596), .ZN(n8439) );
  NAND2_X1 U7054 ( .A1(n8438), .A2(n8439), .ZN(n8912) );
  INV_X1 U7055 ( .A(n8920), .ZN(n9053) );
  AOI22_X1 U7056 ( .A1(n8913), .A2(n8912), .B1(n8596), .B2(n9053), .ZN(n8902)
         );
  AND2_X1 U7057 ( .A1(n5544), .A2(n5543), .ZN(n5546) );
  NAND2_X1 U7058 ( .A1(n7779), .A2(n8297), .ZN(n5548) );
  OR2_X1 U7059 ( .A1(n5377), .A2(n7778), .ZN(n5547) );
  INV_X1 U7060 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U7061 ( .A1(n5550), .A2(n5549), .ZN(n5551) );
  NAND2_X1 U7062 ( .A1(n5552), .A2(n5551), .ZN(n8904) );
  OR2_X1 U7063 ( .A1(n8904), .A2(n5553), .ZN(n5558) );
  INV_X1 U7064 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8905) );
  NAND2_X1 U7065 ( .A1(n5326), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5555) );
  INV_X1 U7066 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n7019) );
  OR2_X1 U7067 ( .A1(n4485), .A2(n7019), .ZN(n5554) );
  OAI211_X1 U7068 ( .C1(n5666), .C2(n8905), .A(n5555), .B(n5554), .ZN(n5556)
         );
  INV_X1 U7069 ( .A(n5556), .ZN(n5557) );
  XNOR2_X1 U7070 ( .A(n8991), .B(n8634), .ZN(n8901) );
  INV_X1 U7071 ( .A(n8991), .ZN(n8445) );
  NAND2_X1 U7072 ( .A1(n8887), .A2(n8605), .ZN(n8332) );
  INV_X1 U7073 ( .A(n5559), .ZN(n5563) );
  INV_X1 U7074 ( .A(n5560), .ZN(n5561) );
  NAND2_X1 U7075 ( .A1(n5561), .A2(SI_24_), .ZN(n5562) );
  INV_X1 U7076 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7952) );
  INV_X1 U7077 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7953) );
  MUX2_X1 U7078 ( .A(n7952), .B(n7953), .S(n4483), .Z(n5566) );
  INV_X1 U7079 ( .A(SI_25_), .ZN(n5565) );
  NAND2_X1 U7080 ( .A1(n5566), .A2(n5565), .ZN(n5579) );
  INV_X1 U7081 ( .A(n5566), .ZN(n5567) );
  NAND2_X1 U7082 ( .A1(n5567), .A2(SI_25_), .ZN(n5568) );
  NAND2_X1 U7083 ( .A1(n5579), .A2(n5568), .ZN(n5580) );
  NAND2_X1 U7084 ( .A1(n7950), .A2(n8297), .ZN(n5570) );
  OR2_X1 U7085 ( .A1(n5377), .A2(n7952), .ZN(n5569) );
  INV_X1 U7086 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8607) );
  NAND2_X1 U7087 ( .A1(n5571), .A2(n8607), .ZN(n5572) );
  NAND2_X1 U7088 ( .A1(n5589), .A2(n5572), .ZN(n8868) );
  INV_X1 U7089 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8869) );
  NAND2_X1 U7090 ( .A1(n5326), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5575) );
  INV_X1 U7091 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n5573) );
  OR2_X1 U7092 ( .A1(n4485), .A2(n5573), .ZN(n5574) );
  OAI211_X1 U7093 ( .C1(n8869), .C2(n5666), .A(n5575), .B(n5574), .ZN(n5576)
         );
  INV_X1 U7094 ( .A(n5576), .ZN(n5577) );
  OAI21_X1 U7095 ( .B1(n8868), .B2(n5578), .A(n5577), .ZN(n8661) );
  INV_X1 U7096 ( .A(n8661), .ZN(n8648) );
  NAND2_X1 U7097 ( .A1(n8980), .A2(n8648), .ZN(n8452) );
  INV_X1 U7098 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7973) );
  INV_X1 U7099 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7975) );
  MUX2_X1 U7100 ( .A(n7973), .B(n7975), .S(n4483), .Z(n5583) );
  INV_X1 U7101 ( .A(SI_26_), .ZN(n5582) );
  NAND2_X1 U7102 ( .A1(n5583), .A2(n5582), .ZN(n5602) );
  INV_X1 U7103 ( .A(n5583), .ZN(n5584) );
  NAND2_X1 U7104 ( .A1(n5584), .A2(SI_26_), .ZN(n5585) );
  AND2_X1 U7105 ( .A1(n5602), .A2(n5585), .ZN(n5600) );
  NAND2_X1 U7106 ( .A1(n7972), .A2(n8297), .ZN(n5587) );
  OR2_X1 U7107 ( .A1(n5377), .A2(n7973), .ZN(n5586) );
  INV_X1 U7108 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U7109 ( .A1(n5589), .A2(n8651), .ZN(n5590) );
  NAND2_X1 U7110 ( .A1(n5623), .A2(n5590), .ZN(n8847) );
  OR2_X1 U7111 ( .A1(n8847), .A2(n5578), .ZN(n5596) );
  INV_X1 U7112 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7113 ( .A1(n5663), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7114 ( .A1(n5326), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5591) );
  OAI211_X1 U7115 ( .C1(n5593), .C2(n5666), .A(n5592), .B(n5591), .ZN(n5594)
         );
  INV_X1 U7116 ( .A(n5594), .ZN(n5595) );
  NAND2_X1 U7117 ( .A1(n5596), .A2(n5595), .ZN(n8660) );
  NAND2_X1 U7118 ( .A1(n9044), .A2(n8660), .ZN(n8451) );
  INV_X1 U7119 ( .A(n8660), .ZN(n5597) );
  NAND2_X1 U7120 ( .A1(n8859), .A2(n5597), .ZN(n8454) );
  NAND2_X1 U7121 ( .A1(n9044), .A2(n5597), .ZN(n5598) );
  NAND2_X1 U7122 ( .A1(n5599), .A2(n5598), .ZN(n8831) );
  INV_X1 U7123 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8067) );
  INV_X1 U7124 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8065) );
  MUX2_X1 U7125 ( .A(n8067), .B(n8065), .S(n4483), .Z(n5605) );
  INV_X1 U7126 ( .A(SI_27_), .ZN(n5604) );
  NAND2_X1 U7127 ( .A1(n5605), .A2(n5604), .ZN(n5618) );
  INV_X1 U7128 ( .A(n5605), .ZN(n5606) );
  NAND2_X1 U7129 ( .A1(n5606), .A2(SI_27_), .ZN(n5607) );
  AND2_X1 U7130 ( .A1(n5618), .A2(n5607), .ZN(n5616) );
  NAND2_X1 U7131 ( .A1(n8064), .A2(n8297), .ZN(n5609) );
  OR2_X1 U7132 ( .A1(n5377), .A2(n8067), .ZN(n5608) );
  XNOR2_X1 U7133 ( .A(n5623), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8839) );
  NAND2_X1 U7134 ( .A1(n8839), .A2(n5668), .ZN(n5614) );
  INV_X1 U7135 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6897) );
  NAND2_X1 U7136 ( .A1(n5326), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5610) );
  OAI211_X1 U7137 ( .C1(n4485), .C2(n6897), .A(n5611), .B(n5610), .ZN(n5612)
         );
  INV_X1 U7138 ( .A(n5612), .ZN(n5613) );
  NAND2_X1 U7139 ( .A1(n5614), .A2(n5613), .ZN(n8659) );
  INV_X1 U7140 ( .A(n8970), .ZN(n8842) );
  NAND2_X1 U7141 ( .A1(n8842), .A2(n8650), .ZN(n5615) );
  MUX2_X1 U7142 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n4483), .Z(n8190) );
  INV_X1 U7143 ( .A(SI_28_), .ZN(n8191) );
  XNOR2_X1 U7144 ( .A(n8190), .B(n8191), .ZN(n8188) );
  NAND2_X1 U7145 ( .A1(n8220), .A2(n8297), .ZN(n5621) );
  INV_X1 U7146 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8117) );
  OR2_X1 U7147 ( .A1(n5377), .A2(n8117), .ZN(n5620) );
  INV_X1 U7148 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6471) );
  INV_X1 U7149 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5622) );
  OAI21_X1 U7150 ( .B1(n5623), .B2(n6471), .A(n5622), .ZN(n5624) );
  NAND2_X1 U7151 ( .A1(n8821), .A2(n5668), .ZN(n5629) );
  INV_X1 U7152 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8822) );
  NAND2_X1 U7153 ( .A1(n5663), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7154 ( .A1(n5326), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5625) );
  OAI211_X1 U7155 ( .C1(n8822), .C2(n5666), .A(n5626), .B(n5625), .ZN(n5627)
         );
  INV_X1 U7156 ( .A(n5627), .ZN(n5628) );
  NAND2_X1 U7157 ( .A1(n5629), .A2(n5628), .ZN(n8815) );
  INV_X1 U7158 ( .A(n8815), .ZN(n8461) );
  NAND2_X1 U7159 ( .A1(n8827), .A2(n8461), .ZN(n8456) );
  XNOR2_X1 U7160 ( .A(n8801), .B(n8800), .ZN(n8820) );
  NAND2_X1 U7161 ( .A1(n5632), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U7162 ( .A1(n5637), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5636) );
  INV_X1 U7163 ( .A(n8330), .ZN(n8517) );
  NAND2_X1 U7164 ( .A1(n8479), .A2(n8517), .ZN(n8524) );
  INV_X1 U7165 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5680) );
  XNOR2_X2 U7166 ( .A(n5681), .B(n5680), .ZN(n5672) );
  INV_X1 U7167 ( .A(n5672), .ZN(n5658) );
  XNOR2_X1 U7168 ( .A(n8524), .B(n5672), .ZN(n5638) );
  OR2_X1 U7169 ( .A1(n5638), .A2(n8327), .ZN(n10266) );
  AND2_X1 U7170 ( .A1(n8479), .A2(n8327), .ZN(n5639) );
  NAND2_X1 U7171 ( .A1(n5639), .A2(n5672), .ZN(n10335) );
  NAND2_X1 U7172 ( .A1(n6328), .A2(n6327), .ZN(n7196) );
  NAND2_X1 U7173 ( .A1(n8361), .A2(n7196), .ZN(n8355) );
  NAND2_X1 U7174 ( .A1(n8355), .A2(n8358), .ZN(n7273) );
  INV_X1 U7175 ( .A(n7273), .ZN(n5641) );
  INV_X1 U7176 ( .A(n8484), .ZN(n5640) );
  NAND2_X1 U7177 ( .A1(n5641), .A2(n5640), .ZN(n5642) );
  NAND2_X1 U7178 ( .A1(n5642), .A2(n8360), .ZN(n7213) );
  INV_X1 U7179 ( .A(n8487), .ZN(n8367) );
  INV_X1 U7180 ( .A(n8348), .ZN(n5643) );
  AOI21_X1 U7181 ( .B1(n7213), .B2(n8367), .A(n5643), .ZN(n8267) );
  INV_X1 U7182 ( .A(n8488), .ZN(n8266) );
  NAND2_X1 U7183 ( .A1(n8267), .A2(n8266), .ZN(n7285) );
  AND2_X1 U7184 ( .A1(n5644), .A2(n8371), .ZN(n8373) );
  NAND2_X1 U7185 ( .A1(n7285), .A2(n8373), .ZN(n5645) );
  NAND2_X1 U7186 ( .A1(n5645), .A2(n8352), .ZN(n10275) );
  XNOR2_X1 U7187 ( .A(n10321), .B(n8677), .ZN(n10287) );
  NAND2_X1 U7188 ( .A1(n10275), .A2(n10287), .ZN(n5646) );
  INV_X1 U7189 ( .A(n8677), .ZN(n8381) );
  NAND2_X1 U7190 ( .A1(n10321), .A2(n8381), .ZN(n8351) );
  NAND2_X1 U7191 ( .A1(n5646), .A2(n8351), .ZN(n7448) );
  INV_X1 U7192 ( .A(n7416), .ZN(n8496) );
  INV_X1 U7193 ( .A(n8392), .ZN(n8337) );
  NOR2_X1 U7194 ( .A1(n8496), .A2(n8337), .ZN(n5647) );
  NAND2_X1 U7195 ( .A1(n7414), .A2(n5647), .ZN(n7415) );
  AND2_X1 U7196 ( .A1(n8399), .A2(n8342), .ZN(n8404) );
  INV_X1 U7197 ( .A(n8410), .ZN(n8500) );
  AND2_X1 U7198 ( .A1(n8404), .A2(n8500), .ZN(n5650) );
  INV_X1 U7199 ( .A(n9919), .ZN(n5651) );
  NOR2_X1 U7200 ( .A1(n5651), .A2(n4914), .ZN(n5652) );
  NAND2_X1 U7201 ( .A1(n9908), .A2(n8412), .ZN(n7932) );
  INV_X1 U7202 ( .A(n7932), .ZN(n5653) );
  INV_X1 U7203 ( .A(n8414), .ZN(n8502) );
  NAND2_X1 U7204 ( .A1(n5653), .A2(n8414), .ZN(n7930) );
  NAND2_X1 U7205 ( .A1(n7930), .A2(n8416), .ZN(n7978) );
  INV_X1 U7206 ( .A(n8418), .ZN(n5654) );
  NOR2_X1 U7207 ( .A1(n8504), .A2(n5654), .ZN(n5655) );
  NOR2_X1 U7208 ( .A1(n9020), .A2(n8243), .ZN(n8425) );
  NAND2_X1 U7209 ( .A1(n9020), .A2(n8243), .ZN(n8430) );
  OR2_X1 U7210 ( .A1(n8248), .A2(n8237), .ZN(n8426) );
  NAND2_X1 U7211 ( .A1(n8248), .A2(n8237), .ZN(n8432) );
  XNOR2_X1 U7212 ( .A(n9002), .B(n8633), .ZN(n8935) );
  NAND2_X1 U7213 ( .A1(n9002), .A2(n8633), .ZN(n8437) );
  INV_X1 U7214 ( .A(n8912), .ZN(n8915) );
  INV_X1 U7215 ( .A(n8901), .ZN(n8894) );
  AND2_X1 U7216 ( .A1(n8991), .A2(n8634), .ZN(n8444) );
  INV_X1 U7217 ( .A(n5656), .ZN(n8447) );
  NOR3_X1 U7218 ( .A1(n8848), .A2(n4818), .A3(n8857), .ZN(n8850) );
  INV_X1 U7219 ( .A(n8454), .ZN(n5657) );
  NAND2_X1 U7220 ( .A1(n8834), .A2(n8833), .ZN(n8832) );
  OR2_X1 U7221 ( .A1(n8970), .A2(n8650), .ZN(n8455) );
  AOI21_X2 U7222 ( .B1(n8832), .B2(n8455), .A(n8800), .ZN(n8313) );
  AND3_X1 U7223 ( .A1(n8832), .A2(n8800), .A3(n8455), .ZN(n5659) );
  OR2_X1 U7224 ( .A1(n8479), .A2(n8330), .ZN(n8328) );
  AND2_X1 U7225 ( .A1(n6323), .A2(n8328), .ZN(n9910) );
  NOR3_X1 U7226 ( .A1(n8313), .A2(n5659), .A3(n9910), .ZN(n5670) );
  OR2_X1 U7227 ( .A1(n5672), .A2(n8330), .ZN(n6602) );
  INV_X1 U7228 ( .A(n6602), .ZN(n7111) );
  INV_X1 U7229 ( .A(n5661), .ZN(n5662) );
  NAND2_X1 U7230 ( .A1(n7111), .A2(n5662), .ZN(n8647) );
  INV_X1 U7231 ( .A(n8808), .ZN(n5669) );
  INV_X1 U7232 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8807) );
  NAND2_X1 U7233 ( .A1(n5663), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U7234 ( .A1(n5326), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5664) );
  OAI211_X1 U7235 ( .C1(n8807), .C2(n5666), .A(n5665), .B(n5664), .ZN(n5667)
         );
  AOI21_X1 U7236 ( .B1(n5669), .B2(n5668), .A(n5667), .ZN(n8314) );
  NAND2_X1 U7237 ( .A1(n7111), .A2(n5661), .ZN(n8649) );
  OAI22_X1 U7238 ( .A1(n8650), .A2(n8647), .B1(n8314), .B2(n8649), .ZN(n6451)
         );
  NOR2_X1 U7239 ( .A1(n5670), .A2(n6451), .ZN(n8830) );
  INV_X1 U7240 ( .A(n8980), .ZN(n8867) );
  NAND2_X1 U7241 ( .A1(n7263), .A2(n7240), .ZN(n7270) );
  OR2_X1 U7242 ( .A1(n7270), .A2(n7493), .ZN(n7271) );
  NAND2_X1 U7243 ( .A1(n8270), .A2(n7465), .ZN(n10288) );
  OR2_X1 U7244 ( .A1(n10288), .A2(n10321), .ZN(n10289) );
  INV_X1 U7245 ( .A(n8588), .ZN(n10336) );
  NAND2_X1 U7246 ( .A1(n10253), .A2(n10336), .ZN(n10252) );
  INV_X1 U7247 ( .A(n8060), .ZN(n7937) );
  NAND2_X1 U7248 ( .A1(n7935), .A2(n7937), .ZN(n7983) );
  INV_X1 U7249 ( .A(n5671), .ZN(n8838) );
  INV_X1 U7250 ( .A(n8295), .ZN(n8805) );
  OAI211_X1 U7251 ( .C1(n8802), .C2(n8838), .A(n8805), .B(n9922), .ZN(n8824)
         );
  NAND2_X1 U7252 ( .A1(n8830), .A2(n8824), .ZN(n5673) );
  AOI21_X1 U7253 ( .B1(n8820), .B2(n10368), .A(n5673), .ZN(n5715) );
  INV_X1 U7254 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U7255 ( .A1(n5674), .A2(n5683), .ZN(n5675) );
  OAI21_X1 U7256 ( .B1(n4504), .B2(n5675), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5677) );
  MUX2_X1 U7257 ( .A(n5677), .B(P2_IR_REG_31__SCAN_IN), .S(n5676), .Z(n5679)
         );
  NAND2_X1 U7258 ( .A1(n5679), .A2(n5686), .ZN(n7951) );
  NAND2_X1 U7259 ( .A1(n5681), .A2(n5680), .ZN(n5682) );
  NAND2_X1 U7260 ( .A1(n5682), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5703) );
  INV_X1 U7261 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U7262 ( .A1(n5703), .A2(n5702), .ZN(n5705) );
  NAND2_X1 U7263 ( .A1(n5705), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5684) );
  XNOR2_X1 U7264 ( .A(n5684), .B(n5683), .ZN(n7826) );
  XNOR2_X1 U7265 ( .A(n7826), .B(P2_B_REG_SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7266 ( .A1(n7951), .A2(n5685), .ZN(n5690) );
  NAND2_X1 U7267 ( .A1(n5686), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5688) );
  XNOR2_X1 U7268 ( .A(n5688), .B(n5687), .ZN(n7974) );
  INV_X1 U7269 ( .A(n7974), .ZN(n5689) );
  INV_X1 U7270 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10311) );
  AND2_X1 U7271 ( .A1(n7974), .A2(n7951), .ZN(n10312) );
  AOI21_X1 U7272 ( .B1(n10297), .B2(n10311), .A(n10312), .ZN(n6425) );
  NOR4_X1 U7273 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5694) );
  NOR4_X1 U7274 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5693) );
  NOR4_X1 U7275 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n5692) );
  NOR4_X1 U7276 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n5691) );
  NAND4_X1 U7277 ( .A1(n5694), .A2(n5693), .A3(n5692), .A4(n5691), .ZN(n5700)
         );
  NOR2_X1 U7278 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .ZN(
        n5698) );
  NOR4_X1 U7279 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5697) );
  NOR4_X1 U7280 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n5696) );
  NOR4_X1 U7281 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5695) );
  NAND4_X1 U7282 ( .A1(n5698), .A2(n5697), .A3(n5696), .A4(n5695), .ZN(n5699)
         );
  OAI21_X1 U7283 ( .B1(n5700), .B2(n5699), .A(n10297), .ZN(n6424) );
  OR2_X1 U7284 ( .A1(n7974), .A2(n7951), .ZN(n5701) );
  OR2_X1 U7285 ( .A1(n7826), .A2(n5701), .ZN(n7114) );
  OR2_X1 U7286 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  NAND2_X1 U7287 ( .A1(n5705), .A2(n5704), .ZN(n6603) );
  NAND2_X1 U7288 ( .A1(n7114), .A2(n10313), .ZN(n7112) );
  INV_X1 U7289 ( .A(n8327), .ZN(n8856) );
  NAND2_X1 U7290 ( .A1(n8479), .A2(n8856), .ZN(n6448) );
  NAND2_X1 U7291 ( .A1(n7111), .A2(n6448), .ZN(n6454) );
  INV_X1 U7292 ( .A(n6454), .ZN(n5706) );
  OR2_X1 U7293 ( .A1(n7112), .A2(n5706), .ZN(n8525) );
  NAND2_X1 U7294 ( .A1(n9922), .A2(n8327), .ZN(n6452) );
  INV_X1 U7295 ( .A(n6452), .ZN(n5707) );
  NOR2_X1 U7296 ( .A1(n8525), .A2(n5707), .ZN(n5708) );
  NAND2_X1 U7297 ( .A1(n6424), .A2(n5708), .ZN(n5709) );
  OR2_X1 U7298 ( .A1(n6425), .A2(n5709), .ZN(n5714) );
  INV_X1 U7299 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10308) );
  AND2_X1 U7300 ( .A1(n10297), .A2(n10308), .ZN(n5710) );
  AND2_X1 U7301 ( .A1(n7826), .A2(n7974), .ZN(n10309) );
  INV_X2 U7302 ( .A(n10380), .ZN(n10382) );
  NAND2_X1 U7303 ( .A1(n5711), .A2(n6448), .ZN(n10362) );
  INV_X1 U7304 ( .A(n10362), .ZN(n9026) );
  NAND2_X1 U7305 ( .A1(n10382), .A2(n9026), .ZN(n9017) );
  INV_X2 U7306 ( .A(n10370), .ZN(n10371) );
  NAND2_X1 U7307 ( .A1(n10371), .A2(n9026), .ZN(n9061) );
  NAND2_X1 U7308 ( .A1(n8827), .A2(n5716), .ZN(n5717) );
  NAND4_X1 U7309 ( .A1(n5720), .A2(n5950), .A3(n5924), .A4(n5719), .ZN(n5721)
         );
  INV_X1 U7310 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5723) );
  NOR2_X1 U7311 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5725) );
  INV_X1 U7312 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5724) );
  NAND2_X1 U7313 ( .A1(n5725), .A2(n5724), .ZN(n5730) );
  NOR2_X1 U7314 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5729) );
  NOR2_X1 U7315 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5728) );
  NOR2_X1 U7316 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5727) );
  NAND2_X1 U7317 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5732) );
  INV_X1 U7318 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U7319 ( .A1(n7779), .A2(n9214), .ZN(n5736) );
  OR2_X1 U7320 ( .A1(n5822), .A2(n7782), .ZN(n5735) );
  INV_X1 U7321 ( .A(n9779), .ZN(n9633) );
  INV_X1 U7322 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n7039) );
  INV_X1 U7323 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5737) );
  INV_X1 U7324 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5781) );
  INV_X1 U7325 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6940) );
  NAND2_X1 U7326 ( .A1(n5776), .A2(n5740), .ZN(n5779) );
  NAND2_X1 U7327 ( .A1(n5743), .A2(n5742), .ZN(n5741) );
  XNOR2_X1 U7328 ( .A(n5743), .B(n5742), .ZN(n5775) );
  INV_X1 U7329 ( .A(n6041), .ZN(n5744) );
  NAND2_X1 U7330 ( .A1(n5059), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5745) );
  OR2_X1 U7331 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5750) );
  OR2_X1 U7332 ( .A1(n5750), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U7333 ( .A1(n4506), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5752) );
  XNOR2_X1 U7334 ( .A(n5752), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6275) );
  NAND2_X1 U7335 ( .A1(n5753), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5754) );
  MUX2_X1 U7336 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5754), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5755) );
  NAND2_X1 U7337 ( .A1(n7625), .A2(n6543), .ZN(n5815) );
  INV_X2 U7338 ( .A(n5815), .ZN(n5802) );
  INV_X2 U7339 ( .A(n5802), .ZN(n6236) );
  NOR3_X1 U7340 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .A3(
        P1_IR_REG_29__SCAN_IN), .ZN(n5760) );
  NAND2_X1 U7341 ( .A1(n5759), .A2(n5760), .ZN(n9848) );
  NAND2_X1 U7342 ( .A1(n9848), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5761) );
  INV_X1 U7343 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9849) );
  XNOR2_X2 U7344 ( .A(n5761), .B(n9849), .ZN(n9855) );
  NAND2_X1 U7345 ( .A1(n5915), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5943) );
  INV_X1 U7346 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5971) );
  INV_X1 U7347 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6029) );
  INV_X1 U7348 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6045) );
  INV_X1 U7349 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7350 ( .A1(n6083), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6102) );
  INV_X1 U7351 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9111) );
  INV_X1 U7352 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6877) );
  NAND2_X1 U7353 ( .A1(n6127), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6128) );
  INV_X1 U7354 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9160) );
  NAND2_X1 U7355 ( .A1(n6190), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6209) );
  OR2_X1 U7356 ( .A1(n6190), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U7357 ( .A1(n6209), .A2(n5762), .ZN(n9630) );
  OR2_X1 U7358 ( .A1(n6527), .A2(n9630), .ZN(n5769) );
  NAND2_X1 U7359 ( .A1(n4482), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U7360 ( .A1(n5764), .A2(n9855), .ZN(n5917) );
  NAND2_X1 U7361 ( .A1(n8555), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5767) );
  NAND2_X4 U7362 ( .A1(n5765), .A2(n9855), .ZN(n8559) );
  NAND2_X1 U7363 ( .A1(n6245), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5766) );
  NAND4_X1 U7364 ( .A1(n5769), .A2(n5768), .A3(n5767), .A4(n5766), .ZN(n9477)
         );
  INV_X1 U7365 ( .A(n9477), .ZN(n9649) );
  INV_X1 U7366 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5771) );
  NAND2_X1 U7367 ( .A1(n5772), .A2(n5771), .ZN(n5773) );
  XNOR2_X2 U7368 ( .A(n5774), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9209) );
  INV_X1 U7369 ( .A(n5776), .ZN(n5777) );
  NAND2_X1 U7370 ( .A1(n5777), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5778) );
  MUX2_X1 U7371 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5778), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5780) );
  NAND2_X1 U7372 ( .A1(n5780), .A2(n5779), .ZN(n9532) );
  AND2_X1 U7373 ( .A1(n5775), .A2(n9532), .ZN(n6292) );
  NAND2_X1 U7374 ( .A1(n6282), .A2(n6292), .ZN(n7627) );
  INV_X1 U7375 ( .A(n5923), .ZN(n6235) );
  OAI22_X1 U7376 ( .A1(n9633), .A2(n6236), .B1(n9649), .B2(n6235), .ZN(n9077)
         );
  NAND2_X1 U7377 ( .A1(n7264), .A2(n9214), .ZN(n5785) );
  OAI21_X1 U7378 ( .B1(n6098), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5782) );
  OR2_X1 U7379 ( .A1(n5782), .A2(n5781), .ZN(n5783) );
  NAND2_X1 U7380 ( .A1(n5782), .A2(n5781), .ZN(n6123) );
  AND2_X1 U7381 ( .A1(n5783), .A2(n6123), .ZN(n9513) );
  AOI22_X1 U7382 ( .A1(n6137), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9986), .B2(
        n9513), .ZN(n5784) );
  INV_X1 U7383 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9498) );
  OR2_X1 U7384 ( .A1(n8559), .A2(n9498), .ZN(n5790) );
  NAND2_X1 U7385 ( .A1(n4482), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5789) );
  AND2_X1 U7386 ( .A1(n6104), .A2(n6877), .ZN(n5786) );
  NOR2_X1 U7387 ( .A1(n6127), .A2(n5786), .ZN(n9739) );
  NAND2_X1 U7388 ( .A1(n5829), .A2(n9739), .ZN(n5788) );
  NAND2_X1 U7389 ( .A1(n8555), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5787) );
  NAND4_X1 U7390 ( .A1(n5790), .A2(n5789), .A3(n5788), .A4(n5787), .ZN(n9719)
         );
  AOI22_X1 U7391 ( .A1(n9809), .A2(n4490), .B1(n6514), .B2(n9719), .ZN(n6122)
         );
  NAND2_X1 U7392 ( .A1(n9809), .A2(n4486), .ZN(n5792) );
  NAND2_X1 U7393 ( .A1(n9719), .A2(n4490), .ZN(n5791) );
  NAND2_X1 U7394 ( .A1(n5792), .A2(n5791), .ZN(n5793) );
  NAND2_X1 U7395 ( .A1(n9209), .A2(n9532), .ZN(n7626) );
  NAND2_X1 U7396 ( .A1(n7626), .A2(n5770), .ZN(n5813) );
  XNOR2_X1 U7397 ( .A(n5793), .B(n7574), .ZN(n6120) );
  INV_X1 U7398 ( .A(n6120), .ZN(n6121) );
  NAND2_X1 U7399 ( .A1(n8555), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5795) );
  INV_X1 U7400 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9991) );
  NAND2_X1 U7401 ( .A1(n5880), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7402 ( .A1(n9492), .A2(n4484), .ZN(n5801) );
  INV_X1 U7403 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5796) );
  AND2_X1 U7404 ( .A1(n5798), .A2(n5797), .ZN(n9860) );
  MUX2_X1 U7405 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9860), .S(n6545), .Z(n7600) );
  NAND2_X1 U7406 ( .A1(n7600), .A2(n4487), .ZN(n5803) );
  NAND2_X1 U7407 ( .A1(n5805), .A2(n5804), .ZN(n5806) );
  NAND2_X1 U7408 ( .A1(n7203), .A2(n5806), .ZN(n5808) );
  INV_X1 U7409 ( .A(n5806), .ZN(n7204) );
  NAND2_X1 U7410 ( .A1(n7204), .A2(n5813), .ZN(n5807) );
  NAND2_X1 U7411 ( .A1(n5808), .A2(n5807), .ZN(n5817) );
  NAND2_X1 U7412 ( .A1(n5880), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7577) );
  INV_X1 U7413 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5809) );
  OR2_X1 U7414 ( .A1(n5917), .A2(n5809), .ZN(n7578) );
  INV_X1 U7415 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6566) );
  INV_X1 U7416 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7639) );
  OR2_X1 U7417 ( .A1(n6301), .A2(n7639), .ZN(n7576) );
  INV_X1 U7418 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7419 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5810) );
  XNOR2_X1 U7420 ( .A(n5810), .B(n5811), .ZN(n6721) );
  INV_X1 U7421 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6594) );
  NAND2_X1 U7422 ( .A1(n7641), .A2(n4486), .ZN(n5812) );
  OAI21_X1 U7423 ( .B1(n7679), .B2(n5815), .A(n5812), .ZN(n5814) );
  INV_X2 U7424 ( .A(n5813), .ZN(n6252) );
  XNOR2_X1 U7425 ( .A(n5814), .B(n6252), .ZN(n5818) );
  NAND2_X1 U7426 ( .A1(n5817), .A2(n5818), .ZN(n7393) );
  NAND2_X1 U7427 ( .A1(n7641), .A2(n5802), .ZN(n5816) );
  OAI21_X1 U7428 ( .B1(n7679), .B2(n6235), .A(n5816), .ZN(n7395) );
  NAND2_X1 U7429 ( .A1(n7393), .A2(n7395), .ZN(n5821) );
  INV_X1 U7430 ( .A(n5817), .ZN(n5820) );
  INV_X1 U7431 ( .A(n5818), .ZN(n5819) );
  NAND2_X1 U7432 ( .A1(n5820), .A2(n5819), .ZN(n7394) );
  OR2_X1 U7433 ( .A1(n5822), .A2(n6590), .ZN(n5828) );
  OR2_X1 U7434 ( .A1(n5823), .A2(n6589), .ZN(n5827) );
  OR2_X1 U7435 ( .A1(n5824), .A2(n5731), .ZN(n5825) );
  INV_X1 U7436 ( .A(n10014), .ZN(n6588) );
  OR2_X1 U7437 ( .A1(n6545), .A2(n6588), .ZN(n5826) );
  AND3_X2 U7438 ( .A1(n5828), .A2(n5827), .A3(n5826), .ZN(n10161) );
  NAND2_X1 U7439 ( .A1(n8555), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5831) );
  INV_X1 U7440 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10220) );
  NAND2_X1 U7441 ( .A1(n9490), .A2(n5802), .ZN(n5832) );
  OAI21_X1 U7442 ( .B1(n10161), .B2(n6216), .A(n5832), .ZN(n5833) );
  XNOR2_X1 U7443 ( .A(n5833), .B(n6252), .ZN(n5838) );
  OR2_X1 U7444 ( .A1(n10161), .A2(n6236), .ZN(n5835) );
  NAND2_X1 U7445 ( .A1(n9490), .A2(n5923), .ZN(n5834) );
  NAND2_X1 U7446 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  XNOR2_X1 U7447 ( .A(n5838), .B(n5836), .ZN(n9167) );
  NAND2_X1 U7448 ( .A1(n9165), .A2(n9167), .ZN(n9166) );
  INV_X1 U7449 ( .A(n5836), .ZN(n5837) );
  NAND2_X1 U7450 ( .A1(n5838), .A2(n5837), .ZN(n5839) );
  OR2_X1 U7451 ( .A1(n5822), .A2(n8253), .ZN(n5843) );
  OR2_X1 U7452 ( .A1(n5823), .A2(n8255), .ZN(n5842) );
  NAND2_X1 U7453 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4516), .ZN(n5840) );
  XNOR2_X1 U7454 ( .A(n5840), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6565) );
  INV_X1 U7455 ( .A(n6565), .ZN(n9862) );
  OR2_X1 U7456 ( .A1(n6545), .A2(n9862), .ZN(n5841) );
  OR2_X1 U7457 ( .A1(n6527), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U7458 ( .A1(n4482), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5846) );
  NAND2_X1 U7459 ( .A1(n8555), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U7460 ( .A1(n6245), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U7461 ( .A1(n7846), .A2(n5802), .ZN(n5848) );
  OAI21_X1 U7462 ( .B1(n10167), .B2(n6216), .A(n5848), .ZN(n5849) );
  XNOR2_X1 U7463 ( .A(n5849), .B(n6252), .ZN(n5852) );
  OR2_X1 U7464 ( .A1(n10167), .A2(n5815), .ZN(n5851) );
  NAND2_X1 U7465 ( .A1(n7846), .A2(n6514), .ZN(n5850) );
  AND2_X1 U7466 ( .A1(n5851), .A2(n5850), .ZN(n5853) );
  AND2_X1 U7467 ( .A1(n5852), .A2(n5853), .ZN(n7292) );
  INV_X1 U7468 ( .A(n5852), .ZN(n5855) );
  INV_X1 U7469 ( .A(n5853), .ZN(n5854) );
  NAND2_X1 U7470 ( .A1(n5855), .A2(n5854), .ZN(n7293) );
  OAI21_X1 U7471 ( .B1(n7296), .B2(n7292), .A(n7293), .ZN(n9138) );
  INV_X1 U7472 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6596) );
  OR2_X1 U7473 ( .A1(n5822), .A2(n6596), .ZN(n5861) );
  OR2_X1 U7474 ( .A1(n5823), .A2(n5856), .ZN(n5860) );
  NAND2_X1 U7475 ( .A1(n5857), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5858) );
  XNOR2_X1 U7476 ( .A(n5858), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10028) );
  INV_X1 U7477 ( .A(n10028), .ZN(n6595) );
  OR2_X1 U7478 ( .A1(n4489), .A2(n6595), .ZN(n5859) );
  NAND2_X1 U7479 ( .A1(n6245), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U7480 ( .A1(n4482), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5865) );
  NOR2_X1 U7481 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5862) );
  NOR2_X1 U7482 ( .A1(n5892), .A2(n5862), .ZN(n9139) );
  NAND2_X1 U7483 ( .A1(n5829), .A2(n9139), .ZN(n5864) );
  NAND2_X1 U7484 ( .A1(n8555), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5863) );
  NAND4_X1 U7485 ( .A1(n5866), .A2(n5865), .A3(n5864), .A4(n5863), .ZN(n9489)
         );
  NAND2_X1 U7486 ( .A1(n9489), .A2(n6255), .ZN(n5867) );
  OAI21_X1 U7487 ( .B1(n10172), .B2(n6216), .A(n5867), .ZN(n5868) );
  XNOR2_X1 U7488 ( .A(n5868), .B(n6252), .ZN(n5871) );
  OR2_X1 U7489 ( .A1(n10172), .A2(n6236), .ZN(n5870) );
  NAND2_X1 U7490 ( .A1(n9489), .A2(n6514), .ZN(n5869) );
  NAND2_X1 U7491 ( .A1(n5870), .A2(n5869), .ZN(n5872) );
  XNOR2_X1 U7492 ( .A(n5871), .B(n5872), .ZN(n9137) );
  NAND2_X1 U7493 ( .A1(n9138), .A2(n9137), .ZN(n9136) );
  INV_X1 U7494 ( .A(n5871), .ZN(n5873) );
  NAND2_X1 U7495 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  INV_X1 U7496 ( .A(n7534), .ZN(n5908) );
  OR2_X1 U7497 ( .A1(n5823), .A2(n8261), .ZN(n5879) );
  OR2_X1 U7498 ( .A1(n5822), .A2(n8258), .ZN(n5878) );
  NOR2_X1 U7499 ( .A1(n5875), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5925) );
  OR2_X1 U7500 ( .A1(n5925), .A2(n5731), .ZN(n5876) );
  XNOR2_X1 U7501 ( .A(n5876), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6732) );
  INV_X1 U7502 ( .A(n6732), .ZN(n8259) );
  OR2_X1 U7503 ( .A1(n6545), .A2(n8259), .ZN(n5877) );
  NAND2_X1 U7504 ( .A1(n6245), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U7505 ( .A1(n4482), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5885) );
  AND2_X1 U7506 ( .A1(n5891), .A2(n5881), .ZN(n5882) );
  NOR2_X1 U7507 ( .A1(n5915), .A2(n5882), .ZN(n7541) );
  NAND2_X1 U7508 ( .A1(n5829), .A2(n7541), .ZN(n5884) );
  NAND2_X1 U7509 ( .A1(n8555), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5883) );
  NAND4_X1 U7510 ( .A1(n5886), .A2(n5885), .A3(n5884), .A4(n5883), .ZN(n9487)
         );
  NAND2_X1 U7511 ( .A1(n9487), .A2(n6255), .ZN(n5887) );
  OAI21_X1 U7512 ( .B1(n7602), .B2(n6216), .A(n5887), .ZN(n5888) );
  XNOR2_X1 U7513 ( .A(n5888), .B(n7574), .ZN(n7537) );
  OR2_X1 U7514 ( .A1(n7602), .A2(n6236), .ZN(n5890) );
  NAND2_X1 U7515 ( .A1(n9487), .A2(n6514), .ZN(n5889) );
  NAND2_X1 U7516 ( .A1(n5890), .A2(n5889), .ZN(n7536) );
  AND2_X1 U7517 ( .A1(n7537), .A2(n7536), .ZN(n5909) );
  OAI21_X1 U7518 ( .B1(n5892), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5891), .ZN(
        n7698) );
  OR2_X1 U7519 ( .A1(n6301), .A2(n7698), .ZN(n5896) );
  NAND2_X1 U7520 ( .A1(n6245), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U7521 ( .A1(n4482), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7522 ( .A1(n8555), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5893) );
  NAND4_X1 U7523 ( .A1(n5896), .A2(n5895), .A3(n5894), .A4(n5893), .ZN(n9488)
         );
  NAND2_X1 U7524 ( .A1(n9488), .A2(n6255), .ZN(n5903) );
  NAND2_X1 U7525 ( .A1(n5875), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5897) );
  MUX2_X1 U7526 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5897), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5899) );
  INV_X1 U7527 ( .A(n5925), .ZN(n5898) );
  INV_X1 U7528 ( .A(n6563), .ZN(n10035) );
  OR2_X1 U7529 ( .A1(n5822), .A2(n6592), .ZN(n5901) );
  OR2_X1 U7530 ( .A1(n5823), .A2(n6591), .ZN(n5900) );
  OAI211_X1 U7531 ( .C1(n4489), .C2(n10035), .A(n5901), .B(n5900), .ZN(n7705)
         );
  NAND2_X1 U7532 ( .A1(n7705), .A2(n4487), .ZN(n5902) );
  NAND2_X1 U7533 ( .A1(n5903), .A2(n5902), .ZN(n5904) );
  XNOR2_X1 U7534 ( .A(n5904), .B(n7574), .ZN(n7535) );
  NAND2_X1 U7535 ( .A1(n9488), .A2(n6514), .ZN(n5906) );
  NAND2_X1 U7536 ( .A1(n7705), .A2(n6255), .ZN(n5905) );
  NAND2_X1 U7537 ( .A1(n5906), .A2(n5905), .ZN(n5910) );
  AND2_X1 U7538 ( .A1(n7535), .A2(n5910), .ZN(n5907) );
  NAND2_X1 U7539 ( .A1(n5908), .A2(n5044), .ZN(n5936) );
  INV_X1 U7540 ( .A(n5909), .ZN(n5914) );
  INV_X1 U7541 ( .A(n7535), .ZN(n7428) );
  INV_X1 U7542 ( .A(n5910), .ZN(n7430) );
  AND2_X1 U7543 ( .A1(n7428), .A2(n7430), .ZN(n5913) );
  INV_X1 U7544 ( .A(n7536), .ZN(n5912) );
  INV_X1 U7545 ( .A(n7537), .ZN(n5911) );
  AOI22_X1 U7546 ( .A1(n5914), .A2(n5913), .B1(n5912), .B2(n5911), .ZN(n5934)
         );
  NAND2_X1 U7547 ( .A1(n5936), .A2(n5934), .ZN(n7437) );
  INV_X1 U7548 ( .A(n7437), .ZN(n5931) );
  NAND2_X1 U7549 ( .A1(n6245), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5922) );
  INV_X1 U7550 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7668) );
  OR2_X1 U7551 ( .A1(n6296), .A2(n7668), .ZN(n5921) );
  OR2_X1 U7552 ( .A1(n5915), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U7553 ( .A1(n5943), .A2(n5916), .ZN(n7667) );
  OR2_X1 U7554 ( .A1(n6527), .A2(n7667), .ZN(n5920) );
  INV_X1 U7555 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5918) );
  OR2_X1 U7556 ( .A1(n6627), .A2(n5918), .ZN(n5919) );
  INV_X1 U7557 ( .A(n7714), .ZN(n9486) );
  NAND2_X1 U7558 ( .A1(n5925), .A2(n5924), .ZN(n5949) );
  NAND2_X1 U7559 ( .A1(n5949), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5926) );
  XNOR2_X1 U7560 ( .A(n5926), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6573) );
  INV_X1 U7561 ( .A(n6573), .ZN(n6706) );
  OR2_X1 U7562 ( .A1(n5823), .A2(n6599), .ZN(n5928) );
  INV_X1 U7563 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6598) );
  OR2_X1 U7564 ( .A1(n5822), .A2(n6598), .ZN(n5927) );
  OAI211_X1 U7565 ( .C1(n4489), .C2(n6706), .A(n5928), .B(n5927), .ZN(n7672)
         );
  AND2_X1 U7566 ( .A1(n7672), .A2(n4490), .ZN(n5929) );
  AOI21_X1 U7567 ( .B1(n9486), .B2(n6514), .A(n5929), .ZN(n7438) );
  INV_X1 U7568 ( .A(n7438), .ZN(n5930) );
  NAND2_X1 U7569 ( .A1(n5931), .A2(n5930), .ZN(n5941) );
  NAND2_X1 U7570 ( .A1(n7672), .A2(n4486), .ZN(n5932) );
  OAI21_X1 U7571 ( .B1(n7714), .B2(n6236), .A(n5932), .ZN(n5933) );
  XNOR2_X1 U7572 ( .A(n5933), .B(n7574), .ZN(n7439) );
  AND2_X1 U7573 ( .A1(n5934), .A2(n7439), .ZN(n5935) );
  NAND2_X1 U7574 ( .A1(n5936), .A2(n5935), .ZN(n5939) );
  INV_X1 U7575 ( .A(n7439), .ZN(n5937) );
  OR2_X1 U7576 ( .A1(n5937), .A2(n7438), .ZN(n5938) );
  AND2_X1 U7577 ( .A1(n5939), .A2(n5938), .ZN(n5940) );
  NAND2_X1 U7578 ( .A1(n6245), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5948) );
  INV_X1 U7579 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7726) );
  OR2_X1 U7580 ( .A1(n6296), .A2(n7726), .ZN(n5947) );
  INV_X1 U7581 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5942) );
  OR2_X1 U7582 ( .A1(n6627), .A2(n5942), .ZN(n5946) );
  NAND2_X1 U7583 ( .A1(n5943), .A2(n7004), .ZN(n5944) );
  NAND2_X1 U7584 ( .A1(n5972), .A2(n5944), .ZN(n7725) );
  OR2_X1 U7585 ( .A1(n6301), .A2(n7725), .ZN(n5945) );
  NAND2_X1 U7586 ( .A1(n5952), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5951) );
  MUX2_X1 U7587 ( .A(n5951), .B(P1_IR_REG_31__SCAN_IN), .S(n5950), .Z(n5953)
         );
  NAND2_X1 U7588 ( .A1(n5953), .A2(n5964), .ZN(n10049) );
  OR2_X1 U7589 ( .A1(n5822), .A2(n6606), .ZN(n5955) );
  OR2_X1 U7590 ( .A1(n5823), .A2(n6607), .ZN(n5954) );
  OAI211_X1 U7591 ( .C1(n6545), .C2(n10049), .A(n5955), .B(n5954), .ZN(n7741)
         );
  NAND2_X1 U7592 ( .A1(n7741), .A2(n4486), .ZN(n5956) );
  OAI21_X1 U7593 ( .B1(n7745), .B2(n6236), .A(n5956), .ZN(n5957) );
  XNOR2_X1 U7594 ( .A(n5957), .B(n6252), .ZN(n7553) );
  AND2_X1 U7595 ( .A1(n7741), .A2(n4490), .ZN(n5958) );
  AOI21_X1 U7596 ( .B1(n9485), .B2(n6514), .A(n5958), .ZN(n7552) );
  NAND2_X1 U7597 ( .A1(n7553), .A2(n7552), .ZN(n5959) );
  INV_X1 U7598 ( .A(n7553), .ZN(n5961) );
  INV_X1 U7599 ( .A(n7552), .ZN(n5960) );
  NAND2_X1 U7600 ( .A1(n5961), .A2(n5960), .ZN(n5962) );
  NAND2_X1 U7601 ( .A1(n5964), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5965) );
  MUX2_X1 U7602 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5965), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n5966) );
  INV_X1 U7603 ( .A(n5966), .ZN(n5968) );
  NOR2_X1 U7604 ( .A1(n5968), .A2(n5967), .ZN(n6741) );
  INV_X1 U7605 ( .A(n6741), .ZN(n6613) );
  NAND2_X1 U7606 ( .A1(n6609), .A2(n9214), .ZN(n5970) );
  OR2_X1 U7607 ( .A1(n5822), .A2(n6611), .ZN(n5969) );
  NAND2_X1 U7608 ( .A1(n7881), .A2(n4486), .ZN(n5979) );
  NAND2_X1 U7609 ( .A1(n4482), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7610 ( .A1(n8555), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5976) );
  AND2_X1 U7611 ( .A1(n5972), .A2(n5971), .ZN(n5973) );
  NOR2_X1 U7612 ( .A1(n5996), .A2(n5973), .ZN(n7749) );
  NAND2_X1 U7613 ( .A1(n5829), .A2(n7749), .ZN(n5975) );
  NAND2_X1 U7614 ( .A1(n6245), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5974) );
  NAND4_X1 U7615 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .ZN(n9484)
         );
  NAND2_X1 U7616 ( .A1(n9484), .A2(n4490), .ZN(n5978) );
  NAND2_X1 U7617 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  XNOR2_X1 U7618 ( .A(n5980), .B(n6252), .ZN(n5983) );
  NAND2_X1 U7619 ( .A1(n7881), .A2(n4490), .ZN(n5982) );
  NAND2_X1 U7620 ( .A1(n9484), .A2(n6514), .ZN(n5981) );
  AND2_X1 U7621 ( .A1(n5982), .A2(n5981), .ZN(n5984) );
  NAND2_X1 U7622 ( .A1(n5983), .A2(n5984), .ZN(n5989) );
  INV_X1 U7623 ( .A(n5983), .ZN(n5986) );
  INV_X1 U7624 ( .A(n5984), .ZN(n5985) );
  NAND2_X1 U7625 ( .A1(n5986), .A2(n5985), .ZN(n5987) );
  NAND2_X1 U7626 ( .A1(n5989), .A2(n5987), .ZN(n7817) );
  NAND2_X1 U7627 ( .A1(n6614), .A2(n9214), .ZN(n5995) );
  NOR2_X1 U7628 ( .A1(n5967), .A2(n5731), .ZN(n5990) );
  MUX2_X1 U7629 ( .A(n5731), .B(n5990), .S(P1_IR_REG_10__SCAN_IN), .Z(n5993)
         );
  OR2_X1 U7630 ( .A1(n5993), .A2(n5992), .ZN(n6742) );
  INV_X1 U7631 ( .A(n6742), .ZN(n6761) );
  AOI22_X1 U7632 ( .A1(n6137), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9986), .B2(
        n6761), .ZN(n5994) );
  NAND2_X1 U7633 ( .A1(n7908), .A2(n4487), .ZN(n6003) );
  NOR2_X1 U7634 ( .A1(n5996), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5997) );
  OR2_X1 U7635 ( .A1(n6011), .A2(n5997), .ZN(n7891) );
  OR2_X1 U7636 ( .A1(n6301), .A2(n7891), .ZN(n6001) );
  NAND2_X1 U7637 ( .A1(n4482), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7638 ( .A1(n8555), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U7639 ( .A1(n6245), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5998) );
  NAND4_X1 U7640 ( .A1(n6001), .A2(n6000), .A3(n5999), .A4(n5998), .ZN(n7899)
         );
  NAND2_X1 U7641 ( .A1(n7899), .A2(n4490), .ZN(n6002) );
  NAND2_X1 U7642 ( .A1(n6003), .A2(n6002), .ZN(n6004) );
  XNOR2_X1 U7643 ( .A(n6004), .B(n6252), .ZN(n6006) );
  AOI22_X1 U7644 ( .A1(n7908), .A2(n4490), .B1(n6514), .B2(n7899), .ZN(n6005)
         );
  OR2_X1 U7645 ( .A1(n6006), .A2(n6005), .ZN(n7830) );
  AND2_X1 U7646 ( .A1(n6006), .A2(n6005), .ZN(n7831) );
  NAND2_X1 U7647 ( .A1(n6618), .A2(n9214), .ZN(n6009) );
  OR2_X1 U7648 ( .A1(n5992), .A2(n5731), .ZN(n6007) );
  XNOR2_X1 U7649 ( .A(n6007), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7253) );
  AOI22_X1 U7650 ( .A1(n6137), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9986), .B2(
        n7253), .ZN(n6008) );
  NAND2_X1 U7651 ( .A1(n4482), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6016) );
  INV_X1 U7652 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6010) );
  OR2_X1 U7653 ( .A1(n8559), .A2(n6010), .ZN(n6015) );
  OR2_X1 U7654 ( .A1(n6011), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U7655 ( .A1(n6030), .A2(n6012), .ZN(n9947) );
  OR2_X1 U7656 ( .A1(n6527), .A2(n9947), .ZN(n6014) );
  OR2_X1 U7657 ( .A1(n6627), .A2(n7915), .ZN(n6013) );
  OAI22_X1 U7658 ( .A1(n9952), .A2(n6216), .B1(n8049), .B2(n6236), .ZN(n6017)
         );
  XNOR2_X1 U7659 ( .A(n6017), .B(n6252), .ZN(n6020) );
  OR2_X1 U7660 ( .A1(n9952), .A2(n6236), .ZN(n6019) );
  NAND2_X1 U7661 ( .A1(n5030), .A2(n6514), .ZN(n6018) );
  NAND2_X1 U7662 ( .A1(n6019), .A2(n6018), .ZN(n6021) );
  XNOR2_X1 U7663 ( .A(n6020), .B(n6021), .ZN(n7923) );
  INV_X1 U7664 ( .A(n6020), .ZN(n6022) );
  NAND2_X1 U7665 ( .A1(n6022), .A2(n6021), .ZN(n6023) );
  NAND2_X1 U7666 ( .A1(n6621), .A2(n9214), .ZN(n6027) );
  NAND2_X1 U7667 ( .A1(n6024), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6025) );
  XNOR2_X1 U7668 ( .A(n6025), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7791) );
  AOI22_X1 U7669 ( .A1(n6137), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9986), .B2(
        n7791), .ZN(n6026) );
  NAND2_X1 U7670 ( .A1(n9972), .A2(n4487), .ZN(n6038) );
  NAND2_X1 U7671 ( .A1(n4482), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6036) );
  INV_X1 U7672 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6028) );
  OR2_X1 U7673 ( .A1(n8559), .A2(n6028), .ZN(n6035) );
  NAND2_X1 U7674 ( .A1(n6030), .A2(n6029), .ZN(n6031) );
  NAND2_X1 U7675 ( .A1(n6046), .A2(n6031), .ZN(n8048) );
  OR2_X1 U7676 ( .A1(n6301), .A2(n8048), .ZN(n6034) );
  INV_X1 U7677 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n6032) );
  OR2_X1 U7678 ( .A1(n6627), .A2(n6032), .ZN(n6033) );
  INV_X1 U7679 ( .A(n7990), .ZN(n9483) );
  NAND2_X1 U7680 ( .A1(n9483), .A2(n4490), .ZN(n6037) );
  NAND2_X1 U7681 ( .A1(n6038), .A2(n6037), .ZN(n6039) );
  XNOR2_X1 U7682 ( .A(n6039), .B(n6252), .ZN(n6059) );
  NOR2_X1 U7683 ( .A1(n7990), .A2(n6235), .ZN(n6040) );
  AOI21_X1 U7684 ( .B1(n9972), .B2(n4490), .A(n6040), .ZN(n6058) );
  XNOR2_X1 U7685 ( .A(n6059), .B(n6058), .ZN(n8045) );
  NAND2_X1 U7686 ( .A1(n6661), .A2(n9214), .ZN(n6044) );
  NAND2_X1 U7687 ( .A1(n6041), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6042) );
  XNOR2_X1 U7688 ( .A(n6042), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10066) );
  AOI22_X1 U7689 ( .A1(n6137), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9986), .B2(
        n10066), .ZN(n6043) );
  NAND2_X1 U7690 ( .A1(n9825), .A2(n4487), .ZN(n6053) );
  NAND2_X1 U7691 ( .A1(n6046), .A2(n6045), .ZN(n6047) );
  NAND2_X1 U7692 ( .A1(n6069), .A2(n6047), .ZN(n8168) );
  OR2_X1 U7693 ( .A1(n6527), .A2(n8168), .ZN(n6051) );
  NAND2_X1 U7694 ( .A1(n4482), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7695 ( .A1(n8555), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7696 ( .A1(n6245), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6048) );
  NAND4_X1 U7697 ( .A1(n6051), .A2(n6050), .A3(n6049), .A4(n6048), .ZN(n9482)
         );
  NAND2_X1 U7698 ( .A1(n9482), .A2(n4490), .ZN(n6052) );
  NAND2_X1 U7699 ( .A1(n6053), .A2(n6052), .ZN(n6054) );
  XNOR2_X1 U7700 ( .A(n6054), .B(n6252), .ZN(n8034) );
  INV_X1 U7701 ( .A(n8034), .ZN(n6057) );
  AND2_X1 U7702 ( .A1(n9482), .A2(n6514), .ZN(n6055) );
  AOI21_X1 U7703 ( .B1(n9825), .B2(n4490), .A(n6055), .ZN(n8033) );
  INV_X1 U7704 ( .A(n8033), .ZN(n6056) );
  OR2_X1 U7705 ( .A1(n8045), .A2(n5051), .ZN(n6061) );
  NAND2_X1 U7706 ( .A1(n6059), .A2(n6058), .ZN(n8032) );
  AND2_X1 U7707 ( .A1(n5057), .A2(n8032), .ZN(n6060) );
  NAND2_X1 U7708 ( .A1(n6679), .A2(n9214), .ZN(n6067) );
  OR2_X1 U7709 ( .A1(n6041), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7710 ( .A1(n6062), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6064) );
  INV_X1 U7711 ( .A(n6064), .ZN(n6063) );
  NAND2_X1 U7712 ( .A1(n6063), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7713 ( .A1(n6064), .A2(n7039), .ZN(n6079) );
  AND2_X1 U7714 ( .A1(n6065), .A2(n6079), .ZN(n7796) );
  AOI22_X1 U7715 ( .A1(n6137), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n9986), .B2(
        n7796), .ZN(n6066) );
  NAND2_X1 U7716 ( .A1(n8131), .A2(n4486), .ZN(n6076) );
  NAND2_X1 U7717 ( .A1(n6245), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7718 ( .A1(n4482), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6073) );
  AND2_X1 U7719 ( .A1(n6069), .A2(n6068), .ZN(n6070) );
  NOR2_X1 U7720 ( .A1(n6083), .A2(n6070), .ZN(n8026) );
  NAND2_X1 U7721 ( .A1(n5829), .A2(n8026), .ZN(n6072) );
  NAND2_X1 U7722 ( .A1(n8555), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6071) );
  NAND4_X1 U7723 ( .A1(n6074), .A2(n6073), .A3(n6072), .A4(n6071), .ZN(n9481)
         );
  NAND2_X1 U7724 ( .A1(n9481), .A2(n4490), .ZN(n6075) );
  NAND2_X1 U7725 ( .A1(n6076), .A2(n6075), .ZN(n6077) );
  XNOR2_X1 U7726 ( .A(n6077), .B(n6252), .ZN(n8023) );
  AND2_X1 U7727 ( .A1(n9481), .A2(n6514), .ZN(n6078) );
  AOI21_X1 U7728 ( .B1(n8131), .B2(n4490), .A(n6078), .ZN(n8022) );
  AND2_X1 U7729 ( .A1(n8023), .A2(n8022), .ZN(n6094) );
  NAND2_X1 U7730 ( .A1(n7192), .A2(n9214), .ZN(n6082) );
  NAND2_X1 U7731 ( .A1(n6079), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6080) );
  XNOR2_X1 U7732 ( .A(n6080), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10080) );
  AOI22_X1 U7733 ( .A1(n6137), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9986), .B2(
        n10080), .ZN(n6081) );
  NAND2_X1 U7734 ( .A1(n8555), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6089) );
  INV_X1 U7735 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8140) );
  OR2_X1 U7736 ( .A1(n6296), .A2(n8140), .ZN(n6088) );
  OR2_X1 U7737 ( .A1(n6083), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7738 ( .A1(n6102), .A2(n6084), .ZN(n9188) );
  OR2_X1 U7739 ( .A1(n6527), .A2(n9188), .ZN(n6087) );
  INV_X1 U7740 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6085) );
  OR2_X1 U7741 ( .A1(n8559), .A2(n6085), .ZN(n6086) );
  OAI22_X1 U7742 ( .A1(n9820), .A2(n6216), .B1(n9113), .B2(n6236), .ZN(n6090)
         );
  XNOR2_X1 U7743 ( .A(n6090), .B(n6252), .ZN(n6093) );
  INV_X1 U7744 ( .A(n8023), .ZN(n6092) );
  INV_X1 U7745 ( .A(n8022), .ZN(n6091) );
  NAND2_X1 U7746 ( .A1(n6092), .A2(n6091), .ZN(n6097) );
  OAI22_X1 U7747 ( .A1(n9820), .A2(n6236), .B1(n9113), .B2(n6235), .ZN(n9196)
         );
  INV_X1 U7748 ( .A(n6093), .ZN(n6095) );
  NAND2_X1 U7749 ( .A1(n6095), .A2(n4853), .ZN(n6096) );
  NAND2_X1 U7750 ( .A1(n7200), .A2(n9214), .ZN(n6101) );
  NAND2_X1 U7751 ( .A1(n6098), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6099) );
  XNOR2_X1 U7752 ( .A(n6099), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10092) );
  AOI22_X1 U7753 ( .A1(n6137), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9986), .B2(
        n10092), .ZN(n6100) );
  NAND2_X1 U7754 ( .A1(n9816), .A2(n4487), .ZN(n6110) );
  NAND2_X1 U7755 ( .A1(n4482), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6108) );
  INV_X1 U7756 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9496) );
  OR2_X1 U7757 ( .A1(n8559), .A2(n9496), .ZN(n6107) );
  NAND2_X1 U7758 ( .A1(n6102), .A2(n9111), .ZN(n6103) );
  NAND2_X1 U7759 ( .A1(n6104), .A2(n6103), .ZN(n9112) );
  OR2_X1 U7760 ( .A1(n6527), .A2(n9112), .ZN(n6106) );
  INV_X1 U7761 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n6886) );
  OR2_X1 U7762 ( .A1(n6627), .A2(n6886), .ZN(n6105) );
  INV_X1 U7763 ( .A(n9193), .ZN(n9734) );
  NAND2_X1 U7764 ( .A1(n9734), .A2(n4490), .ZN(n6109) );
  NAND2_X1 U7765 ( .A1(n6110), .A2(n6109), .ZN(n6111) );
  XNOR2_X1 U7766 ( .A(n6111), .B(n6252), .ZN(n6113) );
  NOR2_X1 U7767 ( .A1(n9193), .A2(n6235), .ZN(n6112) );
  AOI21_X1 U7768 ( .B1(n9816), .B2(n4490), .A(n6112), .ZN(n6114) );
  NAND2_X1 U7769 ( .A1(n6113), .A2(n6114), .ZN(n6118) );
  INV_X1 U7770 ( .A(n6113), .ZN(n6116) );
  INV_X1 U7771 ( .A(n6114), .ZN(n6115) );
  NAND2_X1 U7772 ( .A1(n6116), .A2(n6115), .ZN(n6117) );
  NAND2_X1 U7773 ( .A1(n6118), .A2(n6117), .ZN(n9107) );
  NOR3_X4 U7774 ( .A1(n9201), .A2(n9195), .A3(n9107), .ZN(n9110) );
  INV_X1 U7775 ( .A(n6118), .ZN(n6119) );
  XOR2_X1 U7776 ( .A(n6122), .B(n6120), .Z(n9120) );
  NAND2_X1 U7777 ( .A1(n7318), .A2(n9214), .ZN(n6126) );
  NAND2_X1 U7778 ( .A1(n6123), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6124) );
  XNOR2_X1 U7779 ( .A(n6124), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9521) );
  AOI22_X1 U7780 ( .A1(n6137), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9986), .B2(
        n9521), .ZN(n6125) );
  INV_X1 U7781 ( .A(n9804), .ZN(n9712) );
  NAND2_X1 U7782 ( .A1(n8555), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6133) );
  INV_X1 U7783 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9524) );
  OR2_X1 U7784 ( .A1(n8559), .A2(n9524), .ZN(n6132) );
  INV_X1 U7785 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9503) );
  OR2_X1 U7786 ( .A1(n6296), .A2(n9503), .ZN(n6131) );
  OR2_X1 U7787 ( .A1(n6127), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7788 ( .A1(n6129), .A2(n6128), .ZN(n9709) );
  OR2_X1 U7789 ( .A1(n6527), .A2(n9709), .ZN(n6130) );
  OAI22_X1 U7790 ( .A1(n9712), .A2(n6216), .B1(n9123), .B2(n6236), .ZN(n6134)
         );
  XNOR2_X1 U7791 ( .A(n6134), .B(n7574), .ZN(n6135) );
  INV_X1 U7792 ( .A(n9123), .ZN(n9736) );
  AOI22_X1 U7793 ( .A1(n9804), .A2(n4490), .B1(n6514), .B2(n9736), .ZN(n9179)
         );
  NAND2_X1 U7794 ( .A1(n7402), .A2(n9214), .ZN(n6139) );
  AOI22_X1 U7795 ( .A1(n6137), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9670), .B2(
        n9986), .ZN(n6138) );
  NAND2_X1 U7796 ( .A1(n9800), .A2(n4486), .ZN(n6147) );
  INV_X1 U7797 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n7000) );
  OR2_X1 U7798 ( .A1(n8559), .A2(n7000), .ZN(n6145) );
  NAND2_X1 U7799 ( .A1(n4482), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7800 ( .A1(n8555), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6143) );
  NOR2_X1 U7801 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(n6140), .ZN(n6141) );
  NOR2_X1 U7802 ( .A1(n6155), .A2(n6141), .ZN(n9695) );
  NAND2_X1 U7803 ( .A1(n5829), .A2(n9695), .ZN(n6142) );
  NAND4_X1 U7804 ( .A1(n6145), .A2(n6144), .A3(n6143), .A4(n6142), .ZN(n9718)
         );
  NAND2_X1 U7805 ( .A1(n9718), .A2(n4490), .ZN(n6146) );
  NAND2_X1 U7806 ( .A1(n6147), .A2(n6146), .ZN(n6148) );
  XNOR2_X1 U7807 ( .A(n6148), .B(n6252), .ZN(n6151) );
  AND2_X1 U7808 ( .A1(n9718), .A2(n6514), .ZN(n6149) );
  AOI21_X1 U7809 ( .B1(n9800), .B2(n4490), .A(n6149), .ZN(n6150) );
  NAND2_X1 U7810 ( .A1(n6151), .A2(n6150), .ZN(n6152) );
  OAI21_X1 U7811 ( .B1(n6151), .B2(n6150), .A(n6152), .ZN(n9085) );
  INV_X1 U7812 ( .A(n6152), .ZN(n9148) );
  NAND2_X1 U7813 ( .A1(n7548), .A2(n9214), .ZN(n6154) );
  OR2_X1 U7814 ( .A1(n5822), .A2(n7549), .ZN(n6153) );
  NAND2_X1 U7815 ( .A1(n9796), .A2(n4486), .ZN(n6162) );
  INV_X1 U7816 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n6989) );
  OR2_X1 U7817 ( .A1(n6627), .A2(n6989), .ZN(n6160) );
  NAND2_X1 U7818 ( .A1(n4482), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6159) );
  NAND2_X1 U7819 ( .A1(n6245), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6158) );
  NOR2_X1 U7820 ( .A1(n6155), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6156) );
  NOR2_X1 U7821 ( .A1(n6173), .A2(n6156), .ZN(n9685) );
  NAND2_X1 U7822 ( .A1(n5829), .A2(n9685), .ZN(n6157) );
  NAND4_X1 U7823 ( .A1(n6160), .A2(n6159), .A3(n6158), .A4(n6157), .ZN(n9701)
         );
  NAND2_X1 U7824 ( .A1(n9701), .A2(n4490), .ZN(n6161) );
  NAND2_X1 U7825 ( .A1(n6162), .A2(n6161), .ZN(n6163) );
  XNOR2_X1 U7826 ( .A(n6163), .B(n7574), .ZN(n6167) );
  NAND2_X1 U7827 ( .A1(n9796), .A2(n4490), .ZN(n6165) );
  NAND2_X1 U7828 ( .A1(n9701), .A2(n6514), .ZN(n6164) );
  NAND2_X1 U7829 ( .A1(n6165), .A2(n6164), .ZN(n6166) );
  NOR2_X1 U7830 ( .A1(n6167), .A2(n6166), .ZN(n6168) );
  AOI21_X1 U7831 ( .B1(n6167), .B2(n6166), .A(n6168), .ZN(n9147) );
  INV_X1 U7832 ( .A(n6168), .ZN(n6169) );
  NAND2_X1 U7833 ( .A1(n7620), .A2(n9214), .ZN(n6171) );
  OR2_X1 U7834 ( .A1(n5822), .A2(n7621), .ZN(n6170) );
  NAND2_X1 U7835 ( .A1(n9791), .A2(n4487), .ZN(n6180) );
  NAND2_X1 U7836 ( .A1(n6245), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6178) );
  INV_X1 U7837 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n6172) );
  OR2_X1 U7838 ( .A1(n6296), .A2(n6172), .ZN(n6177) );
  OAI21_X1 U7839 ( .B1(n6173), .B2(P1_REG3_REG_21__SCAN_IN), .A(n6189), .ZN(
        n9668) );
  OR2_X1 U7840 ( .A1(n6301), .A2(n9668), .ZN(n6176) );
  INV_X1 U7841 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n6174) );
  OR2_X1 U7842 ( .A1(n6627), .A2(n6174), .ZN(n6175) );
  NAND2_X1 U7843 ( .A1(n9479), .A2(n4490), .ZN(n6179) );
  NAND2_X1 U7844 ( .A1(n6180), .A2(n6179), .ZN(n6181) );
  XNOR2_X1 U7845 ( .A(n6181), .B(n7574), .ZN(n6184) );
  AOI22_X1 U7846 ( .A1(n9791), .A2(n4490), .B1(n6514), .B2(n9479), .ZN(n6182)
         );
  XNOR2_X1 U7847 ( .A(n6184), .B(n6182), .ZN(n9092) );
  INV_X1 U7848 ( .A(n6182), .ZN(n6183) );
  NAND2_X1 U7849 ( .A1(n7799), .A2(n9214), .ZN(n6187) );
  OR2_X1 U7850 ( .A1(n5822), .A2(n7800), .ZN(n6186) );
  NAND2_X1 U7851 ( .A1(n4482), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6196) );
  INV_X1 U7852 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6188) );
  OR2_X1 U7853 ( .A1(n8559), .A2(n6188), .ZN(n6195) );
  AND2_X1 U7854 ( .A1(n6189), .A2(n9160), .ZN(n6191) );
  OR2_X1 U7855 ( .A1(n6191), .A2(n6190), .ZN(n9651) );
  OR2_X1 U7856 ( .A1(n6527), .A2(n9651), .ZN(n6194) );
  INV_X1 U7857 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n6192) );
  OR2_X1 U7858 ( .A1(n6627), .A2(n6192), .ZN(n6193) );
  INV_X1 U7859 ( .A(n9665), .ZN(n9478) );
  AOI22_X1 U7860 ( .A1(n9786), .A2(n4490), .B1(n5923), .B2(n9478), .ZN(n6202)
         );
  NAND2_X1 U7861 ( .A1(n6201), .A2(n6202), .ZN(n9157) );
  OAI22_X1 U7862 ( .A1(n9655), .A2(n6216), .B1(n9665), .B2(n6236), .ZN(n6197)
         );
  XNOR2_X1 U7863 ( .A(n6197), .B(n7574), .ZN(n9159) );
  NAND2_X1 U7864 ( .A1(n9157), .A2(n9159), .ZN(n6205) );
  NAND2_X1 U7865 ( .A1(n9779), .A2(n4487), .ZN(n6199) );
  NAND2_X1 U7866 ( .A1(n9477), .A2(n4490), .ZN(n6198) );
  NAND2_X1 U7867 ( .A1(n6199), .A2(n6198), .ZN(n6200) );
  XNOR2_X1 U7868 ( .A(n6200), .B(n6252), .ZN(n6204) );
  INV_X1 U7869 ( .A(n6202), .ZN(n6203) );
  NAND2_X1 U7870 ( .A1(n4841), .A2(n6203), .ZN(n9156) );
  NAND3_X1 U7871 ( .A1(n6205), .A2(n6204), .A3(n9156), .ZN(n9074) );
  AOI21_X2 U7872 ( .B1(n6205), .B2(n9156), .A(n6204), .ZN(n9075) );
  NAND2_X1 U7873 ( .A1(n7824), .A2(n9214), .ZN(n6207) );
  OR2_X1 U7874 ( .A1(n5822), .A2(n7827), .ZN(n6206) );
  NAND2_X1 U7875 ( .A1(n6245), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6215) );
  INV_X1 U7876 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6208) );
  OR2_X1 U7877 ( .A1(n6296), .A2(n6208), .ZN(n6214) );
  INV_X1 U7878 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9131) );
  NAND2_X1 U7879 ( .A1(n6209), .A2(n9131), .ZN(n6210) );
  NAND2_X1 U7880 ( .A1(n6227), .A2(n6210), .ZN(n9621) );
  OR2_X1 U7881 ( .A1(n6301), .A2(n9621), .ZN(n6213) );
  INV_X1 U7882 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n6211) );
  OR2_X1 U7883 ( .A1(n6627), .A2(n6211), .ZN(n6212) );
  AND4_X2 U7884 ( .A1(n6215), .A2(n6214), .A3(n6213), .A4(n6212), .ZN(n9638)
         );
  OAI22_X1 U7885 ( .A1(n8539), .A2(n6216), .B1(n9638), .B2(n6236), .ZN(n6217)
         );
  XNOR2_X1 U7886 ( .A(n6217), .B(n7574), .ZN(n6221) );
  OR2_X1 U7887 ( .A1(n8539), .A2(n6236), .ZN(n6219) );
  INV_X1 U7888 ( .A(n9638), .ZN(n9608) );
  NAND2_X1 U7889 ( .A1(n9608), .A2(n6514), .ZN(n6218) );
  NAND2_X1 U7890 ( .A1(n6219), .A2(n6218), .ZN(n6220) );
  NOR2_X1 U7891 ( .A1(n6221), .A2(n6220), .ZN(n6222) );
  AOI21_X1 U7892 ( .B1(n6221), .B2(n6220), .A(n6222), .ZN(n9128) );
  INV_X1 U7893 ( .A(n6222), .ZN(n6223) );
  OR2_X1 U7894 ( .A1(n5822), .A2(n7953), .ZN(n6224) );
  NAND2_X1 U7895 ( .A1(n4482), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6234) );
  INV_X1 U7896 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6226) );
  OR2_X1 U7897 ( .A1(n8559), .A2(n6226), .ZN(n6233) );
  INV_X1 U7898 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U7899 ( .A1(n6227), .A2(n9101), .ZN(n6229) );
  INV_X1 U7900 ( .A(n6244), .ZN(n6228) );
  NAND2_X1 U7901 ( .A1(n6229), .A2(n6228), .ZN(n9599) );
  OR2_X1 U7902 ( .A1(n6301), .A2(n9599), .ZN(n6232) );
  INV_X1 U7903 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n6230) );
  OR2_X1 U7904 ( .A1(n6627), .A2(n6230), .ZN(n6231) );
  OAI22_X1 U7905 ( .A1(n9602), .A2(n6236), .B1(n9618), .B2(n6235), .ZN(n6240)
         );
  NAND2_X1 U7906 ( .A1(n9769), .A2(n4486), .ZN(n6238) );
  INV_X1 U7907 ( .A(n9618), .ZN(n9591) );
  NAND2_X1 U7908 ( .A1(n9591), .A2(n4490), .ZN(n6237) );
  NAND2_X1 U7909 ( .A1(n6238), .A2(n6237), .ZN(n6239) );
  XNOR2_X1 U7910 ( .A(n6239), .B(n7574), .ZN(n6241) );
  XOR2_X1 U7911 ( .A(n6240), .B(n6241), .Z(n9099) );
  INV_X1 U7912 ( .A(n6289), .ZN(n6256) );
  NOR2_X1 U7913 ( .A1(n6241), .A2(n6240), .ZN(n6286) );
  NAND2_X1 U7914 ( .A1(n7972), .A2(n9214), .ZN(n6243) );
  OR2_X1 U7915 ( .A1(n5822), .A2(n7975), .ZN(n6242) );
  NAND2_X1 U7916 ( .A1(n9764), .A2(n4487), .ZN(n6251) );
  INV_X1 U7917 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6977) );
  OR2_X1 U7918 ( .A1(n6296), .A2(n6977), .ZN(n6249) );
  NAND2_X1 U7919 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n6244), .ZN(n6299) );
  OAI21_X1 U7920 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n6244), .A(n6299), .ZN(
        n6307) );
  OR2_X1 U7921 ( .A1(n6527), .A2(n6307), .ZN(n6248) );
  INV_X1 U7922 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n6901) );
  OR2_X1 U7923 ( .A1(n6627), .A2(n6901), .ZN(n6247) );
  NAND2_X1 U7924 ( .A1(n6245), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U7925 ( .A1(n9607), .A2(n4490), .ZN(n6250) );
  NAND2_X1 U7926 ( .A1(n6251), .A2(n6250), .ZN(n6253) );
  XNOR2_X1 U7927 ( .A(n6253), .B(n6252), .ZN(n6477) );
  AND2_X1 U7928 ( .A1(n9607), .A2(n5923), .ZN(n6254) );
  AOI21_X1 U7929 ( .B1(n9764), .B2(n4490), .A(n6254), .ZN(n6478) );
  XNOR2_X1 U7930 ( .A(n6477), .B(n6478), .ZN(n6287) );
  OAI21_X1 U7931 ( .B1(n6256), .B2(n6286), .A(n6287), .ZN(n6290) );
  NOR4_X1 U7932 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6260) );
  NOR4_X1 U7933 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6259) );
  NOR4_X1 U7934 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n6258) );
  NOR4_X1 U7935 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n6257) );
  NAND4_X1 U7936 ( .A1(n6260), .A2(n6259), .A3(n6258), .A4(n6257), .ZN(n6270)
         );
  NOR2_X1 U7937 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .ZN(
        n6264) );
  NOR4_X1 U7938 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n6263) );
  NOR4_X1 U7939 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6262) );
  NOR4_X1 U7940 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6261) );
  NAND4_X1 U7941 ( .A1(n6264), .A2(n6263), .A3(n6262), .A4(n6261), .ZN(n6269)
         );
  INV_X1 U7942 ( .A(n6271), .ZN(n7955) );
  NAND3_X1 U7943 ( .A1(n7955), .A2(P1_B_REG_SCAN_IN), .A3(n7829), .ZN(n6268)
         );
  INV_X1 U7944 ( .A(P1_B_REG_SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7945 ( .A1(n6266), .A2(n6265), .ZN(n6267) );
  OAI21_X1 U7946 ( .B1(n6270), .B2(n6269), .A(n10118), .ZN(n6650) );
  INV_X1 U7947 ( .A(n6650), .ZN(n6273) );
  INV_X1 U7948 ( .A(n10118), .ZN(n6272) );
  OAI22_X1 U7949 ( .A1(n6272), .A2(P1_D_REG_1__SCAN_IN), .B1(n6275), .B2(n6271), .ZN(n6651) );
  NOR2_X1 U7950 ( .A1(n6273), .A2(n6651), .ZN(n7561) );
  INV_X1 U7951 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7952 ( .A1(n10118), .A2(n6274), .ZN(n6277) );
  INV_X1 U7953 ( .A(n6275), .ZN(n7977) );
  NAND2_X1 U7954 ( .A1(n7977), .A2(n7829), .ZN(n6276) );
  NAND2_X1 U7955 ( .A1(n6277), .A2(n6276), .ZN(n7916) );
  INV_X1 U7956 ( .A(n7916), .ZN(n6654) );
  NAND2_X1 U7957 ( .A1(n7561), .A2(n6654), .ZN(n7205) );
  NAND2_X1 U7958 ( .A1(n6278), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6279) );
  MUX2_X1 U7959 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6279), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n6280) );
  NAND2_X1 U7960 ( .A1(n6280), .A2(n5059), .ZN(n7780) );
  AND2_X1 U7961 ( .A1(n7780), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6281) );
  AND2_X1 U7962 ( .A1(n6543), .A2(n6281), .ZN(n7563) );
  INV_X1 U7963 ( .A(n7563), .ZN(n10119) );
  OR2_X1 U7964 ( .A1(n7205), .A2(n10119), .ZN(n6293) );
  INV_X1 U7965 ( .A(n6284), .ZN(n9423) );
  INV_X1 U7966 ( .A(n6292), .ZN(n6285) );
  NAND2_X1 U7967 ( .A1(n9209), .A2(n6284), .ZN(n9368) );
  INV_X1 U7968 ( .A(n9368), .ZN(n7598) );
  OR2_X1 U7969 ( .A1(n9964), .A2(n7598), .ZN(n6308) );
  NOR2_X1 U7970 ( .A1(n6287), .A2(n6286), .ZN(n6288) );
  NAND2_X2 U7971 ( .A1(n6289), .A2(n6288), .ZN(n6495) );
  NAND3_X1 U7972 ( .A1(n6290), .A2(n9168), .A3(n6495), .ZN(n6321) );
  INV_X1 U7973 ( .A(n5775), .ZN(n7588) );
  NAND2_X1 U7974 ( .A1(n7570), .A2(n7588), .ZN(n7568) );
  OR2_X1 U7975 ( .A1(n5770), .A2(n7626), .ZN(n9207) );
  AOI21_X1 U7976 ( .B1(n7568), .B2(n9207), .A(n10119), .ZN(n6291) );
  NAND2_X1 U7977 ( .A1(n7205), .A2(n6291), .ZN(n6313) );
  OR2_X1 U7978 ( .A1(n9368), .A2(n6292), .ZN(n6310) );
  NAND2_X1 U7979 ( .A1(n6310), .A2(n7563), .ZN(n7917) );
  INV_X1 U7980 ( .A(n7917), .ZN(n7562) );
  AND2_X1 U7981 ( .A1(n6313), .A2(n7562), .ZN(n7544) );
  NAND2_X1 U7982 ( .A1(n9764), .A2(n9205), .ZN(n6320) );
  OR2_X1 U7983 ( .A1(n6293), .A2(n9207), .ZN(n6316) );
  INV_X1 U7984 ( .A(n4481), .ZN(n9998) );
  NOR2_X1 U7985 ( .A1(n6316), .A2(n9998), .ZN(n9170) );
  NAND2_X1 U7986 ( .A1(n8555), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6306) );
  INV_X1 U7987 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6295) );
  OR2_X1 U7988 ( .A1(n6296), .A2(n6295), .ZN(n6305) );
  INV_X1 U7989 ( .A(n6299), .ZN(n6297) );
  NAND2_X1 U7990 ( .A1(n6297), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6499) );
  INV_X1 U7991 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U7992 ( .A1(n6299), .A2(n6298), .ZN(n6300) );
  NAND2_X1 U7993 ( .A1(n6499), .A2(n6300), .ZN(n6506) );
  OR2_X1 U7994 ( .A1(n6301), .A2(n6506), .ZN(n6304) );
  INV_X1 U7995 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6302) );
  OR2_X1 U7996 ( .A1(n8559), .A2(n6302), .ZN(n6303) );
  INV_X1 U7997 ( .A(n6307), .ZN(n9584) );
  INV_X1 U7998 ( .A(n6308), .ZN(n6309) );
  NAND2_X1 U7999 ( .A1(n7205), .A2(n6309), .ZN(n6312) );
  AND3_X1 U8000 ( .A1(n6310), .A2(n6543), .A3(n7780), .ZN(n6311) );
  AOI21_X1 U8001 ( .B1(n6312), .B2(n6311), .A(P1_U3084), .ZN(n6315) );
  INV_X1 U8002 ( .A(n6313), .ZN(n6314) );
  AOI22_X1 U8003 ( .A1(n9170), .A2(n9592), .B1(n9584), .B2(n9189), .ZN(n6318)
         );
  NOR2_X2 U8004 ( .A1(n6316), .A2(n4481), .ZN(n9191) );
  AOI22_X1 U8005 ( .A1(n9191), .A2(n9591), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n6317) );
  NAND2_X1 U8006 ( .A1(n6321), .A2(n5061), .ZN(P1_U3238) );
  NAND3_X1 U8007 ( .A1(n6323), .A2(n6322), .A3(n8330), .ZN(n6324) );
  NAND2_X1 U8008 ( .A1(n9922), .A2(n8856), .ZN(n6360) );
  NAND2_X1 U8009 ( .A1(n6398), .A2(n8681), .ZN(n6334) );
  NAND3_X1 U8010 ( .A1(n6360), .A2(n8683), .A3(n6328), .ZN(n6331) );
  NAND2_X1 U8011 ( .A1(n6331), .A2(n6330), .ZN(n6667) );
  INV_X1 U8012 ( .A(n6332), .ZN(n6333) );
  INV_X1 U8013 ( .A(n6334), .ZN(n6335) );
  XNOR2_X1 U8014 ( .A(n4480), .B(n6329), .ZN(n6340) );
  NAND2_X1 U8015 ( .A1(n6398), .A2(n8680), .ZN(n6339) );
  XNOR2_X1 U8016 ( .A(n6340), .B(n6339), .ZN(n6633) );
  XNOR2_X1 U8017 ( .A(n8271), .B(n6329), .ZN(n6342) );
  NAND2_X1 U8018 ( .A1(n6398), .A2(n8679), .ZN(n6341) );
  NAND2_X1 U8019 ( .A1(n6342), .A2(n6341), .ZN(n6343) );
  OAI21_X1 U8020 ( .B1(n6342), .B2(n6341), .A(n6343), .ZN(n6684) );
  XNOR2_X1 U8021 ( .A(n7302), .B(n6422), .ZN(n6345) );
  NAND2_X1 U8022 ( .A1(n6398), .A2(n8678), .ZN(n6344) );
  XNOR2_X1 U8023 ( .A(n6345), .B(n6344), .ZN(n6694) );
  INV_X1 U8024 ( .A(n6344), .ZN(n6346) );
  AND2_X1 U8025 ( .A1(n8329), .A2(n8677), .ZN(n6348) );
  XNOR2_X1 U8026 ( .A(n10321), .B(n6422), .ZN(n6347) );
  NOR2_X1 U8027 ( .A1(n6347), .A2(n6348), .ZN(n6349) );
  AOI21_X1 U8028 ( .B1(n6348), .B2(n6347), .A(n6349), .ZN(n7229) );
  NAND2_X1 U8029 ( .A1(n6398), .A2(n10259), .ZN(n6352) );
  XNOR2_X1 U8030 ( .A(n7458), .B(n6422), .ZN(n6351) );
  XOR2_X1 U8031 ( .A(n6352), .B(n6351), .Z(n7309) );
  INV_X1 U8032 ( .A(n6349), .ZN(n7307) );
  NAND2_X1 U8033 ( .A1(n6351), .A2(n6353), .ZN(n6354) );
  XNOR2_X1 U8034 ( .A(n8588), .B(n6422), .ZN(n6356) );
  NAND2_X1 U8035 ( .A1(n8329), .A2(n8676), .ZN(n6355) );
  XNOR2_X1 U8036 ( .A(n6356), .B(n6355), .ZN(n8580) );
  INV_X1 U8037 ( .A(n6355), .ZN(n6357) );
  XNOR2_X1 U8038 ( .A(n7389), .B(n6422), .ZN(n6359) );
  AND2_X1 U8039 ( .A1(n8329), .A2(n10257), .ZN(n6358) );
  NAND2_X1 U8040 ( .A1(n6359), .A2(n6358), .ZN(n7365) );
  NOR2_X1 U8041 ( .A1(n6359), .A2(n6358), .ZN(n7367) );
  XNOR2_X1 U8042 ( .A(n7425), .B(n6329), .ZN(n6362) );
  NAND2_X1 U8043 ( .A1(n8329), .A2(n8675), .ZN(n6361) );
  NOR2_X1 U8044 ( .A1(n6362), .A2(n6361), .ZN(n6363) );
  AOI21_X1 U8045 ( .B1(n6362), .B2(n6361), .A(n6363), .ZN(n7407) );
  INV_X1 U8046 ( .A(n6363), .ZN(n6364) );
  XNOR2_X1 U8047 ( .A(n7528), .B(n6422), .ZN(n6365) );
  NAND2_X1 U8048 ( .A1(n6398), .A2(n8674), .ZN(n6366) );
  XNOR2_X1 U8049 ( .A(n6365), .B(n6366), .ZN(n7498) );
  NAND2_X1 U8050 ( .A1(n7499), .A2(n7498), .ZN(n7497) );
  INV_X1 U8051 ( .A(n6366), .ZN(n6367) );
  NAND2_X1 U8052 ( .A1(n6365), .A2(n6367), .ZN(n6368) );
  XNOR2_X1 U8053 ( .A(n7479), .B(n6329), .ZN(n6370) );
  NAND2_X1 U8054 ( .A1(n8329), .A2(n8673), .ZN(n6369) );
  NAND2_X1 U8055 ( .A1(n6370), .A2(n6369), .ZN(n7644) );
  NAND2_X1 U8057 ( .A1(n8329), .A2(n8672), .ZN(n6372) );
  XNOR2_X1 U8058 ( .A(n5468), .B(n6422), .ZN(n6371) );
  XOR2_X1 U8059 ( .A(n6372), .B(n6371), .Z(n7734) );
  XNOR2_X1 U8060 ( .A(n9917), .B(n6329), .ZN(n6374) );
  NAND2_X1 U8061 ( .A1(n8329), .A2(n8671), .ZN(n6373) );
  NAND2_X1 U8062 ( .A1(n6374), .A2(n6373), .ZN(n6375) );
  OAI21_X1 U8063 ( .B1(n6374), .B2(n6373), .A(n6375), .ZN(n7855) );
  XOR2_X1 U8064 ( .A(n6422), .B(n8060), .Z(n6377) );
  NAND2_X1 U8065 ( .A1(n6376), .A2(n6377), .ZN(n6381) );
  NOR2_X1 U8066 ( .A1(n8152), .A2(n6673), .ZN(n8055) );
  INV_X1 U8067 ( .A(n6381), .ZN(n8149) );
  XNOR2_X1 U8068 ( .A(n9025), .B(n6422), .ZN(n6384) );
  NAND2_X1 U8069 ( .A1(n8669), .A2(n8329), .ZN(n6382) );
  XNOR2_X1 U8070 ( .A(n6384), .B(n6382), .ZN(n8148) );
  INV_X1 U8071 ( .A(n6382), .ZN(n6383) );
  NAND2_X1 U8072 ( .A1(n8668), .A2(n8329), .ZN(n6387) );
  XNOR2_X1 U8073 ( .A(n8203), .B(n6422), .ZN(n6386) );
  XOR2_X1 U8074 ( .A(n6387), .B(n6386), .Z(n8196) );
  INV_X1 U8075 ( .A(n6386), .ZN(n6388) );
  XNOR2_X1 U8076 ( .A(n9020), .B(n6422), .ZN(n6390) );
  NAND2_X1 U8077 ( .A1(n8667), .A2(n8329), .ZN(n6389) );
  XNOR2_X1 U8078 ( .A(n6390), .B(n6389), .ZN(n8233) );
  INV_X1 U8079 ( .A(n6389), .ZN(n6391) );
  AND2_X1 U8080 ( .A1(n8666), .A2(n8329), .ZN(n6393) );
  XNOR2_X1 U8081 ( .A(n8248), .B(n6422), .ZN(n6392) );
  NOR2_X1 U8082 ( .A1(n6392), .A2(n6393), .ZN(n6394) );
  AOI21_X1 U8083 ( .B1(n6393), .B2(n6392), .A(n6394), .ZN(n8571) );
  NAND2_X1 U8084 ( .A1(n8665), .A2(n8329), .ZN(n6396) );
  XNOR2_X1 U8085 ( .A(n8950), .B(n6422), .ZN(n6395) );
  XOR2_X1 U8086 ( .A(n6396), .B(n6395), .Z(n8621) );
  INV_X1 U8087 ( .A(n6395), .ZN(n6397) );
  NAND2_X1 U8088 ( .A1(n8664), .A2(n6398), .ZN(n6399) );
  XNOR2_X1 U8089 ( .A(n6400), .B(n6399), .ZN(n8593) );
  INV_X1 U8090 ( .A(n6399), .ZN(n6401) );
  XNOR2_X1 U8091 ( .A(n8920), .B(n6422), .ZN(n6402) );
  NAND2_X1 U8092 ( .A1(n8663), .A2(n8329), .ZN(n8629) );
  NAND2_X1 U8093 ( .A1(n8630), .A2(n8629), .ZN(n8628) );
  INV_X1 U8094 ( .A(n6402), .ZN(n6403) );
  NAND2_X1 U8095 ( .A1(n6404), .A2(n6403), .ZN(n6405) );
  NAND2_X1 U8096 ( .A1(n8628), .A2(n6405), .ZN(n6408) );
  XNOR2_X1 U8097 ( .A(n8991), .B(n6422), .ZN(n6406) );
  XNOR2_X1 U8098 ( .A(n6408), .B(n6406), .ZN(n8564) );
  NOR2_X1 U8099 ( .A1(n8634), .A2(n6673), .ZN(n8565) );
  INV_X1 U8100 ( .A(n6406), .ZN(n6407) );
  NOR2_X1 U8101 ( .A1(n6408), .A2(n6407), .ZN(n6409) );
  XNOR2_X1 U8102 ( .A(n8887), .B(n6422), .ZN(n6410) );
  NOR2_X1 U8103 ( .A1(n8605), .A2(n6673), .ZN(n8613) );
  NAND2_X1 U8104 ( .A1(n8612), .A2(n8613), .ZN(n6414) );
  INV_X1 U8105 ( .A(n6410), .ZN(n6411) );
  XNOR2_X1 U8106 ( .A(n8980), .B(n6422), .ZN(n8603) );
  NAND2_X1 U8107 ( .A1(n8601), .A2(n8603), .ZN(n6415) );
  NAND2_X1 U8108 ( .A1(n8661), .A2(n8329), .ZN(n8602) );
  INV_X1 U8109 ( .A(n8601), .ZN(n6417) );
  INV_X1 U8110 ( .A(n8603), .ZN(n6416) );
  XNOR2_X1 U8111 ( .A(n8859), .B(n6422), .ZN(n6419) );
  AND2_X1 U8112 ( .A1(n8660), .A2(n8329), .ZN(n6418) );
  NAND2_X1 U8113 ( .A1(n6419), .A2(n6418), .ZN(n6465) );
  OAI21_X1 U8114 ( .B1(n6419), .B2(n6418), .A(n6465), .ZN(n8643) );
  XNOR2_X1 U8115 ( .A(n8970), .B(n6329), .ZN(n6421) );
  NAND2_X1 U8116 ( .A1(n8659), .A2(n8329), .ZN(n6420) );
  NOR2_X1 U8117 ( .A1(n6421), .A2(n6420), .ZN(n6430) );
  INV_X1 U8118 ( .A(n6467), .ZN(n6431) );
  OR2_X1 U8119 ( .A1(n8643), .A2(n6431), .ZN(n6440) );
  NAND2_X1 U8120 ( .A1(n8815), .A2(n8329), .ZN(n6423) );
  XNOR2_X1 U8121 ( .A(n6423), .B(n6422), .ZN(n6438) );
  AND2_X1 U8122 ( .A1(n6425), .A2(n6424), .ZN(n7346) );
  NOR2_X1 U8123 ( .A1(n6426), .A2(n7112), .ZN(n6427) );
  AND2_X1 U8124 ( .A1(n7346), .A2(n6427), .ZN(n6450) );
  INV_X1 U8125 ( .A(n8479), .ZN(n8516) );
  AND2_X1 U8126 ( .A1(n5711), .A2(n8516), .ZN(n7353) );
  NAND2_X1 U8127 ( .A1(n6450), .A2(n7353), .ZN(n6428) );
  NOR3_X1 U8128 ( .A1(n8802), .A2(n8618), .A3(n6438), .ZN(n6429) );
  AOI21_X1 U8129 ( .B1(n8802), .B2(n6438), .A(n6429), .ZN(n6434) );
  INV_X1 U8130 ( .A(n6430), .ZN(n6432) );
  OR2_X1 U8131 ( .A1(n6431), .A2(n6465), .ZN(n6460) );
  AND2_X1 U8132 ( .A1(n6432), .A2(n6460), .ZN(n6441) );
  NAND2_X1 U8133 ( .A1(n6436), .A2(n6435), .ZN(n6447) );
  NAND3_X1 U8134 ( .A1(n8827), .A2(n8657), .A3(n6438), .ZN(n6437) );
  OAI21_X1 U8135 ( .B1(n8827), .B2(n6438), .A(n6437), .ZN(n6439) );
  INV_X1 U8136 ( .A(n6439), .ZN(n6442) );
  AND2_X1 U8137 ( .A1(n10362), .A2(n6602), .ZN(n6444) );
  NAND2_X1 U8138 ( .A1(n6450), .A2(n6444), .ZN(n8642) );
  OAI21_X1 U8139 ( .B1(n8802), .B2(n8657), .A(n8642), .ZN(n6445) );
  INV_X1 U8140 ( .A(n6448), .ZN(n6449) );
  NAND2_X1 U8141 ( .A1(n7346), .A2(n7344), .ZN(n6453) );
  NAND2_X1 U8142 ( .A1(n6453), .A2(n6452), .ZN(n6644) );
  AND3_X1 U8143 ( .A1(n7114), .A2(n6603), .A3(n6454), .ZN(n6455) );
  NAND2_X1 U8144 ( .A1(n6644), .A2(n6455), .ZN(n6456) );
  AOI22_X1 U8145 ( .A1(n8821), .A2(n8639), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6457) );
  INV_X1 U8146 ( .A(n6460), .ZN(n6461) );
  OR2_X1 U8147 ( .A1(n6461), .A2(n8642), .ZN(n6462) );
  NOR2_X1 U8148 ( .A1(n6463), .A2(n6462), .ZN(n6470) );
  INV_X1 U8149 ( .A(n8643), .ZN(n6464) );
  NAND2_X1 U8150 ( .A1(n6470), .A2(n6469), .ZN(n6476) );
  INV_X1 U8151 ( .A(n8647), .ZN(n10260) );
  AOI22_X1 U8152 ( .A1(n8815), .A2(n10258), .B1(n10260), .B2(n8660), .ZN(n8835) );
  INV_X1 U8153 ( .A(n8654), .ZN(n8637) );
  OAI22_X1 U8154 ( .A1(n8835), .A2(n8637), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6471), .ZN(n6472) );
  AOI21_X1 U8155 ( .B1(n8839), .B2(n8639), .A(n6472), .ZN(n6473) );
  NAND2_X1 U8156 ( .A1(n6476), .A2(n6475), .ZN(P2_U3216) );
  INV_X1 U8157 ( .A(n6477), .ZN(n6480) );
  INV_X1 U8158 ( .A(n6478), .ZN(n6479) );
  NAND2_X1 U8159 ( .A1(n6480), .A2(n6479), .ZN(n6491) );
  OR2_X1 U8160 ( .A1(n5822), .A2(n8065), .ZN(n6481) );
  NAND2_X1 U8161 ( .A1(n9759), .A2(n4487), .ZN(n6484) );
  NAND2_X1 U8162 ( .A1(n9592), .A2(n4490), .ZN(n6483) );
  NAND2_X1 U8163 ( .A1(n6484), .A2(n6483), .ZN(n6485) );
  XNOR2_X1 U8164 ( .A(n6485), .B(n7574), .ZN(n6489) );
  NAND2_X1 U8165 ( .A1(n9759), .A2(n4490), .ZN(n6487) );
  NAND2_X1 U8166 ( .A1(n9592), .A2(n5923), .ZN(n6486) );
  NAND2_X1 U8167 ( .A1(n6487), .A2(n6486), .ZN(n6488) );
  AOI21_X1 U8168 ( .B1(n6489), .B2(n6488), .A(n6523), .ZN(n6490) );
  AOI21_X1 U8169 ( .B1(n6495), .B2(n6491), .A(n6490), .ZN(n6496) );
  INV_X1 U8170 ( .A(n6490), .ZN(n6493) );
  INV_X1 U8171 ( .A(n6491), .ZN(n6492) );
  NOR2_X1 U8172 ( .A1(n6493), .A2(n6492), .ZN(n6494) );
  OAI21_X1 U8173 ( .B1(n6496), .B2(n6539), .A(n9168), .ZN(n6511) );
  NAND2_X1 U8174 ( .A1(n9759), .A2(n9205), .ZN(n6510) );
  NAND2_X1 U8175 ( .A1(n4482), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6505) );
  INV_X1 U8176 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6497) );
  OR2_X1 U8177 ( .A1(n8559), .A2(n6497), .ZN(n6504) );
  INV_X1 U8178 ( .A(n6499), .ZN(n6498) );
  NAND2_X1 U8179 ( .A1(n6498), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8546) );
  INV_X1 U8180 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6525) );
  NAND2_X1 U8181 ( .A1(n6499), .A2(n6525), .ZN(n6500) );
  NAND2_X1 U8182 ( .A1(n8546), .A2(n6500), .ZN(n9553) );
  INV_X1 U8183 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6501) );
  OR2_X1 U8184 ( .A1(n6627), .A2(n6501), .ZN(n6502) );
  INV_X1 U8185 ( .A(n9572), .ZN(n9476) );
  INV_X1 U8186 ( .A(n6506), .ZN(n9569) );
  AOI22_X1 U8187 ( .A1(n9170), .A2(n9476), .B1(n9569), .B2(n9189), .ZN(n6508)
         );
  AOI22_X1 U8188 ( .A1(n9191), .A2(n9607), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n6507) );
  NAND3_X1 U8189 ( .A1(n6511), .A2(n6510), .A3(n6509), .ZN(P1_U3212) );
  INV_X1 U8190 ( .A(n6523), .ZN(n6521) );
  NAND2_X1 U8191 ( .A1(n8220), .A2(n9214), .ZN(n6513) );
  INV_X1 U8192 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8222) );
  OR2_X1 U8193 ( .A1(n5822), .A2(n8222), .ZN(n6512) );
  NAND2_X1 U8194 ( .A1(n9755), .A2(n4490), .ZN(n6516) );
  NAND2_X1 U8195 ( .A1(n9476), .A2(n5923), .ZN(n6515) );
  NAND2_X1 U8196 ( .A1(n6516), .A2(n6515), .ZN(n6517) );
  XNOR2_X1 U8197 ( .A(n6517), .B(n7574), .ZN(n6519) );
  AOI22_X1 U8198 ( .A1(n9755), .A2(n4487), .B1(n5802), .B2(n9476), .ZN(n6518)
         );
  XNOR2_X1 U8199 ( .A(n6519), .B(n6518), .ZN(n6524) );
  INV_X1 U8200 ( .A(n6524), .ZN(n6520) );
  NAND4_X1 U8201 ( .A1(n6522), .A2(n6521), .A3(n6520), .A4(n9168), .ZN(n6541)
         );
  AND2_X1 U8202 ( .A1(n6524), .A2(n9168), .ZN(n6538) );
  NAND3_X1 U8203 ( .A1(n6524), .A2(n9168), .A3(n6523), .ZN(n6536) );
  INV_X1 U8204 ( .A(n9191), .ZN(n9183) );
  OAI22_X1 U8205 ( .A1(n9183), .A2(n8541), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6525), .ZN(n6534) );
  NAND2_X1 U8206 ( .A1(n4482), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6532) );
  INV_X1 U8207 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6526) );
  OR2_X1 U8208 ( .A1(n8559), .A2(n6526), .ZN(n6531) );
  OR2_X1 U8209 ( .A1(n6527), .A2(n8546), .ZN(n6530) );
  INV_X1 U8210 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6528) );
  OR2_X1 U8211 ( .A1(n6627), .A2(n6528), .ZN(n6529) );
  OAI22_X1 U8212 ( .A1(n9194), .A2(n9557), .B1(n9181), .B2(n9553), .ZN(n6533)
         );
  AOI211_X1 U8213 ( .C1(n9755), .C2(n9205), .A(n6534), .B(n6533), .ZN(n6535)
         );
  AOI21_X1 U8214 ( .B1(n6539), .B2(n6538), .A(n6537), .ZN(n6540) );
  NAND2_X1 U8215 ( .A1(n6541), .A2(n6540), .ZN(P1_U3218) );
  INV_X1 U8216 ( .A(n7780), .ZN(n6542) );
  NOR2_X1 U8217 ( .A1(n6543), .A2(n6542), .ZN(n6580) );
  NAND2_X1 U8218 ( .A1(n9368), .A2(n6543), .ZN(n6544) );
  NAND2_X1 U8219 ( .A1(n6544), .A2(n7780), .ZN(n6558) );
  NAND2_X1 U8220 ( .A1(n6558), .A2(n4489), .ZN(n6546) );
  NAND2_X1 U8221 ( .A1(n6546), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8222 ( .A(n10313), .ZN(n10298) );
  NOR2_X1 U8223 ( .A1(n7114), .A2(n10298), .ZN(P2_U3966) );
  AND2_X1 U8224 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7820) );
  NOR2_X1 U8225 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6573), .ZN(n6547) );
  AOI21_X1 U8226 ( .B1(n6573), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6547), .ZN(
        n6702) );
  NOR2_X1 U8227 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6563), .ZN(n6548) );
  AOI21_X1 U8228 ( .B1(n6563), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6548), .ZN(
        n10038) );
  XNOR2_X1 U8229 ( .A(n6721), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n6718) );
  INV_X1 U8230 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10000) );
  INV_X1 U8231 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7573) );
  NOR2_X1 U8232 ( .A1(n10000), .A2(n7573), .ZN(n9996) );
  NAND2_X1 U8233 ( .A1(n6718), .A2(n9996), .ZN(n6717) );
  INV_X1 U8234 ( .A(n6721), .ZN(n6567) );
  NAND2_X1 U8235 ( .A1(n6567), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6549) );
  AND2_X1 U8236 ( .A1(n6717), .A2(n6549), .ZN(n10011) );
  NAND2_X1 U8237 ( .A1(n10014), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6550) );
  OAI21_X1 U8238 ( .B1(n10014), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6550), .ZN(
        n10010) );
  NOR2_X1 U8239 ( .A1(n10011), .A2(n10010), .ZN(n10009) );
  AOI21_X1 U8240 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n10014), .A(n10009), .ZN(
        n9865) );
  INV_X1 U8241 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6551) );
  AOI22_X1 U8242 ( .A1(n6565), .A2(n6551), .B1(P1_REG2_REG_3__SCAN_IN), .B2(
        n9862), .ZN(n9866) );
  AND2_X1 U8243 ( .A1(n6565), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6552) );
  INV_X1 U8244 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6553) );
  MUX2_X1 U8245 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6553), .S(n10028), .Z(n10018) );
  OAI21_X1 U8246 ( .B1(n10028), .B2(P1_REG2_REG_4__SCAN_IN), .A(n10019), .ZN(
        n10039) );
  NAND2_X1 U8247 ( .A1(n10038), .A2(n10039), .ZN(n10037) );
  INV_X1 U8248 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6554) );
  MUX2_X1 U8249 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6554), .S(n6732), .Z(n6555)
         );
  INV_X1 U8250 ( .A(n6555), .ZN(n6728) );
  OAI21_X1 U8251 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6573), .A(n6700), .ZN(
        n10052) );
  XNOR2_X1 U8252 ( .A(n10049), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n10051) );
  NAND2_X1 U8253 ( .A1(n6741), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6556) );
  OAI21_X1 U8254 ( .B1(n6741), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6556), .ZN(
        n6557) );
  INV_X1 U8255 ( .A(n6557), .ZN(n6559) );
  NAND2_X1 U8256 ( .A1(n6558), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9988) );
  OR2_X1 U8257 ( .A1(n9988), .A2(n4491), .ZN(n9522) );
  OR2_X1 U8258 ( .A1(n9522), .A2(n4481), .ZN(n10086) );
  INV_X1 U8259 ( .A(n10086), .ZN(n10104) );
  OAI21_X1 U8260 ( .B1(n6560), .B2(n6559), .A(n10104), .ZN(n6561) );
  NOR2_X1 U8261 ( .A1(n6561), .A2(n6740), .ZN(n6583) );
  INV_X1 U8262 ( .A(n10049), .ZN(n6562) );
  NAND2_X1 U8263 ( .A1(n6562), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6576) );
  NOR2_X1 U8264 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6573), .ZN(n6574) );
  INV_X1 U8265 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10227) );
  NAND2_X1 U8266 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6563), .ZN(n6572) );
  INV_X1 U8267 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6564) );
  MUX2_X1 U8268 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6564), .S(n6563), .Z(n10042)
         );
  INV_X1 U8269 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10224) );
  AOI22_X1 U8270 ( .A1(n10028), .A2(n10224), .B1(P1_REG1_REG_4__SCAN_IN), .B2(
        n6595), .ZN(n10024) );
  INV_X1 U8271 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10222) );
  MUX2_X1 U8272 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10222), .S(n6565), .Z(n9869)
         );
  NAND2_X1 U8273 ( .A1(n10014), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6570) );
  MUX2_X1 U8274 ( .A(n10220), .B(P1_REG1_REG_2__SCAN_IN), .S(n10014), .Z(
        n10005) );
  INV_X1 U8275 ( .A(n10005), .ZN(n6569) );
  MUX2_X1 U8276 ( .A(n6566), .B(P1_REG1_REG_1__SCAN_IN), .S(n6721), .Z(n6713)
         );
  AND2_X1 U8277 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6714) );
  NAND2_X1 U8278 ( .A1(n6713), .A2(n6714), .ZN(n6712) );
  NAND2_X1 U8279 ( .A1(n6567), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6568) );
  NAND2_X1 U8280 ( .A1(n6712), .A2(n6568), .ZN(n10006) );
  NAND2_X1 U8281 ( .A1(n9869), .A2(n9870), .ZN(n9868) );
  OAI21_X1 U8282 ( .B1(n10222), .B2(n9862), .A(n9868), .ZN(n10023) );
  NOR2_X1 U8283 ( .A1(n10024), .A2(n10023), .ZN(n10022) );
  NOR2_X1 U8284 ( .A1(n10028), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U8285 ( .A1(n10042), .A2(n10043), .ZN(n10041) );
  NAND2_X1 U8286 ( .A1(n6572), .A2(n10041), .ZN(n6724) );
  AOI22_X1 U8287 ( .A1(n6732), .A2(n10227), .B1(P1_REG1_REG_6__SCAN_IN), .B2(
        n8259), .ZN(n6723) );
  NOR2_X1 U8288 ( .A1(n6724), .A2(n6723), .ZN(n6722) );
  INV_X1 U8289 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10229) );
  AOI22_X1 U8290 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6706), .B1(n6573), .B2(
        n10229), .ZN(n6704) );
  NOR2_X1 U8291 ( .A1(n6705), .A2(n6704), .ZN(n6703) );
  INV_X1 U8292 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10231) );
  INV_X1 U8293 ( .A(n6576), .ZN(n6575) );
  AOI21_X1 U8294 ( .B1(n10231), .B2(n10049), .A(n6575), .ZN(n10055) );
  NAND2_X1 U8295 ( .A1(n10056), .A2(n10055), .ZN(n10054) );
  NAND2_X1 U8296 ( .A1(n6576), .A2(n10054), .ZN(n6578) );
  INV_X1 U8297 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10234) );
  AOI22_X1 U8298 ( .A1(n6741), .A2(n10234), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6613), .ZN(n6577) );
  NOR2_X1 U8299 ( .A1(n6578), .A2(n6577), .ZN(n6734) );
  AOI21_X1 U8300 ( .B1(n6578), .B2(n6577), .A(n6734), .ZN(n6579) );
  INV_X1 U8301 ( .A(n4491), .ZN(n9995) );
  NOR2_X1 U8302 ( .A1(n6579), .A2(n10070), .ZN(n6582) );
  OR2_X1 U8303 ( .A1(n9522), .A2(n9998), .ZN(n10107) );
  INV_X1 U8304 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10422) );
  OAI22_X1 U8305 ( .A1(n10107), .A2(n6613), .B1(n10116), .B2(n10422), .ZN(
        n6581) );
  OR4_X1 U8306 ( .A1(n7820), .A2(n6583), .A3(n6582), .A4(n6581), .ZN(P1_U3250)
         );
  INV_X2 U8307 ( .A(n8114), .ZN(n9070) );
  OAI222_X1 U8308 ( .A1(P2_U3152), .A2(n7122), .B1(n9070), .B2(n6593), .C1(
        n6584), .C2(n8311), .ZN(P2_U3357) );
  OAI222_X1 U8309 ( .A1(n8311), .A2(n6586), .B1(n9070), .B2(n6589), .C1(
        P2_U3152), .C2(n6585), .ZN(P2_U3356) );
  INV_X1 U8310 ( .A(n7143), .ZN(n7164) );
  OAI222_X1 U8311 ( .A1(n8311), .A2(n6992), .B1(n9070), .B2(n6591), .C1(
        P2_U3152), .C2(n7164), .ZN(P2_U3353) );
  OAI222_X1 U8312 ( .A1(n8311), .A2(n6587), .B1(n9070), .B2(n5856), .C1(
        P2_U3152), .C2(n7146), .ZN(P2_U3354) );
  INV_X1 U8313 ( .A(n8257), .ZN(n7201) );
  INV_X1 U8314 ( .A(n7201), .ZN(n9859) );
  OAI222_X1 U8315 ( .A1(n9859), .A2(n6590), .B1(n9857), .B2(n6589), .C1(n6588), 
        .C2(P1_U3084), .ZN(P1_U3351) );
  OAI222_X1 U8316 ( .A1(n9859), .A2(n6592), .B1(n9857), .B2(n6591), .C1(n10035), .C2(P1_U3084), .ZN(P1_U3348) );
  OAI222_X1 U8317 ( .A1(n9859), .A2(n6594), .B1(n9857), .B2(n6593), .C1(n6721), 
        .C2(P1_U3084), .ZN(P1_U3352) );
  OAI222_X1 U8318 ( .A1(n9859), .A2(n6596), .B1(n9857), .B2(n5856), .C1(n6595), 
        .C2(P1_U3084), .ZN(P1_U3349) );
  NAND2_X1 U8319 ( .A1(n10119), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6597) );
  OAI21_X1 U8320 ( .B1(n6651), .B2(n10119), .A(n6597), .ZN(P1_U3441) );
  OAI222_X1 U8321 ( .A1(n6706), .A2(P1_U3084), .B1(n9857), .B2(n6599), .C1(
        n6598), .C2(n9859), .ZN(P1_U3346) );
  INV_X1 U8322 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6600) );
  INV_X1 U8323 ( .A(n7330), .ZN(n7178) );
  OAI222_X1 U8324 ( .A1(n6600), .A2(n8311), .B1(P2_U3152), .B2(n7178), .C1(
        n9070), .C2(n6599), .ZN(P2_U3351) );
  NAND2_X1 U8325 ( .A1(n6654), .A2(n7563), .ZN(n6601) );
  OAI21_X1 U8326 ( .B1(n7563), .B2(n6274), .A(n6601), .ZN(P1_U3440) );
  OAI21_X1 U8327 ( .B1(n7112), .B2(n6602), .A(n7126), .ZN(n6605) );
  NOR2_X1 U8328 ( .A1(n6603), .A2(P2_U3152), .ZN(n8526) );
  INV_X1 U8329 ( .A(n8526), .ZN(n8530) );
  NAND2_X1 U8330 ( .A1(n7112), .A2(n8530), .ZN(n6604) );
  NAND2_X1 U8331 ( .A1(n6605), .A2(n6604), .ZN(n8791) );
  INV_X1 U8332 ( .A(n8791), .ZN(n10243) );
  NOR2_X1 U8333 ( .A1(n10243), .A2(P2_U3966), .ZN(P2_U3151) );
  OAI222_X1 U8334 ( .A1(n9859), .A2(n6606), .B1(n9857), .B2(n6607), .C1(n10049), .C2(P1_U3084), .ZN(P1_U3345) );
  INV_X1 U8335 ( .A(n7333), .ZN(n8685) );
  OAI222_X1 U8336 ( .A1(n8311), .A2(n6608), .B1(n9070), .B2(n6607), .C1(
        P2_U3152), .C2(n8685), .ZN(P2_U3350) );
  INV_X1 U8337 ( .A(n6609), .ZN(n6612) );
  INV_X1 U8338 ( .A(n8706), .ZN(n7335) );
  OAI222_X1 U8339 ( .A1(n8311), .A2(n6610), .B1(n9070), .B2(n6612), .C1(n7335), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  OAI222_X1 U8340 ( .A1(P1_U3084), .A2(n6613), .B1(n9857), .B2(n6612), .C1(
        n6611), .C2(n9859), .ZN(P1_U3344) );
  INV_X1 U8341 ( .A(n7758), .ZN(n7765) );
  INV_X1 U8342 ( .A(n6614), .ZN(n6617) );
  OAI222_X1 U8343 ( .A1(P2_U3152), .A2(n7765), .B1(n9070), .B2(n6617), .C1(
        n6615), .C2(n8311), .ZN(P2_U3348) );
  OAI222_X1 U8344 ( .A1(P1_U3084), .A2(n6742), .B1(n9857), .B2(n6617), .C1(
        n6616), .C2(n9859), .ZN(P1_U3343) );
  INV_X1 U8345 ( .A(n6618), .ZN(n6620) );
  AOI22_X1 U8346 ( .A1(n8711), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n4568), .ZN(n6619) );
  OAI21_X1 U8347 ( .B1(n6620), .B2(n9070), .A(n6619), .ZN(P2_U3347) );
  INV_X1 U8348 ( .A(n7253), .ZN(n7248) );
  OAI222_X1 U8349 ( .A1(P1_U3084), .A2(n7248), .B1(n9857), .B2(n6620), .C1(
        n6878), .C2(n9859), .ZN(P1_U3342) );
  INV_X1 U8350 ( .A(n6621), .ZN(n6624) );
  INV_X1 U8351 ( .A(n7866), .ZN(n7862) );
  OAI222_X1 U8352 ( .A1(n8311), .A2(n6622), .B1(n9070), .B2(n6624), .C1(
        P2_U3152), .C2(n7862), .ZN(P2_U3346) );
  INV_X1 U8353 ( .A(n7791), .ZN(n7784) );
  OAI222_X1 U8354 ( .A1(n7784), .A2(P1_U3084), .B1(n9857), .B2(n6624), .C1(
        n6623), .C2(n9859), .ZN(P1_U3341) );
  INV_X1 U8355 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U8356 ( .A1(n4482), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6630) );
  INV_X1 U8357 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6625) );
  OR2_X1 U8358 ( .A1(n8559), .A2(n6625), .ZN(n6629) );
  INV_X1 U8359 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6626) );
  OR2_X1 U8360 ( .A1(n6627), .A2(n6626), .ZN(n6628) );
  AND3_X1 U8361 ( .A1(n6630), .A2(n6629), .A3(n6628), .ZN(n9312) );
  INV_X1 U8362 ( .A(n9312), .ZN(n9539) );
  NAND2_X1 U8363 ( .A1(n9539), .A2(P1_U4006), .ZN(n6631) );
  OAI21_X1 U8364 ( .B1(P1_U4006), .B2(n6632), .A(n6631), .ZN(P1_U3586) );
  XNOR2_X1 U8365 ( .A(n6634), .B(n6633), .ZN(n6641) );
  INV_X1 U8366 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7359) );
  NAND2_X1 U8367 ( .A1(n10260), .A2(n8681), .ZN(n6636) );
  NAND2_X1 U8368 ( .A1(n10258), .A2(n8679), .ZN(n6635) );
  NAND2_X1 U8369 ( .A1(n6636), .A2(n6635), .ZN(n7216) );
  AOI22_X1 U8370 ( .A1(n8654), .A2(n7216), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3152), .ZN(n6637) );
  OAI21_X1 U8371 ( .B1(n6638), .B2(n8657), .A(n6637), .ZN(n6639) );
  AOI21_X1 U8372 ( .B1(n8639), .B2(n7359), .A(n6639), .ZN(n6640) );
  OAI21_X1 U8373 ( .B1(n8642), .B2(n6641), .A(n6640), .ZN(P2_U3220) );
  OAI22_X1 U8374 ( .A1(n6642), .A2(n8647), .B1(n6688), .B2(n8649), .ZN(n7274)
         );
  INV_X1 U8375 ( .A(n8525), .ZN(n6643) );
  NAND2_X1 U8376 ( .A1(n6644), .A2(n6643), .ZN(n6671) );
  AOI22_X1 U8377 ( .A1(n8654), .A2(n7274), .B1(n6671), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6649) );
  XOR2_X1 U8378 ( .A(n6646), .B(n6645), .Z(n6647) );
  NAND2_X1 U8379 ( .A1(n8631), .A2(n6647), .ZN(n6648) );
  OAI211_X1 U8380 ( .C1(n7279), .C2(n8657), .A(n6649), .B(n6648), .ZN(P2_U3239) );
  OR2_X1 U8381 ( .A1(n10155), .A2(n6284), .ZN(n6653) );
  AND2_X1 U8382 ( .A1(n6651), .A2(n6650), .ZN(n6652) );
  NOR2_X1 U8383 ( .A1(n7917), .A2(n6654), .ZN(n6655) );
  AND2_X2 U8384 ( .A1(n7919), .A2(n6655), .ZN(n10218) );
  INV_X1 U8385 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6660) );
  INV_X1 U8386 ( .A(n7600), .ZN(n7637) );
  INV_X1 U8387 ( .A(n7570), .ZN(n6658) );
  NAND2_X1 U8388 ( .A1(n7637), .A2(n9492), .ZN(n9429) );
  NAND2_X1 U8389 ( .A1(n7630), .A2(n9429), .ZN(n9335) );
  INV_X1 U8390 ( .A(n9207), .ZN(n6656) );
  NOR2_X1 U8391 ( .A1(n6656), .A2(n7570), .ZN(n6657) );
  INV_X1 U8392 ( .A(n7679), .ZN(n9491) );
  AOI22_X1 U8393 ( .A1(n9335), .A2(n6657), .B1(n9735), .B2(n9491), .ZN(n7565)
         );
  OAI21_X1 U8394 ( .B1(n7637), .B2(n6658), .A(n7565), .ZN(n9830) );
  NAND2_X1 U8395 ( .A1(n9830), .A2(n10218), .ZN(n6659) );
  OAI21_X1 U8396 ( .B1(n10218), .B2(n6660), .A(n6659), .ZN(P1_U3454) );
  INV_X1 U8397 ( .A(n6661), .ZN(n6663) );
  INV_X1 U8398 ( .A(n10066), .ZN(n7785) );
  OAI222_X1 U8399 ( .A1(n9859), .A2(n6662), .B1(n9857), .B2(n6663), .C1(
        P1_U3084), .C2(n7785), .ZN(P1_U3340) );
  INV_X1 U8400 ( .A(n7962), .ZN(n7957) );
  OAI222_X1 U8401 ( .A1(n8311), .A2(n6971), .B1(n9070), .B2(n6663), .C1(n7957), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X2 U8402 ( .A(P2_U3966), .ZN(n8682) );
  NAND2_X1 U8403 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n8682), .ZN(n6664) );
  OAI21_X1 U8404 ( .B1(n8605), .B2(n8682), .A(n6664), .ZN(P2_U3576) );
  AOI21_X1 U8405 ( .B1(n6667), .B2(n6666), .A(n6665), .ZN(n6670) );
  AOI22_X1 U8406 ( .A1(n8618), .A2(n7511), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n6671), .ZN(n6669) );
  OAI22_X1 U8407 ( .A1(n5357), .A2(n8649), .B1(n6327), .B2(n8647), .ZN(n7242)
         );
  NAND2_X1 U8408 ( .A1(n8654), .A2(n7242), .ZN(n6668) );
  OAI211_X1 U8409 ( .C1(n6670), .C2(n8642), .A(n6669), .B(n6668), .ZN(P2_U3224) );
  INV_X1 U8410 ( .A(n6671), .ZN(n6678) );
  NAND2_X1 U8411 ( .A1(n8654), .A2(n10258), .ZN(n8584) );
  INV_X1 U8412 ( .A(n8584), .ZN(n8154) );
  AOI22_X1 U8413 ( .A1(n8154), .A2(n6672), .B1(n8618), .B2(n6328), .ZN(n6677)
         );
  INV_X1 U8414 ( .A(n7196), .ZN(n7241) );
  OR2_X1 U8415 ( .A1(n6327), .A2(n6328), .ZN(n8359) );
  INV_X1 U8416 ( .A(n8359), .ZN(n6674) );
  MUX2_X1 U8417 ( .A(n6674), .B(n6328), .S(n6673), .Z(n6675) );
  OAI21_X1 U8418 ( .B1(n7241), .B2(n6675), .A(n8631), .ZN(n6676) );
  OAI211_X1 U8419 ( .C1(n6678), .C2(n7349), .A(n6677), .B(n6676), .ZN(P2_U3234) );
  INV_X1 U8420 ( .A(n7796), .ZN(n9505) );
  INV_X1 U8421 ( .A(n6679), .ZN(n6681) );
  OAI222_X1 U8422 ( .A1(P1_U3084), .A2(n9505), .B1(n9857), .B2(n6681), .C1(
        n6680), .C2(n9859), .ZN(P1_U3339) );
  INV_X1 U8423 ( .A(n8177), .ZN(n8180) );
  OAI222_X1 U8424 ( .A1(n8311), .A2(n6682), .B1(n9070), .B2(n6681), .C1(n8180), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  AOI21_X1 U8425 ( .B1(n6685), .B2(n6684), .A(n6683), .ZN(n6693) );
  INV_X1 U8426 ( .A(n8272), .ZN(n6691) );
  INV_X1 U8427 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6686) );
  OAI22_X1 U8428 ( .A1(n8657), .A2(n10315), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6686), .ZN(n6690) );
  AND2_X1 U8429 ( .A1(n8654), .A2(n10260), .ZN(n8587) );
  INV_X1 U8430 ( .A(n8587), .ZN(n8200) );
  OAI22_X1 U8431 ( .A1(n8200), .A2(n6688), .B1(n6687), .B2(n8584), .ZN(n6689)
         );
  AOI211_X1 U8432 ( .C1(n6691), .C2(n8639), .A(n6690), .B(n6689), .ZN(n6692)
         );
  OAI21_X1 U8433 ( .B1(n6693), .B2(n8642), .A(n6692), .ZN(P2_U3232) );
  XNOR2_X1 U8434 ( .A(n4566), .B(n6694), .ZN(n6699) );
  AOI22_X1 U8435 ( .A1(n10260), .A2(n8679), .B1(n10258), .B2(n8677), .ZN(n7287) );
  OAI22_X1 U8436 ( .A1(n8637), .A2(n7287), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6695), .ZN(n6697) );
  NOR2_X1 U8437 ( .A1(n8652), .A2(n7463), .ZN(n6696) );
  AOI211_X1 U8438 ( .C1(n7302), .C2(n8618), .A(n6697), .B(n6696), .ZN(n6698)
         );
  OAI21_X1 U8439 ( .B1(n6699), .B2(n8642), .A(n6698), .ZN(P2_U3229) );
  OAI21_X1 U8440 ( .B1(n6702), .B2(n6701), .A(n6700), .ZN(n6710) );
  INV_X1 U8441 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n8100) );
  NAND2_X1 U8442 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7442) );
  OAI21_X1 U8443 ( .B1(n10116), .B2(n8100), .A(n7442), .ZN(n6709) );
  AOI21_X1 U8444 ( .B1(n6705), .B2(n6704), .A(n6703), .ZN(n6707) );
  OAI22_X1 U8445 ( .A1(n6707), .A2(n10070), .B1(n10107), .B2(n6706), .ZN(n6708) );
  AOI211_X1 U8446 ( .C1(n10104), .C2(n6710), .A(n6709), .B(n6708), .ZN(n6711)
         );
  INV_X1 U8447 ( .A(n6711), .ZN(P1_U3248) );
  INV_X1 U8448 ( .A(n10116), .ZN(n9983) );
  OAI21_X1 U8449 ( .B1(n6714), .B2(n6713), .A(n6712), .ZN(n6715) );
  OAI22_X1 U8450 ( .A1(n10070), .A2(n6715), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7639), .ZN(n6716) );
  AOI21_X1 U8451 ( .B1(n9983), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n6716), .ZN(
        n6720) );
  OAI211_X1 U8452 ( .C1(n6718), .C2(n9996), .A(n10104), .B(n6717), .ZN(n6719)
         );
  OAI211_X1 U8453 ( .C1(n10107), .C2(n6721), .A(n6720), .B(n6719), .ZN(
        P1_U3242) );
  INV_X1 U8454 ( .A(n10107), .ZN(n10093) );
  AOI21_X1 U8455 ( .B1(n6724), .B2(n6723), .A(n6722), .ZN(n6726) );
  NAND2_X1 U8456 ( .A1(n9983), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U8457 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7540) );
  OAI211_X1 U8458 ( .C1(n6726), .C2(n10070), .A(n6725), .B(n7540), .ZN(n6731)
         );
  AOI211_X1 U8459 ( .C1(n6729), .C2(n6728), .A(n6727), .B(n10086), .ZN(n6730)
         );
  AOI211_X1 U8460 ( .C1(n10093), .C2(n6732), .A(n6731), .B(n6730), .ZN(n6733)
         );
  INV_X1 U8461 ( .A(n6733), .ZN(P1_U3247) );
  NOR2_X1 U8462 ( .A1(n6741), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6735) );
  INV_X1 U8463 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6736) );
  MUX2_X1 U8464 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6736), .S(n6742), .Z(n6753)
         );
  NAND2_X1 U8465 ( .A1(n6742), .A2(n6736), .ZN(n6737) );
  AOI22_X1 U8466 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n7248), .B1(n7253), .B2(
        n6010), .ZN(n6738) );
  NOR2_X1 U8467 ( .A1(n6739), .A2(n6738), .ZN(n7247) );
  AOI21_X1 U8468 ( .B1(n6739), .B2(n6738), .A(n7247), .ZN(n6750) );
  INV_X1 U8469 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7892) );
  XNOR2_X1 U8470 ( .A(n6742), .B(n7892), .ZN(n6757) );
  AOI21_X1 U8471 ( .B1(n6761), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6756), .ZN(
        n6745) );
  INV_X1 U8472 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6743) );
  AOI22_X1 U8473 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7253), .B1(n7248), .B2(
        n6743), .ZN(n6744) );
  NAND2_X1 U8474 ( .A1(n6744), .A2(n6745), .ZN(n7252) );
  OAI21_X1 U8475 ( .B1(n6745), .B2(n6744), .A(n7252), .ZN(n6748) );
  AND2_X1 U8476 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3084), .ZN(n7927) );
  AOI21_X1 U8477 ( .B1(n9983), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7927), .ZN(
        n6746) );
  OAI21_X1 U8478 ( .B1(n7248), .B2(n10107), .A(n6746), .ZN(n6747) );
  AOI21_X1 U8479 ( .B1(n6748), .B2(n10104), .A(n6747), .ZN(n6749) );
  OAI21_X1 U8480 ( .B1(n6750), .B2(n10070), .A(n6749), .ZN(P1_U3252) );
  INV_X1 U8481 ( .A(n6751), .ZN(n6752) );
  AOI21_X1 U8482 ( .B1(n6754), .B2(n6753), .A(n6752), .ZN(n6763) );
  INV_X1 U8483 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6755) );
  NAND2_X1 U8484 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7836) );
  OAI21_X1 U8485 ( .B1(n10116), .B2(n6755), .A(n7836), .ZN(n6760) );
  AOI211_X1 U8486 ( .C1(n6758), .C2(n6757), .A(n10086), .B(n6756), .ZN(n6759)
         );
  AOI211_X1 U8487 ( .C1(n10093), .C2(n6761), .A(n6760), .B(n6759), .ZN(n6762)
         );
  OAI21_X1 U8488 ( .B1(n6763), .B2(n10070), .A(n6762), .ZN(P1_U3251) );
  MUX2_X1 U8489 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n7899), .S(P1_U4006), .Z(
        n7105) );
  OAI22_X1 U8490 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(keyinput8), .B1(
        P2_IR_REG_14__SCAN_IN), .B2(keyinput96), .ZN(n6764) );
  AOI221_X1 U8491 ( .B1(P1_DATAO_REG_0__SCAN_IN), .B2(keyinput8), .C1(
        keyinput96), .C2(P2_IR_REG_14__SCAN_IN), .A(n6764), .ZN(n6771) );
  OAI22_X1 U8492 ( .A1(P1_D_REG_8__SCAN_IN), .A2(keyinput25), .B1(keyinput89), 
        .B2(P1_REG3_REG_22__SCAN_IN), .ZN(n6765) );
  AOI221_X1 U8493 ( .B1(P1_D_REG_8__SCAN_IN), .B2(keyinput25), .C1(
        P1_REG3_REG_22__SCAN_IN), .C2(keyinput89), .A(n6765), .ZN(n6770) );
  OAI22_X1 U8494 ( .A1(P1_D_REG_14__SCAN_IN), .A2(keyinput49), .B1(keyinput120), .B2(P2_D_REG_1__SCAN_IN), .ZN(n6766) );
  AOI221_X1 U8495 ( .B1(P1_D_REG_14__SCAN_IN), .B2(keyinput49), .C1(
        P2_D_REG_1__SCAN_IN), .C2(keyinput120), .A(n6766), .ZN(n6769) );
  OAI22_X1 U8496 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(keyinput15), .B1(
        keyinput16), .B2(SI_1_), .ZN(n6767) );
  AOI221_X1 U8497 ( .B1(P2_DATAO_REG_3__SCAN_IN), .B2(keyinput15), .C1(SI_1_), 
        .C2(keyinput16), .A(n6767), .ZN(n6768) );
  NAND4_X1 U8498 ( .A1(n6771), .A2(n6770), .A3(n6769), .A4(n6768), .ZN(n6799)
         );
  OAI22_X1 U8499 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput38), .B1(keyinput79), .B2(P2_REG3_REG_4__SCAN_IN), .ZN(n6772) );
  AOI221_X1 U8500 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput38), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput79), .A(n6772), .ZN(n6779) );
  OAI22_X1 U8501 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput18), .B1(
        P1_REG0_REG_26__SCAN_IN), .B2(keyinput40), .ZN(n6773) );
  AOI221_X1 U8502 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput18), .C1(
        keyinput40), .C2(P1_REG0_REG_26__SCAN_IN), .A(n6773), .ZN(n6778) );
  OAI22_X1 U8503 ( .A1(P2_REG0_REG_27__SCAN_IN), .A2(keyinput31), .B1(
        P2_REG0_REG_3__SCAN_IN), .B2(keyinput113), .ZN(n6774) );
  AOI221_X1 U8504 ( .B1(P2_REG0_REG_27__SCAN_IN), .B2(keyinput31), .C1(
        keyinput113), .C2(P2_REG0_REG_3__SCAN_IN), .A(n6774), .ZN(n6777) );
  OAI22_X1 U8505 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput122), .B1(
        P2_REG2_REG_18__SCAN_IN), .B2(keyinput55), .ZN(n6775) );
  AOI221_X1 U8506 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput122), .C1(
        keyinput55), .C2(P2_REG2_REG_18__SCAN_IN), .A(n6775), .ZN(n6776) );
  NAND4_X1 U8507 ( .A1(n6779), .A2(n6778), .A3(n6777), .A4(n6776), .ZN(n6798)
         );
  OAI22_X1 U8508 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(keyinput39), .B1(
        P2_ADDR_REG_7__SCAN_IN), .B2(keyinput115), .ZN(n6780) );
  AOI221_X1 U8509 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(keyinput39), .C1(
        keyinput115), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n6780), .ZN(n6787) );
  OAI22_X1 U8510 ( .A1(P2_D_REG_23__SCAN_IN), .A2(keyinput84), .B1(
        P2_REG0_REG_1__SCAN_IN), .B2(keyinput10), .ZN(n6781) );
  AOI221_X1 U8511 ( .B1(P2_D_REG_23__SCAN_IN), .B2(keyinput84), .C1(keyinput10), .C2(P2_REG0_REG_1__SCAN_IN), .A(n6781), .ZN(n6786) );
  OAI22_X1 U8512 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(keyinput72), .B1(
        keyinput77), .B2(P1_ADDR_REG_16__SCAN_IN), .ZN(n6782) );
  AOI221_X1 U8513 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(keyinput72), .C1(
        P1_ADDR_REG_16__SCAN_IN), .C2(keyinput77), .A(n6782), .ZN(n6785) );
  OAI22_X1 U8514 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput34), .B1(
        keyinput41), .B2(P2_REG3_REG_15__SCAN_IN), .ZN(n6783) );
  AOI221_X1 U8515 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput34), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput41), .A(n6783), .ZN(n6784) );
  NAND4_X1 U8516 ( .A1(n6787), .A2(n6786), .A3(n6785), .A4(n6784), .ZN(n6797)
         );
  OAI22_X1 U8517 ( .A1(SI_28_), .A2(keyinput44), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(keyinput100), .ZN(n6788) );
  AOI221_X1 U8518 ( .B1(SI_28_), .B2(keyinput44), .C1(keyinput100), .C2(
        P2_REG2_REG_23__SCAN_IN), .A(n6788), .ZN(n6795) );
  OAI22_X1 U8519 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(keyinput99), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(keyinput112), .ZN(n6789) );
  AOI221_X1 U8520 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(keyinput99), .C1(
        keyinput112), .C2(P2_REG3_REG_1__SCAN_IN), .A(n6789), .ZN(n6794) );
  OAI22_X1 U8521 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(keyinput4), .B1(keyinput30), .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n6790) );
  AOI221_X1 U8522 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(keyinput4), .C1(
        P2_REG1_REG_0__SCAN_IN), .C2(keyinput30), .A(n6790), .ZN(n6793) );
  OAI22_X1 U8523 ( .A1(SI_4_), .A2(keyinput57), .B1(keyinput43), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n6791) );
  AOI221_X1 U8524 ( .B1(SI_4_), .B2(keyinput57), .C1(P2_REG2_REG_25__SCAN_IN), 
        .C2(keyinput43), .A(n6791), .ZN(n6792) );
  NAND4_X1 U8525 ( .A1(n6795), .A2(n6794), .A3(n6793), .A4(n6792), .ZN(n6796)
         );
  NOR4_X1 U8526 ( .A1(n6799), .A2(n6798), .A3(n6797), .A4(n6796), .ZN(n7103)
         );
  AOI22_X1 U8527 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput173), .B1(
        P1_REG0_REG_20__SCAN_IN), .B2(keyinput245), .ZN(n6800) );
  OAI221_X1 U8528 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput173), .C1(
        P1_REG0_REG_20__SCAN_IN), .C2(keyinput245), .A(n6800), .ZN(n6807) );
  AOI22_X1 U8529 ( .A1(P2_REG0_REG_8__SCAN_IN), .A2(keyinput129), .B1(
        P1_REG1_REG_29__SCAN_IN), .B2(keyinput244), .ZN(n6801) );
  OAI221_X1 U8530 ( .B1(P2_REG0_REG_8__SCAN_IN), .B2(keyinput129), .C1(
        P1_REG1_REG_29__SCAN_IN), .C2(keyinput244), .A(n6801), .ZN(n6806) );
  AOI22_X1 U8531 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(keyinput158), .B1(
        P1_REG2_REG_16__SCAN_IN), .B2(keyinput249), .ZN(n6802) );
  OAI221_X1 U8532 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(keyinput158), .C1(
        P1_REG2_REG_16__SCAN_IN), .C2(keyinput249), .A(n6802), .ZN(n6805) );
  AOI22_X1 U8533 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(keyinput227), .B1(
        P1_REG3_REG_14__SCAN_IN), .B2(keyinput222), .ZN(n6803) );
  OAI221_X1 U8534 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(keyinput227), .C1(
        P1_REG3_REG_14__SCAN_IN), .C2(keyinput222), .A(n6803), .ZN(n6804) );
  NOR4_X1 U8535 ( .A1(n6807), .A2(n6806), .A3(n6805), .A4(n6804), .ZN(n6835)
         );
  AOI22_X1 U8536 ( .A1(P2_REG0_REG_25__SCAN_IN), .A2(keyinput213), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(keyinput136), .ZN(n6808) );
  OAI221_X1 U8537 ( .B1(P2_REG0_REG_25__SCAN_IN), .B2(keyinput213), .C1(
        P1_DATAO_REG_0__SCAN_IN), .C2(keyinput136), .A(n6808), .ZN(n6815) );
  AOI22_X1 U8538 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(keyinput230), .B1(
        P2_D_REG_31__SCAN_IN), .B2(keyinput194), .ZN(n6809) );
  OAI221_X1 U8539 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(keyinput230), .C1(
        P2_D_REG_31__SCAN_IN), .C2(keyinput194), .A(n6809), .ZN(n6814) );
  AOI22_X1 U8540 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(keyinput238), .B1(
        P1_REG2_REG_26__SCAN_IN), .B2(keyinput145), .ZN(n6810) );
  OAI221_X1 U8541 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(keyinput238), .C1(
        P1_REG2_REG_26__SCAN_IN), .C2(keyinput145), .A(n6810), .ZN(n6813) );
  AOI22_X1 U8542 ( .A1(P2_D_REG_28__SCAN_IN), .A2(keyinput211), .B1(
        P1_REG0_REG_7__SCAN_IN), .B2(keyinput215), .ZN(n6811) );
  OAI221_X1 U8543 ( .B1(P2_D_REG_28__SCAN_IN), .B2(keyinput211), .C1(
        P1_REG0_REG_7__SCAN_IN), .C2(keyinput215), .A(n6811), .ZN(n6812) );
  NOR4_X1 U8544 ( .A1(n6815), .A2(n6814), .A3(n6813), .A4(n6812), .ZN(n6834)
         );
  AOI22_X1 U8545 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput207), .B1(
        P1_REG2_REG_0__SCAN_IN), .B2(keyinput235), .ZN(n6816) );
  OAI221_X1 U8546 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput207), .C1(
        P1_REG2_REG_0__SCAN_IN), .C2(keyinput235), .A(n6816), .ZN(n6823) );
  AOI22_X1 U8547 ( .A1(SI_7_), .A2(keyinput170), .B1(P1_D_REG_27__SCAN_IN), 
        .B2(keyinput163), .ZN(n6817) );
  OAI221_X1 U8548 ( .B1(SI_7_), .B2(keyinput170), .C1(P1_D_REG_27__SCAN_IN), 
        .C2(keyinput163), .A(n6817), .ZN(n6822) );
  AOI22_X1 U8549 ( .A1(P2_D_REG_23__SCAN_IN), .A2(keyinput212), .B1(
        P1_IR_REG_1__SCAN_IN), .B2(keyinput254), .ZN(n6818) );
  OAI221_X1 U8550 ( .B1(P2_D_REG_23__SCAN_IN), .B2(keyinput212), .C1(
        P1_IR_REG_1__SCAN_IN), .C2(keyinput254), .A(n6818), .ZN(n6821) );
  AOI22_X1 U8551 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput188), .B1(
        P2_D_REG_12__SCAN_IN), .B2(keyinput140), .ZN(n6819) );
  OAI221_X1 U8552 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput188), .C1(
        P2_D_REG_12__SCAN_IN), .C2(keyinput140), .A(n6819), .ZN(n6820) );
  NOR4_X1 U8553 ( .A1(n6823), .A2(n6822), .A3(n6821), .A4(n6820), .ZN(n6833)
         );
  AOI22_X1 U8554 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(keyinput184), .B1(SI_17_), 
        .B2(keyinput206), .ZN(n6824) );
  OAI221_X1 U8555 ( .B1(P1_DATAO_REG_5__SCAN_IN), .B2(keyinput184), .C1(SI_17_), .C2(keyinput206), .A(n6824), .ZN(n6831) );
  AOI22_X1 U8556 ( .A1(P2_REG0_REG_15__SCAN_IN), .A2(keyinput208), .B1(
        P1_REG2_REG_12__SCAN_IN), .B2(keyinput179), .ZN(n6825) );
  OAI221_X1 U8557 ( .B1(P2_REG0_REG_15__SCAN_IN), .B2(keyinput208), .C1(
        P1_REG2_REG_12__SCAN_IN), .C2(keyinput179), .A(n6825), .ZN(n6830) );
  AOI22_X1 U8558 ( .A1(P2_REG2_REG_7__SCAN_IN), .A2(keyinput139), .B1(SI_28_), 
        .B2(keyinput172), .ZN(n6826) );
  OAI221_X1 U8559 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(keyinput139), .C1(SI_28_), 
        .C2(keyinput172), .A(n6826), .ZN(n6829) );
  AOI22_X1 U8560 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(keyinput191), .B1(SI_13_), 
        .B2(keyinput225), .ZN(n6827) );
  OAI221_X1 U8561 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(keyinput191), .C1(SI_13_), .C2(keyinput225), .A(n6827), .ZN(n6828) );
  NOR4_X1 U8562 ( .A1(n6831), .A2(n6830), .A3(n6829), .A4(n6828), .ZN(n6832)
         );
  NAND4_X1 U8563 ( .A1(n6835), .A2(n6834), .A3(n6833), .A4(n6832), .ZN(n6965)
         );
  AOI22_X1 U8564 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(keyinput242), .B1(SI_4_), 
        .B2(keyinput185), .ZN(n6836) );
  OAI221_X1 U8565 ( .B1(P2_IR_REG_8__SCAN_IN), .B2(keyinput242), .C1(SI_4_), 
        .C2(keyinput185), .A(n6836), .ZN(n6843) );
  AOI22_X1 U8566 ( .A1(P2_D_REG_1__SCAN_IN), .A2(keyinput248), .B1(
        P1_REG1_REG_6__SCAN_IN), .B2(keyinput150), .ZN(n6837) );
  OAI221_X1 U8567 ( .B1(P2_D_REG_1__SCAN_IN), .B2(keyinput248), .C1(
        P1_REG1_REG_6__SCAN_IN), .C2(keyinput150), .A(n6837), .ZN(n6842) );
  AOI22_X1 U8568 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(keyinput198), .B1(
        P2_REG2_REG_21__SCAN_IN), .B2(keyinput226), .ZN(n6838) );
  OAI221_X1 U8569 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(keyinput198), .C1(
        P2_REG2_REG_21__SCAN_IN), .C2(keyinput226), .A(n6838), .ZN(n6841) );
  AOI22_X1 U8570 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(keyinput223), .B1(
        P1_D_REG_23__SCAN_IN), .B2(keyinput201), .ZN(n6839) );
  OAI221_X1 U8571 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(keyinput223), .C1(
        P1_D_REG_23__SCAN_IN), .C2(keyinput201), .A(n6839), .ZN(n6840) );
  NOR4_X1 U8572 ( .A1(n6843), .A2(n6842), .A3(n6841), .A4(n6840), .ZN(n6872)
         );
  AOI22_X1 U8573 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(keyinput196), .B1(
        P1_REG1_REG_3__SCAN_IN), .B2(keyinput219), .ZN(n6844) );
  OAI221_X1 U8574 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(keyinput196), .C1(
        P1_REG1_REG_3__SCAN_IN), .C2(keyinput219), .A(n6844), .ZN(n6851) );
  AOI22_X1 U8575 ( .A1(P2_REG0_REG_23__SCAN_IN), .A2(keyinput210), .B1(
        P2_REG2_REG_18__SCAN_IN), .B2(keyinput183), .ZN(n6845) );
  OAI221_X1 U8576 ( .B1(P2_REG0_REG_23__SCAN_IN), .B2(keyinput210), .C1(
        P2_REG2_REG_18__SCAN_IN), .C2(keyinput183), .A(n6845), .ZN(n6850) );
  AOI22_X1 U8577 ( .A1(P2_REG0_REG_1__SCAN_IN), .A2(keyinput138), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput166), .ZN(n6846) );
  OAI221_X1 U8578 ( .B1(P2_REG0_REG_1__SCAN_IN), .B2(keyinput138), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput166), .A(n6846), .ZN(n6849) );
  AOI22_X1 U8579 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(keyinput243), .B1(
        P2_REG1_REG_6__SCAN_IN), .B2(keyinput132), .ZN(n6847) );
  OAI221_X1 U8580 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(keyinput243), .C1(
        P2_REG1_REG_6__SCAN_IN), .C2(keyinput132), .A(n6847), .ZN(n6848) );
  NOR4_X1 U8581 ( .A1(n6851), .A2(n6850), .A3(n6849), .A4(n6848), .ZN(n6871)
         );
  AOI22_X1 U8582 ( .A1(P2_REG0_REG_24__SCAN_IN), .A2(keyinput134), .B1(
        P1_IR_REG_3__SCAN_IN), .B2(keyinput128), .ZN(n6852) );
  OAI221_X1 U8583 ( .B1(P2_REG0_REG_24__SCAN_IN), .B2(keyinput134), .C1(
        P1_IR_REG_3__SCAN_IN), .C2(keyinput128), .A(n6852), .ZN(n6859) );
  AOI22_X1 U8584 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput135), .B1(
        P1_IR_REG_26__SCAN_IN), .B2(keyinput216), .ZN(n6853) );
  OAI221_X1 U8585 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput135), .C1(
        P1_IR_REG_26__SCAN_IN), .C2(keyinput216), .A(n6853), .ZN(n6858) );
  AOI22_X1 U8586 ( .A1(P2_REG0_REG_12__SCAN_IN), .A2(keyinput130), .B1(
        P2_IR_REG_14__SCAN_IN), .B2(keyinput224), .ZN(n6854) );
  OAI221_X1 U8587 ( .B1(P2_REG0_REG_12__SCAN_IN), .B2(keyinput130), .C1(
        P2_IR_REG_14__SCAN_IN), .C2(keyinput224), .A(n6854), .ZN(n6857) );
  AOI22_X1 U8588 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(keyinput203), .B1(
        P2_D_REG_15__SCAN_IN), .B2(keyinput237), .ZN(n6855) );
  OAI221_X1 U8589 ( .B1(P1_DATAO_REG_29__SCAN_IN), .B2(keyinput203), .C1(
        P2_D_REG_15__SCAN_IN), .C2(keyinput237), .A(n6855), .ZN(n6856) );
  NOR4_X1 U8590 ( .A1(n6859), .A2(n6858), .A3(n6857), .A4(n6856), .ZN(n6870)
         );
  AOI22_X1 U8591 ( .A1(P2_REG2_REG_30__SCAN_IN), .A2(keyinput176), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(keyinput187), .ZN(n6860) );
  OAI221_X1 U8592 ( .B1(P2_REG2_REG_30__SCAN_IN), .B2(keyinput176), .C1(
        P2_DATAO_REG_22__SCAN_IN), .C2(keyinput187), .A(n6860), .ZN(n6868) );
  AOI22_X1 U8593 ( .A1(P2_REG2_REG_19__SCAN_IN), .A2(keyinput186), .B1(
        P1_D_REG_31__SCAN_IN), .B2(keyinput192), .ZN(n6861) );
  OAI221_X1 U8594 ( .B1(P2_REG2_REG_19__SCAN_IN), .B2(keyinput186), .C1(
        P1_D_REG_31__SCAN_IN), .C2(keyinput192), .A(n6861), .ZN(n6867) );
  AOI22_X1 U8595 ( .A1(P2_REG2_REG_25__SCAN_IN), .A2(keyinput171), .B1(SI_20_), 
        .B2(keyinput251), .ZN(n6862) );
  OAI221_X1 U8596 ( .B1(P2_REG2_REG_25__SCAN_IN), .B2(keyinput171), .C1(SI_20_), .C2(keyinput251), .A(n6862), .ZN(n6866) );
  XOR2_X1 U8597 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput165), .Z(n6864) );
  XNOR2_X1 U8598 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput156), .ZN(n6863) );
  NAND2_X1 U8599 ( .A1(n6864), .A2(n6863), .ZN(n6865) );
  NOR4_X1 U8600 ( .A1(n6868), .A2(n6867), .A3(n6866), .A4(n6865), .ZN(n6869)
         );
  NAND4_X1 U8601 ( .A1(n6872), .A2(n6871), .A3(n6870), .A4(n6869), .ZN(n6964)
         );
  INV_X1 U8602 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10300) );
  AOI22_X1 U8603 ( .A1(n8276), .A2(keyinput193), .B1(n10300), .B2(keyinput152), 
        .ZN(n6873) );
  OAI221_X1 U8604 ( .B1(n8276), .B2(keyinput193), .C1(n10300), .C2(keyinput152), .A(n6873), .ZN(n6884) );
  AOI22_X1 U8605 ( .A1(n7614), .A2(keyinput220), .B1(n6875), .B2(keyinput202), 
        .ZN(n6874) );
  OAI221_X1 U8606 ( .B1(n7614), .B2(keyinput220), .C1(n6875), .C2(keyinput202), 
        .A(n6874), .ZN(n6883) );
  AOI22_X1 U8607 ( .A1(n6878), .A2(keyinput146), .B1(keyinput148), .B2(n6877), 
        .ZN(n6876) );
  OAI221_X1 U8608 ( .B1(n6878), .B2(keyinput146), .C1(n6877), .C2(keyinput148), 
        .A(n6876), .ZN(n6882) );
  XNOR2_X1 U8609 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput143), .ZN(n6880) );
  XNOR2_X1 U8610 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput250), .ZN(n6879) );
  NAND2_X1 U8611 ( .A1(n6880), .A2(n6879), .ZN(n6881) );
  NOR4_X1 U8612 ( .A1(n6884), .A2(n6883), .A3(n6882), .A4(n6881), .ZN(n6920)
         );
  INV_X1 U8613 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n8105) );
  AOI22_X1 U8614 ( .A1(n8105), .A2(keyinput229), .B1(n6886), .B2(keyinput236), 
        .ZN(n6885) );
  OAI221_X1 U8615 ( .B1(n8105), .B2(keyinput229), .C1(n6886), .C2(keyinput236), 
        .A(n6885), .ZN(n6894) );
  AOI22_X1 U8616 ( .A1(n10308), .A2(keyinput214), .B1(n7000), .B2(keyinput189), 
        .ZN(n6887) );
  OAI221_X1 U8617 ( .B1(n10308), .B2(keyinput214), .C1(n7000), .C2(keyinput189), .A(n6887), .ZN(n6893) );
  INV_X1 U8618 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10301) );
  AOI22_X1 U8619 ( .A1(n8905), .A2(keyinput228), .B1(n10301), .B2(keyinput253), 
        .ZN(n6888) );
  OAI221_X1 U8620 ( .B1(n8905), .B2(keyinput228), .C1(n10301), .C2(keyinput253), .A(n6888), .ZN(n6892) );
  INV_X1 U8621 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6890) );
  AOI22_X1 U8622 ( .A1(n7227), .A2(keyinput155), .B1(keyinput200), .B2(n6890), 
        .ZN(n6889) );
  OAI221_X1 U8623 ( .B1(n7227), .B2(keyinput155), .C1(n6890), .C2(keyinput200), 
        .A(n6889), .ZN(n6891) );
  NOR4_X1 U8624 ( .A1(n6894), .A2(n6893), .A3(n6892), .A4(n6891), .ZN(n6919)
         );
  INV_X1 U8625 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6896) );
  AOI22_X1 U8626 ( .A1(n6897), .A2(keyinput159), .B1(keyinput255), .B2(n6896), 
        .ZN(n6895) );
  OAI221_X1 U8627 ( .B1(n6897), .B2(keyinput159), .C1(n6896), .C2(keyinput255), 
        .A(n6895), .ZN(n6905) );
  AOI22_X1 U8628 ( .A1(n7039), .A2(keyinput149), .B1(keyinput234), .B2(n7639), 
        .ZN(n6898) );
  OAI221_X1 U8629 ( .B1(n7039), .B2(keyinput149), .C1(n7639), .C2(keyinput234), 
        .A(n6898), .ZN(n6904) );
  AOI22_X1 U8630 ( .A1(n9524), .A2(keyinput218), .B1(n6971), .B2(keyinput239), 
        .ZN(n6899) );
  OAI221_X1 U8631 ( .B1(n9524), .B2(keyinput218), .C1(n6971), .C2(keyinput239), 
        .A(n6899), .ZN(n6903) );
  AOI22_X1 U8632 ( .A1(n7767), .A2(keyinput154), .B1(n6901), .B2(keyinput168), 
        .ZN(n6900) );
  OAI221_X1 U8633 ( .B1(n7767), .B2(keyinput154), .C1(n6901), .C2(keyinput168), 
        .A(n6900), .ZN(n6902) );
  NOR4_X1 U8634 ( .A1(n6905), .A2(n6904), .A3(n6903), .A4(n6902), .ZN(n6918)
         );
  INV_X1 U8635 ( .A(SI_1_), .ZN(n6907) );
  AOI22_X1 U8636 ( .A1(n6295), .A2(keyinput204), .B1(n6907), .B2(keyinput144), 
        .ZN(n6906) );
  OAI221_X1 U8637 ( .B1(n6295), .B2(keyinput204), .C1(n6907), .C2(keyinput144), 
        .A(n6906), .ZN(n6916) );
  INV_X1 U8638 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10137) );
  INV_X1 U8639 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10177) );
  AOI22_X1 U8640 ( .A1(n10137), .A2(keyinput177), .B1(keyinput137), .B2(n10177), .ZN(n6908) );
  OAI221_X1 U8641 ( .B1(n10137), .B2(keyinput177), .C1(n10177), .C2(
        keyinput137), .A(n6908), .ZN(n6915) );
  AOI22_X1 U8642 ( .A1(n6010), .A2(keyinput167), .B1(keyinput175), .B2(n6910), 
        .ZN(n6909) );
  OAI221_X1 U8643 ( .B1(n6010), .B2(keyinput167), .C1(n6910), .C2(keyinput175), 
        .A(n6909), .ZN(n6914) );
  INV_X1 U8644 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6980) );
  XOR2_X1 U8645 ( .A(n6980), .B(keyinput174), .Z(n6912) );
  XNOR2_X1 U8646 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput197), .ZN(n6911) );
  NAND2_X1 U8647 ( .A1(n6912), .A2(n6911), .ZN(n6913) );
  NOR4_X1 U8648 ( .A1(n6916), .A2(n6915), .A3(n6914), .A4(n6913), .ZN(n6917)
         );
  NAND4_X1 U8649 ( .A1(n6920), .A2(n6919), .A3(n6918), .A4(n6917), .ZN(n6963)
         );
  INV_X1 U8650 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10143) );
  AOI22_X1 U8651 ( .A1(n8056), .A2(keyinput169), .B1(n10143), .B2(keyinput153), 
        .ZN(n6921) );
  OAI221_X1 U8652 ( .B1(n8056), .B2(keyinput169), .C1(n10143), .C2(keyinput153), .A(n6921), .ZN(n6929) );
  INV_X1 U8653 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8303) );
  INV_X1 U8654 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10099) );
  AOI22_X1 U8655 ( .A1(n8303), .A2(keyinput164), .B1(keyinput205), .B2(n10099), 
        .ZN(n6922) );
  OAI221_X1 U8656 ( .B1(n8303), .B2(keyinput164), .C1(n10099), .C2(keyinput205), .A(n6922), .ZN(n6928) );
  INV_X1 U8657 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n7020) );
  AOI22_X1 U8658 ( .A1(n7506), .A2(keyinput240), .B1(n7020), .B2(keyinput160), 
        .ZN(n6923) );
  OAI221_X1 U8659 ( .B1(n7506), .B2(keyinput240), .C1(n7020), .C2(keyinput160), 
        .A(n6923), .ZN(n6927) );
  INV_X1 U8660 ( .A(SI_18_), .ZN(n6925) );
  AOI22_X1 U8661 ( .A1(n7825), .A2(keyinput182), .B1(keyinput232), .B2(n6925), 
        .ZN(n6924) );
  OAI221_X1 U8662 ( .B1(n7825), .B2(keyinput182), .C1(n6925), .C2(keyinput232), 
        .A(n6924), .ZN(n6926) );
  NOR4_X1 U8663 ( .A1(n6929), .A2(n6928), .A3(n6927), .A4(n6926), .ZN(n6961)
         );
  INV_X1 U8664 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9980) );
  AOI22_X1 U8665 ( .A1(n9980), .A2(keyinput199), .B1(keyinput141), .B2(n10229), 
        .ZN(n6930) );
  OAI221_X1 U8666 ( .B1(n9980), .B2(keyinput199), .C1(n10229), .C2(keyinput141), .A(n6930), .ZN(n6938) );
  INV_X1 U8667 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10135) );
  INV_X1 U8668 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U8669 ( .A1(n10135), .A2(keyinput157), .B1(keyinput246), .B2(n10304), .ZN(n6931) );
  OAI221_X1 U8670 ( .B1(n10135), .B2(keyinput157), .C1(n10304), .C2(
        keyinput246), .A(n6931), .ZN(n6937) );
  INV_X1 U8671 ( .A(P2_B_REG_SCAN_IN), .ZN(n8528) );
  AOI22_X1 U8672 ( .A1(n7953), .A2(keyinput151), .B1(keyinput178), .B2(n8528), 
        .ZN(n6932) );
  OAI221_X1 U8673 ( .B1(n7953), .B2(keyinput151), .C1(n8528), .C2(keyinput178), 
        .A(n6932), .ZN(n6936) );
  XOR2_X1 U8674 ( .A(n5101), .B(keyinput190), .Z(n6934) );
  XNOR2_X1 U8675 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput131), .ZN(n6933) );
  NAND2_X1 U8676 ( .A1(n6934), .A2(n6933), .ZN(n6935) );
  NOR4_X1 U8677 ( .A1(n6938), .A2(n6937), .A3(n6936), .A4(n6935), .ZN(n6960)
         );
  INV_X1 U8678 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U8679 ( .A1(n6940), .A2(keyinput247), .B1(keyinput195), .B2(n10305), 
        .ZN(n6939) );
  OAI221_X1 U8680 ( .B1(n6940), .B2(keyinput247), .C1(n10305), .C2(keyinput195), .A(n6939), .ZN(n6948) );
  AOI22_X1 U8681 ( .A1(n5942), .A2(keyinput180), .B1(keyinput161), .B2(n7173), 
        .ZN(n6941) );
  OAI221_X1 U8682 ( .B1(n5942), .B2(keyinput180), .C1(n7173), .C2(keyinput161), 
        .A(n6941), .ZN(n6947) );
  AOI22_X1 U8683 ( .A1(n7004), .A2(keyinput231), .B1(keyinput241), .B2(n5363), 
        .ZN(n6942) );
  OAI221_X1 U8684 ( .B1(n7004), .B2(keyinput231), .C1(n5363), .C2(keyinput241), 
        .A(n6942), .ZN(n6946) );
  INV_X1 U8685 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10217) );
  XOR2_X1 U8686 ( .A(n10217), .B(keyinput181), .Z(n6944) );
  XNOR2_X1 U8687 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput221), .ZN(n6943) );
  NAND2_X1 U8688 ( .A1(n6944), .A2(n6943), .ZN(n6945) );
  NOR4_X1 U8689 ( .A1(n6948), .A2(n6947), .A3(n6946), .A4(n6945), .ZN(n6959)
         );
  INV_X1 U8690 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10132) );
  AOI22_X1 U8691 ( .A1(n6028), .A2(keyinput209), .B1(n10132), .B2(keyinput252), 
        .ZN(n6949) );
  OAI221_X1 U8692 ( .B1(n6028), .B2(keyinput209), .C1(n10132), .C2(keyinput252), .A(n6949), .ZN(n6957) );
  AOI22_X1 U8693 ( .A1(n8623), .A2(keyinput162), .B1(n8140), .B2(keyinput233), 
        .ZN(n6950) );
  OAI221_X1 U8694 ( .B1(n8623), .B2(keyinput162), .C1(n8140), .C2(keyinput233), 
        .A(n6950), .ZN(n6956) );
  INV_X1 U8695 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U8696 ( .A1(n10306), .A2(keyinput133), .B1(n9160), .B2(keyinput217), 
        .ZN(n6951) );
  OAI221_X1 U8697 ( .B1(n10306), .B2(keyinput133), .C1(n9160), .C2(keyinput217), .A(n6951), .ZN(n6955) );
  XNOR2_X1 U8698 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput147), .ZN(n6953) );
  XNOR2_X1 U8699 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput142), .ZN(n6952)
         );
  NAND2_X1 U8700 ( .A1(n6953), .A2(n6952), .ZN(n6954) );
  NOR4_X1 U8701 ( .A1(n6957), .A2(n6956), .A3(n6955), .A4(n6954), .ZN(n6958)
         );
  NAND4_X1 U8702 ( .A1(n6961), .A2(n6960), .A3(n6959), .A4(n6958), .ZN(n6962)
         );
  NOR4_X1 U8703 ( .A1(n6965), .A2(n6964), .A3(n6963), .A4(n6962), .ZN(n7064)
         );
  AOI22_X1 U8704 ( .A1(P2_REG0_REG_25__SCAN_IN), .A2(keyinput85), .B1(
        P2_D_REG_7__SCAN_IN), .B2(keyinput67), .ZN(n6966) );
  OAI221_X1 U8705 ( .B1(P2_REG0_REG_25__SCAN_IN), .B2(keyinput85), .C1(
        P2_D_REG_7__SCAN_IN), .C2(keyinput67), .A(n6966), .ZN(n6975) );
  AOI22_X1 U8706 ( .A1(n10304), .A2(keyinput118), .B1(n5101), .B2(keyinput62), 
        .ZN(n6967) );
  OAI221_X1 U8707 ( .B1(n10304), .B2(keyinput118), .C1(n5101), .C2(keyinput62), 
        .A(n6967), .ZN(n6974) );
  INV_X1 U8708 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6969) );
  INV_X1 U8709 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10299) );
  AOI22_X1 U8710 ( .A1(n6969), .A2(keyinput11), .B1(n10299), .B2(keyinput83), 
        .ZN(n6968) );
  OAI221_X1 U8711 ( .B1(n6969), .B2(keyinput11), .C1(n10299), .C2(keyinput83), 
        .A(n6968), .ZN(n6973) );
  AOI22_X1 U8712 ( .A1(n6971), .A2(keyinput111), .B1(keyinput36), .B2(n8303), 
        .ZN(n6970) );
  OAI221_X1 U8713 ( .B1(n6971), .B2(keyinput111), .C1(n8303), .C2(keyinput36), 
        .A(n6970), .ZN(n6972) );
  NOR4_X1 U8714 ( .A1(n6975), .A2(n6974), .A3(n6973), .A4(n6972), .ZN(n7013)
         );
  INV_X1 U8715 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10120) );
  AOI22_X1 U8716 ( .A1(n10120), .A2(keyinput64), .B1(keyinput17), .B2(n6977), 
        .ZN(n6976) );
  OAI221_X1 U8717 ( .B1(n10120), .B2(keyinput64), .C1(n6977), .C2(keyinput17), 
        .A(n6976), .ZN(n6985) );
  AOI22_X1 U8718 ( .A1(n5521), .A2(keyinput98), .B1(keyinput58), .B2(n8778), 
        .ZN(n6978) );
  OAI221_X1 U8719 ( .B1(n5521), .B2(keyinput98), .C1(n8778), .C2(keyinput58), 
        .A(n6978), .ZN(n6984) );
  AOI22_X1 U8720 ( .A1(n6980), .A2(keyinput46), .B1(n7359), .B2(keyinput37), 
        .ZN(n6979) );
  OAI221_X1 U8721 ( .B1(n6980), .B2(keyinput46), .C1(n7359), .C2(keyinput37), 
        .A(n6979), .ZN(n6983) );
  AOI22_X1 U8722 ( .A1(n8105), .A2(keyinput101), .B1(n7953), .B2(keyinput23), 
        .ZN(n6981) );
  OAI221_X1 U8723 ( .B1(n8105), .B2(keyinput101), .C1(n7953), .C2(keyinput23), 
        .A(n6981), .ZN(n6982) );
  NOR4_X1 U8724 ( .A1(n6985), .A2(n6984), .A3(n6983), .A4(n6982), .ZN(n7012)
         );
  AOI22_X1 U8725 ( .A1(n7614), .A2(keyinput92), .B1(keyinput1), .B2(n5321), 
        .ZN(n6986) );
  OAI221_X1 U8726 ( .B1(n7614), .B2(keyinput92), .C1(n5321), .C2(keyinput1), 
        .A(n6986), .ZN(n6998) );
  AOI22_X1 U8727 ( .A1(n6989), .A2(keyinput117), .B1(keyinput80), .B2(n6988), 
        .ZN(n6987) );
  OAI221_X1 U8728 ( .B1(n6989), .B2(keyinput117), .C1(n6988), .C2(keyinput80), 
        .A(n6987), .ZN(n6997) );
  AOI22_X1 U8729 ( .A1(n6992), .A2(keyinput56), .B1(n6991), .B2(keyinput123), 
        .ZN(n6990) );
  OAI221_X1 U8730 ( .B1(n6992), .B2(keyinput56), .C1(n6991), .C2(keyinput123), 
        .A(n6990), .ZN(n6996) );
  XNOR2_X1 U8731 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput88), .ZN(n6994) );
  XNOR2_X1 U8732 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput119), .ZN(n6993) );
  NAND2_X1 U8733 ( .A1(n6994), .A2(n6993), .ZN(n6995) );
  NOR4_X1 U8734 ( .A1(n6998), .A2(n6997), .A3(n6996), .A4(n6995), .ZN(n7011)
         );
  INV_X1 U8735 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U8736 ( .A1(n10303), .A2(keyinput12), .B1(n7000), .B2(keyinput61), 
        .ZN(n6999) );
  OAI221_X1 U8737 ( .B1(n10303), .B2(keyinput12), .C1(n7000), .C2(keyinput61), 
        .A(n6999), .ZN(n7009) );
  INV_X1 U8738 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7002) );
  AOI22_X1 U8739 ( .A1(n7002), .A2(keyinput51), .B1(keyinput60), .B2(n7349), 
        .ZN(n7001) );
  OAI221_X1 U8740 ( .B1(n7002), .B2(keyinput51), .C1(n7349), .C2(keyinput60), 
        .A(n7001), .ZN(n7008) );
  AOI22_X1 U8741 ( .A1(n10177), .A2(keyinput9), .B1(n7004), .B2(keyinput103), 
        .ZN(n7003) );
  OAI221_X1 U8742 ( .B1(n10177), .B2(keyinput9), .C1(n7004), .C2(keyinput103), 
        .A(n7003), .ZN(n7007) );
  AOI22_X1 U8743 ( .A1(n10222), .A2(keyinput91), .B1(n6028), .B2(keyinput81), 
        .ZN(n7005) );
  OAI221_X1 U8744 ( .B1(n10222), .B2(keyinput91), .C1(n6028), .C2(keyinput81), 
        .A(n7005), .ZN(n7006) );
  NOR4_X1 U8745 ( .A1(n7009), .A2(n7008), .A3(n7007), .A4(n7006), .ZN(n7010)
         );
  NAND4_X1 U8746 ( .A1(n7013), .A2(n7012), .A3(n7011), .A4(n7010), .ZN(n7063)
         );
  AOI22_X1 U8747 ( .A1(n8140), .A2(keyinput105), .B1(n10132), .B2(keyinput124), 
        .ZN(n7014) );
  OAI221_X1 U8748 ( .B1(n8140), .B2(keyinput105), .C1(n10132), .C2(keyinput124), .A(n7014), .ZN(n7026) );
  INV_X1 U8749 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7016) );
  AOI22_X1 U8750 ( .A1(n7016), .A2(keyinput102), .B1(n7639), .B2(keyinput106), 
        .ZN(n7015) );
  OAI221_X1 U8751 ( .B1(n7016), .B2(keyinput102), .C1(n7639), .C2(keyinput106), 
        .A(n7015), .ZN(n7025) );
  AOI22_X1 U8752 ( .A1(n7019), .A2(keyinput82), .B1(n7018), .B2(keyinput42), 
        .ZN(n7017) );
  OAI221_X1 U8753 ( .B1(n7019), .B2(keyinput82), .C1(n7018), .C2(keyinput42), 
        .A(n7017), .ZN(n7024) );
  XOR2_X1 U8754 ( .A(n7020), .B(keyinput32), .Z(n7022) );
  XNOR2_X1 U8755 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput126), .ZN(n7021) );
  NAND2_X1 U8756 ( .A1(n7022), .A2(n7021), .ZN(n7023) );
  NOR4_X1 U8757 ( .A1(n7026), .A2(n7025), .A3(n7024), .A4(n7023), .ZN(n7061)
         );
  AOI22_X1 U8758 ( .A1(n10135), .A2(keyinput29), .B1(keyinput107), .B2(n7573), 
        .ZN(n7027) );
  OAI221_X1 U8759 ( .B1(n10135), .B2(keyinput29), .C1(n7573), .C2(keyinput107), 
        .A(n7027), .ZN(n7036) );
  INV_X1 U8760 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n7029) );
  AOI22_X1 U8761 ( .A1(n5918), .A2(keyinput87), .B1(keyinput48), .B2(n7029), 
        .ZN(n7028) );
  OAI221_X1 U8762 ( .B1(n5918), .B2(keyinput87), .C1(n7029), .C2(keyinput48), 
        .A(n7028), .ZN(n7035) );
  XNOR2_X1 U8763 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput93), .ZN(n7032) );
  XNOR2_X1 U8764 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput14), .ZN(n7031) );
  XNOR2_X1 U8765 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput114), .ZN(n7030) );
  NAND3_X1 U8766 ( .A1(n7032), .A2(n7031), .A3(n7030), .ZN(n7034) );
  INV_X1 U8767 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10302) );
  XNOR2_X1 U8768 ( .A(n10302), .B(keyinput109), .ZN(n7033) );
  NOR4_X1 U8769 ( .A1(n7036), .A2(n7035), .A3(n7034), .A4(n7033), .ZN(n7060)
         );
  AOI22_X1 U8770 ( .A1(n10301), .A2(keyinput125), .B1(n10229), .B2(keyinput13), 
        .ZN(n7037) );
  OAI221_X1 U8771 ( .B1(n10301), .B2(keyinput125), .C1(n10229), .C2(keyinput13), .A(n7037), .ZN(n7046) );
  INV_X1 U8772 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10128) );
  AOI22_X1 U8773 ( .A1(n7039), .A2(keyinput21), .B1(keyinput73), .B2(n10128), 
        .ZN(n7038) );
  OAI221_X1 U8774 ( .B1(n7039), .B2(keyinput21), .C1(n10128), .C2(keyinput73), 
        .A(n7038), .ZN(n7045) );
  AOI22_X1 U8775 ( .A1(n9980), .A2(keyinput71), .B1(n8213), .B2(keyinput121), 
        .ZN(n7040) );
  OAI221_X1 U8776 ( .B1(n9980), .B2(keyinput71), .C1(n8213), .C2(keyinput121), 
        .A(n7040), .ZN(n7044) );
  XNOR2_X1 U8777 ( .A(P1_REG1_REG_29__SCAN_IN), .B(keyinput116), .ZN(n7042) );
  XNOR2_X1 U8778 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput69), .ZN(n7041) );
  NAND2_X1 U8779 ( .A1(n7042), .A2(n7041), .ZN(n7043) );
  NOR4_X1 U8780 ( .A1(n7046), .A2(n7045), .A3(n7044), .A4(n7043), .ZN(n7059)
         );
  INV_X1 U8781 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U8782 ( .A1(n10425), .A2(keyinput110), .B1(n10227), .B2(keyinput22), 
        .ZN(n7047) );
  OAI221_X1 U8783 ( .B1(n10425), .B2(keyinput110), .C1(n10227), .C2(keyinput22), .A(n7047), .ZN(n7057) );
  INV_X1 U8784 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7049) );
  AOI22_X1 U8785 ( .A1(n7825), .A2(keyinput54), .B1(keyinput63), .B2(n7049), 
        .ZN(n7048) );
  OAI221_X1 U8786 ( .B1(n7825), .B2(keyinput54), .C1(n7049), .C2(keyinput63), 
        .A(n7048), .ZN(n7056) );
  AOI22_X1 U8787 ( .A1(n7051), .A2(keyinput78), .B1(keyinput90), .B2(n9524), 
        .ZN(n7050) );
  OAI221_X1 U8788 ( .B1(n7051), .B2(keyinput78), .C1(n9524), .C2(keyinput90), 
        .A(n7050), .ZN(n7055) );
  XNOR2_X1 U8789 ( .A(P2_REG0_REG_21__SCAN_IN), .B(keyinput74), .ZN(n7053) );
  XNOR2_X1 U8790 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput19), .ZN(n7052) );
  NAND2_X1 U8791 ( .A1(n7053), .A2(n7052), .ZN(n7054) );
  NOR4_X1 U8792 ( .A1(n7057), .A2(n7056), .A3(n7055), .A4(n7054), .ZN(n7058)
         );
  NAND4_X1 U8793 ( .A1(n7061), .A2(n7060), .A3(n7059), .A4(n7058), .ZN(n7062)
         );
  NOR3_X1 U8794 ( .A1(n7064), .A2(n7063), .A3(n7062), .ZN(n7102) );
  OAI22_X1 U8795 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput45), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(keyinput127), .ZN(n7065) );
  AOI221_X1 U8796 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput45), .C1(
        keyinput127), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n7065), .ZN(n7072) );
  OAI22_X1 U8797 ( .A1(P2_B_REG_SCAN_IN), .A2(keyinput50), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(keyinput75), .ZN(n7066) );
  AOI221_X1 U8798 ( .B1(P2_B_REG_SCAN_IN), .B2(keyinput50), .C1(keyinput75), 
        .C2(P1_DATAO_REG_29__SCAN_IN), .A(n7066), .ZN(n7071) );
  OAI22_X1 U8799 ( .A1(P1_D_REG_27__SCAN_IN), .A2(keyinput35), .B1(SI_29_), 
        .B2(keyinput65), .ZN(n7067) );
  AOI221_X1 U8800 ( .B1(P1_D_REG_27__SCAN_IN), .B2(keyinput35), .C1(keyinput65), .C2(SI_29_), .A(n7067), .ZN(n7070) );
  OAI22_X1 U8801 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput7), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(keyinput59), .ZN(n7068) );
  AOI221_X1 U8802 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput7), .C1(keyinput59), 
        .C2(P2_DATAO_REG_22__SCAN_IN), .A(n7068), .ZN(n7069) );
  NAND4_X1 U8803 ( .A1(n7072), .A2(n7071), .A3(n7070), .A4(n7069), .ZN(n7100)
         );
  OAI22_X1 U8804 ( .A1(P1_REG0_REG_16__SCAN_IN), .A2(keyinput108), .B1(
        P2_REG0_REG_12__SCAN_IN), .B2(keyinput2), .ZN(n7073) );
  AOI221_X1 U8805 ( .B1(P1_REG0_REG_16__SCAN_IN), .B2(keyinput108), .C1(
        keyinput2), .C2(P2_REG0_REG_12__SCAN_IN), .A(n7073), .ZN(n7080) );
  OAI22_X1 U8806 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(keyinput68), .B1(
        P2_ADDR_REG_16__SCAN_IN), .B2(keyinput70), .ZN(n7074) );
  AOI221_X1 U8807 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(keyinput68), .C1(
        keyinput70), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n7074), .ZN(n7079) );
  OAI22_X1 U8808 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(keyinput3), .B1(
        keyinput20), .B2(P1_REG3_REG_17__SCAN_IN), .ZN(n7075) );
  AOI221_X1 U8809 ( .B1(P1_DATAO_REG_2__SCAN_IN), .B2(keyinput3), .C1(
        P1_REG3_REG_17__SCAN_IN), .C2(keyinput20), .A(n7075), .ZN(n7078) );
  OAI22_X1 U8810 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput0), .B1(
        P2_REG1_REG_12__SCAN_IN), .B2(keyinput26), .ZN(n7076) );
  AOI221_X1 U8811 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput0), .C1(keyinput26), 
        .C2(P2_REG1_REG_12__SCAN_IN), .A(n7076), .ZN(n7077) );
  NAND4_X1 U8812 ( .A1(n7080), .A2(n7079), .A3(n7078), .A4(n7077), .ZN(n7099)
         );
  OAI22_X1 U8813 ( .A1(SI_18_), .A2(keyinput104), .B1(P2_REG0_REG_24__SCAN_IN), 
        .B2(keyinput6), .ZN(n7081) );
  AOI221_X1 U8814 ( .B1(SI_18_), .B2(keyinput104), .C1(keyinput6), .C2(
        P2_REG0_REG_24__SCAN_IN), .A(n7081), .ZN(n7088) );
  OAI22_X1 U8815 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(keyinput94), .B1(
        keyinput86), .B2(P2_D_REG_0__SCAN_IN), .ZN(n7082) );
  AOI221_X1 U8816 ( .B1(P1_REG3_REG_14__SCAN_IN), .B2(keyinput94), .C1(
        P2_D_REG_0__SCAN_IN), .C2(keyinput86), .A(n7082), .ZN(n7087) );
  OAI22_X1 U8817 ( .A1(SI_13_), .A2(keyinput97), .B1(P2_D_REG_31__SCAN_IN), 
        .B2(keyinput66), .ZN(n7083) );
  AOI221_X1 U8818 ( .B1(SI_13_), .B2(keyinput97), .C1(keyinput66), .C2(
        P2_D_REG_31__SCAN_IN), .A(n7083), .ZN(n7086) );
  OAI22_X1 U8819 ( .A1(P2_REG1_REG_7__SCAN_IN), .A2(keyinput33), .B1(
        P2_ADDR_REG_12__SCAN_IN), .B2(keyinput95), .ZN(n7084) );
  AOI221_X1 U8820 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(keyinput33), .C1(
        keyinput95), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n7084), .ZN(n7085) );
  NAND4_X1 U8821 ( .A1(n7088), .A2(n7087), .A3(n7086), .A4(n7085), .ZN(n7098)
         );
  OAI22_X1 U8822 ( .A1(P1_REG0_REG_9__SCAN_IN), .A2(keyinput53), .B1(
        keyinput52), .B2(P1_REG0_REG_8__SCAN_IN), .ZN(n7089) );
  AOI221_X1 U8823 ( .B1(P1_REG0_REG_9__SCAN_IN), .B2(keyinput53), .C1(
        P1_REG0_REG_8__SCAN_IN), .C2(keyinput52), .A(n7089), .ZN(n7096) );
  OAI22_X1 U8824 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(keyinput27), .B1(
        P2_IR_REG_3__SCAN_IN), .B2(keyinput47), .ZN(n7090) );
  AOI221_X1 U8825 ( .B1(P1_DATAO_REG_16__SCAN_IN), .B2(keyinput27), .C1(
        keyinput47), .C2(P2_IR_REG_3__SCAN_IN), .A(n7090), .ZN(n7095) );
  OAI22_X1 U8826 ( .A1(P1_REG2_REG_27__SCAN_IN), .A2(keyinput76), .B1(
        keyinput5), .B2(P2_D_REG_4__SCAN_IN), .ZN(n7091) );
  AOI221_X1 U8827 ( .B1(P1_REG2_REG_27__SCAN_IN), .B2(keyinput76), .C1(
        P2_D_REG_4__SCAN_IN), .C2(keyinput5), .A(n7091), .ZN(n7094) );
  OAI22_X1 U8828 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(keyinput28), .B1(
        P2_D_REG_21__SCAN_IN), .B2(keyinput24), .ZN(n7092) );
  AOI221_X1 U8829 ( .B1(P2_DATAO_REG_1__SCAN_IN), .B2(keyinput28), .C1(
        keyinput24), .C2(P2_D_REG_21__SCAN_IN), .A(n7092), .ZN(n7093) );
  NAND4_X1 U8830 ( .A1(n7096), .A2(n7095), .A3(n7094), .A4(n7093), .ZN(n7097)
         );
  NOR4_X1 U8831 ( .A1(n7100), .A2(n7099), .A3(n7098), .A4(n7097), .ZN(n7101)
         );
  NAND3_X1 U8832 ( .A1(n7103), .A2(n7102), .A3(n7101), .ZN(n7104) );
  XNOR2_X1 U8833 ( .A(n7105), .B(n7104), .ZN(P1_U3565) );
  INV_X1 U8834 ( .A(n8254), .ZN(n7109) );
  INV_X1 U8835 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7350) );
  NOR3_X1 U8836 ( .A1(n10246), .A2(n7350), .A3(n9876), .ZN(n9875) );
  AOI21_X1 U8837 ( .B1(n9879), .B2(P2_REG2_REG_1__SCAN_IN), .A(n9875), .ZN(
        n9890) );
  NAND2_X1 U8838 ( .A1(n9892), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7106) );
  OAI21_X1 U8839 ( .B1(n9892), .B2(P2_REG2_REG_2__SCAN_IN), .A(n7106), .ZN(
        n9889) );
  NOR2_X1 U8840 ( .A1(n9890), .A2(n9889), .ZN(n9888) );
  INV_X1 U8841 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7107) );
  MUX2_X1 U8842 ( .A(n7107), .B(P2_REG2_REG_3__SCAN_IN), .S(n8254), .Z(n7108)
         );
  INV_X1 U8843 ( .A(n7108), .ZN(n7182) );
  NOR2_X1 U8844 ( .A1(n7183), .A2(n7182), .ZN(n7181) );
  AOI21_X1 U8845 ( .B1(n7109), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7181), .ZN(
        n7118) );
  INV_X1 U8846 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7110) );
  MUX2_X1 U8847 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7110), .S(n7146), .Z(n7117)
         );
  NOR2_X1 U8848 ( .A1(n7118), .A2(n7117), .ZN(n7135) );
  OR2_X1 U8849 ( .A1(n5661), .A2(P2_U3152), .ZN(n8115) );
  OR2_X1 U8850 ( .A1(n7112), .A2(n7111), .ZN(n7113) );
  OAI211_X1 U8851 ( .C1(n7114), .C2(n8115), .A(n7113), .B(n8530), .ZN(n7128)
         );
  NAND2_X1 U8852 ( .A1(n7128), .A2(n7126), .ZN(n7115) );
  NAND2_X1 U8853 ( .A1(n7115), .A2(n8682), .ZN(n7119) );
  OR2_X1 U8854 ( .A1(n5661), .A2(n8301), .ZN(n8523) );
  INV_X1 U8855 ( .A(n8523), .ZN(n7116) );
  AOI211_X1 U8856 ( .C1(n7118), .C2(n7117), .A(n7135), .B(n9887), .ZN(n7134)
         );
  NAND2_X1 U8857 ( .A1(n7119), .A2(n5661), .ZN(n10239) );
  AND2_X1 U8858 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7120) );
  AOI21_X1 U8859 ( .B1(n10243), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n7120), .ZN(
        n7132) );
  INV_X1 U8860 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7224) );
  MUX2_X1 U8861 ( .A(n7224), .B(P2_REG1_REG_3__SCAN_IN), .S(n8254), .Z(n7186)
         );
  NAND2_X1 U8862 ( .A1(n9892), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7125) );
  MUX2_X1 U8863 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n7121), .S(n9892), .Z(n9895)
         );
  NAND2_X1 U8864 ( .A1(n9879), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7124) );
  INV_X1 U8865 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7123) );
  MUX2_X1 U8866 ( .A(n7123), .B(P2_REG1_REG_1__SCAN_IN), .S(n7122), .Z(n9882)
         );
  NAND3_X1 U8867 ( .A1(n4579), .A2(P2_REG1_REG_0__SCAN_IN), .A3(n9882), .ZN(
        n9881) );
  NAND2_X1 U8868 ( .A1(n7124), .A2(n9881), .ZN(n9896) );
  NAND2_X1 U8869 ( .A1(n9895), .A2(n9896), .ZN(n9894) );
  NAND2_X1 U8870 ( .A1(n7125), .A2(n9894), .ZN(n7187) );
  NAND2_X1 U8871 ( .A1(n7186), .A2(n7187), .ZN(n7185) );
  OAI21_X1 U8872 ( .B1(n8254), .B2(n7224), .A(n7185), .ZN(n7130) );
  MUX2_X1 U8873 ( .A(n5384), .B(P2_REG1_REG_4__SCAN_IN), .S(n7146), .Z(n7129)
         );
  AND2_X1 U8874 ( .A1(n7126), .A2(n8301), .ZN(n7127) );
  NAND2_X1 U8875 ( .A1(n7128), .A2(n7127), .ZN(n10241) );
  INV_X1 U8876 ( .A(n10241), .ZN(n10237) );
  NAND2_X1 U8877 ( .A1(n7129), .A2(n7130), .ZN(n7145) );
  OAI211_X1 U8878 ( .C1(n7130), .C2(n7129), .A(n10237), .B(n7145), .ZN(n7131)
         );
  OAI211_X1 U8879 ( .C1(n10239), .C2(n7146), .A(n7132), .B(n7131), .ZN(n7133)
         );
  OR2_X1 U8880 ( .A1(n7134), .A2(n7133), .ZN(P2_U3249) );
  INV_X1 U8881 ( .A(n7146), .ZN(n7136) );
  NAND2_X1 U8882 ( .A1(n7143), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7137) );
  OAI21_X1 U8883 ( .B1(n7143), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7137), .ZN(
        n7156) );
  NOR2_X1 U8884 ( .A1(n7157), .A2(n7156), .ZN(n7155) );
  INV_X1 U8885 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7138) );
  MUX2_X1 U8886 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7138), .S(n7168), .Z(n7139)
         );
  INV_X1 U8887 ( .A(n7139), .ZN(n7140) );
  AOI211_X1 U8888 ( .C1(n7141), .C2(n7140), .A(n7167), .B(n9887), .ZN(n7154)
         );
  INV_X1 U8889 ( .A(n7168), .ZN(n8260) );
  NOR2_X1 U8890 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7233), .ZN(n7142) );
  AOI21_X1 U8891 ( .B1(n10243), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7142), .ZN(
        n7152) );
  NAND2_X1 U8892 ( .A1(n7143), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7147) );
  MUX2_X1 U8893 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n7144), .S(n7143), .Z(n7160)
         );
  OAI21_X1 U8894 ( .B1(n7146), .B2(n5384), .A(n7145), .ZN(n7161) );
  NAND2_X1 U8895 ( .A1(n7160), .A2(n7161), .ZN(n7159) );
  NAND2_X1 U8896 ( .A1(n7147), .A2(n7159), .ZN(n7150) );
  MUX2_X1 U8897 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7148), .S(n7168), .Z(n7149)
         );
  NAND2_X1 U8898 ( .A1(n7149), .A2(n7150), .ZN(n7172) );
  OAI211_X1 U8899 ( .C1(n7150), .C2(n7149), .A(n10237), .B(n7172), .ZN(n7151)
         );
  OAI211_X1 U8900 ( .C1(n10239), .C2(n8260), .A(n7152), .B(n7151), .ZN(n7153)
         );
  OR2_X1 U8901 ( .A1(n7154), .A2(n7153), .ZN(P2_U3251) );
  AOI211_X1 U8902 ( .C1(n7157), .C2(n7156), .A(n7155), .B(n9887), .ZN(n7166)
         );
  AND2_X1 U8903 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7158) );
  AOI21_X1 U8904 ( .B1(n10243), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7158), .ZN(
        n7163) );
  OAI211_X1 U8905 ( .C1(n7161), .C2(n7160), .A(n10237), .B(n7159), .ZN(n7162)
         );
  OAI211_X1 U8906 ( .C1(n10239), .C2(n7164), .A(n7163), .B(n7162), .ZN(n7165)
         );
  OR2_X1 U8907 ( .A1(n7166), .A2(n7165), .ZN(P2_U3250) );
  NAND2_X1 U8908 ( .A1(n7330), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7169) );
  OAI21_X1 U8909 ( .B1(n7330), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7169), .ZN(
        n7170) );
  AOI211_X1 U8910 ( .C1(n7171), .C2(n7170), .A(n7322), .B(n9887), .ZN(n7180)
         );
  AND2_X1 U8911 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7313) );
  AOI21_X1 U8912 ( .B1(n10243), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7313), .ZN(
        n7177) );
  OAI21_X1 U8913 ( .B1(n8260), .B2(n7148), .A(n7172), .ZN(n7175) );
  MUX2_X1 U8914 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7173), .S(n7330), .Z(n7174)
         );
  NAND2_X1 U8915 ( .A1(n7174), .A2(n7175), .ZN(n7331) );
  OAI211_X1 U8916 ( .C1(n7175), .C2(n7174), .A(n10237), .B(n7331), .ZN(n7176)
         );
  OAI211_X1 U8917 ( .C1(n10239), .C2(n7178), .A(n7177), .B(n7176), .ZN(n7179)
         );
  OR2_X1 U8918 ( .A1(n7180), .A2(n7179), .ZN(P2_U3252) );
  AOI211_X1 U8919 ( .C1(n7183), .C2(n7182), .A(n7181), .B(n9887), .ZN(n7191)
         );
  NOR2_X1 U8920 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7359), .ZN(n7184) );
  AOI21_X1 U8921 ( .B1(n10243), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7184), .ZN(
        n7189) );
  OAI211_X1 U8922 ( .C1(n7187), .C2(n7186), .A(n10237), .B(n7185), .ZN(n7188)
         );
  OAI211_X1 U8923 ( .C1(n10239), .C2(n8254), .A(n7189), .B(n7188), .ZN(n7190)
         );
  OR2_X1 U8924 ( .A1(n7191), .A2(n7190), .ZN(P2_U3248) );
  INV_X1 U8925 ( .A(n7192), .ZN(n7195) );
  INV_X1 U8926 ( .A(n8726), .ZN(n8735) );
  OAI222_X1 U8927 ( .A1(n8311), .A2(n7193), .B1(n9070), .B2(n7195), .C1(
        P2_U3152), .C2(n8735), .ZN(P2_U3343) );
  INV_X1 U8928 ( .A(n10080), .ZN(n9509) );
  OAI222_X1 U8929 ( .A1(n9509), .A2(P1_U3084), .B1(n9857), .B2(n7195), .C1(
        n7194), .C2(n9859), .ZN(P1_U3338) );
  NAND2_X1 U8930 ( .A1(n8359), .A2(n7196), .ZN(n7343) );
  INV_X1 U8931 ( .A(n9910), .ZN(n10278) );
  AND2_X1 U8932 ( .A1(n10258), .A2(n6672), .ZN(n7197) );
  AOI21_X1 U8933 ( .B1(n7343), .B2(n10278), .A(n7197), .ZN(n7348) );
  AOI22_X1 U8934 ( .A1(n7343), .A2(n10368), .B1(n5711), .B2(n6328), .ZN(n7198)
         );
  NAND2_X1 U8935 ( .A1(n7348), .A2(n7198), .ZN(n9031) );
  NAND2_X1 U8936 ( .A1(n10371), .A2(n9031), .ZN(n7199) );
  OAI21_X1 U8937 ( .B1(n10371), .B2(n5341), .A(n7199), .ZN(P2_U3451) );
  INV_X1 U8938 ( .A(n7200), .ZN(n7226) );
  AOI22_X1 U8939 ( .A1(n10092), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n7201), .ZN(n7202) );
  OAI21_X1 U8940 ( .B1(n7226), .B2(n9857), .A(n7202), .ZN(P1_U3337) );
  XNOR2_X1 U8941 ( .A(n7204), .B(n7203), .ZN(n9997) );
  NOR2_X1 U8942 ( .A1(n7205), .A2(n7917), .ZN(n7206) );
  OR2_X1 U8943 ( .A1(n9205), .A2(n7206), .ZN(n9171) );
  INV_X1 U8944 ( .A(n9171), .ZN(n7208) );
  INV_X1 U8945 ( .A(n9205), .ZN(n9117) );
  OAI22_X1 U8946 ( .A1(n9194), .A2(n7679), .B1(n9117), .B2(n7637), .ZN(n7207)
         );
  AOI21_X1 U8947 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n7208), .A(n7207), .ZN(
        n7209) );
  OAI21_X1 U8948 ( .B1(n9199), .B2(n9997), .A(n7209), .ZN(P1_U3230) );
  OR2_X1 U8949 ( .A1(n7211), .A2(n8487), .ZN(n7212) );
  NAND2_X1 U8950 ( .A1(n7210), .A2(n7212), .ZN(n7217) );
  INV_X1 U8951 ( .A(n7217), .ZN(n7364) );
  INV_X1 U8952 ( .A(n10266), .ZN(n7381) );
  XNOR2_X1 U8953 ( .A(n8487), .B(n7213), .ZN(n7214) );
  NOR2_X1 U8954 ( .A1(n7214), .A2(n9910), .ZN(n7215) );
  AOI211_X1 U8955 ( .C1(n7381), .C2(n7217), .A(n7216), .B(n7215), .ZN(n7358)
         );
  NAND2_X1 U8956 ( .A1(n7271), .A2(n4480), .ZN(n7218) );
  INV_X1 U8957 ( .A(n7360), .ZN(n7219) );
  AOI22_X1 U8958 ( .A1(n7219), .A2(n9922), .B1(n9026), .B2(n4480), .ZN(n7220)
         );
  OAI211_X1 U8959 ( .C1(n7364), .C2(n10335), .A(n7358), .B(n7220), .ZN(n7222)
         );
  NAND2_X1 U8960 ( .A1(n7222), .A2(n10371), .ZN(n7221) );
  OAI21_X1 U8961 ( .B1(n10371), .B2(n5363), .A(n7221), .ZN(P2_U3460) );
  NAND2_X1 U8962 ( .A1(n7222), .A2(n10382), .ZN(n7223) );
  OAI21_X1 U8963 ( .B1(n10382), .B2(n7224), .A(n7223), .ZN(P2_U3523) );
  NAND2_X1 U8964 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8682), .ZN(n7225) );
  OAI21_X1 U8965 ( .B1(n8314), .B2(n8682), .A(n7225), .ZN(P2_U3581) );
  INV_X1 U8966 ( .A(n8746), .ZN(n8752) );
  OAI222_X1 U8967 ( .A1(n8311), .A2(n7227), .B1(n9070), .B2(n7226), .C1(n8752), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  OAI21_X1 U8968 ( .B1(n7229), .B2(n7228), .A(n7308), .ZN(n7230) );
  NAND2_X1 U8969 ( .A1(n7230), .A2(n8631), .ZN(n7236) );
  NAND2_X1 U8970 ( .A1(n10260), .A2(n8678), .ZN(n7232) );
  NAND2_X1 U8971 ( .A1(n10258), .A2(n10259), .ZN(n7231) );
  AND2_X1 U8972 ( .A1(n7232), .A2(n7231), .ZN(n10276) );
  OAI22_X1 U8973 ( .A1(n8637), .A2(n10276), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7233), .ZN(n7234) );
  AOI21_X1 U8974 ( .B1(n10321), .B2(n8618), .A(n7234), .ZN(n7235) );
  OAI211_X1 U8975 ( .C1(n8652), .C2(n10280), .A(n7236), .B(n7235), .ZN(
        P2_U3241) );
  OAI21_X1 U8976 ( .B1(n8483), .B2(n7239), .A(n7238), .ZN(n7512) );
  OAI211_X1 U8977 ( .C1(n7263), .C2(n7240), .A(n9922), .B(n7270), .ZN(n7507)
         );
  INV_X1 U8978 ( .A(n7507), .ZN(n7245) );
  XNOR2_X1 U8979 ( .A(n8483), .B(n7241), .ZN(n7244) );
  INV_X1 U8980 ( .A(n7242), .ZN(n7243) );
  OAI21_X1 U8981 ( .B1(n7244), .B2(n9910), .A(n7243), .ZN(n7510) );
  AOI211_X1 U8982 ( .C1(n10368), .C2(n7512), .A(n7245), .B(n7510), .ZN(n7261)
         );
  MUX2_X1 U8983 ( .A(n5327), .B(n7261), .S(n10371), .Z(n7246) );
  OAI21_X1 U8984 ( .B1(n7263), .B2(n9061), .A(n7246), .ZN(P2_U3454) );
  AOI22_X1 U8985 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n7784), .B1(n7791), .B2(
        n6028), .ZN(n7249) );
  NOR2_X1 U8986 ( .A1(n7250), .A2(n7249), .ZN(n7783) );
  AOI21_X1 U8987 ( .B1(n7250), .B2(n7249), .A(n7783), .ZN(n7260) );
  INV_X1 U8988 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7251) );
  NAND2_X1 U8989 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n8046) );
  OAI21_X1 U8990 ( .B1(n10116), .B2(n7251), .A(n8046), .ZN(n7258) );
  OAI21_X1 U8991 ( .B1(n7253), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7252), .ZN(
        n7256) );
  NAND2_X1 U8992 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7791), .ZN(n7254) );
  OAI21_X1 U8993 ( .B1(n7791), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7254), .ZN(
        n7255) );
  NOR2_X1 U8994 ( .A1(n7255), .A2(n7256), .ZN(n7790) );
  AOI211_X1 U8995 ( .C1(n7256), .C2(n7255), .A(n7790), .B(n10086), .ZN(n7257)
         );
  AOI211_X1 U8996 ( .C1(n10093), .C2(n7791), .A(n7258), .B(n7257), .ZN(n7259)
         );
  OAI21_X1 U8997 ( .B1(n7260), .B2(n10070), .A(n7259), .ZN(P1_U3253) );
  MUX2_X1 U8998 ( .A(n7123), .B(n7261), .S(n10382), .Z(n7262) );
  OAI21_X1 U8999 ( .B1(n7263), .B2(n9017), .A(n7262), .ZN(P2_U3521) );
  INV_X1 U9000 ( .A(n9513), .ZN(n10108) );
  INV_X1 U9001 ( .A(n7264), .ZN(n7266) );
  INV_X1 U9002 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7265) );
  OAI222_X1 U9003 ( .A1(P1_U3084), .A2(n10108), .B1(n9857), .B2(n7266), .C1(
        n7265), .C2(n8257), .ZN(P1_U3336) );
  INV_X1 U9004 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7267) );
  INV_X1 U9005 ( .A(n8767), .ZN(n8760) );
  OAI222_X1 U9006 ( .A1(n8311), .A2(n7267), .B1(n9070), .B2(n7266), .C1(n8760), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  OAI21_X1 U9007 ( .B1(n7269), .B2(n8484), .A(n7268), .ZN(n7494) );
  INV_X1 U9008 ( .A(n9922), .ZN(n10364) );
  AOI21_X1 U9009 ( .B1(n7270), .B2(n7493), .A(n10364), .ZN(n7272) );
  NAND2_X1 U9010 ( .A1(n7272), .A2(n7271), .ZN(n7490) );
  INV_X1 U9011 ( .A(n7490), .ZN(n7277) );
  XNOR2_X1 U9012 ( .A(n8484), .B(n7273), .ZN(n7275) );
  AOI21_X1 U9013 ( .B1(n7275), .B2(n10278), .A(n7274), .ZN(n7487) );
  INV_X1 U9014 ( .A(n7487), .ZN(n7276) );
  AOI211_X1 U9015 ( .C1(n10368), .C2(n7494), .A(n7277), .B(n7276), .ZN(n7306)
         );
  INV_X1 U9016 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7278) );
  OAI22_X1 U9017 ( .A1(n9061), .A2(n7279), .B1(n10371), .B2(n7278), .ZN(n7280)
         );
  INV_X1 U9018 ( .A(n7280), .ZN(n7281) );
  OAI21_X1 U9019 ( .B1(n7306), .B2(n10370), .A(n7281), .ZN(P2_U3457) );
  NAND2_X1 U9020 ( .A1(n7282), .A2(n8489), .ZN(n10285) );
  OAI21_X1 U9021 ( .B1(n7282), .B2(n8489), .A(n10285), .ZN(n7469) );
  INV_X1 U9022 ( .A(n8270), .ZN(n7284) );
  INV_X1 U9023 ( .A(n10288), .ZN(n7283) );
  AOI211_X1 U9024 ( .C1(n7302), .C2(n7284), .A(n10364), .B(n7283), .ZN(n7468)
         );
  NAND2_X1 U9025 ( .A1(n7285), .A2(n5644), .ZN(n7286) );
  XOR2_X1 U9026 ( .A(n8489), .B(n7286), .Z(n7288) );
  OAI21_X1 U9027 ( .B1(n7288), .B2(n9910), .A(n7287), .ZN(n7462) );
  AOI211_X1 U9028 ( .C1(n10368), .C2(n7469), .A(n7468), .B(n7462), .ZN(n7304)
         );
  INV_X1 U9029 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7289) );
  OAI22_X1 U9030 ( .A1(n9061), .A2(n7465), .B1(n10371), .B2(n7289), .ZN(n7290)
         );
  INV_X1 U9031 ( .A(n7290), .ZN(n7291) );
  OAI21_X1 U9032 ( .B1(n7304), .B2(n10370), .A(n7291), .ZN(P2_U3466) );
  INV_X1 U9033 ( .A(n7292), .ZN(n7294) );
  NAND2_X1 U9034 ( .A1(n7294), .A2(n7293), .ZN(n7295) );
  XNOR2_X1 U9035 ( .A(n7296), .B(n7295), .ZN(n7301) );
  INV_X1 U9036 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7808) );
  AOI22_X1 U9037 ( .A1(n9170), .A2(n9489), .B1(n7808), .B2(n9189), .ZN(n7300)
         );
  NAND2_X1 U9038 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9873) );
  INV_X1 U9039 ( .A(n9873), .ZN(n7298) );
  NOR2_X1 U9040 ( .A1(n9117), .A2(n10167), .ZN(n7297) );
  AOI211_X1 U9041 ( .C1(n9191), .C2(n9490), .A(n7298), .B(n7297), .ZN(n7299)
         );
  OAI211_X1 U9042 ( .C1(n7301), .C2(n9199), .A(n7300), .B(n7299), .ZN(P1_U3216) );
  AOI22_X1 U9043 ( .A1(n5712), .A2(n7302), .B1(n10380), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n7303) );
  OAI21_X1 U9044 ( .B1(n7304), .B2(n10380), .A(n7303), .ZN(P2_U3525) );
  AOI22_X1 U9045 ( .A1(n5712), .A2(n7493), .B1(n10380), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n7305) );
  OAI21_X1 U9046 ( .B1(n7306), .B2(n10380), .A(n7305), .ZN(P2_U3522) );
  XOR2_X1 U9047 ( .A(n7309), .B(n4562), .Z(n7310) );
  NAND2_X1 U9048 ( .A1(n7310), .A2(n8631), .ZN(n7317) );
  INV_X1 U9049 ( .A(n7458), .ZN(n10331) );
  NAND2_X1 U9050 ( .A1(n10260), .A2(n8677), .ZN(n7312) );
  NAND2_X1 U9051 ( .A1(n10258), .A2(n8676), .ZN(n7311) );
  NAND2_X1 U9052 ( .A1(n7312), .A2(n7311), .ZN(n7449) );
  AOI21_X1 U9053 ( .B1(n8654), .B2(n7449), .A(n7313), .ZN(n7314) );
  OAI21_X1 U9054 ( .B1(n8657), .B2(n10331), .A(n7314), .ZN(n7315) );
  INV_X1 U9055 ( .A(n7315), .ZN(n7316) );
  OAI211_X1 U9056 ( .C1(n8652), .C2(n7452), .A(n7317), .B(n7316), .ZN(P2_U3215) );
  INV_X1 U9057 ( .A(n9521), .ZN(n9525) );
  INV_X1 U9058 ( .A(n7318), .ZN(n7320) );
  INV_X1 U9059 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7319) );
  OAI222_X1 U9060 ( .A1(n9525), .A2(P1_U3084), .B1(n9857), .B2(n7320), .C1(
        n7319), .C2(n8257), .ZN(P1_U3335) );
  INV_X1 U9061 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7321) );
  INV_X1 U9062 ( .A(n8769), .ZN(n8781) );
  OAI222_X1 U9063 ( .A1(n8311), .A2(n7321), .B1(n9070), .B2(n7320), .C1(
        P2_U3152), .C2(n8781), .ZN(P2_U3340) );
  XNOR2_X1 U9064 ( .A(n7333), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U9065 ( .A1(n7333), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7323) );
  NAND2_X1 U9066 ( .A1(n8691), .A2(n7323), .ZN(n8704) );
  OR2_X1 U9067 ( .A1(n8706), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7325) );
  NAND2_X1 U9068 ( .A1(n8706), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7324) );
  AND2_X1 U9069 ( .A1(n7325), .A2(n7324), .ZN(n8705) );
  NAND2_X1 U9070 ( .A1(n8704), .A2(n8705), .ZN(n8703) );
  INV_X1 U9071 ( .A(n8703), .ZN(n7326) );
  NAND2_X1 U9072 ( .A1(n7758), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7327) );
  OAI21_X1 U9073 ( .B1(n7758), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7327), .ZN(
        n7328) );
  AOI211_X1 U9074 ( .C1(n7329), .C2(n7328), .A(n7757), .B(n9887), .ZN(n7342)
         );
  AND2_X1 U9075 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7410) );
  AOI21_X1 U9076 ( .B1(n10243), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7410), .ZN(
        n7340) );
  INV_X1 U9077 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10376) );
  MUX2_X1 U9078 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10376), .S(n8706), .Z(n8699)
         );
  INV_X1 U9079 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7334) );
  NAND2_X1 U9080 ( .A1(n7330), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7332) );
  NAND2_X1 U9081 ( .A1(n7332), .A2(n7331), .ZN(n8694) );
  MUX2_X1 U9082 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7334), .S(n7333), .Z(n8693)
         );
  NAND2_X1 U9083 ( .A1(n8694), .A2(n8693), .ZN(n8692) );
  OAI21_X1 U9084 ( .B1(n7334), .B2(n8685), .A(n8692), .ZN(n8700) );
  NAND2_X1 U9085 ( .A1(n8699), .A2(n8700), .ZN(n8698) );
  OAI21_X1 U9086 ( .B1(n7335), .B2(n10376), .A(n8698), .ZN(n7338) );
  INV_X1 U9087 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7336) );
  MUX2_X1 U9088 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7336), .S(n7758), .Z(n7337)
         );
  NAND2_X1 U9089 ( .A1(n7337), .A2(n7338), .ZN(n7764) );
  OAI211_X1 U9090 ( .C1(n7338), .C2(n7337), .A(n10237), .B(n7764), .ZN(n7339)
         );
  OAI211_X1 U9091 ( .C1(n10239), .C2(n7765), .A(n7340), .B(n7339), .ZN(n7341)
         );
  OR2_X1 U9092 ( .A1(n7342), .A2(n7341), .ZN(P2_U3255) );
  INV_X1 U9093 ( .A(n7343), .ZN(n8485) );
  NOR2_X1 U9094 ( .A1(n7344), .A2(n8525), .ZN(n7345) );
  NAND2_X1 U9095 ( .A1(n7346), .A2(n7345), .ZN(n7455) );
  OR2_X1 U9096 ( .A1(n8524), .A2(n8856), .ZN(n7356) );
  NAND2_X1 U9097 ( .A1(n10266), .A2(n7356), .ZN(n7347) );
  NAND2_X1 U9098 ( .A1(n10272), .A2(n7347), .ZN(n8956) );
  OAI21_X1 U9099 ( .B1(n7349), .B2(n8903), .A(n7348), .ZN(n7352) );
  NOR2_X1 U9100 ( .A1(n10272), .A2(n7350), .ZN(n7351) );
  AOI21_X1 U9101 ( .B1(n10272), .B2(n7352), .A(n7351), .ZN(n7355) );
  OR2_X1 U9102 ( .A1(n7455), .A2(n8329), .ZN(n7476) );
  INV_X1 U9103 ( .A(n7476), .ZN(n10255) );
  OAI21_X1 U9104 ( .B1(n10283), .B2(n10255), .A(n6328), .ZN(n7354) );
  OAI211_X1 U9105 ( .C1(n8485), .C2(n8956), .A(n7355), .B(n7354), .ZN(P2_U3296) );
  INV_X1 U9106 ( .A(n7356), .ZN(n7357) );
  NAND2_X1 U9107 ( .A1(n10272), .A2(n7357), .ZN(n10251) );
  MUX2_X1 U9108 ( .A(n7107), .B(n7358), .S(n10272), .Z(n7363) );
  OAI22_X1 U9109 ( .A1(n7476), .A2(n7360), .B1(n8903), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n7361) );
  AOI21_X1 U9110 ( .B1(n10283), .B2(n4480), .A(n7361), .ZN(n7362) );
  OAI211_X1 U9111 ( .C1(n7364), .C2(n10251), .A(n7363), .B(n7362), .ZN(
        P2_U3293) );
  INV_X1 U9112 ( .A(n7389), .ZN(n10341) );
  INV_X1 U9113 ( .A(n7365), .ZN(n7366) );
  NOR2_X1 U9114 ( .A1(n7367), .A2(n7366), .ZN(n7368) );
  XNOR2_X1 U9115 ( .A(n7369), .B(n7368), .ZN(n7370) );
  NAND2_X1 U9116 ( .A1(n7370), .A2(n8631), .ZN(n7375) );
  NAND2_X1 U9117 ( .A1(n8587), .A2(n8676), .ZN(n7371) );
  OAI21_X1 U9118 ( .B1(n8652), .B2(n7384), .A(n7371), .ZN(n7373) );
  NAND2_X1 U9119 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8701) );
  OAI21_X1 U9120 ( .B1(n8584), .B2(n7500), .A(n8701), .ZN(n7372) );
  NOR2_X1 U9121 ( .A1(n7373), .A2(n7372), .ZN(n7374) );
  OAI211_X1 U9122 ( .C1(n10341), .C2(n8657), .A(n7375), .B(n7374), .ZN(
        P2_U3233) );
  OAI21_X1 U9123 ( .B1(n7377), .B2(n8495), .A(n7376), .ZN(n10345) );
  INV_X1 U9124 ( .A(n10345), .ZN(n7392) );
  XNOR2_X1 U9125 ( .A(n7378), .B(n8495), .ZN(n7383) );
  OAI22_X1 U9126 ( .A1(n7379), .A2(n8647), .B1(n7500), .B2(n8649), .ZN(n7380)
         );
  AOI21_X1 U9127 ( .B1(n10345), .B2(n7381), .A(n7380), .ZN(n7382) );
  OAI21_X1 U9128 ( .B1(n9910), .B2(n7383), .A(n7382), .ZN(n10343) );
  NAND2_X1 U9129 ( .A1(n10343), .A2(n10272), .ZN(n7391) );
  INV_X1 U9130 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7385) );
  OAI22_X1 U9131 ( .A1(n10272), .A2(n7385), .B1(n7384), .B2(n8903), .ZN(n7388)
         );
  NAND2_X1 U9132 ( .A1(n10252), .A2(n7389), .ZN(n7386) );
  NAND2_X1 U9133 ( .A1(n7421), .A2(n7386), .ZN(n10342) );
  NOR2_X1 U9134 ( .A1(n10342), .A2(n7476), .ZN(n7387) );
  AOI211_X1 U9135 ( .C1(n10283), .C2(n7389), .A(n7388), .B(n7387), .ZN(n7390)
         );
  OAI211_X1 U9136 ( .C1(n7392), .C2(n10251), .A(n7391), .B(n7390), .ZN(
        P2_U3287) );
  NAND2_X1 U9137 ( .A1(n7393), .A2(n7394), .ZN(n7396) );
  XNOR2_X1 U9138 ( .A(n7396), .B(n7395), .ZN(n7400) );
  AND2_X1 U9139 ( .A1(n7641), .A2(n9964), .ZN(n10152) );
  AOI22_X1 U9140 ( .A1(n9191), .A2(n9492), .B1(n10152), .B2(n7544), .ZN(n7398)
         );
  NAND2_X1 U9141 ( .A1(n9170), .A2(n9490), .ZN(n7397) );
  OAI211_X1 U9142 ( .C1(n9171), .C2(n7639), .A(n7398), .B(n7397), .ZN(n7399)
         );
  AOI21_X1 U9143 ( .B1(n7400), .B2(n9168), .A(n7399), .ZN(n7401) );
  INV_X1 U9144 ( .A(n7401), .ZN(P1_U3220) );
  INV_X1 U9145 ( .A(n7402), .ZN(n7404) );
  OAI222_X1 U9146 ( .A1(P1_U3084), .A2(n9532), .B1(n9857), .B2(n7404), .C1(
        n7403), .C2(n8257), .ZN(P1_U3334) );
  OAI222_X1 U9147 ( .A1(n8311), .A2(n7405), .B1(n9070), .B2(n7404), .C1(n8856), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI211_X1 U9148 ( .C1(n7408), .C2(n7407), .A(n7406), .B(n8631), .ZN(n7412)
         );
  OAI22_X1 U9149 ( .A1(n8200), .A2(n8583), .B1(n8652), .B2(n7420), .ZN(n7409)
         );
  AOI211_X1 U9150 ( .C1(n8154), .C2(n8674), .A(n7410), .B(n7409), .ZN(n7411)
         );
  OAI211_X1 U9151 ( .C1(n10348), .C2(n8657), .A(n7412), .B(n7411), .ZN(
        P2_U3219) );
  XNOR2_X1 U9152 ( .A(n7413), .B(n7416), .ZN(n10347) );
  AOI22_X1 U9153 ( .A1(n10258), .A2(n8674), .B1(n10260), .B2(n10257), .ZN(
        n7419) );
  AND2_X1 U9154 ( .A1(n7414), .A2(n8392), .ZN(n7417) );
  OAI211_X1 U9155 ( .C1(n7417), .C2(n7416), .A(n10278), .B(n7415), .ZN(n7418)
         );
  OAI211_X1 U9156 ( .C1(n10347), .C2(n10266), .A(n7419), .B(n7418), .ZN(n10350) );
  NAND2_X1 U9157 ( .A1(n10350), .A2(n10272), .ZN(n7427) );
  OAI22_X1 U9158 ( .A1(n10272), .A2(n7049), .B1(n7420), .B2(n8903), .ZN(n7424)
         );
  AND2_X1 U9159 ( .A1(n7421), .A2(n7425), .ZN(n7422) );
  OR2_X1 U9160 ( .A1(n7422), .A2(n7522), .ZN(n10349) );
  NOR2_X1 U9161 ( .A1(n10349), .A2(n7476), .ZN(n7423) );
  AOI211_X1 U9162 ( .C1(n10283), .C2(n7425), .A(n7424), .B(n7423), .ZN(n7426)
         );
  OAI211_X1 U9163 ( .C1(n10347), .C2(n10251), .A(n7427), .B(n7426), .ZN(
        P2_U3286) );
  XNOR2_X1 U9164 ( .A(n7534), .B(n7428), .ZN(n7429) );
  NAND2_X1 U9165 ( .A1(n7429), .A2(n7430), .ZN(n7533) );
  OAI21_X1 U9166 ( .B1(n7430), .B2(n7429), .A(n7533), .ZN(n7435) );
  AOI22_X1 U9167 ( .A1(n9191), .A2(n9489), .B1(n9170), .B2(n9487), .ZN(n7433)
         );
  INV_X1 U9168 ( .A(n7705), .ZN(n7701) );
  INV_X1 U9169 ( .A(n9964), .ZN(n10208) );
  NOR2_X1 U9170 ( .A1(n7701), .A2(n10208), .ZN(n10178) );
  NAND2_X1 U9171 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10046) );
  INV_X1 U9172 ( .A(n10046), .ZN(n7431) );
  AOI21_X1 U9173 ( .B1(n10178), .B2(n7544), .A(n7431), .ZN(n7432) );
  OAI211_X1 U9174 ( .C1(n9181), .C2(n7698), .A(n7433), .B(n7432), .ZN(n7434)
         );
  AOI21_X1 U9175 ( .B1(n7435), .B2(n9168), .A(n7434), .ZN(n7436) );
  INV_X1 U9176 ( .A(n7436), .ZN(P1_U3225) );
  INV_X1 U9177 ( .A(n7544), .ZN(n7447) );
  NAND2_X1 U9178 ( .A1(n7672), .A2(n9964), .ZN(n10196) );
  XNOR2_X1 U9179 ( .A(n7439), .B(n7438), .ZN(n7440) );
  XNOR2_X1 U9180 ( .A(n7437), .B(n7440), .ZN(n7441) );
  NAND2_X1 U9181 ( .A1(n7441), .A2(n9168), .ZN(n7446) );
  INV_X1 U9182 ( .A(n7442), .ZN(n7444) );
  OAI22_X1 U9183 ( .A1(n9194), .A2(n7745), .B1(n9181), .B2(n7667), .ZN(n7443)
         );
  AOI211_X1 U9184 ( .C1(n9191), .C2(n9487), .A(n7444), .B(n7443), .ZN(n7445)
         );
  OAI211_X1 U9185 ( .C1(n7447), .C2(n10196), .A(n7446), .B(n7445), .ZN(
        P1_U3211) );
  AOI21_X1 U9186 ( .B1(n7448), .B2(n8380), .A(n9910), .ZN(n7451) );
  AOI21_X1 U9187 ( .B1(n7451), .B2(n7450), .A(n7449), .ZN(n10330) );
  OAI22_X1 U9188 ( .A1(n10272), .A2(n6969), .B1(n7452), .B2(n8903), .ZN(n7457)
         );
  INV_X1 U9189 ( .A(n10289), .ZN(n7454) );
  INV_X1 U9190 ( .A(n10253), .ZN(n7453) );
  OAI211_X1 U9191 ( .C1(n10331), .C2(n7454), .A(n7453), .B(n9922), .ZN(n10329)
         );
  OR2_X1 U9192 ( .A1(n7455), .A2(n8327), .ZN(n8909) );
  NOR2_X1 U9193 ( .A1(n10329), .A2(n8909), .ZN(n7456) );
  AOI211_X1 U9194 ( .C1(n10283), .C2(n7458), .A(n7457), .B(n7456), .ZN(n7461)
         );
  XNOR2_X1 U9195 ( .A(n8380), .B(n7459), .ZN(n10333) );
  NAND2_X1 U9196 ( .A1(n10333), .A2(n10293), .ZN(n7460) );
  OAI211_X1 U9197 ( .C1(n10296), .C2(n10330), .A(n7461), .B(n7460), .ZN(
        P2_U3289) );
  INV_X1 U9198 ( .A(n7462), .ZN(n7472) );
  INV_X1 U9199 ( .A(n8909), .ZN(n10292) );
  INV_X1 U9200 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7464) );
  OAI22_X1 U9201 ( .A1(n10272), .A2(n7464), .B1(n7463), .B2(n8903), .ZN(n7467)
         );
  NOR2_X1 U9202 ( .A1(n10270), .A2(n7465), .ZN(n7466) );
  AOI211_X1 U9203 ( .C1(n7468), .C2(n10292), .A(n7467), .B(n7466), .ZN(n7471)
         );
  NAND2_X1 U9204 ( .A1(n7469), .A2(n10293), .ZN(n7470) );
  OAI211_X1 U9205 ( .C1(n10296), .C2(n7472), .A(n7471), .B(n7470), .ZN(
        P2_U3291) );
  AOI21_X1 U9206 ( .B1(n8499), .B2(n7474), .A(n7473), .ZN(n10361) );
  OAI22_X1 U9207 ( .A1(n10272), .A2(n7475), .B1(n7649), .B2(n8903), .ZN(n7478)
         );
  OAI21_X1 U9208 ( .B1(n7523), .B2(n10363), .A(n7615), .ZN(n10365) );
  NOR2_X1 U9209 ( .A1(n10365), .A2(n7476), .ZN(n7477) );
  AOI211_X1 U9210 ( .C1(n10283), .C2(n7479), .A(n7478), .B(n7477), .ZN(n7486)
         );
  NAND2_X1 U9211 ( .A1(n7606), .A2(n8342), .ZN(n7481) );
  INV_X1 U9212 ( .A(n8499), .ZN(n7480) );
  XNOR2_X1 U9213 ( .A(n7481), .B(n7480), .ZN(n7482) );
  NAND2_X1 U9214 ( .A1(n7482), .A2(n10278), .ZN(n7484) );
  AOI22_X1 U9215 ( .A1(n10260), .A2(n8674), .B1(n10258), .B2(n8672), .ZN(n7483) );
  NAND2_X1 U9216 ( .A1(n7484), .A2(n7483), .ZN(n10367) );
  NAND2_X1 U9217 ( .A1(n10367), .A2(n10272), .ZN(n7485) );
  OAI211_X1 U9218 ( .C1(n10361), .C2(n8956), .A(n7486), .B(n7485), .ZN(
        P2_U3284) );
  INV_X1 U9219 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7488) );
  OAI21_X1 U9220 ( .B1(n7488), .B2(n8903), .A(n7487), .ZN(n7492) );
  INV_X1 U9221 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7489) );
  OAI22_X1 U9222 ( .A1(n8909), .A2(n7490), .B1(n10272), .B2(n7489), .ZN(n7491)
         );
  AOI21_X1 U9223 ( .B1(n10272), .B2(n7492), .A(n7491), .ZN(n7496) );
  AOI22_X1 U9224 ( .A1(n10293), .A2(n7494), .B1(n10283), .B2(n7493), .ZN(n7495) );
  NAND2_X1 U9225 ( .A1(n7496), .A2(n7495), .ZN(P2_U3294) );
  OAI211_X1 U9226 ( .C1(n7499), .C2(n7498), .A(n7497), .B(n8631), .ZN(n7504)
         );
  OAI22_X1 U9227 ( .A1(n8584), .A2(n7736), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8712), .ZN(n7502) );
  OAI22_X1 U9228 ( .A1(n8200), .A2(n7500), .B1(n8652), .B2(n7525), .ZN(n7501)
         );
  AOI211_X1 U9229 ( .C1(n7528), .C2(n8618), .A(n7502), .B(n7501), .ZN(n7503)
         );
  NAND2_X1 U9230 ( .A1(n7504), .A2(n7503), .ZN(P2_U3238) );
  INV_X1 U9231 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7505) );
  NOR2_X1 U9232 ( .A1(n10272), .A2(n7505), .ZN(n7509) );
  OAI22_X1 U9233 ( .A1(n8909), .A2(n7507), .B1(n7506), .B2(n8903), .ZN(n7508)
         );
  AOI211_X1 U9234 ( .C1(n10272), .C2(n7510), .A(n7509), .B(n7508), .ZN(n7514)
         );
  AOI22_X1 U9235 ( .A1(n10293), .A2(n7512), .B1(n10283), .B2(n7511), .ZN(n7513) );
  NAND2_X1 U9236 ( .A1(n7514), .A2(n7513), .ZN(P2_U3295) );
  XNOR2_X1 U9237 ( .A(n7515), .B(n8497), .ZN(n7516) );
  NAND2_X1 U9238 ( .A1(n7516), .A2(n10278), .ZN(n7518) );
  AOI22_X1 U9239 ( .A1(n10260), .A2(n8675), .B1(n10258), .B2(n8673), .ZN(n7517) );
  NAND2_X1 U9240 ( .A1(n7518), .A2(n7517), .ZN(n10358) );
  INV_X1 U9241 ( .A(n10358), .ZN(n7532) );
  OAI21_X1 U9242 ( .B1(n7520), .B2(n8497), .A(n7519), .ZN(n7521) );
  INV_X1 U9243 ( .A(n7521), .ZN(n10359) );
  OAI21_X1 U9244 ( .B1(n7522), .B2(n10356), .A(n9922), .ZN(n7524) );
  OR2_X1 U9245 ( .A1(n7524), .A2(n7523), .ZN(n10355) );
  OAI22_X1 U9246 ( .A1(n10272), .A2(n7526), .B1(n7525), .B2(n8903), .ZN(n7527)
         );
  AOI21_X1 U9247 ( .B1(n10283), .B2(n7528), .A(n7527), .ZN(n7529) );
  OAI21_X1 U9248 ( .B1(n10355), .B2(n8909), .A(n7529), .ZN(n7530) );
  AOI21_X1 U9249 ( .B1(n10359), .B2(n10293), .A(n7530), .ZN(n7531) );
  OAI21_X1 U9250 ( .B1(n10296), .B2(n7532), .A(n7531), .ZN(P2_U3285) );
  OAI21_X1 U9251 ( .B1(n7535), .B2(n7534), .A(n7533), .ZN(n7539) );
  XNOR2_X1 U9252 ( .A(n7537), .B(n7536), .ZN(n7538) );
  XNOR2_X1 U9253 ( .A(n7539), .B(n7538), .ZN(n7547) );
  INV_X1 U9254 ( .A(n7540), .ZN(n7543) );
  INV_X1 U9255 ( .A(n7541), .ZN(n7601) );
  OAI22_X1 U9256 ( .A1(n9194), .A2(n7714), .B1(n9181), .B2(n7601), .ZN(n7542)
         );
  AOI211_X1 U9257 ( .C1(n9191), .C2(n9488), .A(n7543), .B(n7542), .ZN(n7546)
         );
  NOR2_X1 U9258 ( .A1(n7602), .A2(n10208), .ZN(n10186) );
  NAND2_X1 U9259 ( .A1(n10186), .A2(n7544), .ZN(n7545) );
  OAI211_X1 U9260 ( .C1(n7547), .C2(n9199), .A(n7546), .B(n7545), .ZN(P1_U3237) );
  INV_X1 U9261 ( .A(n7548), .ZN(n7550) );
  OAI222_X1 U9262 ( .A1(n5775), .A2(P1_U3084), .B1(n9857), .B2(n7550), .C1(
        n7549), .C2(n9859), .ZN(P1_U3333) );
  OAI222_X1 U9263 ( .A1(n8311), .A2(n7551), .B1(P2_U3152), .B2(n8479), .C1(
        n9070), .C2(n7550), .ZN(P2_U3338) );
  XNOR2_X1 U9264 ( .A(n7553), .B(n7552), .ZN(n7554) );
  XNOR2_X1 U9265 ( .A(n7555), .B(n7554), .ZN(n7556) );
  NAND2_X1 U9266 ( .A1(n7556), .A2(n9168), .ZN(n7560) );
  NAND2_X1 U9267 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10059) );
  INV_X1 U9268 ( .A(n10059), .ZN(n7558) );
  INV_X1 U9269 ( .A(n9484), .ZN(n7887) );
  OAI22_X1 U9270 ( .A1(n9194), .A2(n7887), .B1(n9181), .B2(n7725), .ZN(n7557)
         );
  AOI211_X1 U9271 ( .C1(n9191), .C2(n9486), .A(n7558), .B(n7557), .ZN(n7559)
         );
  OAI211_X1 U9272 ( .C1(n10202), .C2(n9117), .A(n7560), .B(n7559), .ZN(
        P1_U3219) );
  NAND3_X1 U9273 ( .A1(n7562), .A2(n7561), .A3(n7916), .ZN(n7569) );
  NAND2_X1 U9274 ( .A1(n7563), .A2(n9423), .ZN(n7564) );
  INV_X1 U9275 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7566) );
  OAI21_X1 U9276 ( .B1(n7566), .B2(n9669), .A(n7565), .ZN(n7567) );
  NAND2_X1 U9277 ( .A1(n7567), .A2(n9728), .ZN(n7572) );
  OR2_X1 U9278 ( .A1(n7569), .A2(n9670), .ZN(n8212) );
  OR2_X1 U9279 ( .A1(n8212), .A2(n10210), .ZN(n9549) );
  INV_X1 U9280 ( .A(n9549), .ZN(n9743) );
  OAI21_X1 U9281 ( .B1(n9660), .B2(n9743), .A(n7600), .ZN(n7571) );
  OAI211_X1 U9282 ( .C1(n7573), .C2(n9728), .A(n7572), .B(n7571), .ZN(P1_U3291) );
  NAND2_X1 U9283 ( .A1(n9207), .A2(n7574), .ZN(n7575) );
  OR2_X1 U9284 ( .A1(n9487), .A2(n7602), .ZN(n9220) );
  NAND2_X1 U9285 ( .A1(n7602), .A2(n9487), .ZN(n9228) );
  OR2_X1 U9286 ( .A1(n9490), .A2(n10161), .ZN(n7592) );
  NAND2_X1 U9287 ( .A1(n10161), .A2(n9490), .ZN(n9435) );
  AND2_X1 U9288 ( .A1(n7592), .A2(n9435), .ZN(n7591) );
  NAND2_X1 U9289 ( .A1(n7679), .A2(n7641), .ZN(n7590) );
  INV_X1 U9290 ( .A(n7641), .ZN(n7638) );
  NAND4_X1 U9291 ( .A1(n7579), .A2(n7578), .A3(n7577), .A4(n7576), .ZN(n7580)
         );
  NAND2_X1 U9292 ( .A1(n7638), .A2(n7580), .ZN(n9430) );
  AND2_X1 U9293 ( .A1(n9492), .A2(n7600), .ZN(n7623) );
  NAND2_X1 U9294 ( .A1(n7580), .A2(n7641), .ZN(n7581) );
  INV_X1 U9295 ( .A(n10161), .ZN(n9172) );
  OR2_X1 U9296 ( .A1(n9490), .A2(n9172), .ZN(n7582) );
  NAND2_X1 U9297 ( .A1(n7802), .A2(n7803), .ZN(n7584) );
  INV_X1 U9298 ( .A(n7846), .ZN(n9438) );
  NAND2_X1 U9299 ( .A1(n9438), .A2(n10167), .ZN(n7583) );
  NAND2_X1 U9300 ( .A1(n7584), .A2(n7583), .ZN(n7841) );
  OR2_X1 U9301 ( .A1(n9489), .A2(n10172), .ZN(n7691) );
  NAND2_X1 U9302 ( .A1(n10172), .A2(n9489), .ZN(n7693) );
  NAND2_X1 U9303 ( .A1(n7691), .A2(n7693), .ZN(n9334) );
  NAND2_X1 U9304 ( .A1(n7841), .A2(n9334), .ZN(n7586) );
  INV_X1 U9305 ( .A(n10172), .ZN(n9142) );
  OR2_X1 U9306 ( .A1(n9489), .A2(n9142), .ZN(n7585) );
  XNOR2_X1 U9307 ( .A(n9488), .B(n7705), .ZN(n9339) );
  NAND2_X1 U9308 ( .A1(n9488), .A2(n7705), .ZN(n7587) );
  XOR2_X1 U9309 ( .A(n9340), .B(n7666), .Z(n10191) );
  NAND2_X1 U9310 ( .A1(n9209), .A2(n9670), .ZN(n7589) );
  NAND2_X1 U9311 ( .A1(n6284), .A2(n7588), .ZN(n9464) );
  NAND2_X1 U9312 ( .A1(n7589), .A2(n9464), .ZN(n9738) );
  OR2_X1 U9313 ( .A1(n9336), .A2(n7630), .ZN(n7631) );
  NAND2_X1 U9314 ( .A1(n7631), .A2(n7590), .ZN(n9431) );
  INV_X1 U9315 ( .A(n7591), .ZN(n9337) );
  NAND2_X1 U9316 ( .A1(n9431), .A2(n7591), .ZN(n7678) );
  INV_X1 U9317 ( .A(n7592), .ZN(n7593) );
  INV_X1 U9318 ( .A(n7803), .ZN(n9338) );
  INV_X1 U9319 ( .A(n10167), .ZN(n9437) );
  NAND2_X1 U9320 ( .A1(n9438), .A2(n9437), .ZN(n9439) );
  INV_X1 U9321 ( .A(n9488), .ZN(n9140) );
  NAND2_X1 U9322 ( .A1(n9140), .A2(n7705), .ZN(n7594) );
  AND2_X1 U9323 ( .A1(n7594), .A2(n7691), .ZN(n7654) );
  NAND2_X1 U9324 ( .A1(n7595), .A2(n7654), .ZN(n7597) );
  AND2_X1 U9325 ( .A1(n7701), .A2(n9488), .ZN(n7656) );
  INV_X1 U9326 ( .A(n7656), .ZN(n7596) );
  NAND2_X1 U9327 ( .A1(n7597), .A2(n7596), .ZN(n9218) );
  XNOR2_X1 U9328 ( .A(n9219), .B(n9340), .ZN(n7599) );
  AOI222_X1 U9329 ( .A1(n9738), .A2(n7599), .B1(n9488), .B2(n9733), .C1(n9486), 
        .C2(n9735), .ZN(n10190) );
  MUX2_X1 U9330 ( .A(n6554), .B(n10190), .S(n9728), .Z(n7605) );
  INV_X1 U9331 ( .A(n7602), .ZN(n7665) );
  OR2_X1 U9332 ( .A1(n7641), .A2(n7600), .ZN(n7684) );
  NAND2_X1 U9333 ( .A1(n7807), .A2(n10167), .ZN(n7842) );
  AOI21_X1 U9334 ( .B1(n7665), .B2(n7700), .A(n7669), .ZN(n10188) );
  OAI22_X1 U9335 ( .A1(n9951), .A2(n7602), .B1(n7601), .B2(n9669), .ZN(n7603)
         );
  AOI21_X1 U9336 ( .B1(n10188), .B2(n9743), .A(n7603), .ZN(n7604) );
  OAI211_X1 U9337 ( .C1(n9745), .C2(n10191), .A(n7605), .B(n7604), .ZN(
        P1_U3285) );
  NAND2_X1 U9338 ( .A1(n7606), .A2(n8404), .ZN(n7607) );
  NAND2_X1 U9339 ( .A1(n7607), .A2(n8402), .ZN(n7609) );
  OAI21_X1 U9340 ( .B1(n8500), .B2(n7609), .A(n7608), .ZN(n7610) );
  AOI222_X1 U9341 ( .A1(n10278), .A2(n7610), .B1(n8671), .B2(n10258), .C1(
        n8673), .C2(n10260), .ZN(n9935) );
  OAI21_X1 U9342 ( .B1(n7612), .B2(n8410), .A(n7611), .ZN(n7613) );
  INV_X1 U9343 ( .A(n7613), .ZN(n9938) );
  NAND2_X1 U9344 ( .A1(n9938), .A2(n10293), .ZN(n7619) );
  OAI22_X1 U9345 ( .A1(n10272), .A2(n7614), .B1(n7735), .B2(n8903), .ZN(n7617)
         );
  OAI211_X1 U9346 ( .C1(n4746), .C2(n9936), .A(n9922), .B(n9921), .ZN(n9934)
         );
  NOR2_X1 U9347 ( .A1(n9934), .A2(n8909), .ZN(n7616) );
  AOI211_X1 U9348 ( .C1(n10283), .C2(n5468), .A(n7617), .B(n7616), .ZN(n7618)
         );
  OAI211_X1 U9349 ( .C1(n10296), .C2(n9935), .A(n7619), .B(n7618), .ZN(
        P2_U3283) );
  INV_X1 U9350 ( .A(n7620), .ZN(n7710) );
  OAI222_X1 U9351 ( .A1(n9423), .A2(P1_U3084), .B1(n9857), .B2(n7710), .C1(
        n7621), .C2(n9859), .ZN(P1_U3332) );
  OAI21_X1 U9352 ( .B1(n9336), .B2(n7623), .A(n7622), .ZN(n10156) );
  NAND2_X1 U9353 ( .A1(n7625), .A2(n9670), .ZN(n7624) );
  OR2_X1 U9354 ( .A1(n7626), .A2(n7625), .ZN(n7629) );
  OR2_X1 U9355 ( .A1(n7627), .A2(n9423), .ZN(n7628) );
  AND2_X1 U9356 ( .A1(n7629), .A2(n7628), .ZN(n7998) );
  AOI22_X1 U9357 ( .A1(n9733), .A2(n9492), .B1(n9490), .B2(n9735), .ZN(n7636)
         );
  INV_X1 U9358 ( .A(n9336), .ZN(n7633) );
  INV_X1 U9359 ( .A(n7630), .ZN(n7632) );
  OAI21_X1 U9360 ( .B1(n7633), .B2(n7632), .A(n7631), .ZN(n7634) );
  NAND2_X1 U9361 ( .A1(n7634), .A2(n9738), .ZN(n7635) );
  OAI211_X1 U9362 ( .C1(n10156), .C2(n7998), .A(n7636), .B(n7635), .ZN(n10158)
         );
  OAI211_X1 U9363 ( .C1(n7638), .C2(n7637), .A(n10187), .B(n7684), .ZN(n10153)
         );
  OAI22_X1 U9364 ( .A1(n10153), .A2(n9670), .B1(n9669), .B2(n7639), .ZN(n7640)
         );
  OAI21_X1 U9365 ( .B1(n10158), .B2(n7640), .A(n9728), .ZN(n7643) );
  AOI22_X1 U9366 ( .A1(n9660), .A2(n7641), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n9703), .ZN(n7642) );
  OAI211_X1 U9367 ( .C1(n10156), .C2(n9953), .A(n7643), .B(n7642), .ZN(
        P1_U3290) );
  NAND2_X1 U9368 ( .A1(n4564), .A2(n7644), .ZN(n7645) );
  XNOR2_X1 U9369 ( .A(n7646), .B(n7645), .ZN(n7647) );
  NAND2_X1 U9370 ( .A1(n7647), .A2(n8631), .ZN(n7653) );
  NAND2_X1 U9371 ( .A1(n8587), .A2(n8674), .ZN(n7648) );
  OAI21_X1 U9372 ( .B1(n8652), .B2(n7649), .A(n7648), .ZN(n7651) );
  NAND2_X1 U9373 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7770) );
  OAI21_X1 U9374 ( .B1(n8584), .B2(n7856), .A(n7770), .ZN(n7650) );
  NOR2_X1 U9375 ( .A1(n7651), .A2(n7650), .ZN(n7652) );
  OAI211_X1 U9376 ( .C1(n10363), .C2(n8657), .A(n7653), .B(n7652), .ZN(
        P2_U3226) );
  NAND2_X1 U9377 ( .A1(n7654), .A2(n9220), .ZN(n7655) );
  INV_X1 U9378 ( .A(n7655), .ZN(n9440) );
  INV_X1 U9379 ( .A(n7693), .ZN(n7659) );
  NAND2_X1 U9380 ( .A1(n7656), .A2(n9220), .ZN(n7657) );
  NAND2_X1 U9381 ( .A1(n7657), .A2(n9228), .ZN(n7658) );
  AOI21_X1 U9382 ( .B1(n9440), .B2(n7659), .A(n7658), .ZN(n9443) );
  NAND2_X1 U9383 ( .A1(n7714), .A2(n7672), .ZN(n9231) );
  INV_X1 U9384 ( .A(n7672), .ZN(n7713) );
  NAND2_X1 U9385 ( .A1(n7713), .A2(n9486), .ZN(n9442) );
  NAND2_X1 U9386 ( .A1(n9231), .A2(n9442), .ZN(n9342) );
  INV_X1 U9387 ( .A(n9342), .ZN(n7661) );
  XNOR2_X1 U9388 ( .A(n7718), .B(n7661), .ZN(n7664) );
  NAND2_X1 U9389 ( .A1(n9487), .A2(n9733), .ZN(n7662) );
  OAI21_X1 U9390 ( .B1(n7745), .B2(n9683), .A(n7662), .ZN(n7663) );
  AOI21_X1 U9391 ( .B1(n7664), .B2(n9738), .A(n7663), .ZN(n10197) );
  XNOR2_X1 U9392 ( .A(n7712), .B(n9342), .ZN(n10200) );
  INV_X1 U9393 ( .A(n9745), .ZN(n7707) );
  NAND2_X1 U9394 ( .A1(n10200), .A2(n7707), .ZN(n7674) );
  OAI22_X1 U9395 ( .A1(n9728), .A2(n7668), .B1(n7667), .B2(n9669), .ZN(n7671)
         );
  OAI211_X1 U9396 ( .C1(n7669), .C2(n7713), .A(n7727), .B(n10187), .ZN(n10195)
         );
  NOR2_X1 U9397 ( .A1(n10195), .A2(n8212), .ZN(n7670) );
  AOI211_X1 U9398 ( .C1(n9660), .C2(n7672), .A(n7671), .B(n7670), .ZN(n7673)
         );
  OAI211_X1 U9399 ( .C1(n9703), .C2(n10197), .A(n7674), .B(n7673), .ZN(
        P1_U3284) );
  INV_X1 U9400 ( .A(n7675), .ZN(n7676) );
  AOI21_X1 U9401 ( .B1(n7591), .B2(n7677), .A(n7676), .ZN(n10159) );
  OAI21_X1 U9402 ( .B1(n7591), .B2(n9431), .A(n7678), .ZN(n7681) );
  INV_X1 U9403 ( .A(n9733), .ZN(n9681) );
  OAI22_X1 U9404 ( .A1(n9438), .A2(n9683), .B1(n7679), .B2(n9681), .ZN(n7680)
         );
  AOI21_X1 U9405 ( .B1(n7681), .B2(n9738), .A(n7680), .ZN(n7682) );
  OAI21_X1 U9406 ( .B1(n10159), .B2(n7998), .A(n7682), .ZN(n10162) );
  NAND2_X1 U9407 ( .A1(n10162), .A2(n9728), .ZN(n7690) );
  INV_X1 U9408 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7683) );
  INV_X1 U9409 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10007) );
  OAI22_X1 U9410 ( .A1(n9728), .A2(n7683), .B1(n10007), .B2(n9669), .ZN(n7688)
         );
  INV_X1 U9411 ( .A(n7684), .ZN(n7686) );
  INV_X1 U9412 ( .A(n7807), .ZN(n7685) );
  OAI211_X1 U9413 ( .C1(n10161), .C2(n7686), .A(n7685), .B(n10187), .ZN(n10160) );
  NOR2_X1 U9414 ( .A1(n10160), .A2(n8212), .ZN(n7687) );
  AOI211_X1 U9415 ( .C1(n9660), .C2(n9172), .A(n7688), .B(n7687), .ZN(n7689)
         );
  OAI211_X1 U9416 ( .C1(n10159), .C2(n9953), .A(n7690), .B(n7689), .ZN(
        P1_U3289) );
  INV_X1 U9417 ( .A(n7691), .ZN(n7692) );
  OR2_X1 U9418 ( .A1(n7845), .A2(n7692), .ZN(n7694) );
  AND2_X1 U9419 ( .A1(n7694), .A2(n7693), .ZN(n7696) );
  NAND2_X1 U9420 ( .A1(n7696), .A2(n9339), .ZN(n7695) );
  OAI21_X1 U9421 ( .B1(n7696), .B2(n9339), .A(n7695), .ZN(n7697) );
  AOI222_X1 U9422 ( .A1(n9738), .A2(n7697), .B1(n9487), .B2(n9735), .C1(n9489), 
        .C2(n9733), .ZN(n10184) );
  INV_X1 U9423 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7699) );
  OAI22_X1 U9424 ( .A1(n9728), .A2(n7699), .B1(n7698), .B2(n9669), .ZN(n7704)
         );
  INV_X1 U9425 ( .A(n7843), .ZN(n7702) );
  OAI211_X1 U9426 ( .C1(n7702), .C2(n7701), .A(n10187), .B(n7700), .ZN(n10182)
         );
  NOR2_X1 U9427 ( .A1(n10182), .A2(n8212), .ZN(n7703) );
  AOI211_X1 U9428 ( .C1(n9660), .C2(n7705), .A(n7704), .B(n7703), .ZN(n7709)
         );
  NAND2_X1 U9429 ( .A1(n7706), .A2(n9339), .ZN(n10179) );
  NAND3_X1 U9430 ( .A1(n10180), .A2(n10179), .A3(n7707), .ZN(n7708) );
  OAI211_X1 U9431 ( .C1(n10184), .C2(n9703), .A(n7709), .B(n7708), .ZN(
        P1_U3286) );
  OAI222_X1 U9432 ( .A1(n8311), .A2(n7711), .B1(P2_U3152), .B2(n8330), .C1(
        n9070), .C2(n7710), .ZN(P2_U3337) );
  NAND2_X1 U9433 ( .A1(n7712), .A2(n9342), .ZN(n7716) );
  NAND2_X1 U9434 ( .A1(n7714), .A2(n7713), .ZN(n7715) );
  NAND2_X1 U9435 ( .A1(n7745), .A2(n7741), .ZN(n9230) );
  OR2_X1 U9436 ( .A1(n7877), .A2(n7878), .ZN(n7742) );
  NAND2_X1 U9437 ( .A1(n7877), .A2(n7878), .ZN(n7717) );
  NAND2_X1 U9438 ( .A1(n7742), .A2(n7717), .ZN(n10201) );
  AOI22_X1 U9439 ( .A1(n9486), .A2(n9733), .B1(n9735), .B2(n9484), .ZN(n7724)
         );
  NAND2_X1 U9440 ( .A1(n7718), .A2(n9442), .ZN(n7721) );
  INV_X1 U9441 ( .A(n7721), .ZN(n9376) );
  INV_X1 U9442 ( .A(n9231), .ZN(n7719) );
  OAI21_X1 U9443 ( .B1(n9376), .B2(n7719), .A(n9343), .ZN(n7722) );
  NOR2_X1 U9444 ( .A1(n9343), .A2(n7719), .ZN(n7720) );
  NAND2_X1 U9445 ( .A1(n7721), .A2(n7720), .ZN(n7744) );
  NAND3_X1 U9446 ( .A1(n7722), .A2(n9738), .A3(n7744), .ZN(n7723) );
  OAI211_X1 U9447 ( .C1(n10201), .C2(n7998), .A(n7724), .B(n7723), .ZN(n10204)
         );
  NAND2_X1 U9448 ( .A1(n10204), .A2(n9728), .ZN(n7732) );
  OAI22_X1 U9449 ( .A1(n9728), .A2(n7726), .B1(n7725), .B2(n9669), .ZN(n7730)
         );
  NAND2_X1 U9450 ( .A1(n7727), .A2(n7741), .ZN(n7728) );
  NAND2_X1 U9451 ( .A1(n7751), .A2(n7728), .ZN(n10203) );
  NOR2_X1 U9452 ( .A1(n10203), .A2(n9549), .ZN(n7729) );
  AOI211_X1 U9453 ( .C1(n9660), .C2(n7741), .A(n7730), .B(n7729), .ZN(n7731)
         );
  OAI211_X1 U9454 ( .C1(n10201), .C2(n9953), .A(n7732), .B(n7731), .ZN(
        P1_U3283) );
  XNOR2_X1 U9455 ( .A(n7733), .B(n7734), .ZN(n7740) );
  NAND2_X1 U9456 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7871) );
  OAI21_X1 U9457 ( .B1(n8584), .B2(n8058), .A(n7871), .ZN(n7738) );
  OAI22_X1 U9458 ( .A1(n8200), .A2(n7736), .B1(n8652), .B2(n7735), .ZN(n7737)
         );
  AOI211_X1 U9459 ( .C1(n5468), .C2(n8618), .A(n7738), .B(n7737), .ZN(n7739)
         );
  OAI21_X1 U9460 ( .B1(n7740), .B2(n8642), .A(n7739), .ZN(P2_U3236) );
  NAND2_X1 U9461 ( .A1(n9485), .A2(n7741), .ZN(n7879) );
  NAND2_X1 U9462 ( .A1(n7742), .A2(n7879), .ZN(n7743) );
  AND2_X1 U9463 ( .A1(n7887), .A2(n7881), .ZN(n7906) );
  INV_X1 U9464 ( .A(n7906), .ZN(n9222) );
  INV_X1 U9465 ( .A(n7881), .ZN(n10209) );
  NAND2_X1 U9466 ( .A1(n10209), .A2(n9484), .ZN(n7905) );
  NAND2_X1 U9467 ( .A1(n9222), .A2(n7905), .ZN(n9344) );
  XNOR2_X1 U9468 ( .A(n7743), .B(n9344), .ZN(n10207) );
  XNOR2_X1 U9469 ( .A(n7910), .B(n9344), .ZN(n7747) );
  INV_X1 U9470 ( .A(n7899), .ZN(n7925) );
  OAI22_X1 U9471 ( .A1(n7925), .A2(n9683), .B1(n7745), .B2(n9681), .ZN(n7746)
         );
  AOI21_X1 U9472 ( .B1(n7747), .B2(n9738), .A(n7746), .ZN(n7748) );
  OAI21_X1 U9473 ( .B1(n10207), .B2(n7998), .A(n7748), .ZN(n10212) );
  NAND2_X1 U9474 ( .A1(n10212), .A2(n9728), .ZN(n7756) );
  INV_X1 U9475 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7750) );
  INV_X1 U9476 ( .A(n7749), .ZN(n7818) );
  OAI22_X1 U9477 ( .A1(n9728), .A2(n7750), .B1(n7818), .B2(n9669), .ZN(n7754)
         );
  AND2_X1 U9478 ( .A1(n7751), .A2(n7881), .ZN(n7752) );
  OR2_X1 U9479 ( .A1(n7752), .A2(n7893), .ZN(n10211) );
  NOR2_X1 U9480 ( .A1(n10211), .A2(n9549), .ZN(n7753) );
  AOI211_X1 U9481 ( .C1(n9660), .C2(n7881), .A(n7754), .B(n7753), .ZN(n7755)
         );
  OAI211_X1 U9482 ( .C1(n10207), .C2(n9953), .A(n7756), .B(n7755), .ZN(
        P1_U3282) );
  MUX2_X1 U9483 ( .A(n7526), .B(P2_REG2_REG_11__SCAN_IN), .S(n8711), .Z(n7759)
         );
  INV_X1 U9484 ( .A(n7759), .ZN(n8716) );
  NAND2_X1 U9485 ( .A1(n7866), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7760) );
  OAI21_X1 U9486 ( .B1(n7866), .B2(P2_REG2_REG_12__SCAN_IN), .A(n7760), .ZN(
        n7761) );
  NOR2_X1 U9487 ( .A1(n7761), .A2(n7762), .ZN(n7865) );
  AOI211_X1 U9488 ( .C1(n7762), .C2(n7761), .A(n7865), .B(n9887), .ZN(n7776)
         );
  NAND2_X1 U9489 ( .A1(n8711), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7766) );
  INV_X1 U9490 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7763) );
  MUX2_X1 U9491 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7763), .S(n8711), .Z(n8719)
         );
  OAI21_X1 U9492 ( .B1(n7765), .B2(n7336), .A(n7764), .ZN(n8720) );
  NAND2_X1 U9493 ( .A1(n8719), .A2(n8720), .ZN(n8718) );
  NAND2_X1 U9494 ( .A1(n7766), .A2(n8718), .ZN(n7769) );
  MUX2_X1 U9495 ( .A(n7767), .B(P2_REG1_REG_12__SCAN_IN), .S(n7866), .Z(n7768)
         );
  NOR2_X1 U9496 ( .A1(n7769), .A2(n7768), .ZN(n7861) );
  AOI21_X1 U9497 ( .B1(n7769), .B2(n7768), .A(n7861), .ZN(n7774) );
  INV_X1 U9498 ( .A(n10239), .ZN(n9893) );
  NAND2_X1 U9499 ( .A1(n9893), .A2(n7866), .ZN(n7773) );
  INV_X1 U9500 ( .A(n7770), .ZN(n7771) );
  AOI21_X1 U9501 ( .B1(n10243), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7771), .ZN(
        n7772) );
  OAI211_X1 U9502 ( .C1(n7774), .C2(n10241), .A(n7773), .B(n7772), .ZN(n7775)
         );
  OR2_X1 U9503 ( .A1(n7776), .A2(n7775), .ZN(P2_U3257) );
  NAND2_X1 U9504 ( .A1(n7779), .A2(n8114), .ZN(n7777) );
  OAI211_X1 U9505 ( .C1(n7778), .C2(n8311), .A(n7777), .B(n8530), .ZN(P2_U3335) );
  NAND2_X1 U9506 ( .A1(n7779), .A2(n4567), .ZN(n7781) );
  NOR2_X1 U9507 ( .A1(n7780), .A2(P1_U3084), .ZN(n9468) );
  INV_X1 U9508 ( .A(n9468), .ZN(n9208) );
  OAI211_X1 U9509 ( .C1(n7782), .C2(n9859), .A(n7781), .B(n9208), .ZN(P1_U3330) );
  INV_X1 U9510 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7786) );
  MUX2_X1 U9511 ( .A(n7786), .B(P1_REG1_REG_13__SCAN_IN), .S(n10066), .Z(
        n10068) );
  NOR2_X1 U9512 ( .A1(n10069), .A2(n10068), .ZN(n10067) );
  INV_X1 U9513 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9970) );
  AOI22_X1 U9514 ( .A1(n7796), .A2(n9970), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n9505), .ZN(n7787) );
  NOR2_X1 U9515 ( .A1(n7788), .A2(n7787), .ZN(n9493) );
  AOI21_X1 U9516 ( .B1(n7788), .B2(n7787), .A(n9493), .ZN(n7798) );
  INV_X1 U9517 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7789) );
  NAND2_X1 U9518 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n8027) );
  OAI21_X1 U9519 ( .B1(n10116), .B2(n7789), .A(n8027), .ZN(n7795) );
  XNOR2_X1 U9520 ( .A(n10066), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n10062) );
  INV_X1 U9521 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7792) );
  NOR2_X1 U9522 ( .A1(n7792), .A2(n7793), .ZN(n9507) );
  AOI211_X1 U9523 ( .C1(n7793), .C2(n7792), .A(n9507), .B(n10086), .ZN(n7794)
         );
  AOI211_X1 U9524 ( .C1(n10093), .C2(n7796), .A(n7795), .B(n7794), .ZN(n7797)
         );
  OAI21_X1 U9525 ( .B1(n7798), .B2(n10070), .A(n7797), .ZN(P1_U3255) );
  INV_X1 U9526 ( .A(n7799), .ZN(n8309) );
  OAI222_X1 U9527 ( .A1(P1_U3084), .A2(n6282), .B1(n9857), .B2(n8309), .C1(
        n7800), .C2(n9859), .ZN(P1_U3331) );
  INV_X1 U9528 ( .A(n9738), .ZN(n9678) );
  XNOR2_X1 U9529 ( .A(n7801), .B(n7803), .ZN(n7806) );
  XNOR2_X1 U9530 ( .A(n7802), .B(n7803), .ZN(n10170) );
  INV_X1 U9531 ( .A(n7998), .ZN(n9945) );
  NAND2_X1 U9532 ( .A1(n10170), .A2(n9945), .ZN(n7805) );
  AOI22_X1 U9533 ( .A1(n9733), .A2(n9490), .B1(n9489), .B2(n9735), .ZN(n7804)
         );
  OAI211_X1 U9534 ( .C1(n9678), .C2(n7806), .A(n7805), .B(n7804), .ZN(n10168)
         );
  INV_X1 U9535 ( .A(n10168), .ZN(n7813) );
  INV_X1 U9536 ( .A(n9953), .ZN(n7852) );
  OAI211_X1 U9537 ( .C1(n7807), .C2(n10167), .A(n7842), .B(n10187), .ZN(n10166) );
  INV_X1 U9538 ( .A(n9669), .ZN(n9948) );
  AOI22_X1 U9539 ( .A1(n9703), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9948), .B2(
        n7808), .ZN(n7810) );
  NAND2_X1 U9540 ( .A1(n9660), .A2(n9437), .ZN(n7809) );
  OAI211_X1 U9541 ( .C1(n10166), .C2(n8212), .A(n7810), .B(n7809), .ZN(n7811)
         );
  AOI21_X1 U9542 ( .B1(n10170), .B2(n7852), .A(n7811), .ZN(n7812) );
  OAI21_X1 U9543 ( .B1(n7813), .B2(n9703), .A(n7812), .ZN(P1_U3288) );
  INV_X1 U9544 ( .A(n7815), .ZN(n7816) );
  AOI21_X1 U9545 ( .B1(n7817), .B2(n7814), .A(n7816), .ZN(n7823) );
  OAI22_X1 U9546 ( .A1(n9194), .A2(n7925), .B1(n9181), .B2(n7818), .ZN(n7819)
         );
  AOI211_X1 U9547 ( .C1(n9191), .C2(n9485), .A(n7820), .B(n7819), .ZN(n7822)
         );
  NAND2_X1 U9548 ( .A1(n9205), .A2(n7881), .ZN(n7821) );
  OAI211_X1 U9549 ( .C1(n7823), .C2(n9199), .A(n7822), .B(n7821), .ZN(P1_U3229) );
  INV_X1 U9550 ( .A(n7824), .ZN(n7828) );
  OAI222_X1 U9551 ( .A1(n7826), .A2(P2_U3152), .B1(n9070), .B2(n7828), .C1(
        n7825), .C2(n8311), .ZN(P2_U3334) );
  OAI222_X1 U9552 ( .A1(n7829), .A2(P1_U3084), .B1(n9857), .B2(n7828), .C1(
        n7827), .C2(n9859), .ZN(P1_U3329) );
  INV_X1 U9553 ( .A(n7908), .ZN(n9901) );
  INV_X1 U9554 ( .A(n7830), .ZN(n7832) );
  NOR2_X1 U9555 ( .A1(n7832), .A2(n7831), .ZN(n7833) );
  XNOR2_X1 U9556 ( .A(n7834), .B(n7833), .ZN(n7835) );
  NAND2_X1 U9557 ( .A1(n7835), .A2(n9168), .ZN(n7840) );
  INV_X1 U9558 ( .A(n7836), .ZN(n7838) );
  OAI22_X1 U9559 ( .A1(n9194), .A2(n8049), .B1(n9181), .B2(n7891), .ZN(n7837)
         );
  AOI211_X1 U9560 ( .C1(n9191), .C2(n9484), .A(n7838), .B(n7837), .ZN(n7839)
         );
  OAI211_X1 U9561 ( .C1(n9901), .C2(n9117), .A(n7840), .B(n7839), .ZN(P1_U3215) );
  XNOR2_X1 U9562 ( .A(n7841), .B(n9334), .ZN(n10176) );
  OAI21_X1 U9563 ( .B1(n4762), .B2(n10172), .A(n7843), .ZN(n10173) );
  AOI22_X1 U9564 ( .A1(n9660), .A2(n9142), .B1(n9139), .B2(n9948), .ZN(n7844)
         );
  OAI21_X1 U9565 ( .B1(n10173), .B2(n9549), .A(n7844), .ZN(n7851) );
  XNOR2_X1 U9566 ( .A(n7845), .B(n9334), .ZN(n7849) );
  NAND2_X1 U9567 ( .A1(n10176), .A2(n9945), .ZN(n7848) );
  AOI22_X1 U9568 ( .A1(n9733), .A2(n7846), .B1(n9488), .B2(n9735), .ZN(n7847)
         );
  OAI211_X1 U9569 ( .C1(n7849), .C2(n9678), .A(n7848), .B(n7847), .ZN(n10174)
         );
  MUX2_X1 U9570 ( .A(n10174), .B(P1_REG2_REG_4__SCAN_IN), .S(n9703), .Z(n7850)
         );
  AOI211_X1 U9571 ( .C1(n7852), .C2(n10176), .A(n7851), .B(n7850), .ZN(n7853)
         );
  INV_X1 U9572 ( .A(n7853), .ZN(P1_U3287) );
  AOI21_X1 U9573 ( .B1(n7855), .B2(n7854), .A(n4563), .ZN(n7860) );
  NAND2_X1 U9574 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7966) );
  OAI22_X1 U9575 ( .A1(n8152), .A2(n8649), .B1(n7856), .B2(n8647), .ZN(n9913)
         );
  NAND2_X1 U9576 ( .A1(n8654), .A2(n9913), .ZN(n7857) );
  OAI211_X1 U9577 ( .C1(n8652), .C2(n9915), .A(n7966), .B(n7857), .ZN(n7858)
         );
  AOI21_X1 U9578 ( .B1(n9917), .B2(n8618), .A(n7858), .ZN(n7859) );
  OAI21_X1 U9579 ( .B1(n7860), .B2(n8642), .A(n7859), .ZN(P2_U3217) );
  AOI21_X1 U9580 ( .B1(n7862), .B2(n7767), .A(n7861), .ZN(n7864) );
  INV_X1 U9581 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9939) );
  AOI22_X1 U9582 ( .A1(n7962), .A2(n9939), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7957), .ZN(n7863) );
  NOR2_X1 U9583 ( .A1(n7864), .A2(n7863), .ZN(n7956) );
  AOI21_X1 U9584 ( .B1(n7864), .B2(n7863), .A(n7956), .ZN(n7876) );
  NOR2_X1 U9585 ( .A1(n7962), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7867) );
  AOI21_X1 U9586 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7962), .A(n7867), .ZN(
        n7868) );
  NAND2_X1 U9587 ( .A1(n7869), .A2(n7868), .ZN(n7961) );
  OAI21_X1 U9588 ( .B1(n7869), .B2(n7868), .A(n7961), .ZN(n7870) );
  NAND2_X1 U9589 ( .A1(n7870), .A2(n10238), .ZN(n7875) );
  INV_X1 U9590 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7872) );
  OAI21_X1 U9591 ( .B1(n8791), .B2(n7872), .A(n7871), .ZN(n7873) );
  AOI21_X1 U9592 ( .B1(n9893), .B2(n7962), .A(n7873), .ZN(n7874) );
  OAI211_X1 U9593 ( .C1(n7876), .C2(n10241), .A(n7875), .B(n7874), .ZN(
        P2_U3258) );
  XNOR2_X1 U9594 ( .A(n7908), .B(n7899), .ZN(n9346) );
  NOR2_X1 U9595 ( .A1(n9484), .A2(n7881), .ZN(n7880) );
  OR2_X1 U9596 ( .A1(n7880), .A2(n7879), .ZN(n7883) );
  NAND2_X1 U9597 ( .A1(n7881), .A2(n9484), .ZN(n7882) );
  OR2_X2 U9598 ( .A1(n7885), .A2(n9346), .ZN(n7901) );
  INV_X1 U9599 ( .A(n7901), .ZN(n7884) );
  AOI21_X1 U9600 ( .B1(n9346), .B2(n7885), .A(n7884), .ZN(n9900) );
  OAI21_X1 U9601 ( .B1(n4881), .B2(n9344), .A(n7905), .ZN(n7886) );
  XOR2_X1 U9602 ( .A(n9346), .B(n7886), .Z(n7889) );
  OAI22_X1 U9603 ( .A1(n7887), .A2(n9681), .B1(n8049), .B2(n9683), .ZN(n7888)
         );
  AOI21_X1 U9604 ( .B1(n7889), .B2(n9738), .A(n7888), .ZN(n7890) );
  OAI21_X1 U9605 ( .B1(n9900), .B2(n7998), .A(n7890), .ZN(n9903) );
  NAND2_X1 U9606 ( .A1(n9903), .A2(n9728), .ZN(n7898) );
  OAI22_X1 U9607 ( .A1(n9728), .A2(n7892), .B1(n7891), .B2(n9669), .ZN(n7896)
         );
  NOR2_X1 U9608 ( .A1(n7893), .A2(n9901), .ZN(n7894) );
  OR2_X1 U9609 ( .A1(n7902), .A2(n7894), .ZN(n9902) );
  NOR2_X1 U9610 ( .A1(n9902), .A2(n9549), .ZN(n7895) );
  AOI211_X1 U9611 ( .C1(n9660), .C2(n7908), .A(n7896), .B(n7895), .ZN(n7897)
         );
  OAI211_X1 U9612 ( .C1(n9900), .C2(n9953), .A(n7898), .B(n7897), .ZN(P1_U3281) );
  INV_X1 U9613 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7915) );
  OR2_X1 U9614 ( .A1(n7899), .A2(n7908), .ZN(n7900) );
  NAND2_X2 U9615 ( .A1(n7901), .A2(n7900), .ZN(n7989) );
  INV_X1 U9616 ( .A(n9952), .ZN(n7912) );
  AND2_X1 U9617 ( .A1(n7912), .A2(n8049), .ZN(n7992) );
  OR2_X1 U9618 ( .A1(n7912), .A2(n8049), .ZN(n8009) );
  AND2_X1 U9619 ( .A1(n4874), .A2(n8009), .ZN(n9347) );
  XNOR2_X1 U9620 ( .A(n7989), .B(n9347), .ZN(n9954) );
  INV_X1 U9621 ( .A(n7902), .ZN(n7904) );
  NAND2_X1 U9622 ( .A1(n7902), .A2(n9952), .ZN(n7999) );
  INV_X1 U9623 ( .A(n7999), .ZN(n7903) );
  AOI211_X1 U9624 ( .C1(n7912), .C2(n7904), .A(n10210), .B(n7903), .ZN(n9958)
         );
  OR2_X1 U9625 ( .A1(n7925), .A2(n7908), .ZN(n7907) );
  NAND2_X1 U9626 ( .A1(n7907), .A2(n7905), .ZN(n9235) );
  NAND2_X1 U9627 ( .A1(n7907), .A2(n7906), .ZN(n7909) );
  NAND2_X1 U9628 ( .A1(n7908), .A2(n7925), .ZN(n9224) );
  AND2_X1 U9629 ( .A1(n7909), .A2(n9224), .ZN(n9370) );
  XOR2_X1 U9630 ( .A(n9347), .B(n7993), .Z(n7911) );
  OAI222_X1 U9631 ( .A1(n9683), .A2(n7990), .B1(n9681), .B2(n7925), .C1(n7911), 
        .C2(n9678), .ZN(n9944) );
  AOI211_X1 U9632 ( .C1(n9964), .C2(n7912), .A(n9958), .B(n9944), .ZN(n7913)
         );
  OAI21_X1 U9633 ( .B1(n10192), .B2(n9954), .A(n7913), .ZN(n7920) );
  NAND2_X1 U9634 ( .A1(n7920), .A2(n10218), .ZN(n7914) );
  OAI21_X1 U9635 ( .B1(n10218), .B2(n7915), .A(n7914), .ZN(P1_U3487) );
  NOR2_X1 U9636 ( .A1(n7917), .A2(n7916), .ZN(n7918) );
  AND2_X2 U9637 ( .A1(n7919), .A2(n7918), .ZN(n10236) );
  NAND2_X1 U9638 ( .A1(n7920), .A2(n10236), .ZN(n7921) );
  OAI21_X1 U9639 ( .B1(n10236), .B2(n6010), .A(n7921), .ZN(P1_U3534) );
  OAI211_X1 U9640 ( .C1(n7924), .C2(n7923), .A(n7922), .B(n9168), .ZN(n7929)
         );
  OAI22_X1 U9641 ( .A1(n9183), .A2(n7925), .B1(n9181), .B2(n9947), .ZN(n7926)
         );
  AOI211_X1 U9642 ( .C1(n9170), .C2(n9483), .A(n7927), .B(n7926), .ZN(n7928)
         );
  OAI211_X1 U9643 ( .C1(n9952), .C2(n9117), .A(n7929), .B(n7928), .ZN(P1_U3234) );
  INV_X1 U9644 ( .A(n7930), .ZN(n7931) );
  AOI21_X1 U9645 ( .B1(n8502), .B2(n7932), .A(n7931), .ZN(n7933) );
  OAI222_X1 U9646 ( .A1(n8647), .A2(n8058), .B1(n8649), .B2(n8199), .C1(n9910), 
        .C2(n7933), .ZN(n7944) );
  INV_X1 U9647 ( .A(n7944), .ZN(n7943) );
  XNOR2_X1 U9648 ( .A(n7934), .B(n8414), .ZN(n7946) );
  NAND2_X1 U9649 ( .A1(n7946), .A2(n10293), .ZN(n7942) );
  INV_X1 U9650 ( .A(n7935), .ZN(n9923) );
  INV_X1 U9651 ( .A(n7983), .ZN(n7936) );
  AOI211_X1 U9652 ( .C1(n8060), .C2(n9923), .A(n10364), .B(n7936), .ZN(n7945)
         );
  NOR2_X1 U9653 ( .A1(n7937), .A2(n10270), .ZN(n7940) );
  OAI22_X1 U9654 ( .A1(n10272), .A2(n7938), .B1(n8057), .B2(n8903), .ZN(n7939)
         );
  AOI211_X1 U9655 ( .C1(n7945), .C2(n10292), .A(n7940), .B(n7939), .ZN(n7941)
         );
  OAI211_X1 U9656 ( .C1(n10296), .C2(n7943), .A(n7942), .B(n7941), .ZN(
        P2_U3281) );
  AOI211_X1 U9657 ( .C1(n7946), .C2(n10368), .A(n7945), .B(n7944), .ZN(n7949)
         );
  AOI22_X1 U9658 ( .A1(n8060), .A2(n5716), .B1(P2_REG0_REG_15__SCAN_IN), .B2(
        n10370), .ZN(n7947) );
  OAI21_X1 U9659 ( .B1(n7949), .B2(n10370), .A(n7947), .ZN(P2_U3496) );
  AOI22_X1 U9660 ( .A1(n8060), .A2(n5712), .B1(P2_REG1_REG_15__SCAN_IN), .B2(
        n10380), .ZN(n7948) );
  OAI21_X1 U9661 ( .B1(n7949), .B2(n10380), .A(n7948), .ZN(P2_U3535) );
  INV_X1 U9662 ( .A(n7950), .ZN(n7954) );
  OAI222_X1 U9663 ( .A1(n8311), .A2(n7952), .B1(n9070), .B2(n7954), .C1(n7951), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U9664 ( .A1(P1_U3084), .A2(n7955), .B1(n9857), .B2(n7954), .C1(
        n7953), .C2(n8257), .ZN(P1_U3328) );
  AOI21_X1 U9665 ( .B1(n7957), .B2(n9939), .A(n7956), .ZN(n7959) );
  INV_X1 U9666 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9933) );
  AOI22_X1 U9667 ( .A1(n8177), .A2(n9933), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n8180), .ZN(n7958) );
  NOR2_X1 U9668 ( .A1(n7959), .A2(n7958), .ZN(n8179) );
  AOI21_X1 U9669 ( .B1(n7959), .B2(n7958), .A(n8179), .ZN(n7971) );
  INV_X1 U9670 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7960) );
  AOI22_X1 U9671 ( .A1(n8177), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7960), .B2(
        n8180), .ZN(n7964) );
  OAI21_X1 U9672 ( .B1(n7964), .B2(n7963), .A(n8176), .ZN(n7965) );
  NAND2_X1 U9673 ( .A1(n7965), .A2(n10238), .ZN(n7970) );
  INV_X1 U9674 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7967) );
  OAI21_X1 U9675 ( .B1(n8791), .B2(n7967), .A(n7966), .ZN(n7968) );
  AOI21_X1 U9676 ( .B1(n9893), .B2(n8177), .A(n7968), .ZN(n7969) );
  OAI211_X1 U9677 ( .C1(n7971), .C2(n10241), .A(n7970), .B(n7969), .ZN(
        P2_U3259) );
  INV_X1 U9678 ( .A(n7972), .ZN(n7976) );
  OAI222_X1 U9679 ( .A1(n7974), .A2(P2_U3152), .B1(n9070), .B2(n7976), .C1(
        n7973), .C2(n8311), .ZN(P2_U3332) );
  OAI222_X1 U9680 ( .A1(n7977), .A2(P1_U3084), .B1(n9857), .B2(n7976), .C1(
        n7975), .C2(n8257), .ZN(P1_U3327) );
  OAI21_X1 U9681 ( .B1(n8482), .B2(n7978), .A(n8068), .ZN(n7979) );
  AOI222_X1 U9682 ( .A1(n10278), .A2(n7979), .B1(n8668), .B2(n10258), .C1(
        n8670), .C2(n10260), .ZN(n9028) );
  AOI21_X1 U9683 ( .B1(n8482), .B2(n7981), .A(n7980), .ZN(n9023) );
  NAND2_X1 U9684 ( .A1(n9023), .A2(n10293), .ZN(n7988) );
  INV_X1 U9685 ( .A(n8073), .ZN(n7982) );
  AOI211_X1 U9686 ( .C1(n9025), .C2(n7983), .A(n10364), .B(n7982), .ZN(n9024)
         );
  INV_X1 U9687 ( .A(n9025), .ZN(n8157) );
  NOR2_X1 U9688 ( .A1(n8157), .A2(n10270), .ZN(n7986) );
  OAI22_X1 U9689 ( .A1(n10272), .A2(n7984), .B1(n8151), .B2(n8903), .ZN(n7985)
         );
  AOI211_X1 U9690 ( .C1(n9024), .C2(n10292), .A(n7986), .B(n7985), .ZN(n7987)
         );
  OAI211_X1 U9691 ( .C1(n10296), .C2(n9028), .A(n7988), .B(n7987), .ZN(
        P2_U3280) );
  OR2_X1 U9692 ( .A1(n9972), .A2(n7990), .ZN(n9242) );
  NAND2_X1 U9693 ( .A1(n9972), .A2(n7990), .ZN(n9244) );
  OR2_X1 U9694 ( .A1(n8008), .A2(n9348), .ZN(n8159) );
  NAND2_X1 U9695 ( .A1(n8008), .A2(n9348), .ZN(n7991) );
  NAND2_X1 U9696 ( .A1(n8159), .A2(n7991), .ZN(n9971) );
  NAND2_X1 U9697 ( .A1(n8010), .A2(n8009), .ZN(n7994) );
  XOR2_X1 U9698 ( .A(n9348), .B(n7994), .Z(n7996) );
  INV_X1 U9699 ( .A(n9482), .ZN(n8047) );
  OAI22_X1 U9700 ( .A1(n8047), .A2(n9683), .B1(n8049), .B2(n9681), .ZN(n7995)
         );
  AOI21_X1 U9701 ( .B1(n7996), .B2(n9738), .A(n7995), .ZN(n7997) );
  OAI21_X1 U9702 ( .B1(n9971), .B2(n7998), .A(n7997), .ZN(n9975) );
  NAND2_X1 U9703 ( .A1(n9975), .A2(n9728), .ZN(n8004) );
  OAI22_X1 U9704 ( .A1(n9728), .A2(n7002), .B1(n8048), .B2(n9669), .ZN(n8002)
         );
  NAND2_X1 U9705 ( .A1(n7999), .A2(n9972), .ZN(n8000) );
  NAND2_X1 U9706 ( .A1(n8167), .A2(n8000), .ZN(n9974) );
  NOR2_X1 U9707 ( .A1(n9974), .A2(n9549), .ZN(n8001) );
  AOI211_X1 U9708 ( .C1(n9660), .C2(n9972), .A(n8002), .B(n8001), .ZN(n8003)
         );
  OAI211_X1 U9709 ( .C1(n9971), .C2(n9953), .A(n8004), .B(n8003), .ZN(P1_U3279) );
  NAND2_X1 U9710 ( .A1(n9972), .A2(n9483), .ZN(n8158) );
  NAND2_X1 U9711 ( .A1(n9825), .A2(n9482), .ZN(n8005) );
  AND2_X1 U9712 ( .A1(n8158), .A2(n8005), .ZN(n8006) );
  INV_X1 U9713 ( .A(n9481), .ZN(n8037) );
  OR2_X1 U9714 ( .A1(n8131), .A2(n8037), .ZN(n9255) );
  NAND2_X1 U9715 ( .A1(n8131), .A2(n8037), .ZN(n9253) );
  XNOR2_X1 U9716 ( .A(n8132), .B(n9333), .ZN(n9969) );
  INV_X1 U9717 ( .A(n9969), .ZN(n8021) );
  AND2_X1 U9718 ( .A1(n9242), .A2(n8009), .ZN(n9245) );
  OR2_X1 U9719 ( .A1(n9825), .A2(n8047), .ZN(n9252) );
  NAND2_X1 U9720 ( .A1(n9825), .A2(n8047), .ZN(n9241) );
  INV_X1 U9721 ( .A(n9241), .ZN(n8011) );
  OAI21_X1 U9722 ( .B1(n8012), .B2(n9333), .A(n9738), .ZN(n8013) );
  OR2_X1 U9723 ( .A1(n8013), .A2(n8216), .ZN(n8015) );
  INV_X1 U9724 ( .A(n9113), .ZN(n9480) );
  AOI22_X1 U9725 ( .A1(n9480), .A2(n9735), .B1(n9733), .B2(n9482), .ZN(n8014)
         );
  NAND2_X1 U9726 ( .A1(n8015), .A2(n8014), .ZN(n9968) );
  INV_X1 U9727 ( .A(n8131), .ZN(n9966) );
  INV_X1 U9728 ( .A(n8141), .ZN(n8016) );
  OAI211_X1 U9729 ( .C1(n9966), .C2(n8166), .A(n8016), .B(n10187), .ZN(n9965)
         );
  AOI22_X1 U9730 ( .A1(n9703), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8026), .B2(
        n9948), .ZN(n8018) );
  NAND2_X1 U9731 ( .A1(n8131), .A2(n9660), .ZN(n8017) );
  OAI211_X1 U9732 ( .C1(n9965), .C2(n8212), .A(n8018), .B(n8017), .ZN(n8019)
         );
  AOI21_X1 U9733 ( .B1(n9968), .B2(n9728), .A(n8019), .ZN(n8020) );
  OAI21_X1 U9734 ( .B1(n8021), .B2(n9745), .A(n8020), .ZN(P1_U3277) );
  XNOR2_X1 U9735 ( .A(n8023), .B(n8022), .ZN(n8024) );
  XNOR2_X1 U9736 ( .A(n8025), .B(n8024), .ZN(n8031) );
  AOI22_X1 U9737 ( .A1(n9191), .A2(n9482), .B1(n8026), .B2(n9189), .ZN(n8028)
         );
  OAI211_X1 U9738 ( .C1(n9194), .C2(n9113), .A(n8028), .B(n8027), .ZN(n8029)
         );
  AOI21_X1 U9739 ( .B1(n8131), .B2(n9205), .A(n8029), .ZN(n8030) );
  OAI21_X1 U9740 ( .B1(n8031), .B2(n9199), .A(n8030), .ZN(P1_U3213) );
  OR2_X1 U9741 ( .A1(n8044), .A2(n8045), .ZN(n8042) );
  NAND2_X1 U9742 ( .A1(n8042), .A2(n8032), .ZN(n8036) );
  XNOR2_X1 U9743 ( .A(n8034), .B(n8033), .ZN(n8035) );
  XNOR2_X1 U9744 ( .A(n8036), .B(n8035), .ZN(n8041) );
  AND2_X1 U9745 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10065) );
  OAI22_X1 U9746 ( .A1(n9194), .A2(n8037), .B1(n9181), .B2(n8168), .ZN(n8038)
         );
  AOI211_X1 U9747 ( .C1(n9191), .C2(n9483), .A(n10065), .B(n8038), .ZN(n8040)
         );
  NAND2_X1 U9748 ( .A1(n9825), .A2(n9205), .ZN(n8039) );
  OAI211_X1 U9749 ( .C1(n8041), .C2(n9199), .A(n8040), .B(n8039), .ZN(P1_U3232) );
  INV_X1 U9750 ( .A(n8042), .ZN(n8043) );
  AOI21_X1 U9751 ( .B1(n8045), .B2(n8044), .A(n8043), .ZN(n8053) );
  OAI21_X1 U9752 ( .B1(n9194), .B2(n8047), .A(n8046), .ZN(n8051) );
  OAI22_X1 U9753 ( .A1(n9183), .A2(n8049), .B1(n9181), .B2(n8048), .ZN(n8050)
         );
  AOI211_X1 U9754 ( .C1(n9205), .C2(n9972), .A(n8051), .B(n8050), .ZN(n8052)
         );
  OAI21_X1 U9755 ( .B1(n8053), .B2(n9199), .A(n8052), .ZN(P1_U3222) );
  AOI21_X1 U9756 ( .B1(n8055), .B2(n8054), .A(n4554), .ZN(n8063) );
  NOR2_X1 U9757 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8056), .ZN(n8182) );
  OAI22_X1 U9758 ( .A1(n8200), .A2(n8058), .B1(n8652), .B2(n8057), .ZN(n8059)
         );
  AOI211_X1 U9759 ( .C1(n8154), .C2(n8669), .A(n8182), .B(n8059), .ZN(n8062)
         );
  NAND2_X1 U9760 ( .A1(n8060), .A2(n8618), .ZN(n8061) );
  OAI211_X1 U9761 ( .C1(n8063), .C2(n8642), .A(n8062), .B(n8061), .ZN(P2_U3243) );
  INV_X1 U9762 ( .A(n8064), .ZN(n8066) );
  OAI222_X1 U9763 ( .A1(n8311), .A2(n8067), .B1(n9070), .B2(n8066), .C1(n8301), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  NAND2_X1 U9764 ( .A1(n8068), .A2(n8418), .ZN(n8069) );
  XNOR2_X1 U9765 ( .A(n8069), .B(n8504), .ZN(n8070) );
  OAI222_X1 U9766 ( .A1(n8649), .A2(n8243), .B1(n8647), .B2(n8199), .C1(n8070), 
        .C2(n9910), .ZN(n8223) );
  INV_X1 U9767 ( .A(n8223), .ZN(n8079) );
  OAI21_X1 U9768 ( .B1(n8072), .B2(n8504), .A(n8071), .ZN(n8225) );
  NAND2_X1 U9769 ( .A1(n8225), .A2(n10293), .ZN(n8078) );
  AOI211_X1 U9770 ( .C1(n8203), .C2(n8073), .A(n10364), .B(n8123), .ZN(n8224)
         );
  INV_X1 U9771 ( .A(n8203), .ZN(n8230) );
  NOR2_X1 U9772 ( .A1(n8230), .A2(n10270), .ZN(n8076) );
  OAI22_X1 U9773 ( .A1(n10272), .A2(n8074), .B1(n8198), .B2(n8903), .ZN(n8075)
         );
  AOI211_X1 U9774 ( .C1(n8224), .C2(n10292), .A(n8076), .B(n8075), .ZN(n8077)
         );
  OAI211_X1 U9775 ( .C1(n10296), .C2(n8079), .A(n8078), .B(n8077), .ZN(
        P2_U3279) );
  INV_X1 U9776 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10418) );
  NOR2_X1 U9777 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n8080) );
  AOI21_X1 U9778 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n8080), .ZN(n10388) );
  NOR2_X1 U9779 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8081) );
  AOI21_X1 U9780 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n8081), .ZN(n10391) );
  NOR2_X1 U9781 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8082) );
  AOI21_X1 U9782 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n8082), .ZN(n10394) );
  NOR2_X1 U9783 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8083) );
  AOI21_X1 U9784 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n8083), .ZN(n10397) );
  NOR2_X1 U9785 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8084) );
  AOI21_X1 U9786 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n8084), .ZN(n10400) );
  NOR2_X1 U9787 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8093) );
  INV_X1 U9788 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10034) );
  XOR2_X1 U9789 ( .A(n10034), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10430) );
  NAND2_X1 U9790 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n8091) );
  XOR2_X1 U9791 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10428) );
  NAND2_X1 U9792 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n8089) );
  AOI21_X1 U9793 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10383) );
  INV_X1 U9794 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n8086) );
  NAND2_X1 U9795 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n8085) );
  NOR2_X1 U9796 ( .A1(n8086), .A2(n8085), .ZN(n10384) );
  NOR2_X1 U9797 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10384), .ZN(n8087) );
  NOR2_X1 U9798 ( .A1(n10383), .A2(n8087), .ZN(n10412) );
  INV_X1 U9799 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10017) );
  XNOR2_X1 U9800 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n10017), .ZN(n10411) );
  NAND2_X1 U9801 ( .A1(n10412), .A2(n10411), .ZN(n8088) );
  NAND2_X1 U9802 ( .A1(n8089), .A2(n8088), .ZN(n10427) );
  NAND2_X1 U9803 ( .A1(n10428), .A2(n10427), .ZN(n8090) );
  NAND2_X1 U9804 ( .A1(n8091), .A2(n8090), .ZN(n10429) );
  NOR2_X1 U9805 ( .A1(n10430), .A2(n10429), .ZN(n8092) );
  NOR2_X1 U9806 ( .A1(n8093), .A2(n8092), .ZN(n8094) );
  NOR2_X1 U9807 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n8094), .ZN(n10413) );
  AND2_X1 U9808 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n8094), .ZN(n10414) );
  NOR2_X1 U9809 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10414), .ZN(n8095) );
  NOR2_X1 U9810 ( .A1(n10413), .A2(n8095), .ZN(n8096) );
  NAND2_X1 U9811 ( .A1(n8096), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n8098) );
  XOR2_X1 U9812 ( .A(n8096), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10410) );
  NAND2_X1 U9813 ( .A1(n10410), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n8097) );
  NAND2_X1 U9814 ( .A1(n8098), .A2(n8097), .ZN(n8099) );
  NAND2_X1 U9815 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n8099), .ZN(n8102) );
  XNOR2_X1 U9816 ( .A(n8100), .B(n8099), .ZN(n10426) );
  NAND2_X1 U9817 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10426), .ZN(n8101) );
  NAND2_X1 U9818 ( .A1(n8102), .A2(n8101), .ZN(n8103) );
  AND2_X1 U9819 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n8103), .ZN(n8104) );
  XNOR2_X1 U9820 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n8103), .ZN(n10424) );
  NOR2_X1 U9821 ( .A1(n10425), .A2(n10424), .ZN(n10423) );
  NOR2_X1 U9822 ( .A1(n8106), .A2(n8105), .ZN(n8107) );
  XOR2_X1 U9823 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n8106), .Z(n10421) );
  NAND2_X1 U9824 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n8108) );
  OAI21_X1 U9825 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n8108), .ZN(n10408) );
  AOI21_X1 U9826 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10407), .ZN(n10406) );
  NAND2_X1 U9827 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n8109) );
  OAI21_X1 U9828 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n8109), .ZN(n10405) );
  NOR2_X1 U9829 ( .A1(n10406), .A2(n10405), .ZN(n10404) );
  AOI21_X1 U9830 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10404), .ZN(n10403) );
  NOR2_X1 U9831 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8110) );
  AOI21_X1 U9832 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n8110), .ZN(n10402) );
  NAND2_X1 U9833 ( .A1(n10403), .A2(n10402), .ZN(n10401) );
  OAI21_X1 U9834 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10401), .ZN(n10399) );
  NAND2_X1 U9835 ( .A1(n10400), .A2(n10399), .ZN(n10398) );
  OAI21_X1 U9836 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10398), .ZN(n10396) );
  NAND2_X1 U9837 ( .A1(n10397), .A2(n10396), .ZN(n10395) );
  OAI21_X1 U9838 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10395), .ZN(n10393) );
  NAND2_X1 U9839 ( .A1(n10394), .A2(n10393), .ZN(n10392) );
  OAI21_X1 U9840 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10392), .ZN(n10390) );
  NAND2_X1 U9841 ( .A1(n10391), .A2(n10390), .ZN(n10389) );
  OAI21_X1 U9842 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10389), .ZN(n10387) );
  NAND2_X1 U9843 ( .A1(n10388), .A2(n10387), .ZN(n10386) );
  OAI21_X1 U9844 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10386), .ZN(n10417) );
  NOR2_X1 U9845 ( .A1(n10418), .A2(n10417), .ZN(n8111) );
  NAND2_X1 U9846 ( .A1(n10418), .A2(n10417), .ZN(n10416) );
  OAI21_X1 U9847 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n8111), .A(n10416), .ZN(
        n8113) );
  XNOR2_X1 U9848 ( .A(n4822), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n8112) );
  XNOR2_X1 U9849 ( .A(n8113), .B(n8112), .ZN(ADD_1071_U4) );
  NAND2_X1 U9850 ( .A1(n8220), .A2(n8114), .ZN(n8116) );
  OAI211_X1 U9851 ( .C1(n8311), .C2(n8117), .A(n8116), .B(n8115), .ZN(P2_U3330) );
  INV_X1 U9852 ( .A(n8430), .ZN(n8118) );
  XNOR2_X1 U9853 ( .A(n8119), .B(n4503), .ZN(n9022) );
  XNOR2_X1 U9854 ( .A(n8120), .B(n4503), .ZN(n8121) );
  OAI222_X1 U9855 ( .A1(n8649), .A2(n8237), .B1(n8647), .B2(n8122), .C1(n9910), 
        .C2(n8121), .ZN(n9018) );
  INV_X1 U9856 ( .A(n8123), .ZN(n8125) );
  INV_X1 U9857 ( .A(n8247), .ZN(n8124) );
  AOI211_X1 U9858 ( .C1(n9020), .C2(n8125), .A(n10364), .B(n8124), .ZN(n9019)
         );
  NAND2_X1 U9859 ( .A1(n9019), .A2(n10292), .ZN(n8127) );
  INV_X1 U9860 ( .A(n8903), .ZN(n10282) );
  AOI22_X1 U9861 ( .A1(n10296), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8235), .B2(
        n10282), .ZN(n8126) );
  OAI211_X1 U9862 ( .C1(n8128), .C2(n10270), .A(n8127), .B(n8126), .ZN(n8129)
         );
  AOI21_X1 U9863 ( .B1(n9018), .B2(n10272), .A(n8129), .ZN(n8130) );
  OAI21_X1 U9864 ( .B1(n9022), .B2(n8956), .A(n8130), .ZN(P2_U3278) );
  OR2_X1 U9865 ( .A1(n9204), .A2(n9113), .ZN(n9260) );
  NAND2_X1 U9866 ( .A1(n9204), .A2(n9113), .ZN(n9386) );
  NAND2_X1 U9867 ( .A1(n9260), .A2(n9386), .ZN(n9353) );
  XNOR2_X1 U9868 ( .A(n8206), .B(n9353), .ZN(n9819) );
  INV_X1 U9869 ( .A(n9819), .ZN(n8147) );
  NAND2_X1 U9870 ( .A1(n9819), .A2(n9945), .ZN(n8139) );
  INV_X1 U9871 ( .A(n9255), .ZN(n8133) );
  OR2_X1 U9872 ( .A1(n8216), .A2(n8133), .ZN(n8134) );
  XNOR2_X1 U9873 ( .A(n8134), .B(n9353), .ZN(n8137) );
  NAND2_X1 U9874 ( .A1(n9481), .A2(n9733), .ZN(n8135) );
  OAI21_X1 U9875 ( .B1(n9193), .B2(n9683), .A(n8135), .ZN(n8136) );
  AOI21_X1 U9876 ( .B1(n8137), .B2(n9738), .A(n8136), .ZN(n8138) );
  NAND2_X1 U9877 ( .A1(n8139), .A2(n8138), .ZN(n9824) );
  NAND2_X1 U9878 ( .A1(n9824), .A2(n9728), .ZN(n8146) );
  OAI22_X1 U9879 ( .A1(n9728), .A2(n8140), .B1(n9188), .B2(n9669), .ZN(n8144)
         );
  OR2_X1 U9880 ( .A1(n8141), .A2(n9820), .ZN(n8142) );
  NAND2_X1 U9881 ( .A1(n8211), .A2(n8142), .ZN(n9821) );
  NOR2_X1 U9882 ( .A1(n9821), .A2(n9549), .ZN(n8143) );
  AOI211_X1 U9883 ( .C1(n9660), .C2(n9204), .A(n8144), .B(n8143), .ZN(n8145)
         );
  OAI211_X1 U9884 ( .C1(n8147), .C2(n9953), .A(n8146), .B(n8145), .ZN(P1_U3276) );
  NOR3_X1 U9885 ( .A1(n4554), .A2(n8149), .A3(n8148), .ZN(n8150) );
  OAI21_X1 U9886 ( .B1(n4557), .B2(n8150), .A(n8631), .ZN(n8156) );
  AND2_X1 U9887 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8731) );
  OAI22_X1 U9888 ( .A1(n8200), .A2(n8152), .B1(n8652), .B2(n8151), .ZN(n8153)
         );
  AOI211_X1 U9889 ( .C1(n8154), .C2(n8668), .A(n8731), .B(n8153), .ZN(n8155)
         );
  OAI211_X1 U9890 ( .C1(n8157), .C2(n8657), .A(n8156), .B(n8155), .ZN(P2_U3228) );
  NAND2_X1 U9891 ( .A1(n8159), .A2(n8158), .ZN(n8160) );
  XNOR2_X1 U9892 ( .A(n8160), .B(n8161), .ZN(n8172) );
  INV_X1 U9893 ( .A(n8161), .ZN(n9350) );
  XNOR2_X1 U9894 ( .A(n8162), .B(n9350), .ZN(n8164) );
  AOI22_X1 U9895 ( .A1(n9483), .A2(n9733), .B1(n9735), .B2(n9481), .ZN(n8163)
         );
  OAI21_X1 U9896 ( .B1(n8164), .B2(n9678), .A(n8163), .ZN(n8165) );
  AOI21_X1 U9897 ( .B1(n8172), .B2(n9945), .A(n8165), .ZN(n9828) );
  AOI21_X1 U9898 ( .B1(n9825), .B2(n8167), .A(n8166), .ZN(n9826) );
  INV_X1 U9899 ( .A(n9825), .ZN(n8171) );
  INV_X1 U9900 ( .A(n8168), .ZN(n8169) );
  AOI22_X1 U9901 ( .A1(n9703), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8169), .B2(
        n9948), .ZN(n8170) );
  OAI21_X1 U9902 ( .B1(n8171), .B2(n9951), .A(n8170), .ZN(n8174) );
  INV_X1 U9903 ( .A(n8172), .ZN(n9829) );
  NOR2_X1 U9904 ( .A1(n9829), .A2(n9953), .ZN(n8173) );
  AOI211_X1 U9905 ( .C1(n9826), .C2(n9743), .A(n8174), .B(n8173), .ZN(n8175)
         );
  OAI21_X1 U9906 ( .B1(n9703), .B2(n9828), .A(n8175), .ZN(P1_U3278) );
  NAND2_X1 U9907 ( .A1(n8178), .A2(n7938), .ZN(n8736) );
  OAI21_X1 U9908 ( .B1(n8178), .B2(n7938), .A(n8736), .ZN(n8186) );
  AOI21_X1 U9909 ( .B1(n8180), .B2(n9933), .A(n8179), .ZN(n8725) );
  XNOR2_X1 U9910 ( .A(n8725), .B(n8735), .ZN(n8181) );
  NAND2_X1 U9911 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8181), .ZN(n8727) );
  OAI211_X1 U9912 ( .C1(n8181), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10237), .B(
        n8727), .ZN(n8184) );
  AOI21_X1 U9913 ( .B1(n10243), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8182), .ZN(
        n8183) );
  OAI211_X1 U9914 ( .C1(n10239), .C2(n8735), .A(n8184), .B(n8183), .ZN(n8185)
         );
  AOI21_X1 U9915 ( .B1(n10238), .B2(n8186), .A(n8185), .ZN(n8187) );
  INV_X1 U9916 ( .A(n8187), .ZN(P2_U3260) );
  INV_X1 U9917 ( .A(n8190), .ZN(n8192) );
  NAND2_X1 U9918 ( .A1(n8192), .A2(n8191), .ZN(n8193) );
  INV_X1 U9919 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8292) );
  INV_X1 U9920 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8543) );
  MUX2_X1 U9921 ( .A(n8292), .B(n8543), .S(n4483), .Z(n8277) );
  XNOR2_X1 U9922 ( .A(n8277), .B(SI_29_), .ZN(n8195) );
  INV_X1 U9923 ( .A(n8542), .ZN(n8232) );
  XNOR2_X1 U9924 ( .A(n8197), .B(n8196), .ZN(n8205) );
  OAI22_X1 U9925 ( .A1(n8584), .A2(n8243), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8748), .ZN(n8202) );
  OAI22_X1 U9926 ( .A1(n8200), .A2(n8199), .B1(n8652), .B2(n8198), .ZN(n8201)
         );
  AOI211_X1 U9927 ( .C1(n8203), .C2(n8618), .A(n8202), .B(n8201), .ZN(n8204)
         );
  OAI21_X1 U9928 ( .B1(n8205), .B2(n8642), .A(n8204), .ZN(P2_U3230) );
  NAND2_X1 U9929 ( .A1(n9816), .A2(n9193), .ZN(n9385) );
  OAI21_X1 U9930 ( .B1(n9113), .B2(n9820), .A(n8206), .ZN(n8207) );
  OAI21_X1 U9931 ( .B1(n9204), .B2(n9480), .A(n8207), .ZN(n8208) );
  AOI21_X1 U9932 ( .B1(n9355), .B2(n8208), .A(n8533), .ZN(n8209) );
  INV_X1 U9933 ( .A(n8209), .ZN(n9818) );
  INV_X1 U9934 ( .A(n9725), .ZN(n8210) );
  AOI211_X1 U9935 ( .C1(n9816), .C2(n8211), .A(n10210), .B(n8210), .ZN(n9815)
         );
  INV_X1 U9936 ( .A(n8212), .ZN(n9957) );
  INV_X1 U9937 ( .A(n9816), .ZN(n9118) );
  NOR2_X1 U9938 ( .A1(n9118), .A2(n9951), .ZN(n8215) );
  INV_X1 U9939 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8213) );
  OAI22_X1 U9940 ( .A1(n9728), .A2(n8213), .B1(n9112), .B2(n9669), .ZN(n8214)
         );
  AOI211_X1 U9941 ( .C1(n9815), .C2(n9957), .A(n8215), .B(n8214), .ZN(n8219)
         );
  INV_X1 U9942 ( .A(n9719), .ZN(n9182) );
  NAND2_X1 U9943 ( .A1(n9260), .A2(n9255), .ZN(n9377) );
  OAI21_X1 U9944 ( .B1(n8216), .B2(n9377), .A(n9386), .ZN(n8551) );
  XOR2_X1 U9945 ( .A(n9355), .B(n8551), .Z(n8217) );
  OAI222_X1 U9946 ( .A1(n9683), .A2(n9182), .B1(n9681), .B2(n9113), .C1(n8217), 
        .C2(n9678), .ZN(n9814) );
  NAND2_X1 U9947 ( .A1(n9814), .A2(n9728), .ZN(n8218) );
  OAI211_X1 U9948 ( .C1(n9818), .C2(n9745), .A(n8219), .B(n8218), .ZN(P1_U3275) );
  INV_X1 U9949 ( .A(n8220), .ZN(n8221) );
  OAI222_X1 U9950 ( .A1(n9859), .A2(n8222), .B1(P1_U3084), .B2(n4481), .C1(
        n8221), .C2(n9857), .ZN(P1_U3325) );
  INV_X1 U9951 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8761) );
  AOI211_X1 U9952 ( .C1(n8225), .C2(n10368), .A(n8224), .B(n8223), .ZN(n8227)
         );
  MUX2_X1 U9953 ( .A(n8761), .B(n8227), .S(n10382), .Z(n8226) );
  OAI21_X1 U9954 ( .B1(n8230), .B2(n9017), .A(n8226), .ZN(P2_U3537) );
  INV_X1 U9955 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8228) );
  MUX2_X1 U9956 ( .A(n8228), .B(n8227), .S(n10371), .Z(n8229) );
  OAI21_X1 U9957 ( .B1(n8230), .B2(n9061), .A(n8229), .ZN(P2_U3502) );
  OAI222_X1 U9958 ( .A1(n9070), .A2(n8232), .B1(P2_U3152), .B2(n8231), .C1(
        n8292), .C2(n8311), .ZN(P2_U3329) );
  XNOR2_X1 U9959 ( .A(n8234), .B(n8233), .ZN(n8240) );
  AOI22_X1 U9960 ( .A1(n8587), .A2(n8668), .B1(n8639), .B2(n8235), .ZN(n8236)
         );
  NAND2_X1 U9961 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8764) );
  OAI211_X1 U9962 ( .C1(n8237), .C2(n8584), .A(n8236), .B(n8764), .ZN(n8238)
         );
  AOI21_X1 U9963 ( .B1(n9020), .B2(n8618), .A(n8238), .ZN(n8239) );
  OAI21_X1 U9964 ( .B1(n8240), .B2(n8642), .A(n8239), .ZN(P2_U3240) );
  OAI21_X1 U9965 ( .B1(n8506), .B2(n8242), .A(n8241), .ZN(n8244) );
  OAI22_X1 U9966 ( .A1(n8595), .A2(n8649), .B1(n8243), .B2(n8647), .ZN(n8577)
         );
  AOI21_X1 U9967 ( .B1(n8244), .B2(n10278), .A(n8577), .ZN(n9011) );
  XNOR2_X1 U9968 ( .A(n8245), .B(n8506), .ZN(n9014) );
  NAND2_X1 U9969 ( .A1(n9014), .A2(n10293), .ZN(n8252) );
  INV_X1 U9970 ( .A(n8949), .ZN(n8246) );
  AOI211_X1 U9971 ( .C1(n8248), .C2(n8247), .A(n10364), .B(n8246), .ZN(n9013)
         );
  NOR2_X1 U9972 ( .A1(n9062), .A2(n10270), .ZN(n8250) );
  OAI22_X1 U9973 ( .A1(n10272), .A2(n8778), .B1(n8574), .B2(n8903), .ZN(n8249)
         );
  AOI211_X1 U9974 ( .C1(n9013), .C2(n10292), .A(n8250), .B(n8249), .ZN(n8251)
         );
  OAI211_X1 U9975 ( .C1(n10296), .C2(n9011), .A(n8252), .B(n8251), .ZN(
        P2_U3277) );
  OAI222_X1 U9976 ( .A1(n9859), .A2(n8253), .B1(n9857), .B2(n8255), .C1(n9862), 
        .C2(P1_U3084), .ZN(P1_U3350) );
  OAI222_X1 U9977 ( .A1(n8311), .A2(n8256), .B1(n9070), .B2(n8255), .C1(
        P2_U3152), .C2(n8254), .ZN(P2_U3355) );
  OAI222_X1 U9978 ( .A1(n8259), .A2(P1_U3084), .B1(n9857), .B2(n8261), .C1(
        n8258), .C2(n8257), .ZN(P1_U3347) );
  OAI222_X1 U9979 ( .A1(n8311), .A2(n8262), .B1(n9070), .B2(n8261), .C1(
        P2_U3152), .C2(n8260), .ZN(P2_U3352) );
  NAND2_X1 U9980 ( .A1(n7210), .A2(n8263), .ZN(n8265) );
  NAND2_X1 U9981 ( .A1(n8265), .A2(n8488), .ZN(n8264) );
  OAI21_X1 U9982 ( .B1(n8265), .B2(n8488), .A(n8264), .ZN(n10319) );
  OAI211_X1 U9983 ( .C1(n8267), .C2(n8266), .A(n7285), .B(n10278), .ZN(n8269)
         );
  AOI22_X1 U9984 ( .A1(n10260), .A2(n8680), .B1(n10258), .B2(n8678), .ZN(n8268) );
  NAND2_X1 U9985 ( .A1(n8269), .A2(n8268), .ZN(n10318) );
  AOI22_X1 U9986 ( .A1(n10293), .A2(n10319), .B1(n10272), .B2(n10318), .ZN(
        n8275) );
  OAI22_X1 U9987 ( .A1(n8903), .A2(n8272), .B1(n7110), .B2(n10272), .ZN(n8273)
         );
  AOI21_X1 U9988 ( .B1(n10255), .B2(n10314), .A(n8273), .ZN(n8274) );
  OAI211_X1 U9989 ( .C1(n10315), .C2(n10270), .A(n8275), .B(n8274), .ZN(
        P2_U3292) );
  INV_X1 U9990 ( .A(SI_29_), .ZN(n8276) );
  AND2_X1 U9991 ( .A1(n8277), .A2(n8276), .ZN(n8280) );
  INV_X1 U9992 ( .A(n8277), .ZN(n8278) );
  NAND2_X1 U9993 ( .A1(n8278), .A2(SI_29_), .ZN(n8279) );
  INV_X1 U9994 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9858) );
  INV_X1 U9995 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9071) );
  NAND2_X1 U9996 ( .A1(n8296), .A2(SI_30_), .ZN(n8286) );
  INV_X1 U9997 ( .A(n8282), .ZN(n8283) );
  NAND2_X1 U9998 ( .A1(n8284), .A2(n8283), .ZN(n8285) );
  XNOR2_X1 U9999 ( .A(n8287), .B(SI_31_), .ZN(n8288) );
  OR2_X1 U10000 ( .A1(n5377), .A2(n6632), .ZN(n8290) );
  INV_X1 U10001 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8307) );
  NAND2_X1 U10002 ( .A1(n8542), .A2(n8297), .ZN(n8294) );
  OR2_X1 U10003 ( .A1(n5377), .A2(n8292), .ZN(n8293) );
  INV_X1 U10004 ( .A(n8965), .ZN(n8806) );
  OR2_X1 U10005 ( .A1(n5377), .A2(n9071), .ZN(n8298) );
  NOR2_X1 U10006 ( .A1(n8301), .A2(n8528), .ZN(n8302) );
  NOR2_X1 U10007 ( .A1(n8649), .A2(n8302), .ZN(n8814) );
  OR2_X1 U10008 ( .A1(n4485), .A2(n8303), .ZN(n8305) );
  OR2_X1 U10009 ( .A1(n8318), .A2(n8307), .ZN(n8304) );
  AND3_X1 U10010 ( .A1(n8306), .A2(n8305), .A3(n8304), .ZN(n8322) );
  INV_X1 U10011 ( .A(n8322), .ZN(n8658) );
  NAND2_X1 U10012 ( .A1(n8814), .A2(n8658), .ZN(n8958) );
  OAI21_X1 U10013 ( .B1(n9035), .B2(n9017), .A(n8308), .ZN(P2_U3551) );
  OAI222_X1 U10014 ( .A1(n8311), .A2(n8310), .B1(n9070), .B2(n8309), .C1(n5672), .C2(P2_U3152), .ZN(P2_U3336) );
  INV_X1 U10015 ( .A(n8312), .ZN(n8460) );
  NAND2_X1 U10016 ( .A1(n8965), .A2(n8314), .ZN(n8467) );
  INV_X1 U10017 ( .A(n8467), .ZN(n8315) );
  AOI21_X1 U10018 ( .B1(n8812), .B2(n8466), .A(n8315), .ZN(n8319) );
  INV_X1 U10019 ( .A(n8319), .ZN(n8321) );
  INV_X1 U10020 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8960) );
  INV_X1 U10021 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9036) );
  OR2_X1 U10022 ( .A1(n4485), .A2(n9036), .ZN(n8316) );
  OAI211_X1 U10023 ( .C1(n8318), .C2(n8960), .A(n8317), .B(n8316), .ZN(n8813)
         );
  INV_X1 U10024 ( .A(n8813), .ZN(n8324) );
  NOR2_X1 U10025 ( .A1(n8795), .A2(n8324), .ZN(n8473) );
  OAI22_X1 U10026 ( .A1(n8319), .A2(n8473), .B1(n8330), .B2(n8658), .ZN(n8320)
         );
  OAI21_X1 U10027 ( .B1(n8321), .B2(n8795), .A(n8320), .ZN(n8326) );
  AND2_X1 U10028 ( .A1(n8795), .A2(n8324), .ZN(n8468) );
  INV_X1 U10029 ( .A(n8468), .ZN(n8325) );
  NAND2_X1 U10030 ( .A1(n8477), .A2(n8325), .ZN(n8472) );
  INV_X1 U10031 ( .A(n8472), .ZN(n8513) );
  NAND2_X1 U10032 ( .A1(n8329), .A2(n8328), .ZN(n8522) );
  NOR2_X1 U10033 ( .A1(n8856), .A2(n8330), .ZN(n8331) );
  INV_X1 U10034 ( .A(n8332), .ZN(n8443) );
  INV_X1 U10035 ( .A(n8438), .ZN(n8333) );
  NOR3_X1 U10036 ( .A1(n8333), .A2(n8434), .A3(n8465), .ZN(n8442) );
  AND2_X1 U10037 ( .A1(n8430), .A2(n8334), .ZN(n8335) );
  MUX2_X1 U10038 ( .A(n8336), .B(n8335), .S(n8478), .Z(n8424) );
  AND2_X1 U10039 ( .A1(n8398), .A2(n8338), .ZN(n8346) );
  INV_X1 U10040 ( .A(n8338), .ZN(n8339) );
  INV_X1 U10041 ( .A(n8340), .ZN(n8344) );
  NAND2_X1 U10042 ( .A1(n8342), .A2(n8341), .ZN(n8343) );
  AOI21_X1 U10043 ( .B1(n8395), .B2(n8344), .A(n8343), .ZN(n8345) );
  MUX2_X1 U10044 ( .A(n8346), .B(n8345), .S(n8465), .Z(n8397) );
  AND2_X1 U10045 ( .A1(n8352), .A2(n8349), .ZN(n8347) );
  MUX2_X1 U10046 ( .A(n8373), .B(n8347), .S(n8478), .Z(n8376) );
  NAND2_X1 U10047 ( .A1(n8349), .A2(n8348), .ZN(n8350) );
  NAND2_X1 U10048 ( .A1(n8376), .A2(n8350), .ZN(n8353) );
  NAND3_X1 U10049 ( .A1(n8353), .A2(n8352), .A3(n8351), .ZN(n8354) );
  NAND2_X1 U10050 ( .A1(n8354), .A2(n8465), .ZN(n8370) );
  AND2_X1 U10051 ( .A1(n8359), .A2(n8517), .ZN(n8356) );
  OAI211_X1 U10052 ( .C1(n8356), .C2(n8355), .A(n8358), .B(n8363), .ZN(n8357)
         );
  NAND2_X1 U10053 ( .A1(n8357), .A2(n8360), .ZN(n8366) );
  NAND2_X1 U10054 ( .A1(n8359), .A2(n8358), .ZN(n8362) );
  NAND3_X1 U10055 ( .A1(n8362), .A2(n8361), .A3(n8360), .ZN(n8364) );
  NAND2_X1 U10056 ( .A1(n8364), .A2(n8363), .ZN(n8365) );
  MUX2_X1 U10057 ( .A(n8366), .B(n8365), .S(n8478), .Z(n8368) );
  NAND3_X1 U10058 ( .A1(n8368), .A2(n8376), .A3(n8367), .ZN(n8369) );
  NOR2_X1 U10059 ( .A1(n10321), .A2(n8381), .ZN(n8377) );
  AOI21_X1 U10060 ( .B1(n8370), .B2(n8369), .A(n8377), .ZN(n8384) );
  INV_X1 U10061 ( .A(n8371), .ZN(n8375) );
  NAND2_X1 U10062 ( .A1(n8373), .A2(n8372), .ZN(n8374) );
  OAI21_X1 U10063 ( .B1(n8376), .B2(n8375), .A(n8374), .ZN(n8379) );
  INV_X1 U10064 ( .A(n8377), .ZN(n8378) );
  AOI21_X1 U10065 ( .B1(n8379), .B2(n8378), .A(n8465), .ZN(n8383) );
  INV_X1 U10066 ( .A(n8380), .ZN(n8492) );
  NAND3_X1 U10067 ( .A1(n10321), .A2(n8381), .A3(n8478), .ZN(n8382) );
  OAI211_X1 U10068 ( .C1(n8384), .C2(n8383), .A(n8492), .B(n8382), .ZN(n8388)
         );
  INV_X1 U10069 ( .A(n10261), .ZN(n8493) );
  MUX2_X1 U10070 ( .A(n8386), .B(n8385), .S(n8465), .Z(n8387) );
  NAND3_X1 U10071 ( .A1(n8388), .A2(n8493), .A3(n8387), .ZN(n8393) );
  MUX2_X1 U10072 ( .A(n8390), .B(n8389), .S(n8478), .Z(n8391) );
  NAND3_X1 U10073 ( .A1(n8393), .A2(n8392), .A3(n8391), .ZN(n8394) );
  NAND2_X1 U10074 ( .A1(n8395), .A2(n8394), .ZN(n8396) );
  NAND2_X1 U10075 ( .A1(n8397), .A2(n8396), .ZN(n8405) );
  AND2_X1 U10076 ( .A1(n8402), .A2(n8398), .ZN(n8401) );
  INV_X1 U10077 ( .A(n8399), .ZN(n8400) );
  AOI21_X1 U10078 ( .B1(n8405), .B2(n8401), .A(n8400), .ZN(n8407) );
  INV_X1 U10079 ( .A(n8402), .ZN(n8403) );
  AOI21_X1 U10080 ( .B1(n8405), .B2(n8404), .A(n8403), .ZN(n8406) );
  MUX2_X1 U10081 ( .A(n8408), .B(n9909), .S(n8478), .Z(n8409) );
  MUX2_X1 U10082 ( .A(n8412), .B(n8411), .S(n8465), .Z(n8413) );
  MUX2_X1 U10083 ( .A(n8416), .B(n8415), .S(n8465), .Z(n8417) );
  INV_X1 U10084 ( .A(n8504), .ZN(n8421) );
  MUX2_X1 U10085 ( .A(n8419), .B(n8418), .S(n8465), .Z(n8420) );
  NAND3_X1 U10086 ( .A1(n8422), .A2(n8421), .A3(n8420), .ZN(n8423) );
  NAND2_X1 U10087 ( .A1(n8424), .A2(n8423), .ZN(n8431) );
  INV_X1 U10088 ( .A(n8425), .ZN(n8427) );
  INV_X1 U10089 ( .A(n8432), .ZN(n8428) );
  AOI21_X1 U10090 ( .B1(n8431), .B2(n4527), .A(n8428), .ZN(n8429) );
  OAI211_X1 U10091 ( .C1(n8429), .C2(n4908), .A(n8437), .B(n8433), .ZN(n8441)
         );
  INV_X1 U10092 ( .A(n8434), .ZN(n8435) );
  INV_X1 U10093 ( .A(n8439), .ZN(n8440) );
  INV_X1 U10094 ( .A(n8634), .ZN(n8662) );
  AOI21_X1 U10095 ( .B1(n8445), .B2(n8662), .A(n8447), .ZN(n8446) );
  OAI22_X1 U10096 ( .A1(n8448), .A2(n8447), .B1(n8446), .B2(n8465), .ZN(n8450)
         );
  NAND3_X1 U10097 ( .A1(n8887), .A2(n8605), .A3(n8478), .ZN(n8449) );
  NAND2_X1 U10098 ( .A1(n8454), .A2(n8452), .ZN(n8453) );
  INV_X1 U10099 ( .A(n8455), .ZN(n8458) );
  OAI21_X1 U10100 ( .B1(n8842), .B2(n8659), .A(n8456), .ZN(n8457) );
  MUX2_X1 U10101 ( .A(n8458), .B(n8457), .S(n8465), .Z(n8459) );
  MUX2_X1 U10102 ( .A(n8802), .B(n8461), .S(n8465), .Z(n8462) );
  AOI21_X1 U10103 ( .B1(n8827), .B2(n8815), .A(n8462), .ZN(n8463) );
  NAND2_X1 U10104 ( .A1(n8466), .A2(n8467), .ZN(n8811) );
  INV_X1 U10105 ( .A(n8811), .ZN(n8512) );
  OAI21_X1 U10106 ( .B1(n8464), .B2(n8463), .A(n8512), .ZN(n8470) );
  MUX2_X1 U10107 ( .A(n8467), .B(n8466), .S(n8465), .Z(n8469) );
  AOI211_X1 U10108 ( .C1(n8470), .C2(n8469), .A(n8473), .B(n8468), .ZN(n8471)
         );
  AOI21_X1 U10109 ( .B1(n8478), .B2(n8472), .A(n8471), .ZN(n8475) );
  NOR2_X1 U10110 ( .A1(n8474), .A2(n8473), .ZN(n8514) );
  OAI22_X1 U10111 ( .A1(n8475), .A2(n8474), .B1(n8514), .B2(n8478), .ZN(n8476)
         );
  OAI21_X1 U10112 ( .B1(n8478), .B2(n8477), .A(n8476), .ZN(n8480) );
  INV_X1 U10113 ( .A(n6323), .ZN(n8481) );
  INV_X1 U10114 ( .A(n8482), .ZN(n8503) );
  INV_X1 U10115 ( .A(n8483), .ZN(n8486) );
  NAND4_X1 U10116 ( .A1(n8486), .A2(n8485), .A3(n5640), .A4(n8516), .ZN(n8490)
         );
  NOR4_X1 U10117 ( .A1(n8490), .A2(n8489), .A3(n8488), .A4(n8487), .ZN(n8491)
         );
  NAND4_X1 U10118 ( .A1(n8493), .A2(n8492), .A3(n8491), .A4(n10287), .ZN(n8494) );
  NOR4_X1 U10119 ( .A1(n8497), .A2(n8496), .A3(n8495), .A4(n8494), .ZN(n8498)
         );
  NAND4_X1 U10120 ( .A1(n9919), .A2(n8500), .A3(n8499), .A4(n8498), .ZN(n8501)
         );
  NOR4_X1 U10121 ( .A1(n8504), .A2(n8503), .A3(n8502), .A4(n8501), .ZN(n8505)
         );
  NAND3_X1 U10122 ( .A1(n8506), .A2(n8505), .A3(n4503), .ZN(n8507) );
  NOR4_X1 U10123 ( .A1(n8912), .A2(n8935), .A3(n8944), .A4(n8507), .ZN(n8508)
         );
  NAND4_X1 U10124 ( .A1(n8875), .A2(n8881), .A3(n8508), .A4(n8894), .ZN(n8509)
         );
  NOR4_X1 U10125 ( .A1(n8800), .A2(n8510), .A3(n8857), .A4(n8509), .ZN(n8511)
         );
  NAND4_X1 U10126 ( .A1(n8514), .A2(n8513), .A3(n8512), .A4(n8511), .ZN(n8515)
         );
  XNOR2_X1 U10127 ( .A(n8515), .B(n8856), .ZN(n8518) );
  OAI22_X1 U10128 ( .A1(n8518), .A2(n8517), .B1(n8516), .B2(n6323), .ZN(n8519)
         );
  NOR3_X1 U10129 ( .A1(n8525), .A2(n8524), .A3(n8523), .ZN(n8527) );
  MUX2_X1 U10130 ( .A(n8527), .B(n8526), .S(n5672), .Z(n8529) );
  OAI22_X1 U10131 ( .A1(n8531), .A2(n8530), .B1(n8529), .B2(n8528), .ZN(
        P2_U3244) );
  INV_X1 U10132 ( .A(n9755), .ZN(n9556) );
  INV_X1 U10133 ( .A(n9701), .ZN(n9664) );
  INV_X1 U10134 ( .A(n9796), .ZN(n9688) );
  NOR2_X1 U10135 ( .A1(n9809), .A2(n9719), .ZN(n8534) );
  INV_X1 U10136 ( .A(n9809), .ZN(n9730) );
  OR2_X1 U10137 ( .A1(n9804), .A2(n9123), .ZN(n9269) );
  NAND2_X1 U10138 ( .A1(n9804), .A2(n9123), .ZN(n9272) );
  NAND2_X1 U10139 ( .A1(n9269), .A2(n9272), .ZN(n9717) );
  NAND2_X1 U10140 ( .A1(n9800), .A2(n9718), .ZN(n8537) );
  INV_X1 U10141 ( .A(n9718), .ZN(n9680) );
  NAND2_X1 U10142 ( .A1(n9791), .A2(n9682), .ZN(n9279) );
  AOI22_X2 U10143 ( .A1(n9659), .A2(n9658), .B1(n9479), .B2(n9791), .ZN(n9645)
         );
  OAI21_X1 U10144 ( .B1(n9665), .B2(n9655), .A(n9645), .ZN(n8538) );
  OAI21_X1 U10145 ( .B1(n9786), .B2(n9478), .A(n8538), .ZN(n9626) );
  NAND2_X1 U10146 ( .A1(n9779), .A2(n9477), .ZN(n9285) );
  OAI21_X2 U10147 ( .B1(n9626), .B2(n8552), .A(n9285), .ZN(n9613) );
  NOR2_X1 U10148 ( .A1(n8539), .A2(n9638), .ZN(n8540) );
  NAND2_X1 U10149 ( .A1(n9769), .A2(n9618), .ZN(n9298) );
  NAND2_X1 U10150 ( .A1(n9759), .A2(n8541), .ZN(n9411) );
  NAND2_X1 U10151 ( .A1(n9755), .A2(n9572), .ZN(n9412) );
  NAND2_X1 U10152 ( .A1(n9550), .A2(n9559), .ZN(n9551) );
  NAND2_X1 U10153 ( .A1(n8542), .A2(n9214), .ZN(n8545) );
  OR2_X1 U10154 ( .A1(n5822), .A2(n8543), .ZN(n8544) );
  NAND2_X1 U10155 ( .A1(n9749), .A2(n9557), .ZN(n9455) );
  NAND2_X1 U10156 ( .A1(n9708), .A2(n9697), .ZN(n9692) );
  INV_X1 U10157 ( .A(n9759), .ZN(n9571) );
  AOI21_X1 U10158 ( .B1(n9749), .B2(n9552), .A(n9544), .ZN(n9750) );
  INV_X1 U10159 ( .A(n9749), .ZN(n8549) );
  INV_X1 U10160 ( .A(n8546), .ZN(n8547) );
  AOI22_X1 U10161 ( .A1(n9703), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8547), .B2(
        n9948), .ZN(n8548) );
  OAI21_X1 U10162 ( .B1(n8549), .B2(n9951), .A(n8548), .ZN(n8562) );
  INV_X1 U10163 ( .A(n9385), .ZN(n8550) );
  NAND2_X1 U10164 ( .A1(n9809), .A2(n9182), .ZN(n9715) );
  AND2_X1 U10165 ( .A1(n9272), .A2(n9715), .ZN(n9391) );
  OR2_X1 U10166 ( .A1(n9809), .A2(n9182), .ZN(n9713) );
  NAND2_X1 U10167 ( .A1(n9269), .A2(n9713), .ZN(n9266) );
  AOI22_X1 U10168 ( .A1(n9731), .A2(n9391), .B1(n9266), .B2(n9272), .ZN(n9699)
         );
  OR2_X1 U10169 ( .A1(n9800), .A2(n9680), .ZN(n9273) );
  NAND2_X1 U10170 ( .A1(n9800), .A2(n9680), .ZN(n9369) );
  NAND2_X1 U10171 ( .A1(n9699), .A2(n9700), .ZN(n9698) );
  NAND2_X1 U10172 ( .A1(n9698), .A2(n9369), .ZN(n9677) );
  AND2_X1 U10173 ( .A1(n9796), .A2(n9664), .ZN(n9330) );
  OR2_X1 U10174 ( .A1(n9796), .A2(n9664), .ZN(n9331) );
  OAI21_X1 U10175 ( .B1(n9662), .B2(n9658), .A(n9279), .ZN(n9646) );
  INV_X1 U10176 ( .A(n8552), .ZN(n8553) );
  NAND2_X1 U10177 ( .A1(n8553), .A2(n9285), .ZN(n9635) );
  NAND2_X1 U10178 ( .A1(n9634), .A2(n9635), .ZN(n9640) );
  OR2_X1 U10179 ( .A1(n9779), .A2(n9649), .ZN(n9406) );
  NAND2_X1 U10180 ( .A1(n9640), .A2(n9406), .ZN(n9615) );
  NAND2_X1 U10181 ( .A1(n9776), .A2(n9638), .ZN(n9603) );
  NAND2_X2 U10182 ( .A1(n9407), .A2(n9603), .ZN(n9616) );
  NOR2_X2 U10183 ( .A1(n9615), .A2(n9616), .ZN(n9614) );
  NAND2_X1 U10184 ( .A1(n9298), .A2(n9603), .ZN(n9409) );
  OAI21_X1 U10185 ( .B1(n9764), .B2(n9102), .A(n9293), .ZN(n9417) );
  NAND2_X1 U10186 ( .A1(n9764), .A2(n9102), .ZN(n9413) );
  INV_X1 U10187 ( .A(n9416), .ZN(n9414) );
  INV_X1 U10188 ( .A(n9419), .ZN(n8554) );
  INV_X1 U10189 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U10190 ( .A1(n4482), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U10191 ( .A1(n8555), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8556) );
  OAI211_X1 U10192 ( .C1(n8559), .C2(n8558), .A(n8557), .B(n8556), .ZN(n9474)
         );
  AND2_X1 U10193 ( .A1(n9995), .A2(P1_B_REG_SCAN_IN), .ZN(n8560) );
  NOR2_X1 U10194 ( .A1(n9683), .A2(n8560), .ZN(n9538) );
  NOR2_X1 U10195 ( .A1(n9752), .A2(n9703), .ZN(n8561) );
  AOI211_X1 U10196 ( .C1(n9750), .C2(n9743), .A(n8562), .B(n8561), .ZN(n8563)
         );
  OAI21_X1 U10197 ( .B1(n9753), .B2(n9745), .A(n8563), .ZN(P1_U3355) );
  XNOR2_X1 U10198 ( .A(n8564), .B(n8565), .ZN(n8569) );
  OAI22_X1 U10199 ( .A1(n8605), .A2(n8649), .B1(n8596), .B2(n8647), .ZN(n8896)
         );
  AOI22_X1 U10200 ( .A1(n8896), .A2(n8654), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8566) );
  OAI21_X1 U10201 ( .B1(n8904), .B2(n8652), .A(n8566), .ZN(n8567) );
  AOI21_X1 U10202 ( .B1(n8991), .B2(n8618), .A(n8567), .ZN(n8568) );
  OAI21_X1 U10203 ( .B1(n8569), .B2(n8642), .A(n8568), .ZN(P2_U3218) );
  OAI21_X1 U10204 ( .B1(n8572), .B2(n8571), .A(n8570), .ZN(n8573) );
  NAND2_X1 U10205 ( .A1(n8573), .A2(n8631), .ZN(n8579) );
  NAND2_X1 U10206 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8789) );
  INV_X1 U10207 ( .A(n8789), .ZN(n8576) );
  NOR2_X1 U10208 ( .A1(n8652), .A2(n8574), .ZN(n8575) );
  AOI211_X1 U10209 ( .C1(n8654), .C2(n8577), .A(n8576), .B(n8575), .ZN(n8578)
         );
  OAI211_X1 U10210 ( .C1(n9062), .C2(n8657), .A(n8579), .B(n8578), .ZN(
        P2_U3221) );
  XOR2_X1 U10211 ( .A(n8581), .B(n8580), .Z(n8582) );
  NAND2_X1 U10212 ( .A1(n8582), .A2(n8631), .ZN(n8592) );
  NAND2_X1 U10213 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8684) );
  OAI21_X1 U10214 ( .B1(n8584), .B2(n8583), .A(n8684), .ZN(n8585) );
  INV_X1 U10215 ( .A(n8585), .ZN(n8591) );
  INV_X1 U10216 ( .A(n8586), .ZN(n10268) );
  AOI22_X1 U10217 ( .A1(n8587), .A2(n10259), .B1(n8639), .B2(n10268), .ZN(
        n8590) );
  NAND2_X1 U10218 ( .A1(n8618), .A2(n8588), .ZN(n8589) );
  NAND4_X1 U10219 ( .A1(n8592), .A2(n8591), .A3(n8590), .A4(n8589), .ZN(
        P2_U3223) );
  XNOR2_X1 U10220 ( .A(n8594), .B(n8593), .ZN(n8600) );
  OAI22_X1 U10221 ( .A1(n8596), .A2(n8649), .B1(n8595), .B2(n8647), .ZN(n8937)
         );
  AOI22_X1 U10222 ( .A1(n8654), .A2(n8937), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8597) );
  OAI21_X1 U10223 ( .B1(n8652), .B2(n8931), .A(n8597), .ZN(n8598) );
  AOI21_X1 U10224 ( .B1(n9002), .B2(n8618), .A(n8598), .ZN(n8599) );
  OAI21_X1 U10225 ( .B1(n8600), .B2(n8642), .A(n8599), .ZN(P2_U3225) );
  XNOR2_X1 U10226 ( .A(n8603), .B(n8602), .ZN(n8604) );
  XNOR2_X1 U10227 ( .A(n8601), .B(n8604), .ZN(n8611) );
  NOR2_X1 U10228 ( .A1(n8652), .A2(n8868), .ZN(n8609) );
  NOR2_X1 U10229 ( .A1(n8605), .A2(n8647), .ZN(n8606) );
  AOI21_X1 U10230 ( .B1(n8660), .B2(n10258), .A(n8606), .ZN(n8876) );
  OAI22_X1 U10231 ( .A1(n8876), .A2(n8637), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8607), .ZN(n8608) );
  AOI211_X1 U10232 ( .C1(n8980), .C2(n8618), .A(n8609), .B(n8608), .ZN(n8610)
         );
  OAI21_X1 U10233 ( .B1(n8611), .B2(n8642), .A(n8610), .ZN(P2_U3227) );
  XNOR2_X1 U10234 ( .A(n8612), .B(n8613), .ZN(n8620) );
  NOR2_X1 U10235 ( .A1(n8652), .A2(n8888), .ZN(n8617) );
  NOR2_X1 U10236 ( .A1(n8634), .A2(n8647), .ZN(n8614) );
  AOI21_X1 U10237 ( .B1(n8661), .B2(n10258), .A(n8614), .ZN(n8884) );
  OAI22_X1 U10238 ( .A1(n8884), .A2(n8637), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8615), .ZN(n8616) );
  AOI211_X1 U10239 ( .C1(n8887), .C2(n8618), .A(n8617), .B(n8616), .ZN(n8619)
         );
  OAI21_X1 U10240 ( .B1(n8620), .B2(n8642), .A(n8619), .ZN(P2_U3231) );
  XNOR2_X1 U10241 ( .A(n8622), .B(n8621), .ZN(n8627) );
  AOI22_X1 U10242 ( .A1(n8664), .A2(n10258), .B1(n10260), .B2(n8666), .ZN(
        n8946) );
  OAI22_X1 U10243 ( .A1(n8637), .A2(n8946), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8623), .ZN(n8625) );
  NOR2_X1 U10244 ( .A1(n4739), .A2(n8657), .ZN(n8624) );
  AOI211_X1 U10245 ( .C1(n8639), .C2(n8951), .A(n8625), .B(n8624), .ZN(n8626)
         );
  OAI21_X1 U10246 ( .B1(n8627), .B2(n8642), .A(n8626), .ZN(P2_U3235) );
  OAI21_X1 U10247 ( .B1(n8630), .B2(n8629), .A(n8628), .ZN(n8632) );
  NAND2_X1 U10248 ( .A1(n8632), .A2(n8631), .ZN(n8641) );
  OAI22_X1 U10249 ( .A1(n8634), .A2(n8649), .B1(n8633), .B2(n8647), .ZN(n8635)
         );
  INV_X1 U10250 ( .A(n8635), .ZN(n8917) );
  OAI22_X1 U10251 ( .A1(n8917), .A2(n8637), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8636), .ZN(n8638) );
  AOI21_X1 U10252 ( .B1(n8921), .B2(n8639), .A(n8638), .ZN(n8640) );
  OAI211_X1 U10253 ( .C1(n9053), .C2(n8657), .A(n8641), .B(n8640), .ZN(
        P2_U3237) );
  AOI21_X1 U10254 ( .B1(n8644), .B2(n8643), .A(n8642), .ZN(n8646) );
  NAND2_X1 U10255 ( .A1(n8646), .A2(n8645), .ZN(n8656) );
  OAI22_X1 U10256 ( .A1(n8650), .A2(n8649), .B1(n8648), .B2(n8647), .ZN(n8852)
         );
  OAI22_X1 U10257 ( .A1(n8652), .A2(n8847), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8651), .ZN(n8653) );
  AOI21_X1 U10258 ( .B1(n8852), .B2(n8654), .A(n8653), .ZN(n8655) );
  OAI211_X1 U10259 ( .C1(n9044), .C2(n8657), .A(n8656), .B(n8655), .ZN(
        P2_U3242) );
  MUX2_X1 U10260 ( .A(n8658), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8682), .Z(
        P2_U3583) );
  MUX2_X1 U10261 ( .A(n8813), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8682), .Z(
        P2_U3582) );
  MUX2_X1 U10262 ( .A(n8815), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8682), .Z(
        P2_U3580) );
  MUX2_X1 U10263 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8659), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10264 ( .A(n8660), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8682), .Z(
        P2_U3578) );
  MUX2_X1 U10265 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8661), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U10266 ( .A(n8662), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8682), .Z(
        P2_U3575) );
  MUX2_X1 U10267 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8663), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10268 ( .A(n8664), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8682), .Z(
        P2_U3573) );
  MUX2_X1 U10269 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8665), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10270 ( .A(n8666), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8682), .Z(
        P2_U3571) );
  MUX2_X1 U10271 ( .A(n8667), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8682), .Z(
        P2_U3570) );
  MUX2_X1 U10272 ( .A(n8668), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8682), .Z(
        P2_U3569) );
  MUX2_X1 U10273 ( .A(n8669), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8682), .Z(
        P2_U3568) );
  MUX2_X1 U10274 ( .A(n8670), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8682), .Z(
        P2_U3567) );
  MUX2_X1 U10275 ( .A(n8671), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8682), .Z(
        P2_U3566) );
  MUX2_X1 U10276 ( .A(n8672), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8682), .Z(
        P2_U3565) );
  MUX2_X1 U10277 ( .A(n8673), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8682), .Z(
        P2_U3564) );
  MUX2_X1 U10278 ( .A(n8674), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8682), .Z(
        P2_U3563) );
  MUX2_X1 U10279 ( .A(n8675), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8682), .Z(
        P2_U3562) );
  MUX2_X1 U10280 ( .A(n10257), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8682), .Z(
        P2_U3561) );
  MUX2_X1 U10281 ( .A(n8676), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8682), .Z(
        P2_U3560) );
  MUX2_X1 U10282 ( .A(n10259), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8682), .Z(
        P2_U3559) );
  MUX2_X1 U10283 ( .A(n8677), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8682), .Z(
        P2_U3558) );
  MUX2_X1 U10284 ( .A(n8678), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8682), .Z(
        P2_U3557) );
  MUX2_X1 U10285 ( .A(n8679), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8682), .Z(
        P2_U3556) );
  MUX2_X1 U10286 ( .A(n8680), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8682), .Z(
        P2_U3555) );
  MUX2_X1 U10287 ( .A(n8681), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8682), .Z(
        P2_U3554) );
  MUX2_X1 U10288 ( .A(n6672), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8682), .Z(
        P2_U3553) );
  MUX2_X1 U10289 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8683), .S(P2_U3966), .Z(
        P2_U3552) );
  INV_X1 U10290 ( .A(n8684), .ZN(n8687) );
  NOR2_X1 U10291 ( .A1(n10239), .A2(n8685), .ZN(n8686) );
  AOI211_X1 U10292 ( .C1(n10243), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n8687), .B(
        n8686), .ZN(n8697) );
  NAND2_X1 U10293 ( .A1(n8689), .A2(n8688), .ZN(n8690) );
  NAND3_X1 U10294 ( .A1(n10238), .A2(n8691), .A3(n8690), .ZN(n8696) );
  OAI211_X1 U10295 ( .C1(n8694), .C2(n8693), .A(n8692), .B(n10237), .ZN(n8695)
         );
  NAND3_X1 U10296 ( .A1(n8697), .A2(n8696), .A3(n8695), .ZN(P2_U3253) );
  OAI211_X1 U10297 ( .C1(n8700), .C2(n8699), .A(n10237), .B(n8698), .ZN(n8710)
         );
  INV_X1 U10298 ( .A(n8701), .ZN(n8702) );
  AOI21_X1 U10299 ( .B1(n10243), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8702), .ZN(
        n8709) );
  OAI211_X1 U10300 ( .C1(n8705), .C2(n8704), .A(n10238), .B(n8703), .ZN(n8708)
         );
  NAND2_X1 U10301 ( .A1(n9893), .A2(n8706), .ZN(n8707) );
  NAND4_X1 U10302 ( .A1(n8710), .A2(n8709), .A3(n8708), .A4(n8707), .ZN(
        P2_U3254) );
  NAND2_X1 U10303 ( .A1(n9893), .A2(n8711), .ZN(n8724) );
  NOR2_X1 U10304 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8712), .ZN(n8713) );
  AOI21_X1 U10305 ( .B1(n10243), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8713), .ZN(
        n8723) );
  OAI21_X1 U10306 ( .B1(n8716), .B2(n8715), .A(n8714), .ZN(n8717) );
  NAND2_X1 U10307 ( .A1(n10238), .A2(n8717), .ZN(n8722) );
  OAI211_X1 U10308 ( .C1(n8720), .C2(n8719), .A(n10237), .B(n8718), .ZN(n8721)
         );
  NAND4_X1 U10309 ( .A1(n8724), .A2(n8723), .A3(n8722), .A4(n8721), .ZN(
        P2_U3256) );
  NAND2_X1 U10310 ( .A1(n8726), .A2(n8725), .ZN(n8728) );
  NAND2_X1 U10311 ( .A1(n8728), .A2(n8727), .ZN(n8730) );
  XNOR2_X1 U10312 ( .A(n8746), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8729) );
  NOR2_X1 U10313 ( .A1(n8729), .A2(n8730), .ZN(n8750) );
  AOI21_X1 U10314 ( .B1(n8730), .B2(n8729), .A(n8750), .ZN(n8744) );
  INV_X1 U10315 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8733) );
  INV_X1 U10316 ( .A(n8731), .ZN(n8732) );
  OAI21_X1 U10317 ( .B1(n8791), .B2(n8733), .A(n8732), .ZN(n8742) );
  NAND2_X1 U10318 ( .A1(n8735), .A2(n8734), .ZN(n8737) );
  NAND2_X1 U10319 ( .A1(n8746), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8738) );
  OAI21_X1 U10320 ( .B1(n8746), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8738), .ZN(
        n8739) );
  AOI211_X1 U10321 ( .C1(n8740), .C2(n8739), .A(n8745), .B(n9887), .ZN(n8741)
         );
  AOI211_X1 U10322 ( .C1(n9893), .C2(n8746), .A(n8742), .B(n8741), .ZN(n8743)
         );
  OAI21_X1 U10323 ( .B1(n8744), .B2(n10241), .A(n8743), .ZN(P2_U3261) );
  XNOR2_X1 U10324 ( .A(n8767), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n8747) );
  AOI211_X1 U10325 ( .C1(n4556), .C2(n8747), .A(n8766), .B(n9887), .ZN(n8758)
         );
  NOR2_X1 U10326 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8748), .ZN(n8749) );
  AOI21_X1 U10327 ( .B1(n10243), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8749), .ZN(
        n8756) );
  INV_X1 U10328 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8751) );
  AOI21_X1 U10329 ( .B1(n8752), .B2(n8751), .A(n8750), .ZN(n8754) );
  XNOR2_X1 U10330 ( .A(n8767), .B(n8761), .ZN(n8753) );
  NAND2_X1 U10331 ( .A1(n8753), .A2(n8754), .ZN(n8759) );
  OAI211_X1 U10332 ( .C1(n8754), .C2(n8753), .A(n10237), .B(n8759), .ZN(n8755)
         );
  OAI211_X1 U10333 ( .C1(n10239), .C2(n8760), .A(n8756), .B(n8755), .ZN(n8757)
         );
  OR2_X1 U10334 ( .A1(n8758), .A2(n8757), .ZN(P2_U3262) );
  OAI21_X1 U10335 ( .B1(n8761), .B2(n8760), .A(n8759), .ZN(n8763) );
  AOI22_X1 U10336 ( .A1(n8769), .A2(n8780), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8781), .ZN(n8762) );
  NOR2_X1 U10337 ( .A1(n8763), .A2(n8762), .ZN(n8779) );
  AOI21_X1 U10338 ( .B1(n8763), .B2(n8762), .A(n8779), .ZN(n8774) );
  OAI21_X1 U10339 ( .B1(n8791), .B2(n10418), .A(n8764), .ZN(n8765) );
  AOI21_X1 U10340 ( .B1(n9893), .B2(n8769), .A(n8765), .ZN(n8773) );
  INV_X1 U10341 ( .A(n8775), .ZN(n8768) );
  AOI21_X1 U10342 ( .B1(n8770), .B2(n5496), .A(n8776), .ZN(n8771) );
  NAND2_X1 U10343 ( .A1(n10238), .A2(n8771), .ZN(n8772) );
  OAI211_X1 U10344 ( .C1(n8774), .C2(n10241), .A(n8773), .B(n8772), .ZN(
        P2_U3263) );
  NOR2_X1 U10345 ( .A1(n8775), .A2(n8781), .ZN(n8777) );
  INV_X1 U10346 ( .A(n8786), .ZN(n8784) );
  AOI21_X1 U10347 ( .B1(n8781), .B2(n8780), .A(n8779), .ZN(n8782) );
  XOR2_X1 U10348 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8782), .Z(n8785) );
  OAI21_X1 U10349 ( .B1(n8785), .B2(n10241), .A(n10239), .ZN(n8783) );
  AOI21_X1 U10350 ( .B1(n8784), .B2(n10238), .A(n8783), .ZN(n8788) );
  AOI22_X1 U10351 ( .A1(n8786), .A2(n10238), .B1(n10237), .B2(n8785), .ZN(
        n8787) );
  OAI211_X1 U10352 ( .C1(n4822), .C2(n8791), .A(n8790), .B(n8789), .ZN(
        P2_U3264) );
  NOR2_X1 U10353 ( .A1(n10296), .A2(n8958), .ZN(n8798) );
  NOR2_X1 U10354 ( .A1(n9035), .A2(n10270), .ZN(n8792) );
  AOI211_X1 U10355 ( .C1(n10296), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8798), .B(
        n8792), .ZN(n8793) );
  OAI21_X1 U10356 ( .B1(n8794), .B2(n8909), .A(n8793), .ZN(P2_U3265) );
  OAI211_X1 U10357 ( .C1(n8300), .C2(n8804), .A(n9922), .B(n8796), .ZN(n8959)
         );
  NOR2_X1 U10358 ( .A1(n8300), .A2(n10270), .ZN(n8797) );
  AOI211_X1 U10359 ( .C1(n10296), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8798), .B(
        n8797), .ZN(n8799) );
  OAI21_X1 U10360 ( .B1(n8959), .B2(n8909), .A(n8799), .ZN(P2_U3266) );
  XNOR2_X1 U10361 ( .A(n8803), .B(n8811), .ZN(n8962) );
  INV_X1 U10362 ( .A(n8962), .ZN(n8819) );
  AOI211_X1 U10363 ( .C1(n8965), .C2(n8805), .A(n10364), .B(n8804), .ZN(n8964)
         );
  NOR2_X1 U10364 ( .A1(n8806), .A2(n10270), .ZN(n8810) );
  OAI22_X1 U10365 ( .A1(n8808), .A2(n8903), .B1(n8807), .B2(n10272), .ZN(n8809) );
  AOI211_X1 U10366 ( .C1(n8964), .C2(n10292), .A(n8810), .B(n8809), .ZN(n8818)
         );
  AOI22_X1 U10367 ( .A1(n8815), .A2(n10260), .B1(n8814), .B2(n8813), .ZN(n8816) );
  NAND2_X1 U10368 ( .A1(n8963), .A2(n10272), .ZN(n8817) );
  OAI211_X1 U10369 ( .C1(n8819), .C2(n8956), .A(n8818), .B(n8817), .ZN(
        P2_U3267) );
  NAND2_X1 U10370 ( .A1(n8820), .A2(n10293), .ZN(n8829) );
  INV_X1 U10371 ( .A(n8821), .ZN(n8823) );
  OAI22_X1 U10372 ( .A1(n8823), .A2(n8903), .B1(n8822), .B2(n10272), .ZN(n8826) );
  NOR2_X1 U10373 ( .A1(n8824), .A2(n8909), .ZN(n8825) );
  AOI211_X1 U10374 ( .C1(n10283), .C2(n8827), .A(n8826), .B(n8825), .ZN(n8828)
         );
  OAI211_X1 U10375 ( .C1(n8830), .C2(n10296), .A(n8829), .B(n8828), .ZN(
        P2_U3268) );
  XNOR2_X1 U10376 ( .A(n8831), .B(n8833), .ZN(n8972) );
  OAI211_X1 U10377 ( .C1(n8834), .C2(n8833), .A(n8832), .B(n10278), .ZN(n8836)
         );
  NAND2_X1 U10378 ( .A1(n8836), .A2(n8835), .ZN(n8968) );
  AOI211_X1 U10379 ( .C1(n8970), .C2(n8845), .A(n10364), .B(n8838), .ZN(n8969)
         );
  NAND2_X1 U10380 ( .A1(n8969), .A2(n10292), .ZN(n8841) );
  AOI22_X1 U10381 ( .A1(n8839), .A2(n10282), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n10296), .ZN(n8840) );
  OAI211_X1 U10382 ( .C1(n8842), .C2(n10270), .A(n8841), .B(n8840), .ZN(n8843)
         );
  AOI21_X1 U10383 ( .B1(n8968), .B2(n10272), .A(n8843), .ZN(n8844) );
  OAI21_X1 U10384 ( .B1(n8972), .B2(n8956), .A(n8844), .ZN(P2_U3269) );
  AOI21_X1 U10385 ( .B1(n8859), .B2(n8865), .A(n10364), .ZN(n8846) );
  AND2_X1 U10386 ( .A1(n8846), .A2(n8845), .ZN(n8974) );
  NOR2_X1 U10387 ( .A1(n8847), .A2(n8903), .ZN(n8855) );
  INV_X1 U10388 ( .A(n8848), .ZN(n8873) );
  NAND2_X1 U10389 ( .A1(n8873), .A2(n8849), .ZN(n8851) );
  AOI21_X1 U10390 ( .B1(n8857), .B2(n8851), .A(n8850), .ZN(n8854) );
  INV_X1 U10391 ( .A(n8852), .ZN(n8853) );
  OAI21_X1 U10392 ( .B1(n8854), .B2(n9910), .A(n8853), .ZN(n8973) );
  AOI211_X1 U10393 ( .C1(n8974), .C2(n8856), .A(n8855), .B(n8973), .ZN(n8862)
         );
  XNOR2_X1 U10394 ( .A(n8858), .B(n8857), .ZN(n8975) );
  NAND2_X1 U10395 ( .A1(n8975), .A2(n10293), .ZN(n8861) );
  AOI22_X1 U10396 ( .A1(n8859), .A2(n10283), .B1(n10296), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8860) );
  OAI211_X1 U10397 ( .C1(n10296), .C2(n8862), .A(n8861), .B(n8860), .ZN(
        P2_U3270) );
  XNOR2_X1 U10398 ( .A(n8864), .B(n8863), .ZN(n8982) );
  INV_X1 U10399 ( .A(n8865), .ZN(n8866) );
  AOI211_X1 U10400 ( .C1(n8980), .C2(n4735), .A(n10364), .B(n8866), .ZN(n8979)
         );
  NOR2_X1 U10401 ( .A1(n8867), .A2(n10270), .ZN(n8871) );
  OAI22_X1 U10402 ( .A1(n10272), .A2(n8869), .B1(n8868), .B2(n8903), .ZN(n8870) );
  AOI211_X1 U10403 ( .C1(n8979), .C2(n10292), .A(n8871), .B(n8870), .ZN(n8879)
         );
  INV_X1 U10404 ( .A(n8872), .ZN(n8874) );
  OAI211_X1 U10405 ( .C1(n8875), .C2(n8874), .A(n8873), .B(n10278), .ZN(n8877)
         );
  NAND2_X1 U10406 ( .A1(n8877), .A2(n8876), .ZN(n8978) );
  NAND2_X1 U10407 ( .A1(n8978), .A2(n10272), .ZN(n8878) );
  OAI211_X1 U10408 ( .C1(n8982), .C2(n8956), .A(n8879), .B(n8878), .ZN(
        P2_U3271) );
  OAI21_X1 U10409 ( .B1(n8882), .B2(n8881), .A(n10278), .ZN(n8883) );
  OR2_X1 U10410 ( .A1(n4553), .A2(n8883), .ZN(n8885) );
  NAND2_X1 U10411 ( .A1(n8885), .A2(n8884), .ZN(n8984) );
  AOI211_X1 U10412 ( .C1(n8887), .C2(n8899), .A(n10364), .B(n8886), .ZN(n8985)
         );
  NAND2_X1 U10413 ( .A1(n8985), .A2(n10292), .ZN(n8891) );
  INV_X1 U10414 ( .A(n8888), .ZN(n8889) );
  AOI22_X1 U10415 ( .A1(n10296), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8889), 
        .B2(n10282), .ZN(n8890) );
  OAI211_X1 U10416 ( .C1(n4734), .C2(n10270), .A(n8891), .B(n8890), .ZN(n8892)
         );
  AOI21_X1 U10417 ( .B1(n8984), .B2(n10272), .A(n8892), .ZN(n8893) );
  OAI21_X1 U10418 ( .B1(n8983), .B2(n8956), .A(n8893), .ZN(P2_U3272) );
  XNOR2_X1 U10419 ( .A(n8895), .B(n8894), .ZN(n8897) );
  AOI21_X1 U10420 ( .B1(n8897), .B2(n10278), .A(n8896), .ZN(n8994) );
  AOI21_X1 U10421 ( .B1(n8991), .B2(n8919), .A(n10364), .ZN(n8900) );
  NAND2_X1 U10422 ( .A1(n8900), .A2(n8899), .ZN(n8993) );
  OR2_X1 U10423 ( .A1(n8902), .A2(n8901), .ZN(n8990) );
  NAND3_X1 U10424 ( .A1(n8990), .A2(n8989), .A3(n10293), .ZN(n8908) );
  OAI22_X1 U10425 ( .A1(n10272), .A2(n8905), .B1(n8904), .B2(n8903), .ZN(n8906) );
  AOI21_X1 U10426 ( .B1(n8991), .B2(n10283), .A(n8906), .ZN(n8907) );
  OAI211_X1 U10427 ( .C1(n8993), .C2(n8909), .A(n8908), .B(n8907), .ZN(n8910)
         );
  INV_X1 U10428 ( .A(n8910), .ZN(n8911) );
  OAI21_X1 U10429 ( .B1(n10296), .B2(n8994), .A(n8911), .ZN(P2_U3273) );
  XNOR2_X1 U10430 ( .A(n8913), .B(n8912), .ZN(n8998) );
  INV_X1 U10431 ( .A(n8998), .ZN(n8926) );
  OAI211_X1 U10432 ( .C1(n8916), .C2(n8915), .A(n8914), .B(n10278), .ZN(n8918)
         );
  NAND2_X1 U10433 ( .A1(n8918), .A2(n8917), .ZN(n8996) );
  AOI211_X1 U10434 ( .C1(n8920), .C2(n8929), .A(n10364), .B(n8898), .ZN(n8997)
         );
  NAND2_X1 U10435 ( .A1(n8997), .A2(n10292), .ZN(n8923) );
  AOI22_X1 U10436 ( .A1(n10296), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8921), 
        .B2(n10282), .ZN(n8922) );
  OAI211_X1 U10437 ( .C1(n9053), .C2(n10270), .A(n8923), .B(n8922), .ZN(n8924)
         );
  AOI21_X1 U10438 ( .B1(n10272), .B2(n8996), .A(n8924), .ZN(n8925) );
  OAI21_X1 U10439 ( .B1(n8926), .B2(n8956), .A(n8925), .ZN(P2_U3274) );
  XOR2_X1 U10440 ( .A(n8928), .B(n8935), .Z(n9005) );
  INV_X1 U10441 ( .A(n8929), .ZN(n8930) );
  AOI211_X1 U10442 ( .C1(n9002), .C2(n4741), .A(n10364), .B(n8930), .ZN(n9001)
         );
  INV_X1 U10443 ( .A(n8931), .ZN(n8932) );
  AOI22_X1 U10444 ( .A1(n10296), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8932), 
        .B2(n10282), .ZN(n8933) );
  OAI21_X1 U10445 ( .B1(n8934), .B2(n10270), .A(n8933), .ZN(n8940) );
  XNOR2_X1 U10446 ( .A(n8936), .B(n8935), .ZN(n8938) );
  AOI21_X1 U10447 ( .B1(n8938), .B2(n10278), .A(n8937), .ZN(n9004) );
  NOR2_X1 U10448 ( .A1(n9004), .A2(n10296), .ZN(n8939) );
  AOI211_X1 U10449 ( .C1(n9001), .C2(n10292), .A(n8940), .B(n8939), .ZN(n8941)
         );
  OAI21_X1 U10450 ( .B1(n9005), .B2(n8956), .A(n8941), .ZN(P2_U3275) );
  XOR2_X1 U10451 ( .A(n8942), .B(n8944), .Z(n9008) );
  INV_X1 U10452 ( .A(n9008), .ZN(n8957) );
  OAI211_X1 U10453 ( .C1(n4906), .C2(n4907), .A(n10278), .B(n8945), .ZN(n8947)
         );
  NAND2_X1 U10454 ( .A1(n8947), .A2(n8946), .ZN(n9006) );
  AOI211_X1 U10455 ( .C1(n8950), .C2(n8949), .A(n10364), .B(n8948), .ZN(n9007)
         );
  NAND2_X1 U10456 ( .A1(n9007), .A2(n10292), .ZN(n8953) );
  AOI22_X1 U10457 ( .A1(n10296), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8951), 
        .B2(n10282), .ZN(n8952) );
  OAI211_X1 U10458 ( .C1(n4739), .C2(n10270), .A(n8953), .B(n8952), .ZN(n8954)
         );
  AOI21_X1 U10459 ( .B1(n10272), .B2(n9006), .A(n8954), .ZN(n8955) );
  OAI21_X1 U10460 ( .B1(n8957), .B2(n8956), .A(n8955), .ZN(P2_U3276) );
  AND2_X1 U10461 ( .A1(n8959), .A2(n8958), .ZN(n9037) );
  MUX2_X1 U10462 ( .A(n9037), .B(n8960), .S(n10380), .Z(n8961) );
  OAI21_X1 U10463 ( .B1(n8300), .B2(n9017), .A(n8961), .ZN(P2_U3550) );
  NAND2_X1 U10464 ( .A1(n8962), .A2(n10368), .ZN(n8967) );
  NAND2_X1 U10465 ( .A1(n8967), .A2(n8966), .ZN(n9039) );
  MUX2_X1 U10466 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9039), .S(n10382), .Z(
        P2_U3549) );
  INV_X1 U10467 ( .A(n10368), .ZN(n9029) );
  AOI211_X1 U10468 ( .C1(n9026), .C2(n8970), .A(n8969), .B(n8968), .ZN(n8971)
         );
  OAI21_X1 U10469 ( .B1(n8972), .B2(n9029), .A(n8971), .ZN(n9040) );
  MUX2_X1 U10470 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9040), .S(n10382), .Z(
        P2_U3547) );
  INV_X1 U10471 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8976) );
  AOI211_X1 U10472 ( .C1(n8975), .C2(n10368), .A(n8974), .B(n8973), .ZN(n9041)
         );
  MUX2_X1 U10473 ( .A(n8976), .B(n9041), .S(n10382), .Z(n8977) );
  AOI211_X1 U10474 ( .C1(n9026), .C2(n8980), .A(n8979), .B(n8978), .ZN(n8981)
         );
  OAI21_X1 U10475 ( .B1(n8982), .B2(n9029), .A(n8981), .ZN(n9045) );
  MUX2_X1 U10476 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9045), .S(n10382), .Z(
        P2_U3545) );
  INV_X1 U10477 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8987) );
  INV_X1 U10478 ( .A(n8983), .ZN(n8986) );
  MUX2_X1 U10479 ( .A(n8987), .B(n9046), .S(n10382), .Z(n8988) );
  OAI21_X1 U10480 ( .B1(n4734), .B2(n9017), .A(n8988), .ZN(P2_U3544) );
  NAND3_X1 U10481 ( .A1(n8990), .A2(n8989), .A3(n10368), .ZN(n8995) );
  NAND2_X1 U10482 ( .A1(n8991), .A2(n9026), .ZN(n8992) );
  NAND4_X1 U10483 ( .A1(n8995), .A2(n8994), .A3(n8993), .A4(n8992), .ZN(n9049)
         );
  MUX2_X1 U10484 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9049), .S(n10382), .Z(
        P2_U3543) );
  INV_X1 U10485 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8999) );
  AOI211_X1 U10486 ( .C1(n8998), .C2(n10368), .A(n8997), .B(n8996), .ZN(n9050)
         );
  MUX2_X1 U10487 ( .A(n8999), .B(n9050), .S(n10382), .Z(n9000) );
  OAI21_X1 U10488 ( .B1(n9053), .B2(n9017), .A(n9000), .ZN(P2_U3542) );
  AOI21_X1 U10489 ( .B1(n9026), .B2(n9002), .A(n9001), .ZN(n9003) );
  OAI211_X1 U10490 ( .C1(n9005), .C2(n9029), .A(n9004), .B(n9003), .ZN(n9054)
         );
  MUX2_X1 U10491 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9054), .S(n10382), .Z(
        P2_U3541) );
  INV_X1 U10492 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9009) );
  AOI211_X1 U10493 ( .C1(n9008), .C2(n10368), .A(n9007), .B(n9006), .ZN(n9055)
         );
  MUX2_X1 U10494 ( .A(n9009), .B(n9055), .S(n10382), .Z(n9010) );
  OAI21_X1 U10495 ( .B1(n4739), .B2(n9017), .A(n9010), .ZN(P2_U3540) );
  INV_X1 U10496 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9015) );
  INV_X1 U10497 ( .A(n9011), .ZN(n9012) );
  AOI211_X1 U10498 ( .C1(n9014), .C2(n10368), .A(n9013), .B(n9012), .ZN(n9058)
         );
  MUX2_X1 U10499 ( .A(n9015), .B(n9058), .S(n10382), .Z(n9016) );
  OAI21_X1 U10500 ( .B1(n9062), .B2(n9017), .A(n9016), .ZN(P2_U3539) );
  AOI211_X1 U10501 ( .C1(n9026), .C2(n9020), .A(n9019), .B(n9018), .ZN(n9021)
         );
  OAI21_X1 U10502 ( .B1(n9022), .B2(n9029), .A(n9021), .ZN(n9063) );
  MUX2_X1 U10503 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9063), .S(n10382), .Z(
        P2_U3538) );
  INV_X1 U10504 ( .A(n9023), .ZN(n9030) );
  AOI21_X1 U10505 ( .B1(n9026), .B2(n9025), .A(n9024), .ZN(n9027) );
  OAI211_X1 U10506 ( .C1(n9030), .C2(n9029), .A(n9028), .B(n9027), .ZN(n9064)
         );
  MUX2_X1 U10507 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9064), .S(n10382), .Z(
        P2_U3536) );
  MUX2_X1 U10508 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n9031), .S(n10382), .Z(
        P2_U3520) );
  MUX2_X1 U10509 ( .A(n9032), .B(P2_REG0_REG_31__SCAN_IN), .S(n10370), .Z(
        n9033) );
  INV_X1 U10510 ( .A(n9033), .ZN(n9034) );
  OAI21_X1 U10511 ( .B1(n9035), .B2(n9061), .A(n9034), .ZN(P2_U3519) );
  MUX2_X1 U10512 ( .A(n9037), .B(n9036), .S(n10370), .Z(n9038) );
  OAI21_X1 U10513 ( .B1(n8300), .B2(n9061), .A(n9038), .ZN(P2_U3518) );
  MUX2_X1 U10514 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9039), .S(n10371), .Z(
        P2_U3517) );
  MUX2_X1 U10515 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9040), .S(n10371), .Z(
        P2_U3515) );
  INV_X1 U10516 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9042) );
  MUX2_X1 U10517 ( .A(n9042), .B(n9041), .S(n10371), .Z(n9043) );
  MUX2_X1 U10518 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9045), .S(n10371), .Z(
        P2_U3513) );
  MUX2_X1 U10519 ( .A(n9047), .B(n9046), .S(n10371), .Z(n9048) );
  OAI21_X1 U10520 ( .B1(n4734), .B2(n9061), .A(n9048), .ZN(P2_U3512) );
  MUX2_X1 U10521 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9049), .S(n10371), .Z(
        P2_U3511) );
  INV_X1 U10522 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9051) );
  MUX2_X1 U10523 ( .A(n9051), .B(n9050), .S(n10371), .Z(n9052) );
  OAI21_X1 U10524 ( .B1(n9053), .B2(n9061), .A(n9052), .ZN(P2_U3510) );
  MUX2_X1 U10525 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9054), .S(n10371), .Z(
        P2_U3509) );
  INV_X1 U10526 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9056) );
  MUX2_X1 U10527 ( .A(n9056), .B(n9055), .S(n10371), .Z(n9057) );
  OAI21_X1 U10528 ( .B1(n4739), .B2(n9061), .A(n9057), .ZN(P2_U3508) );
  INV_X1 U10529 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9059) );
  MUX2_X1 U10530 ( .A(n9059), .B(n9058), .S(n10371), .Z(n9060) );
  OAI21_X1 U10531 ( .B1(n9062), .B2(n9061), .A(n9060), .ZN(P2_U3507) );
  MUX2_X1 U10532 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9063), .S(n10371), .Z(
        P2_U3505) );
  MUX2_X1 U10533 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9064), .S(n10371), .Z(
        P2_U3499) );
  INV_X1 U10534 ( .A(n9853), .ZN(n9069) );
  NOR4_X1 U10535 ( .A1(n9066), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9065), .A4(
        P2_U3152), .ZN(n9067) );
  AOI21_X1 U10536 ( .B1(n4568), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9067), .ZN(
        n9068) );
  OAI21_X1 U10537 ( .B1(n9069), .B2(n9070), .A(n9068), .ZN(P2_U3327) );
  INV_X1 U10538 ( .A(n9210), .ZN(n9856) );
  OAI222_X1 U10539 ( .A1(n8311), .A2(n9071), .B1(n9070), .B2(n9856), .C1(n5093), .C2(P2_U3152), .ZN(P2_U3328) );
  INV_X1 U10540 ( .A(n9072), .ZN(n9073) );
  MUX2_X1 U10541 ( .A(n9073), .B(n4579), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10542 ( .A(n9074), .ZN(n9076) );
  NOR2_X1 U10543 ( .A1(n9076), .A2(n9075), .ZN(n9078) );
  XNOR2_X1 U10544 ( .A(n9078), .B(n9077), .ZN(n9083) );
  INV_X1 U10545 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9079) );
  OAI22_X1 U10546 ( .A1(n9183), .A2(n9665), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9079), .ZN(n9081) );
  OAI22_X1 U10547 ( .A1(n9194), .A2(n9638), .B1(n9181), .B2(n9630), .ZN(n9080)
         );
  AOI211_X1 U10548 ( .C1(n9779), .C2(n9205), .A(n9081), .B(n9080), .ZN(n9082)
         );
  OAI21_X1 U10549 ( .B1(n9083), .B2(n9199), .A(n9082), .ZN(P1_U3214) );
  AOI21_X1 U10550 ( .B1(n9085), .B2(n9084), .A(n9149), .ZN(n9089) );
  AOI22_X1 U10551 ( .A1(n9191), .A2(n9736), .B1(n9695), .B2(n9189), .ZN(n9086)
         );
  NAND2_X1 U10552 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9535) );
  OAI211_X1 U10553 ( .C1(n9194), .C2(n9664), .A(n9086), .B(n9535), .ZN(n9087)
         );
  AOI21_X1 U10554 ( .B1(n9800), .B2(n9205), .A(n9087), .ZN(n9088) );
  OAI21_X1 U10555 ( .B1(n9089), .B2(n9199), .A(n9088), .ZN(P1_U3217) );
  OAI21_X1 U10556 ( .B1(n9092), .B2(n9091), .A(n9090), .ZN(n9093) );
  NAND2_X1 U10557 ( .A1(n9093), .A2(n9168), .ZN(n9097) );
  NOR2_X1 U10558 ( .A1(n9183), .A2(n9664), .ZN(n9095) );
  OAI22_X1 U10559 ( .A1(n9194), .A2(n9665), .B1(n9181), .B2(n9668), .ZN(n9094)
         );
  AOI211_X1 U10560 ( .C1(P1_REG3_REG_21__SCAN_IN), .C2(P1_U3084), .A(n9095), 
        .B(n9094), .ZN(n9096) );
  OAI211_X1 U10561 ( .C1(n4753), .C2(n9117), .A(n9097), .B(n9096), .ZN(
        P1_U3221) );
  OAI21_X1 U10562 ( .B1(n9099), .B2(n9098), .A(n6289), .ZN(n9100) );
  NAND2_X1 U10563 ( .A1(n9100), .A2(n9168), .ZN(n9106) );
  OAI22_X1 U10564 ( .A1(n9194), .A2(n9102), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9101), .ZN(n9104) );
  OAI22_X1 U10565 ( .A1(n9183), .A2(n9638), .B1(n9181), .B2(n9599), .ZN(n9103)
         );
  AOI211_X1 U10566 ( .C1(n9769), .C2(n9205), .A(n9104), .B(n9103), .ZN(n9105)
         );
  NAND2_X1 U10567 ( .A1(n9106), .A2(n9105), .ZN(P1_U3223) );
  OAI21_X1 U10568 ( .B1(n9201), .B2(n9195), .A(n9107), .ZN(n9108) );
  INV_X1 U10569 ( .A(n9108), .ZN(n9109) );
  OAI21_X1 U10570 ( .B1(n9110), .B2(n9109), .A(n9168), .ZN(n9116) );
  NOR2_X1 U10571 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9111), .ZN(n10091) );
  OAI22_X1 U10572 ( .A1(n9183), .A2(n9113), .B1(n9181), .B2(n9112), .ZN(n9114)
         );
  AOI211_X1 U10573 ( .C1(n9170), .C2(n9719), .A(n10091), .B(n9114), .ZN(n9115)
         );
  OAI211_X1 U10574 ( .C1(n9118), .C2(n9117), .A(n9116), .B(n9115), .ZN(
        P1_U3224) );
  AOI21_X1 U10575 ( .B1(n9121), .B2(n9120), .A(n9119), .ZN(n9126) );
  AOI22_X1 U10576 ( .A1(n9191), .A2(n9734), .B1(n9739), .B2(n9189), .ZN(n9122)
         );
  NAND2_X1 U10577 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10105)
         );
  OAI211_X1 U10578 ( .C1(n9194), .C2(n9123), .A(n9122), .B(n10105), .ZN(n9124)
         );
  AOI21_X1 U10579 ( .B1(n9809), .B2(n9205), .A(n9124), .ZN(n9125) );
  OAI21_X1 U10580 ( .B1(n9126), .B2(n9199), .A(n9125), .ZN(P1_U3226) );
  OAI21_X1 U10581 ( .B1(n9129), .B2(n9128), .A(n9127), .ZN(n9130) );
  NAND2_X1 U10582 ( .A1(n9130), .A2(n9168), .ZN(n9135) );
  OAI22_X1 U10583 ( .A1(n9194), .A2(n9618), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9131), .ZN(n9133) );
  OAI22_X1 U10584 ( .A1(n9183), .A2(n9649), .B1(n9181), .B2(n9621), .ZN(n9132)
         );
  AOI211_X1 U10585 ( .C1(n9776), .C2(n9205), .A(n9133), .B(n9132), .ZN(n9134)
         );
  NAND2_X1 U10586 ( .A1(n9135), .A2(n9134), .ZN(P1_U3227) );
  OAI211_X1 U10587 ( .C1(n9138), .C2(n9137), .A(n9136), .B(n9168), .ZN(n9145)
         );
  AOI22_X1 U10588 ( .A1(n9191), .A2(n7846), .B1(n9139), .B2(n9189), .ZN(n9144)
         );
  NAND2_X1 U10589 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n10025) );
  OAI21_X1 U10590 ( .B1(n9194), .B2(n9140), .A(n10025), .ZN(n9141) );
  AOI21_X1 U10591 ( .B1(n9205), .B2(n9142), .A(n9141), .ZN(n9143) );
  NAND3_X1 U10592 ( .A1(n9145), .A2(n9144), .A3(n9143), .ZN(P1_U3228) );
  INV_X1 U10593 ( .A(n9146), .ZN(n9151) );
  NOR3_X1 U10594 ( .A1(n9149), .A2(n9148), .A3(n9147), .ZN(n9150) );
  OAI21_X1 U10595 ( .B1(n9151), .B2(n9150), .A(n9168), .ZN(n9155) );
  AOI22_X1 U10596 ( .A1(n9170), .A2(n9479), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9154) );
  AOI22_X1 U10597 ( .A1(n9191), .A2(n9718), .B1(n9685), .B2(n9189), .ZN(n9153)
         );
  NAND2_X1 U10598 ( .A1(n9796), .A2(n9205), .ZN(n9152) );
  NAND4_X1 U10599 ( .A1(n9155), .A2(n9154), .A3(n9153), .A4(n9152), .ZN(
        P1_U3231) );
  NAND2_X1 U10600 ( .A1(n9157), .A2(n9156), .ZN(n9158) );
  XOR2_X1 U10601 ( .A(n9159), .B(n9158), .Z(n9164) );
  OAI22_X1 U10602 ( .A1(n9183), .A2(n9682), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9160), .ZN(n9162) );
  OAI22_X1 U10603 ( .A1(n9194), .A2(n9649), .B1(n9181), .B2(n9651), .ZN(n9161)
         );
  AOI211_X1 U10604 ( .C1(n9786), .C2(n9205), .A(n9162), .B(n9161), .ZN(n9163)
         );
  OAI21_X1 U10605 ( .B1(n9164), .B2(n9199), .A(n9163), .ZN(P1_U3233) );
  OAI21_X1 U10606 ( .B1(n9165), .B2(n9167), .A(n9166), .ZN(n9169) );
  NAND2_X1 U10607 ( .A1(n9169), .A2(n9168), .ZN(n9176) );
  AOI22_X1 U10608 ( .A1(n9170), .A2(n7846), .B1(n9191), .B2(n9491), .ZN(n9175)
         );
  OR2_X1 U10609 ( .A1(n9171), .A2(n10007), .ZN(n9174) );
  NAND2_X1 U10610 ( .A1(n9205), .A2(n9172), .ZN(n9173) );
  NAND4_X1 U10611 ( .A1(n9176), .A2(n9175), .A3(n9174), .A4(n9173), .ZN(
        P1_U3235) );
  NAND2_X1 U10612 ( .A1(n4864), .A2(n9178), .ZN(n9180) );
  XNOR2_X1 U10613 ( .A(n9180), .B(n9179), .ZN(n9187) );
  NAND2_X1 U10614 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9501) );
  OAI21_X1 U10615 ( .B1(n9194), .B2(n9680), .A(n9501), .ZN(n9185) );
  OAI22_X1 U10616 ( .A1(n9183), .A2(n9182), .B1(n9181), .B2(n9709), .ZN(n9184)
         );
  AOI211_X1 U10617 ( .C1(n9804), .C2(n9205), .A(n9185), .B(n9184), .ZN(n9186)
         );
  OAI21_X1 U10618 ( .B1(n9187), .B2(n9199), .A(n9186), .ZN(P1_U3236) );
  INV_X1 U10619 ( .A(n9188), .ZN(n9190) );
  AOI22_X1 U10620 ( .A1(n9191), .A2(n9481), .B1(n9190), .B2(n9189), .ZN(n9192)
         );
  NAND2_X1 U10621 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3084), .ZN(n10075)
         );
  OAI211_X1 U10622 ( .C1(n9194), .C2(n9193), .A(n9192), .B(n10075), .ZN(n9203)
         );
  INV_X1 U10623 ( .A(n9195), .ZN(n9200) );
  AOI21_X1 U10624 ( .B1(n9200), .B2(n9197), .A(n9196), .ZN(n9198) );
  AOI211_X1 U10625 ( .C1(n9201), .C2(n9200), .A(n9199), .B(n9198), .ZN(n9202)
         );
  AOI211_X1 U10626 ( .C1(n9205), .C2(n9204), .A(n9203), .B(n9202), .ZN(n9206)
         );
  INV_X1 U10627 ( .A(n9206), .ZN(P1_U3239) );
  NOR4_X1 U10628 ( .A1(n9207), .A2(n10119), .A3(n4481), .A4(n4491), .ZN(n9473)
         );
  OAI21_X1 U10629 ( .B1(n9209), .B2(n9208), .A(P1_B_REG_SCAN_IN), .ZN(n9472)
         );
  NAND2_X1 U10630 ( .A1(n9210), .A2(n9214), .ZN(n9212) );
  OR2_X1 U10631 ( .A1(n5822), .A2(n9858), .ZN(n9211) );
  INV_X1 U10632 ( .A(n9474), .ZN(n9365) );
  INV_X1 U10633 ( .A(n9454), .ZN(n9213) );
  NAND2_X1 U10634 ( .A1(n9213), .A2(n9539), .ZN(n9217) );
  NAND2_X1 U10635 ( .A1(n9853), .A2(n9214), .ZN(n9216) );
  INV_X1 U10636 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9850) );
  OR2_X1 U10637 ( .A1(n5822), .A2(n9850), .ZN(n9215) );
  INV_X1 U10638 ( .A(n9425), .ZN(n9315) );
  NAND3_X1 U10639 ( .A1(n9229), .A2(n9220), .A3(n9231), .ZN(n9221) );
  NAND3_X1 U10640 ( .A1(n9221), .A2(n9233), .A3(n9442), .ZN(n9223) );
  NAND3_X1 U10641 ( .A1(n9223), .A2(n9230), .A3(n9222), .ZN(n9227) );
  INV_X1 U10642 ( .A(n9235), .ZN(n9226) );
  NAND2_X1 U10643 ( .A1(n9244), .A2(n9224), .ZN(n9225) );
  AOI21_X1 U10644 ( .B1(n9227), .B2(n9226), .A(n9225), .ZN(n9240) );
  NAND3_X1 U10645 ( .A1(n9229), .A2(n9228), .A3(n9442), .ZN(n9232) );
  AND2_X1 U10646 ( .A1(n9231), .A2(n9230), .ZN(n9373) );
  NAND2_X1 U10647 ( .A1(n9232), .A2(n9373), .ZN(n9236) );
  INV_X1 U10648 ( .A(n9233), .ZN(n9234) );
  NOR2_X1 U10649 ( .A1(n9235), .A2(n9234), .ZN(n9384) );
  NAND2_X1 U10650 ( .A1(n9236), .A2(n9384), .ZN(n9238) );
  INV_X1 U10651 ( .A(n9242), .ZN(n9237) );
  AOI21_X1 U10652 ( .B1(n9238), .B2(n9370), .A(n9237), .ZN(n9239) );
  MUX2_X1 U10653 ( .A(n9240), .B(n9239), .S(n4673), .Z(n9251) );
  NAND2_X1 U10654 ( .A1(n9253), .A2(n9241), .ZN(n9378) );
  NAND2_X1 U10655 ( .A1(n9244), .A2(n4874), .ZN(n9371) );
  AND2_X1 U10656 ( .A1(n9371), .A2(n9242), .ZN(n9243) );
  OR2_X1 U10657 ( .A1(n9378), .A2(n9243), .ZN(n9249) );
  OR2_X1 U10658 ( .A1(n9245), .A2(n4875), .ZN(n9246) );
  NAND2_X1 U10659 ( .A1(n9246), .A2(n9252), .ZN(n9379) );
  INV_X1 U10660 ( .A(n9379), .ZN(n9247) );
  NAND2_X1 U10661 ( .A1(n9247), .A2(n9255), .ZN(n9248) );
  MUX2_X1 U10662 ( .A(n9249), .B(n9248), .S(n9318), .Z(n9250) );
  AOI21_X1 U10663 ( .B1(n9251), .B2(n9347), .A(n9250), .ZN(n9263) );
  INV_X1 U10664 ( .A(n9353), .ZN(n9259) );
  NAND2_X1 U10665 ( .A1(n9255), .A2(n9252), .ZN(n9254) );
  NAND2_X1 U10666 ( .A1(n9254), .A2(n9253), .ZN(n9257) );
  NAND2_X1 U10667 ( .A1(n9378), .A2(n9255), .ZN(n9256) );
  MUX2_X1 U10668 ( .A(n9257), .B(n9256), .S(n9318), .Z(n9258) );
  NAND2_X1 U10669 ( .A1(n9259), .A2(n9258), .ZN(n9262) );
  MUX2_X1 U10670 ( .A(n9260), .B(n9386), .S(n4673), .Z(n9261) );
  OAI211_X1 U10671 ( .C1(n9263), .C2(n9262), .A(n9355), .B(n9261), .ZN(n9265)
         );
  MUX2_X1 U10672 ( .A(n9388), .B(n9385), .S(n9318), .Z(n9264) );
  NAND3_X1 U10673 ( .A1(n9265), .A2(n9732), .A3(n9264), .ZN(n9268) );
  INV_X1 U10674 ( .A(n9266), .ZN(n9398) );
  MUX2_X1 U10675 ( .A(n9398), .B(n9391), .S(n4673), .Z(n9267) );
  INV_X1 U10676 ( .A(n9369), .ZN(n9270) );
  OR2_X1 U10677 ( .A1(n9330), .A2(n9270), .ZN(n9271) );
  NAND2_X1 U10678 ( .A1(n9369), .A2(n9272), .ZN(n9397) );
  INV_X1 U10679 ( .A(n9397), .ZN(n9275) );
  AND2_X1 U10680 ( .A1(n9331), .A2(n9273), .ZN(n9395) );
  INV_X1 U10681 ( .A(n9395), .ZN(n9274) );
  NAND3_X1 U10682 ( .A1(n9276), .A2(n9400), .A3(n9396), .ZN(n9277) );
  NAND2_X1 U10683 ( .A1(n9278), .A2(n9396), .ZN(n9282) );
  NAND2_X1 U10684 ( .A1(n9396), .A2(n9330), .ZN(n9280) );
  NAND2_X1 U10685 ( .A1(n9280), .A2(n9279), .ZN(n9281) );
  NOR2_X1 U10686 ( .A1(n9328), .A2(n9281), .ZN(n9394) );
  NAND2_X1 U10687 ( .A1(n9282), .A2(n9394), .ZN(n9283) );
  MUX2_X1 U10688 ( .A(n9477), .B(n9779), .S(n9318), .Z(n9284) );
  OR2_X1 U10689 ( .A1(n9616), .A2(n9284), .ZN(n9288) );
  OAI21_X1 U10690 ( .B1(n9616), .B2(n9285), .A(n9288), .ZN(n9286) );
  OAI211_X1 U10691 ( .C1(n9288), .C2(n9649), .A(n9293), .B(n9407), .ZN(n9287)
         );
  INV_X1 U10692 ( .A(n9287), .ZN(n9291) );
  INV_X1 U10693 ( .A(n9288), .ZN(n9289) );
  AOI21_X1 U10694 ( .B1(n9289), .B2(n9779), .A(n9409), .ZN(n9290) );
  MUX2_X1 U10695 ( .A(n9291), .B(n9290), .S(n4673), .Z(n9292) );
  INV_X1 U10696 ( .A(n9293), .ZN(n9587) );
  OAI21_X1 U10697 ( .B1(n9587), .B2(n9586), .A(n9411), .ZN(n9296) );
  NAND2_X1 U10698 ( .A1(n9298), .A2(n9607), .ZN(n9294) );
  NAND2_X1 U10699 ( .A1(n9416), .A2(n9294), .ZN(n9295) );
  MUX2_X1 U10700 ( .A(n9296), .B(n9295), .S(n9318), .Z(n9297) );
  OAI21_X1 U10701 ( .B1(n9303), .B2(n9575), .A(n9297), .ZN(n9305) );
  NOR2_X1 U10702 ( .A1(n9298), .A2(n9607), .ZN(n9299) );
  NOR2_X1 U10703 ( .A1(n9299), .A2(n9764), .ZN(n9301) );
  OAI21_X1 U10704 ( .B1(n9587), .B2(n9607), .A(n9413), .ZN(n9300) );
  MUX2_X1 U10705 ( .A(n9301), .B(n9300), .S(n4673), .Z(n9302) );
  OAI21_X1 U10706 ( .B1(n9303), .B2(n9325), .A(n9302), .ZN(n9304) );
  NAND2_X1 U10707 ( .A1(n9305), .A2(n9304), .ZN(n9307) );
  INV_X1 U10708 ( .A(n9559), .ZN(n9362) );
  MUX2_X1 U10709 ( .A(n9411), .B(n9416), .S(n4673), .Z(n9306) );
  NAND3_X1 U10710 ( .A1(n9307), .A2(n9362), .A3(n9306), .ZN(n9309) );
  MUX2_X1 U10711 ( .A(n9412), .B(n9419), .S(n9318), .Z(n9308) );
  NAND3_X1 U10712 ( .A1(n9425), .A2(n9319), .A3(n9749), .ZN(n9313) );
  NAND2_X1 U10713 ( .A1(n9474), .A2(n9539), .ZN(n9311) );
  NAND2_X1 U10714 ( .A1(n9310), .A2(n9311), .ZN(n9420) );
  AND2_X1 U10715 ( .A1(n9746), .A2(n9312), .ZN(n9458) );
  AOI21_X1 U10716 ( .B1(n9313), .B2(n9420), .A(n9458), .ZN(n9314) );
  MUX2_X1 U10717 ( .A(n9315), .B(n9314), .S(n9318), .Z(n9324) );
  INV_X1 U10718 ( .A(n9557), .ZN(n9475) );
  NAND2_X1 U10719 ( .A1(n9749), .A2(n4673), .ZN(n9316) );
  OAI21_X1 U10720 ( .B1(n4673), .B2(n9557), .A(n9316), .ZN(n9317) );
  NOR2_X1 U10721 ( .A1(n9557), .A2(n9318), .ZN(n9320) );
  INV_X1 U10722 ( .A(n9420), .ZN(n9321) );
  INV_X1 U10723 ( .A(n9746), .ZN(n9540) );
  INV_X1 U10724 ( .A(n9422), .ZN(n9465) );
  OAI21_X1 U10725 ( .B1(n9322), .B2(n9321), .A(n9465), .ZN(n9323) );
  INV_X1 U10726 ( .A(n9325), .ZN(n9327) );
  INV_X1 U10727 ( .A(n9575), .ZN(n9361) );
  INV_X1 U10728 ( .A(n9400), .ZN(n9329) );
  NOR2_X1 U10729 ( .A1(n9329), .A2(n9328), .ZN(n9647) );
  INV_X1 U10730 ( .A(n9658), .ZN(n9661) );
  INV_X1 U10731 ( .A(n9330), .ZN(n9332) );
  NAND2_X1 U10732 ( .A1(n9332), .A2(n9331), .ZN(n9676) );
  INV_X1 U10733 ( .A(n9700), .ZN(n9357) );
  INV_X1 U10734 ( .A(n9333), .ZN(n9352) );
  NOR4_X1 U10735 ( .A1(n9337), .A2(n9336), .A3(n9335), .A4(n9334), .ZN(n9341)
         );
  NAND4_X1 U10736 ( .A1(n9341), .A2(n9340), .A3(n9339), .A4(n9338), .ZN(n9345)
         );
  NOR4_X1 U10737 ( .A1(n9345), .A2(n9344), .A3(n9343), .A4(n9342), .ZN(n9349)
         );
  NAND4_X1 U10738 ( .A1(n9349), .A2(n9348), .A3(n9347), .A4(n9346), .ZN(n9351)
         );
  NOR4_X1 U10739 ( .A1(n9353), .A2(n9352), .A3(n9351), .A4(n9350), .ZN(n9354)
         );
  NAND3_X1 U10740 ( .A1(n9732), .A2(n9355), .A3(n9354), .ZN(n9356) );
  NOR4_X1 U10741 ( .A1(n9676), .A2(n9357), .A3(n9717), .A4(n9356), .ZN(n9358)
         );
  NAND4_X1 U10742 ( .A1(n9635), .A2(n9647), .A3(n9661), .A4(n9358), .ZN(n9359)
         );
  NOR3_X1 U10743 ( .A1(n9605), .A2(n9616), .A3(n9359), .ZN(n9360) );
  NAND4_X1 U10744 ( .A1(n9589), .A2(n9362), .A3(n9361), .A4(n9360), .ZN(n9363)
         );
  NOR4_X1 U10745 ( .A1(n9458), .A2(n9454), .A3(n9364), .A4(n9363), .ZN(n9366)
         );
  AOI21_X1 U10746 ( .B1(n9365), .B2(n9310), .A(n9422), .ZN(n9457) );
  AOI21_X1 U10747 ( .B1(n9366), .B2(n9457), .A(n6284), .ZN(n9427) );
  INV_X1 U10748 ( .A(n9427), .ZN(n9367) );
  NAND2_X1 U10749 ( .A1(n9779), .A2(n9649), .ZN(n9403) );
  NAND3_X1 U10750 ( .A1(n9394), .A2(n9369), .A3(n9403), .ZN(n9393) );
  INV_X1 U10751 ( .A(n9391), .ZN(n9375) );
  OR3_X1 U10752 ( .A1(n9378), .A2(n9371), .A3(n4876), .ZN(n9383) );
  INV_X1 U10753 ( .A(n9383), .ZN(n9372) );
  NAND4_X1 U10754 ( .A1(n9385), .A2(n9373), .A3(n9372), .A4(n9386), .ZN(n9374)
         );
  OR3_X1 U10755 ( .A1(n9393), .A2(n9375), .A3(n9374), .ZN(n9447) );
  NOR2_X1 U10756 ( .A1(n9447), .A2(n9376), .ZN(n9410) );
  INV_X1 U10757 ( .A(n9377), .ZN(n9382) );
  INV_X1 U10758 ( .A(n9378), .ZN(n9380) );
  NAND2_X1 U10759 ( .A1(n9380), .A2(n9379), .ZN(n9381) );
  OAI211_X1 U10760 ( .C1(n9384), .C2(n9383), .A(n9382), .B(n9381), .ZN(n9387)
         );
  NAND3_X1 U10761 ( .A1(n9387), .A2(n9386), .A3(n9385), .ZN(n9389) );
  NAND2_X1 U10762 ( .A1(n9389), .A2(n9388), .ZN(n9390) );
  NAND2_X1 U10763 ( .A1(n9391), .A2(n9390), .ZN(n9392) );
  OR2_X1 U10764 ( .A1(n9393), .A2(n9392), .ZN(n9408) );
  INV_X1 U10765 ( .A(n9394), .ZN(n9402) );
  OAI211_X1 U10766 ( .C1(n9398), .C2(n9397), .A(n9396), .B(n9395), .ZN(n9399)
         );
  INV_X1 U10767 ( .A(n9399), .ZN(n9401) );
  OAI21_X1 U10768 ( .B1(n9402), .B2(n9401), .A(n9400), .ZN(n9404) );
  NAND2_X1 U10769 ( .A1(n9404), .A2(n9403), .ZN(n9405) );
  NAND4_X1 U10770 ( .A1(n9408), .A2(n9407), .A3(n9406), .A4(n9405), .ZN(n9445)
         );
  OAI21_X1 U10771 ( .B1(n9410), .B2(n9445), .A(n4890), .ZN(n9415) );
  OAI211_X1 U10772 ( .C1(n9414), .C2(n9413), .A(n9412), .B(n9411), .ZN(n9452)
         );
  AOI21_X1 U10773 ( .B1(n9416), .B2(n9415), .A(n9452), .ZN(n9421) );
  OAI211_X1 U10774 ( .C1(n9452), .C2(n4891), .A(n9419), .B(n9418), .ZN(n9450)
         );
  OAI211_X1 U10775 ( .C1(n9421), .C2(n9450), .A(n9420), .B(n9455), .ZN(n9424)
         );
  AOI211_X1 U10776 ( .C1(n9425), .C2(n9424), .A(n9423), .B(n9422), .ZN(n9426)
         );
  NOR2_X1 U10777 ( .A1(n9427), .A2(n9426), .ZN(n9428) );
  INV_X1 U10778 ( .A(n9429), .ZN(n9434) );
  NAND2_X1 U10779 ( .A1(n9430), .A2(n6284), .ZN(n9433) );
  INV_X1 U10780 ( .A(n9431), .ZN(n9432) );
  OAI211_X1 U10781 ( .C1(n9434), .C2(n9433), .A(n9432), .B(n7592), .ZN(n9436)
         );
  OAI211_X1 U10782 ( .C1(n9438), .C2(n9437), .A(n9436), .B(n9435), .ZN(n9441)
         );
  NAND3_X1 U10783 ( .A1(n9441), .A2(n9440), .A3(n9439), .ZN(n9444) );
  AND3_X1 U10784 ( .A1(n9444), .A2(n9443), .A3(n9442), .ZN(n9448) );
  INV_X1 U10785 ( .A(n9445), .ZN(n9446) );
  OAI21_X1 U10786 ( .B1(n9448), .B2(n9447), .A(n9446), .ZN(n9449) );
  AOI21_X1 U10787 ( .B1(n4890), .B2(n9449), .A(n9575), .ZN(n9453) );
  INV_X1 U10788 ( .A(n9450), .ZN(n9451) );
  OAI21_X1 U10789 ( .B1(n9453), .B2(n9452), .A(n9451), .ZN(n9456) );
  AOI21_X1 U10790 ( .B1(n9456), .B2(n9455), .A(n9454), .ZN(n9461) );
  INV_X1 U10791 ( .A(n9457), .ZN(n9460) );
  INV_X1 U10792 ( .A(n9458), .ZN(n9459) );
  OAI21_X1 U10793 ( .B1(n9461), .B2(n9460), .A(n9459), .ZN(n9462) );
  XNOR2_X1 U10794 ( .A(n9462), .B(n9670), .ZN(n9463) );
  INV_X1 U10795 ( .A(n9464), .ZN(n9466) );
  OAI21_X1 U10796 ( .B1(n9470), .B2(n9469), .A(n9468), .ZN(n9471) );
  OAI21_X1 U10797 ( .B1(n9473), .B2(n9472), .A(n9471), .ZN(P1_U3240) );
  MUX2_X1 U10798 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9474), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10799 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9475), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10800 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9476), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10801 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9592), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10802 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9607), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10803 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9591), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10804 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9608), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10805 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9477), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10806 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9478), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10807 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9479), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10808 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9701), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10809 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9718), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10810 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9736), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10811 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9719), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10812 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9734), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10813 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9480), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10814 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9481), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10815 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9482), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10816 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9483), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10817 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n5030), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10818 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9484), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10819 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9485), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10820 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9486), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10821 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9487), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10822 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9488), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10823 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9489), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10824 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n7846), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10825 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9490), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10826 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9491), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10827 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9492), .S(P1_U4006), .Z(
        P1_U3555) );
  AOI22_X1 U10828 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n9525), .B1(n9521), .B2(
        n9524), .ZN(n9500) );
  XNOR2_X1 U10829 ( .A(n10108), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10113) );
  INV_X1 U10830 ( .A(n10092), .ZN(n9497) );
  XOR2_X1 U10831 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10092), .Z(n10095) );
  NAND2_X1 U10832 ( .A1(n10080), .A2(n9494), .ZN(n9495) );
  XNOR2_X1 U10833 ( .A(n9494), .B(n9509), .ZN(n10082) );
  NAND2_X1 U10834 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n10082), .ZN(n10081) );
  NAND2_X1 U10835 ( .A1(n10095), .A2(n10096), .ZN(n10094) );
  NAND2_X1 U10836 ( .A1(n10113), .A2(n10112), .ZN(n10110) );
  OAI21_X1 U10837 ( .B1(n10108), .B2(n9498), .A(n10110), .ZN(n9499) );
  NOR2_X1 U10838 ( .A1(n9500), .A2(n9499), .ZN(n9523) );
  AOI21_X1 U10839 ( .B1(n9500), .B2(n9499), .A(n9523), .ZN(n9519) );
  INV_X1 U10840 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9502) );
  OAI21_X1 U10841 ( .B1(n10116), .B2(n9502), .A(n9501), .ZN(n9517) );
  NOR2_X1 U10842 ( .A1(n9521), .A2(n9503), .ZN(n9504) );
  AOI21_X1 U10843 ( .B1(n9521), .B2(n9503), .A(n9504), .ZN(n9515) );
  NOR2_X1 U10844 ( .A1(n9506), .A2(n9505), .ZN(n9508) );
  NAND2_X1 U10845 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n10092), .ZN(n9511) );
  OAI21_X1 U10846 ( .B1(n10092), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9511), .ZN(
        n10088) );
  NOR2_X1 U10847 ( .A1(n10089), .A2(n10088), .ZN(n10087) );
  AOI21_X1 U10848 ( .B1(n10092), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10087), 
        .ZN(n10101) );
  NAND2_X1 U10849 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9513), .ZN(n9512) );
  OAI21_X1 U10850 ( .B1(n9513), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9512), .ZN(
        n10102) );
  NOR2_X1 U10851 ( .A1(n10101), .A2(n10102), .ZN(n10100) );
  AOI211_X1 U10852 ( .C1(n9515), .C2(n9514), .A(n9520), .B(n10086), .ZN(n9516)
         );
  AOI211_X1 U10853 ( .C1(n10093), .C2(n9521), .A(n9517), .B(n9516), .ZN(n9518)
         );
  OAI21_X1 U10854 ( .B1(n9519), .B2(n10070), .A(n9518), .ZN(P1_U3259) );
  INV_X1 U10855 ( .A(n9531), .ZN(n9529) );
  INV_X1 U10856 ( .A(n9522), .ZN(n9528) );
  XOR2_X1 U10857 ( .A(n9526), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9530) );
  OAI21_X1 U10858 ( .B1(n9530), .B2(n10070), .A(n10107), .ZN(n9527) );
  AOI21_X1 U10859 ( .B1(n9529), .B2(n9528), .A(n9527), .ZN(n9534) );
  INV_X1 U10860 ( .A(n10070), .ZN(n10111) );
  AOI22_X1 U10861 ( .A1(n9531), .A2(n10104), .B1(n10111), .B2(n9530), .ZN(
        n9533) );
  MUX2_X1 U10862 ( .A(n9534), .B(n9533), .S(n9532), .Z(n9536) );
  OAI211_X1 U10863 ( .C1(n9537), .C2(n10116), .A(n9536), .B(n9535), .ZN(
        P1_U3260) );
  XNOR2_X1 U10864 ( .A(n9543), .B(n9746), .ZN(n9748) );
  NAND2_X1 U10865 ( .A1(n9539), .A2(n9538), .ZN(n9961) );
  NOR2_X1 U10866 ( .A1(n9961), .A2(n9703), .ZN(n9547) );
  NOR2_X1 U10867 ( .A1(n9540), .A2(n9951), .ZN(n9541) );
  AOI211_X1 U10868 ( .C1(n9703), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9547), .B(
        n9541), .ZN(n9542) );
  OAI21_X1 U10869 ( .B1(n9549), .B2(n9748), .A(n9542), .ZN(P1_U3261) );
  NOR2_X1 U10870 ( .A1(n9545), .A2(n9951), .ZN(n9546) );
  AOI211_X1 U10871 ( .C1(n9703), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9547), .B(
        n9546), .ZN(n9548) );
  OAI21_X1 U10872 ( .B1(n9549), .B2(n9962), .A(n9548), .ZN(P1_U3262) );
  OAI21_X1 U10873 ( .B1(n9550), .B2(n9559), .A(n9551), .ZN(n9758) );
  AOI211_X1 U10874 ( .C1(n9755), .C2(n9567), .A(n10210), .B(n4763), .ZN(n9754)
         );
  INV_X1 U10875 ( .A(n9553), .ZN(n9554) );
  AOI22_X1 U10876 ( .A1(n9703), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9554), .B2(
        n9948), .ZN(n9555) );
  OAI21_X1 U10877 ( .B1(n9556), .B2(n9951), .A(n9555), .ZN(n9564) );
  NOR2_X1 U10878 ( .A1(n9557), .A2(n9683), .ZN(n9562) );
  AOI211_X1 U10879 ( .C1(n9560), .C2(n9559), .A(n9678), .B(n9558), .ZN(n9561)
         );
  NOR2_X1 U10880 ( .A1(n9757), .A2(n9703), .ZN(n9563) );
  AOI211_X1 U10881 ( .C1(n9754), .C2(n9957), .A(n9564), .B(n9563), .ZN(n9565)
         );
  OAI21_X1 U10882 ( .B1(n9745), .B2(n9758), .A(n9565), .ZN(P1_U3263) );
  XOR2_X1 U10883 ( .A(n9575), .B(n9566), .Z(n9763) );
  INV_X1 U10884 ( .A(n9582), .ZN(n9568) );
  AOI21_X1 U10885 ( .B1(n9759), .B2(n9568), .A(n4764), .ZN(n9760) );
  AOI22_X1 U10886 ( .A1(n9703), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9569), .B2(
        n9948), .ZN(n9570) );
  OAI21_X1 U10887 ( .B1(n9571), .B2(n9951), .A(n9570), .ZN(n9579) );
  NOR2_X1 U10888 ( .A1(n9572), .A2(n9683), .ZN(n9577) );
  AOI211_X1 U10889 ( .C1(n9575), .C2(n9574), .A(n9678), .B(n9573), .ZN(n9576)
         );
  AOI211_X1 U10890 ( .C1(n9733), .C2(n9607), .A(n9577), .B(n9576), .ZN(n9762)
         );
  NOR2_X1 U10891 ( .A1(n9762), .A2(n9703), .ZN(n9578) );
  AOI211_X1 U10892 ( .C1(n9743), .C2(n9760), .A(n9579), .B(n9578), .ZN(n9580)
         );
  OAI21_X1 U10893 ( .B1(n9763), .B2(n9745), .A(n9580), .ZN(P1_U3264) );
  XOR2_X1 U10894 ( .A(n9589), .B(n9581), .Z(n9768) );
  INV_X1 U10895 ( .A(n9598), .ZN(n9583) );
  AOI21_X1 U10896 ( .B1(n9764), .B2(n9583), .A(n9582), .ZN(n9765) );
  AOI22_X1 U10897 ( .A1(n9703), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9584), .B2(
        n9948), .ZN(n9585) );
  OAI21_X1 U10898 ( .B1(n9586), .B2(n9951), .A(n9585), .ZN(n9595) );
  NOR2_X1 U10899 ( .A1(n9588), .A2(n9587), .ZN(n9590) );
  XNOR2_X1 U10900 ( .A(n9590), .B(n9589), .ZN(n9593) );
  AOI222_X1 U10901 ( .A1(n9738), .A2(n9593), .B1(n9592), .B2(n9735), .C1(n9591), .C2(n9733), .ZN(n9767) );
  NOR2_X1 U10902 ( .A1(n9767), .A2(n9703), .ZN(n9594) );
  AOI211_X1 U10903 ( .C1(n9765), .C2(n9743), .A(n9595), .B(n9594), .ZN(n9596)
         );
  OAI21_X1 U10904 ( .B1(n9768), .B2(n9745), .A(n9596), .ZN(P1_U3265) );
  XOR2_X1 U10905 ( .A(n9605), .B(n9597), .Z(n9773) );
  AOI21_X1 U10906 ( .B1(n9769), .B2(n9619), .A(n9598), .ZN(n9770) );
  INV_X1 U10907 ( .A(n9599), .ZN(n9600) );
  AOI22_X1 U10908 ( .A1(n9703), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9600), .B2(
        n9948), .ZN(n9601) );
  OAI21_X1 U10909 ( .B1(n9602), .B2(n9951), .A(n9601), .ZN(n9611) );
  INV_X1 U10910 ( .A(n9603), .ZN(n9604) );
  NOR2_X1 U10911 ( .A1(n9614), .A2(n9604), .ZN(n9606) );
  XNOR2_X1 U10912 ( .A(n9606), .B(n9605), .ZN(n9609) );
  AOI222_X1 U10913 ( .A1(n9738), .A2(n9609), .B1(n9608), .B2(n9733), .C1(n9607), .C2(n9735), .ZN(n9772) );
  NOR2_X1 U10914 ( .A1(n9772), .A2(n9703), .ZN(n9610) );
  AOI211_X1 U10915 ( .C1(n9770), .C2(n9743), .A(n9611), .B(n9610), .ZN(n9612)
         );
  OAI21_X1 U10916 ( .B1(n9773), .B2(n9745), .A(n9612), .ZN(P1_U3266) );
  XNOR2_X1 U10917 ( .A(n9613), .B(n9616), .ZN(n9778) );
  AOI22_X1 U10918 ( .A1(n9776), .A2(n9660), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9703), .ZN(n9625) );
  AOI21_X1 U10919 ( .B1(n9616), .B2(n9615), .A(n9614), .ZN(n9617) );
  OAI222_X1 U10920 ( .A1(n9681), .A2(n9649), .B1(n9683), .B2(n9618), .C1(n9678), .C2(n9617), .ZN(n9774) );
  INV_X1 U10921 ( .A(n9619), .ZN(n9620) );
  AOI211_X1 U10922 ( .C1(n9776), .C2(n9627), .A(n10210), .B(n9620), .ZN(n9775)
         );
  INV_X1 U10923 ( .A(n9775), .ZN(n9622) );
  OAI22_X1 U10924 ( .A1(n9622), .A2(n9670), .B1(n9669), .B2(n9621), .ZN(n9623)
         );
  OAI21_X1 U10925 ( .B1(n9774), .B2(n9623), .A(n9728), .ZN(n9624) );
  OAI211_X1 U10926 ( .C1(n9778), .C2(n9745), .A(n9625), .B(n9624), .ZN(
        P1_U3267) );
  XNOR2_X1 U10927 ( .A(n9626), .B(n9635), .ZN(n9783) );
  INV_X1 U10928 ( .A(n9650), .ZN(n9629) );
  INV_X1 U10929 ( .A(n9627), .ZN(n9628) );
  AOI21_X1 U10930 ( .B1(n9779), .B2(n9629), .A(n9628), .ZN(n9780) );
  INV_X1 U10931 ( .A(n9630), .ZN(n9631) );
  AOI22_X1 U10932 ( .A1(n9703), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9631), .B2(
        n9948), .ZN(n9632) );
  OAI21_X1 U10933 ( .B1(n9633), .B2(n9951), .A(n9632), .ZN(n9643) );
  INV_X1 U10934 ( .A(n9634), .ZN(n9637) );
  INV_X1 U10935 ( .A(n9635), .ZN(n9636) );
  AOI21_X1 U10936 ( .B1(n9637), .B2(n9636), .A(n9678), .ZN(n9641) );
  OAI22_X1 U10937 ( .A1(n9665), .A2(n9681), .B1(n9638), .B2(n9683), .ZN(n9639)
         );
  AOI21_X1 U10938 ( .B1(n9641), .B2(n9640), .A(n9639), .ZN(n9782) );
  NOR2_X1 U10939 ( .A1(n9782), .A2(n9703), .ZN(n9642) );
  AOI211_X1 U10940 ( .C1(n9780), .C2(n9743), .A(n9643), .B(n9642), .ZN(n9644)
         );
  OAI21_X1 U10941 ( .B1(n9783), .B2(n9745), .A(n9644), .ZN(P1_U3268) );
  XNOR2_X1 U10942 ( .A(n9645), .B(n9647), .ZN(n9788) );
  XOR2_X1 U10943 ( .A(n9647), .B(n9646), .Z(n9648) );
  OAI222_X1 U10944 ( .A1(n9683), .A2(n9649), .B1(n9681), .B2(n9682), .C1(n9648), .C2(n9678), .ZN(n9784) );
  AOI211_X1 U10945 ( .C1(n9786), .C2(n9666), .A(n10210), .B(n9650), .ZN(n9785)
         );
  NAND2_X1 U10946 ( .A1(n9785), .A2(n9957), .ZN(n9654) );
  INV_X1 U10947 ( .A(n9651), .ZN(n9652) );
  AOI22_X1 U10948 ( .A1(n9703), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9652), .B2(
        n9948), .ZN(n9653) );
  OAI211_X1 U10949 ( .C1(n9655), .C2(n9951), .A(n9654), .B(n9653), .ZN(n9656)
         );
  AOI21_X1 U10950 ( .B1(n9784), .B2(n9728), .A(n9656), .ZN(n9657) );
  OAI21_X1 U10951 ( .B1(n9788), .B2(n9745), .A(n9657), .ZN(P1_U3269) );
  XNOR2_X1 U10952 ( .A(n9659), .B(n9658), .ZN(n9793) );
  AOI22_X1 U10953 ( .A1(n9791), .A2(n9660), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9703), .ZN(n9674) );
  XNOR2_X1 U10954 ( .A(n9662), .B(n9661), .ZN(n9663) );
  OAI222_X1 U10955 ( .A1(n9683), .A2(n9665), .B1(n9681), .B2(n9664), .C1(n9678), .C2(n9663), .ZN(n9789) );
  INV_X1 U10956 ( .A(n9666), .ZN(n9667) );
  AOI211_X1 U10957 ( .C1(n9791), .C2(n9684), .A(n10210), .B(n9667), .ZN(n9790)
         );
  INV_X1 U10958 ( .A(n9790), .ZN(n9671) );
  OAI22_X1 U10959 ( .A1(n9671), .A2(n9670), .B1(n9669), .B2(n9668), .ZN(n9672)
         );
  OAI21_X1 U10960 ( .B1(n9789), .B2(n9672), .A(n9728), .ZN(n9673) );
  OAI211_X1 U10961 ( .C1(n9793), .C2(n9745), .A(n9674), .B(n9673), .ZN(
        P1_U3270) );
  XNOR2_X1 U10962 ( .A(n9675), .B(n9676), .ZN(n9798) );
  XNOR2_X1 U10963 ( .A(n9677), .B(n9676), .ZN(n9679) );
  OAI222_X1 U10964 ( .A1(n9683), .A2(n9682), .B1(n9681), .B2(n9680), .C1(n9679), .C2(n9678), .ZN(n9794) );
  AOI211_X1 U10965 ( .C1(n9796), .C2(n9692), .A(n10210), .B(n4754), .ZN(n9795)
         );
  NAND2_X1 U10966 ( .A1(n9795), .A2(n9957), .ZN(n9687) );
  AOI22_X1 U10967 ( .A1(n9703), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9685), .B2(
        n9948), .ZN(n9686) );
  OAI211_X1 U10968 ( .C1(n9688), .C2(n9951), .A(n9687), .B(n9686), .ZN(n9689)
         );
  AOI21_X1 U10969 ( .B1(n9794), .B2(n9728), .A(n9689), .ZN(n9690) );
  OAI21_X1 U10970 ( .B1(n9798), .B2(n9745), .A(n9690), .ZN(P1_U3271) );
  XNOR2_X1 U10971 ( .A(n9691), .B(n9700), .ZN(n9803) );
  INV_X1 U10972 ( .A(n9708), .ZN(n9694) );
  INV_X1 U10973 ( .A(n9692), .ZN(n9693) );
  AOI211_X1 U10974 ( .C1(n9800), .C2(n9694), .A(n10210), .B(n9693), .ZN(n9799)
         );
  AOI22_X1 U10975 ( .A1(n9703), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9695), .B2(
        n9948), .ZN(n9696) );
  OAI21_X1 U10976 ( .B1(n9697), .B2(n9951), .A(n9696), .ZN(n9705) );
  OAI21_X1 U10977 ( .B1(n9700), .B2(n9699), .A(n9698), .ZN(n9702) );
  AOI222_X1 U10978 ( .A1(n9738), .A2(n9702), .B1(n9736), .B2(n9733), .C1(n9701), .C2(n9735), .ZN(n9802) );
  NOR2_X1 U10979 ( .A1(n9802), .A2(n9703), .ZN(n9704) );
  AOI211_X1 U10980 ( .C1(n9799), .C2(n9957), .A(n9705), .B(n9704), .ZN(n9706)
         );
  OAI21_X1 U10981 ( .B1(n9803), .B2(n9745), .A(n9706), .ZN(P1_U3272) );
  XNOR2_X1 U10982 ( .A(n9707), .B(n9717), .ZN(n9808) );
  AOI21_X1 U10983 ( .B1(n9804), .B2(n4760), .A(n9708), .ZN(n9805) );
  INV_X1 U10984 ( .A(n9709), .ZN(n9710) );
  AOI22_X1 U10985 ( .A1(n9703), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9710), .B2(
        n9948), .ZN(n9711) );
  OAI21_X1 U10986 ( .B1(n9712), .B2(n9951), .A(n9711), .ZN(n9722) );
  INV_X1 U10987 ( .A(n9713), .ZN(n9714) );
  AOI21_X1 U10988 ( .B1(n9731), .B2(n9715), .A(n9714), .ZN(n9716) );
  XOR2_X1 U10989 ( .A(n9717), .B(n9716), .Z(n9720) );
  AOI222_X1 U10990 ( .A1(n9738), .A2(n9720), .B1(n9719), .B2(n9733), .C1(n9718), .C2(n9735), .ZN(n9807) );
  NOR2_X1 U10991 ( .A1(n9807), .A2(n9703), .ZN(n9721) );
  AOI211_X1 U10992 ( .C1(n9805), .C2(n9743), .A(n9722), .B(n9721), .ZN(n9723)
         );
  OAI21_X1 U10993 ( .B1(n9808), .B2(n9745), .A(n9723), .ZN(P1_U3273) );
  XNOR2_X1 U10994 ( .A(n9724), .B(n9732), .ZN(n9813) );
  AND2_X1 U10995 ( .A1(n9725), .A2(n9809), .ZN(n9726) );
  NOR2_X1 U10996 ( .A1(n9727), .A2(n9726), .ZN(n9810) );
  INV_X1 U10997 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9729) );
  OAI22_X1 U10998 ( .A1(n9730), .A2(n9951), .B1(n9729), .B2(n9728), .ZN(n9742)
         );
  XOR2_X1 U10999 ( .A(n9732), .B(n9731), .Z(n9737) );
  AOI222_X1 U11000 ( .A1(n9738), .A2(n9737), .B1(n9736), .B2(n9735), .C1(n9734), .C2(n9733), .ZN(n9812) );
  NAND2_X1 U11001 ( .A1(n9948), .A2(n9739), .ZN(n9740) );
  AOI21_X1 U11002 ( .B1(n9812), .B2(n9740), .A(n9703), .ZN(n9741) );
  AOI211_X1 U11003 ( .C1(n9810), .C2(n9743), .A(n9742), .B(n9741), .ZN(n9744)
         );
  OAI21_X1 U11004 ( .B1(n9813), .B2(n9745), .A(n9744), .ZN(P1_U3274) );
  NAND2_X1 U11005 ( .A1(n9746), .A2(n9964), .ZN(n9747) );
  OAI211_X1 U11006 ( .C1(n9748), .C2(n10210), .A(n9961), .B(n9747), .ZN(n9831)
         );
  MUX2_X1 U11007 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9831), .S(n10236), .Z(
        P1_U3554) );
  AOI22_X1 U11008 ( .A1(n9750), .A2(n10187), .B1(n9964), .B2(n9749), .ZN(n9751) );
  AOI21_X1 U11009 ( .B1(n9964), .B2(n9755), .A(n9754), .ZN(n9756) );
  OAI211_X1 U11010 ( .C1(n9758), .C2(n10192), .A(n9757), .B(n9756), .ZN(n9833)
         );
  MUX2_X1 U11011 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9833), .S(n10236), .Z(
        P1_U3551) );
  AOI22_X1 U11012 ( .A1(n9760), .A2(n10187), .B1(n9964), .B2(n9759), .ZN(n9761) );
  OAI211_X1 U11013 ( .C1(n9763), .C2(n10192), .A(n9762), .B(n9761), .ZN(n9834)
         );
  MUX2_X1 U11014 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9834), .S(n10236), .Z(
        P1_U3550) );
  AOI22_X1 U11015 ( .A1(n9765), .A2(n10187), .B1(n9964), .B2(n9764), .ZN(n9766) );
  OAI211_X1 U11016 ( .C1(n9768), .C2(n10192), .A(n9767), .B(n9766), .ZN(n9835)
         );
  MUX2_X1 U11017 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9835), .S(n10236), .Z(
        P1_U3549) );
  AOI22_X1 U11018 ( .A1(n9770), .A2(n10187), .B1(n9964), .B2(n9769), .ZN(n9771) );
  OAI211_X1 U11019 ( .C1(n9773), .C2(n10192), .A(n9772), .B(n9771), .ZN(n9836)
         );
  MUX2_X1 U11020 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9836), .S(n10236), .Z(
        P1_U3548) );
  AOI211_X1 U11021 ( .C1(n9964), .C2(n9776), .A(n9775), .B(n9774), .ZN(n9777)
         );
  OAI21_X1 U11022 ( .B1(n9778), .B2(n10192), .A(n9777), .ZN(n9837) );
  MUX2_X1 U11023 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9837), .S(n10236), .Z(
        P1_U3547) );
  AOI22_X1 U11024 ( .A1(n9780), .A2(n10187), .B1(n9964), .B2(n9779), .ZN(n9781) );
  OAI211_X1 U11025 ( .C1(n9783), .C2(n10192), .A(n9782), .B(n9781), .ZN(n9838)
         );
  MUX2_X1 U11026 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9838), .S(n10236), .Z(
        P1_U3546) );
  AOI211_X1 U11027 ( .C1(n9964), .C2(n9786), .A(n9785), .B(n9784), .ZN(n9787)
         );
  OAI21_X1 U11028 ( .B1(n9788), .B2(n10192), .A(n9787), .ZN(n9839) );
  MUX2_X1 U11029 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9839), .S(n10236), .Z(
        P1_U3545) );
  AOI211_X1 U11030 ( .C1(n9964), .C2(n9791), .A(n9790), .B(n9789), .ZN(n9792)
         );
  OAI21_X1 U11031 ( .B1(n9793), .B2(n10192), .A(n9792), .ZN(n9840) );
  MUX2_X1 U11032 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9840), .S(n10236), .Z(
        P1_U3544) );
  AOI211_X1 U11033 ( .C1(n9964), .C2(n9796), .A(n9795), .B(n9794), .ZN(n9797)
         );
  OAI21_X1 U11034 ( .B1(n9798), .B2(n10192), .A(n9797), .ZN(n9841) );
  MUX2_X1 U11035 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9841), .S(n10236), .Z(
        P1_U3543) );
  AOI21_X1 U11036 ( .B1(n9964), .B2(n9800), .A(n9799), .ZN(n9801) );
  OAI211_X1 U11037 ( .C1(n9803), .C2(n10192), .A(n9802), .B(n9801), .ZN(n9842)
         );
  MUX2_X1 U11038 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9842), .S(n10236), .Z(
        P1_U3542) );
  AOI22_X1 U11039 ( .A1(n9805), .A2(n10187), .B1(n9964), .B2(n9804), .ZN(n9806) );
  OAI211_X1 U11040 ( .C1(n9808), .C2(n10192), .A(n9807), .B(n9806), .ZN(n9843)
         );
  MUX2_X1 U11041 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9843), .S(n10236), .Z(
        P1_U3541) );
  AOI22_X1 U11042 ( .A1(n9810), .A2(n10187), .B1(n9964), .B2(n9809), .ZN(n9811) );
  OAI211_X1 U11043 ( .C1(n9813), .C2(n10192), .A(n9812), .B(n9811), .ZN(n9844)
         );
  MUX2_X1 U11044 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9844), .S(n10236), .Z(
        P1_U3540) );
  AOI211_X1 U11045 ( .C1(n9964), .C2(n9816), .A(n9815), .B(n9814), .ZN(n9817)
         );
  OAI21_X1 U11046 ( .B1(n9818), .B2(n10192), .A(n9817), .ZN(n9845) );
  MUX2_X1 U11047 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9845), .S(n10236), .Z(
        P1_U3539) );
  INV_X1 U11048 ( .A(n10155), .ZN(n10215) );
  AND2_X1 U11049 ( .A1(n9819), .A2(n10215), .ZN(n9823) );
  OAI22_X1 U11050 ( .A1(n9821), .A2(n10210), .B1(n9820), .B2(n10208), .ZN(
        n9822) );
  MUX2_X1 U11051 ( .A(n9846), .B(P1_REG1_REG_15__SCAN_IN), .S(n10233), .Z(
        P1_U3538) );
  AOI22_X1 U11052 ( .A1(n9826), .A2(n10187), .B1(n9964), .B2(n9825), .ZN(n9827) );
  OAI211_X1 U11053 ( .C1(n10155), .C2(n9829), .A(n9828), .B(n9827), .ZN(n9847)
         );
  MUX2_X1 U11054 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9847), .S(n10236), .Z(
        P1_U3536) );
  MUX2_X1 U11055 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9830), .S(n10236), .Z(
        P1_U3523) );
  MUX2_X1 U11056 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9831), .S(n10218), .Z(
        P1_U3522) );
  MUX2_X1 U11057 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9832), .S(n10218), .Z(
        P1_U3520) );
  MUX2_X1 U11058 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9833), .S(n10218), .Z(
        P1_U3519) );
  MUX2_X1 U11059 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9834), .S(n10218), .Z(
        P1_U3518) );
  MUX2_X1 U11060 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9835), .S(n10218), .Z(
        P1_U3517) );
  MUX2_X1 U11061 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9836), .S(n10218), .Z(
        P1_U3516) );
  MUX2_X1 U11062 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9837), .S(n10218), .Z(
        P1_U3515) );
  MUX2_X1 U11063 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9838), .S(n10218), .Z(
        P1_U3514) );
  MUX2_X1 U11064 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9839), .S(n10218), .Z(
        P1_U3513) );
  MUX2_X1 U11065 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9840), .S(n10218), .Z(
        P1_U3512) );
  MUX2_X1 U11066 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9841), .S(n10218), .Z(
        P1_U3511) );
  MUX2_X1 U11067 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9842), .S(n10218), .Z(
        P1_U3510) );
  MUX2_X1 U11068 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9843), .S(n10218), .Z(
        P1_U3508) );
  MUX2_X1 U11069 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9844), .S(n10218), .Z(
        P1_U3505) );
  MUX2_X1 U11070 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9845), .S(n10218), .Z(
        P1_U3502) );
  MUX2_X1 U11071 ( .A(n9846), .B(P1_REG0_REG_15__SCAN_IN), .S(n10216), .Z(
        P1_U3499) );
  MUX2_X1 U11072 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9847), .S(n10218), .Z(
        P1_U3493) );
  NAND3_X1 U11073 ( .A1(n9849), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9851) );
  OAI22_X1 U11074 ( .A1(n9848), .A2(n9851), .B1(n9850), .B2(n9859), .ZN(n9852)
         );
  AOI21_X1 U11075 ( .B1(n9853), .B2(n4567), .A(n9852), .ZN(n9854) );
  INV_X1 U11076 ( .A(n9854), .ZN(P1_U3322) );
  OAI222_X1 U11077 ( .A1(n9859), .A2(n9858), .B1(n9857), .B2(n9856), .C1(
        P1_U3084), .C2(n9855), .ZN(P1_U3323) );
  MUX2_X1 U11078 ( .A(n9860), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U11079 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9861) );
  OAI22_X1 U11080 ( .A1(n10107), .A2(n9862), .B1(n10116), .B2(n9861), .ZN(
        n9863) );
  INV_X1 U11081 ( .A(n9863), .ZN(n9874) );
  AOI21_X1 U11082 ( .B1(n9866), .B2(n9865), .A(n9864), .ZN(n9867) );
  NAND2_X1 U11083 ( .A1(n10104), .A2(n9867), .ZN(n9872) );
  OAI211_X1 U11084 ( .C1(n9870), .C2(n9869), .A(n10111), .B(n9868), .ZN(n9871)
         );
  NAND4_X1 U11085 ( .A1(n9874), .A2(n9873), .A3(n9872), .A4(n9871), .ZN(
        P1_U3244) );
  AOI22_X1 U11086 ( .A1(n10243), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9886) );
  NAND2_X1 U11087 ( .A1(n4579), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9877) );
  AOI211_X1 U11088 ( .C1(n9877), .C2(n9876), .A(n9875), .B(n9887), .ZN(n9878)
         );
  AOI21_X1 U11089 ( .B1(n9893), .B2(n9879), .A(n9878), .ZN(n9885) );
  NOR2_X1 U11090 ( .A1(n10246), .A2(n9880), .ZN(n9883) );
  OAI211_X1 U11091 ( .C1(n9883), .C2(n9882), .A(n10237), .B(n9881), .ZN(n9884)
         );
  NAND3_X1 U11092 ( .A1(n9886), .A2(n9885), .A3(n9884), .ZN(P2_U3246) );
  AOI22_X1 U11093 ( .A1(n10243), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9899) );
  AOI211_X1 U11094 ( .C1(n9890), .C2(n9889), .A(n9888), .B(n9887), .ZN(n9891)
         );
  AOI21_X1 U11095 ( .B1(n9893), .B2(n9892), .A(n9891), .ZN(n9898) );
  OAI211_X1 U11096 ( .C1(n9896), .C2(n9895), .A(n10237), .B(n9894), .ZN(n9897)
         );
  NAND3_X1 U11097 ( .A1(n9899), .A2(n9898), .A3(n9897), .ZN(P2_U3247) );
  INV_X1 U11098 ( .A(n9900), .ZN(n9905) );
  OAI22_X1 U11099 ( .A1(n9902), .A2(n10210), .B1(n9901), .B2(n10208), .ZN(
        n9904) );
  AOI211_X1 U11100 ( .C1(n10215), .C2(n9905), .A(n9904), .B(n9903), .ZN(n9907)
         );
  INV_X1 U11101 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9906) );
  AOI22_X1 U11102 ( .A1(n10218), .A2(n9907), .B1(n9906), .B2(n10216), .ZN(
        P1_U3484) );
  AOI22_X1 U11103 ( .A1(n10236), .A2(n9907), .B1(n6736), .B2(n10233), .ZN(
        P1_U3533) );
  INV_X1 U11104 ( .A(n9908), .ZN(n9912) );
  AOI21_X1 U11105 ( .B1(n7608), .B2(n9909), .A(n9919), .ZN(n9911) );
  NOR3_X1 U11106 ( .A1(n9912), .A2(n9911), .A3(n9910), .ZN(n9914) );
  NOR2_X1 U11107 ( .A1(n9914), .A2(n9913), .ZN(n9929) );
  INV_X1 U11108 ( .A(n9915), .ZN(n9916) );
  AOI222_X1 U11109 ( .A1(n9917), .A2(n10283), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n10296), .C1(n10282), .C2(n9916), .ZN(n9927) );
  AOI21_X1 U11110 ( .B1(n9919), .B2(n9918), .A(n4561), .ZN(n9920) );
  INV_X1 U11111 ( .A(n9920), .ZN(n9932) );
  INV_X1 U11112 ( .A(n9921), .ZN(n9924) );
  OAI211_X1 U11113 ( .C1(n9930), .C2(n9924), .A(n9923), .B(n9922), .ZN(n9928)
         );
  INV_X1 U11114 ( .A(n9928), .ZN(n9925) );
  AOI22_X1 U11115 ( .A1(n9932), .A2(n10293), .B1(n10292), .B2(n9925), .ZN(
        n9926) );
  OAI211_X1 U11116 ( .C1(n10296), .C2(n9929), .A(n9927), .B(n9926), .ZN(
        P2_U3282) );
  OAI211_X1 U11117 ( .C1(n9930), .C2(n10362), .A(n9929), .B(n9928), .ZN(n9931)
         );
  AOI21_X1 U11118 ( .B1(n9932), .B2(n10368), .A(n9931), .ZN(n9941) );
  AOI22_X1 U11119 ( .A1(n10382), .A2(n9941), .B1(n9933), .B2(n10380), .ZN(
        P2_U3534) );
  OAI211_X1 U11120 ( .C1(n9936), .C2(n10362), .A(n9935), .B(n9934), .ZN(n9937)
         );
  AOI21_X1 U11121 ( .B1(n9938), .B2(n10368), .A(n9937), .ZN(n9943) );
  AOI22_X1 U11122 ( .A1(n10382), .A2(n9943), .B1(n9939), .B2(n10380), .ZN(
        P2_U3533) );
  INV_X1 U11123 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9940) );
  AOI22_X1 U11124 ( .A1(n10371), .A2(n9941), .B1(n9940), .B2(n10370), .ZN(
        P2_U3493) );
  INV_X1 U11125 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9942) );
  AOI22_X1 U11126 ( .A1(n10371), .A2(n9943), .B1(n9942), .B2(n10370), .ZN(
        P2_U3490) );
  INV_X1 U11127 ( .A(n9954), .ZN(n9946) );
  AOI21_X1 U11128 ( .B1(n9946), .B2(n9945), .A(n9944), .ZN(n9960) );
  INV_X1 U11129 ( .A(n9947), .ZN(n9949) );
  AOI22_X1 U11130 ( .A1(n9703), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9949), .B2(
        n9948), .ZN(n9950) );
  OAI21_X1 U11131 ( .B1(n9952), .B2(n9951), .A(n9950), .ZN(n9956) );
  NOR2_X1 U11132 ( .A1(n9954), .A2(n9953), .ZN(n9955) );
  AOI211_X1 U11133 ( .C1(n9958), .C2(n9957), .A(n9956), .B(n9955), .ZN(n9959)
         );
  OAI21_X1 U11134 ( .B1(n9703), .B2(n9960), .A(n9959), .ZN(P1_U3280) );
  INV_X1 U11135 ( .A(n9961), .ZN(n9963) );
  AOI22_X1 U11136 ( .A1(n10236), .A2(n9979), .B1(n8558), .B2(n10233), .ZN(
        P1_U3553) );
  INV_X1 U11137 ( .A(n10192), .ZN(n10199) );
  OAI21_X1 U11138 ( .B1(n9966), .B2(n10208), .A(n9965), .ZN(n9967) );
  AOI211_X1 U11139 ( .C1(n9969), .C2(n10199), .A(n9968), .B(n9967), .ZN(n9981)
         );
  AOI22_X1 U11140 ( .A1(n10236), .A2(n9981), .B1(n9970), .B2(n10233), .ZN(
        P1_U3537) );
  INV_X1 U11141 ( .A(n9971), .ZN(n9977) );
  INV_X1 U11142 ( .A(n9972), .ZN(n9973) );
  OAI22_X1 U11143 ( .A1(n9974), .A2(n10210), .B1(n9973), .B2(n10208), .ZN(
        n9976) );
  AOI211_X1 U11144 ( .C1(n10215), .C2(n9977), .A(n9976), .B(n9975), .ZN(n9982)
         );
  AOI22_X1 U11145 ( .A1(n10236), .A2(n9982), .B1(n6028), .B2(n10233), .ZN(
        P1_U3535) );
  INV_X1 U11146 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9978) );
  AOI22_X1 U11147 ( .A1(n10218), .A2(n9979), .B1(n9978), .B2(n10216), .ZN(
        P1_U3521) );
  AOI22_X1 U11148 ( .A1(n10218), .A2(n9981), .B1(n9980), .B2(n10216), .ZN(
        P1_U3496) );
  AOI22_X1 U11149 ( .A1(n10218), .A2(n9982), .B1(n6032), .B2(n10216), .ZN(
        P1_U3490) );
  XNOR2_X1 U11150 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XOR2_X1 U11151 ( .A(n5101), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  AOI22_X1 U11152 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9983), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n9994) );
  NOR2_X1 U11153 ( .A1(n4491), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9984) );
  OR2_X1 U11154 ( .A1(n9984), .A2(n4481), .ZN(n10001) );
  XNOR2_X1 U11155 ( .A(n10001), .B(n10000), .ZN(n9985) );
  INV_X1 U11156 ( .A(n9988), .ZN(n9989) );
  NAND2_X1 U11157 ( .A1(n9990), .A2(n9989), .ZN(n9993) );
  NAND3_X1 U11158 ( .A1(n10111), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9991), .ZN(
        n9992) );
  NAND3_X1 U11159 ( .A1(n9994), .A2(n9993), .A3(n9992), .ZN(P1_U3241) );
  MUX2_X1 U11160 ( .A(n9997), .B(n9996), .S(n9995), .Z(n9999) );
  NAND2_X1 U11161 ( .A1(n9999), .A2(n9998), .ZN(n10004) );
  NAND2_X1 U11162 ( .A1(n10001), .A2(n10000), .ZN(n10002) );
  AND2_X1 U11163 ( .A1(n10002), .A2(P1_U4006), .ZN(n10003) );
  NAND2_X1 U11164 ( .A1(n10004), .A2(n10003), .ZN(n10030) );
  XOR2_X1 U11165 ( .A(n10006), .B(n10005), .Z(n10008) );
  OAI22_X1 U11166 ( .A1(n10070), .A2(n10008), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10007), .ZN(n10013) );
  AOI211_X1 U11167 ( .C1(n10011), .C2(n10010), .A(n10009), .B(n10086), .ZN(
        n10012) );
  AOI211_X1 U11168 ( .C1(n10093), .C2(n10014), .A(n10013), .B(n10012), .ZN(
        n10015) );
  AND2_X1 U11169 ( .A1(n10030), .A2(n10015), .ZN(n10016) );
  OAI21_X1 U11170 ( .B1(n10116), .B2(n10017), .A(n10016), .ZN(P1_U3243) );
  INV_X1 U11171 ( .A(n10019), .ZN(n10020) );
  AOI21_X1 U11172 ( .B1(n10021), .B2(n4712), .A(n10020), .ZN(n10031) );
  AOI21_X1 U11173 ( .B1(n10024), .B2(n10023), .A(n10022), .ZN(n10026) );
  OAI21_X1 U11174 ( .B1(n10070), .B2(n10026), .A(n10025), .ZN(n10027) );
  AOI21_X1 U11175 ( .B1(n10093), .B2(n10028), .A(n10027), .ZN(n10029) );
  OAI211_X1 U11176 ( .C1(n10031), .C2(n10086), .A(n10030), .B(n10029), .ZN(
        n10032) );
  INV_X1 U11177 ( .A(n10032), .ZN(n10033) );
  OAI21_X1 U11178 ( .B1(n10116), .B2(n10034), .A(n10033), .ZN(P1_U3245) );
  OAI22_X1 U11179 ( .A1(n10107), .A2(n10035), .B1(n10116), .B2(n7016), .ZN(
        n10036) );
  INV_X1 U11180 ( .A(n10036), .ZN(n10047) );
  OAI21_X1 U11181 ( .B1(n10039), .B2(n10038), .A(n10037), .ZN(n10040) );
  NAND2_X1 U11182 ( .A1(n10104), .A2(n10040), .ZN(n10045) );
  OAI211_X1 U11183 ( .C1(n10043), .C2(n10042), .A(n10111), .B(n10041), .ZN(
        n10044) );
  NAND4_X1 U11184 ( .A1(n10047), .A2(n10046), .A3(n10045), .A4(n10044), .ZN(
        P1_U3246) );
  INV_X1 U11185 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10048) );
  OAI22_X1 U11186 ( .A1(n10107), .A2(n10049), .B1(n10116), .B2(n10048), .ZN(
        n10050) );
  INV_X1 U11187 ( .A(n10050), .ZN(n10060) );
  XNOR2_X1 U11188 ( .A(n10052), .B(n10051), .ZN(n10053) );
  NAND2_X1 U11189 ( .A1(n10053), .A2(n10104), .ZN(n10058) );
  OAI211_X1 U11190 ( .C1(n10056), .C2(n10055), .A(n10054), .B(n10111), .ZN(
        n10057) );
  NAND4_X1 U11191 ( .A1(n10060), .A2(n10059), .A3(n10058), .A4(n10057), .ZN(
        P1_U3249) );
  INV_X1 U11192 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10074) );
  AOI211_X1 U11193 ( .C1(n10063), .C2(n10062), .A(n10061), .B(n10086), .ZN(
        n10064) );
  AOI211_X1 U11194 ( .C1(n10093), .C2(n10066), .A(n10065), .B(n10064), .ZN(
        n10073) );
  AOI21_X1 U11195 ( .B1(n10069), .B2(n10068), .A(n10067), .ZN(n10071) );
  OR2_X1 U11196 ( .A1(n10071), .A2(n10070), .ZN(n10072) );
  OAI211_X1 U11197 ( .C1(n10074), .C2(n10116), .A(n10073), .B(n10072), .ZN(
        P1_U3254) );
  INV_X1 U11198 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10085) );
  INV_X1 U11199 ( .A(n10075), .ZN(n10079) );
  AOI211_X1 U11200 ( .C1(n10077), .C2(n8140), .A(n10076), .B(n10086), .ZN(
        n10078) );
  AOI211_X1 U11201 ( .C1(n10093), .C2(n10080), .A(n10079), .B(n10078), .ZN(
        n10084) );
  OAI211_X1 U11202 ( .C1(n10082), .C2(P1_REG1_REG_15__SCAN_IN), .A(n10111), 
        .B(n10081), .ZN(n10083) );
  OAI211_X1 U11203 ( .C1(n10085), .C2(n10116), .A(n10084), .B(n10083), .ZN(
        P1_U3256) );
  AOI211_X1 U11204 ( .C1(n10089), .C2(n10088), .A(n10087), .B(n10086), .ZN(
        n10090) );
  AOI211_X1 U11205 ( .C1(n10093), .C2(n10092), .A(n10091), .B(n10090), .ZN(
        n10098) );
  OAI211_X1 U11206 ( .C1(n10096), .C2(n10095), .A(n10111), .B(n10094), .ZN(
        n10097) );
  OAI211_X1 U11207 ( .C1(n10099), .C2(n10116), .A(n10098), .B(n10097), .ZN(
        P1_U3257) );
  INV_X1 U11208 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10117) );
  AOI21_X1 U11209 ( .B1(n10102), .B2(n10101), .A(n10100), .ZN(n10103) );
  NAND2_X1 U11210 ( .A1(n10104), .A2(n10103), .ZN(n10106) );
  OAI211_X1 U11211 ( .C1(n10108), .C2(n10107), .A(n10106), .B(n10105), .ZN(
        n10109) );
  INV_X1 U11212 ( .A(n10109), .ZN(n10115) );
  OAI211_X1 U11213 ( .C1(n10113), .C2(n10112), .A(n10111), .B(n10110), .ZN(
        n10114) );
  OAI211_X1 U11214 ( .C1(n10117), .C2(n10116), .A(n10115), .B(n10114), .ZN(
        P1_U3258) );
  NOR2_X1 U11215 ( .A1(n10119), .A2(n10118), .ZN(n10144) );
  NOR2_X1 U11216 ( .A1(n10151), .A2(n10120), .ZN(P1_U3292) );
  INV_X1 U11217 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10121) );
  NOR2_X1 U11218 ( .A1(n10151), .A2(n10121), .ZN(P1_U3293) );
  INV_X1 U11219 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10122) );
  NOR2_X1 U11220 ( .A1(n10151), .A2(n10122), .ZN(P1_U3294) );
  INV_X1 U11221 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10123) );
  NOR2_X1 U11222 ( .A1(n10151), .A2(n10123), .ZN(P1_U3295) );
  INV_X1 U11223 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10124) );
  NOR2_X1 U11224 ( .A1(n10151), .A2(n10124), .ZN(P1_U3296) );
  INV_X1 U11225 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10125) );
  NOR2_X1 U11226 ( .A1(n10151), .A2(n10125), .ZN(P1_U3297) );
  INV_X1 U11227 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10126) );
  NOR2_X1 U11228 ( .A1(n10151), .A2(n10126), .ZN(P1_U3298) );
  INV_X1 U11229 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10127) );
  NOR2_X1 U11230 ( .A1(n10151), .A2(n10127), .ZN(P1_U3299) );
  NOR2_X1 U11231 ( .A1(n10151), .A2(n10128), .ZN(P1_U3300) );
  INV_X1 U11232 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10129) );
  NOR2_X1 U11233 ( .A1(n10151), .A2(n10129), .ZN(P1_U3301) );
  INV_X1 U11234 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10130) );
  NOR2_X1 U11235 ( .A1(n10151), .A2(n10130), .ZN(P1_U3302) );
  INV_X1 U11236 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10131) );
  NOR2_X1 U11237 ( .A1(n10144), .A2(n10131), .ZN(P1_U3303) );
  NOR2_X1 U11238 ( .A1(n10144), .A2(n10132), .ZN(P1_U3304) );
  INV_X1 U11239 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10133) );
  NOR2_X1 U11240 ( .A1(n10144), .A2(n10133), .ZN(P1_U3305) );
  INV_X1 U11241 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10134) );
  NOR2_X1 U11242 ( .A1(n10144), .A2(n10134), .ZN(P1_U3306) );
  NOR2_X1 U11243 ( .A1(n10144), .A2(n10135), .ZN(P1_U3307) );
  INV_X1 U11244 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10136) );
  NOR2_X1 U11245 ( .A1(n10144), .A2(n10136), .ZN(P1_U3308) );
  NOR2_X1 U11246 ( .A1(n10144), .A2(n10137), .ZN(P1_U3309) );
  INV_X1 U11247 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10138) );
  NOR2_X1 U11248 ( .A1(n10151), .A2(n10138), .ZN(P1_U3310) );
  INV_X1 U11249 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10139) );
  NOR2_X1 U11250 ( .A1(n10151), .A2(n10139), .ZN(P1_U3311) );
  INV_X1 U11251 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10140) );
  NOR2_X1 U11252 ( .A1(n10144), .A2(n10140), .ZN(P1_U3312) );
  INV_X1 U11253 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10141) );
  NOR2_X1 U11254 ( .A1(n10144), .A2(n10141), .ZN(P1_U3313) );
  INV_X1 U11255 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10142) );
  NOR2_X1 U11256 ( .A1(n10144), .A2(n10142), .ZN(P1_U3314) );
  NOR2_X1 U11257 ( .A1(n10144), .A2(n10143), .ZN(P1_U3315) );
  INV_X1 U11258 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10145) );
  NOR2_X1 U11259 ( .A1(n10151), .A2(n10145), .ZN(P1_U3316) );
  INV_X1 U11260 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10146) );
  NOR2_X1 U11261 ( .A1(n10151), .A2(n10146), .ZN(P1_U3317) );
  INV_X1 U11262 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10147) );
  NOR2_X1 U11263 ( .A1(n10151), .A2(n10147), .ZN(P1_U3318) );
  INV_X1 U11264 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10148) );
  NOR2_X1 U11265 ( .A1(n10151), .A2(n10148), .ZN(P1_U3319) );
  INV_X1 U11266 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10149) );
  NOR2_X1 U11267 ( .A1(n10151), .A2(n10149), .ZN(P1_U3320) );
  INV_X1 U11268 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10150) );
  NOR2_X1 U11269 ( .A1(n10151), .A2(n10150), .ZN(P1_U3321) );
  INV_X1 U11270 ( .A(n10152), .ZN(n10154) );
  OAI211_X1 U11271 ( .C1(n10156), .C2(n10155), .A(n10154), .B(n10153), .ZN(
        n10157) );
  NOR2_X1 U11272 ( .A1(n10158), .A2(n10157), .ZN(n10219) );
  AOI22_X1 U11273 ( .A1(n10218), .A2(n10219), .B1(n5809), .B2(n10216), .ZN(
        P1_U3457) );
  INV_X1 U11274 ( .A(n10159), .ZN(n10164) );
  OAI21_X1 U11275 ( .B1(n10161), .B2(n10208), .A(n10160), .ZN(n10163) );
  AOI211_X1 U11276 ( .C1(n10215), .C2(n10164), .A(n10163), .B(n10162), .ZN(
        n10221) );
  INV_X1 U11277 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U11278 ( .A1(n10218), .A2(n10221), .B1(n10165), .B2(n10216), .ZN(
        P1_U3460) );
  OAI21_X1 U11279 ( .B1(n10167), .B2(n10208), .A(n10166), .ZN(n10169) );
  AOI211_X1 U11280 ( .C1(n10215), .C2(n10170), .A(n10169), .B(n10168), .ZN(
        n10223) );
  INV_X1 U11281 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10171) );
  AOI22_X1 U11282 ( .A1(n10218), .A2(n10223), .B1(n10171), .B2(n10216), .ZN(
        P1_U3463) );
  OAI22_X1 U11283 ( .A1(n10173), .A2(n10210), .B1(n10172), .B2(n10208), .ZN(
        n10175) );
  AOI211_X1 U11284 ( .C1(n10215), .C2(n10176), .A(n10175), .B(n10174), .ZN(
        n10225) );
  AOI22_X1 U11285 ( .A1(n10218), .A2(n10225), .B1(n10177), .B2(n10216), .ZN(
        P1_U3466) );
  INV_X1 U11286 ( .A(n10178), .ZN(n10183) );
  NAND3_X1 U11287 ( .A1(n10180), .A2(n10179), .A3(n10199), .ZN(n10181) );
  AND4_X1 U11288 ( .A1(n10184), .A2(n10183), .A3(n10182), .A4(n10181), .ZN(
        n10226) );
  INV_X1 U11289 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U11290 ( .A1(n10218), .A2(n10226), .B1(n10185), .B2(n10216), .ZN(
        P1_U3469) );
  AOI21_X1 U11291 ( .B1(n10188), .B2(n10187), .A(n10186), .ZN(n10189) );
  OAI211_X1 U11292 ( .C1(n10192), .C2(n10191), .A(n10190), .B(n10189), .ZN(
        n10193) );
  INV_X1 U11293 ( .A(n10193), .ZN(n10228) );
  INV_X1 U11294 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10194) );
  AOI22_X1 U11295 ( .A1(n10218), .A2(n10228), .B1(n10194), .B2(n10216), .ZN(
        P1_U3472) );
  NAND3_X1 U11296 ( .A1(n10197), .A2(n10196), .A3(n10195), .ZN(n10198) );
  AOI21_X1 U11297 ( .B1(n10200), .B2(n10199), .A(n10198), .ZN(n10230) );
  AOI22_X1 U11298 ( .A1(n10218), .A2(n10230), .B1(n5918), .B2(n10216), .ZN(
        P1_U3475) );
  INV_X1 U11299 ( .A(n10201), .ZN(n10206) );
  OAI22_X1 U11300 ( .A1(n10203), .A2(n10210), .B1(n10202), .B2(n10208), .ZN(
        n10205) );
  AOI211_X1 U11301 ( .C1(n10215), .C2(n10206), .A(n10205), .B(n10204), .ZN(
        n10232) );
  AOI22_X1 U11302 ( .A1(n10218), .A2(n10232), .B1(n5942), .B2(n10216), .ZN(
        P1_U3478) );
  INV_X1 U11303 ( .A(n10207), .ZN(n10214) );
  OAI22_X1 U11304 ( .A1(n10211), .A2(n10210), .B1(n10209), .B2(n10208), .ZN(
        n10213) );
  AOI211_X1 U11305 ( .C1(n10215), .C2(n10214), .A(n10213), .B(n10212), .ZN(
        n10235) );
  AOI22_X1 U11306 ( .A1(n10218), .A2(n10235), .B1(n10217), .B2(n10216), .ZN(
        P1_U3481) );
  AOI22_X1 U11307 ( .A1(n10236), .A2(n10219), .B1(n6566), .B2(n10233), .ZN(
        P1_U3524) );
  AOI22_X1 U11308 ( .A1(n10236), .A2(n10221), .B1(n10220), .B2(n10233), .ZN(
        P1_U3525) );
  AOI22_X1 U11309 ( .A1(n10236), .A2(n10223), .B1(n10222), .B2(n10233), .ZN(
        P1_U3526) );
  AOI22_X1 U11310 ( .A1(n10236), .A2(n10225), .B1(n10224), .B2(n10233), .ZN(
        P1_U3527) );
  AOI22_X1 U11311 ( .A1(n10236), .A2(n10226), .B1(n6564), .B2(n10233), .ZN(
        P1_U3528) );
  AOI22_X1 U11312 ( .A1(n10236), .A2(n10228), .B1(n10227), .B2(n10233), .ZN(
        P1_U3529) );
  AOI22_X1 U11313 ( .A1(n10236), .A2(n10230), .B1(n10229), .B2(n10233), .ZN(
        P1_U3530) );
  AOI22_X1 U11314 ( .A1(n10236), .A2(n10232), .B1(n10231), .B2(n10233), .ZN(
        P1_U3531) );
  AOI22_X1 U11315 ( .A1(n10236), .A2(n10235), .B1(n10234), .B2(n10233), .ZN(
        P1_U3532) );
  AOI22_X1 U11316 ( .A1(n10238), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10237), .ZN(n10247) );
  NAND2_X1 U11317 ( .A1(n10238), .A2(n7350), .ZN(n10240) );
  OAI211_X1 U11318 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n10241), .A(n10240), .B(
        n10239), .ZN(n10242) );
  INV_X1 U11319 ( .A(n10242), .ZN(n10245) );
  AOI22_X1 U11320 ( .A1(n10243), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10244) );
  OAI221_X1 U11321 ( .B1(n4579), .B2(n10247), .C1(n10246), .C2(n10245), .A(
        n10244), .ZN(P2_U3245) );
  NOR2_X1 U11322 ( .A1(n10248), .A2(n10261), .ZN(n10249) );
  OR2_X1 U11323 ( .A1(n10250), .A2(n10249), .ZN(n10267) );
  INV_X1 U11324 ( .A(n10267), .ZN(n10340) );
  INV_X1 U11325 ( .A(n10251), .ZN(n10256) );
  OAI21_X1 U11326 ( .B1(n10253), .B2(n10336), .A(n10252), .ZN(n10337) );
  INV_X1 U11327 ( .A(n10337), .ZN(n10254) );
  AOI22_X1 U11328 ( .A1(n10340), .A2(n10256), .B1(n10255), .B2(n10254), .ZN(
        n10274) );
  AOI22_X1 U11329 ( .A1(n10260), .A2(n10259), .B1(n10258), .B2(n10257), .ZN(
        n10265) );
  XNOR2_X1 U11330 ( .A(n10262), .B(n10261), .ZN(n10263) );
  NAND2_X1 U11331 ( .A1(n10263), .A2(n10278), .ZN(n10264) );
  OAI211_X1 U11332 ( .C1(n10267), .C2(n10266), .A(n10265), .B(n10264), .ZN(
        n10338) );
  AOI22_X1 U11333 ( .A1(n10296), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n10268), 
        .B2(n10282), .ZN(n10269) );
  OAI21_X1 U11334 ( .B1(n10336), .B2(n10270), .A(n10269), .ZN(n10271) );
  AOI21_X1 U11335 ( .B1(n10338), .B2(n10272), .A(n10271), .ZN(n10273) );
  NAND2_X1 U11336 ( .A1(n10274), .A2(n10273), .ZN(P2_U3288) );
  XNOR2_X1 U11337 ( .A(n10275), .B(n10287), .ZN(n10279) );
  INV_X1 U11338 ( .A(n10276), .ZN(n10277) );
  AOI21_X1 U11339 ( .B1(n10279), .B2(n10278), .A(n10277), .ZN(n10324) );
  INV_X1 U11340 ( .A(n10280), .ZN(n10281) );
  AOI222_X1 U11341 ( .A1(n10321), .A2(n10283), .B1(P2_REG2_REG_6__SCAN_IN), 
        .B2(n10296), .C1(n10282), .C2(n10281), .ZN(n10295) );
  NAND2_X1 U11342 ( .A1(n10285), .A2(n10284), .ZN(n10286) );
  XOR2_X1 U11343 ( .A(n10287), .B(n10286), .Z(n10327) );
  AOI21_X1 U11344 ( .B1(n10288), .B2(n10321), .A(n10364), .ZN(n10290) );
  NAND2_X1 U11345 ( .A1(n10290), .A2(n10289), .ZN(n10322) );
  INV_X1 U11346 ( .A(n10322), .ZN(n10291) );
  AOI22_X1 U11347 ( .A1(n10327), .A2(n10293), .B1(n10292), .B2(n10291), .ZN(
        n10294) );
  OAI211_X1 U11348 ( .C1(n10296), .C2(n10324), .A(n10295), .B(n10294), .ZN(
        P2_U3290) );
  NOR2_X1 U11349 ( .A1(n10298), .A2(n10297), .ZN(n10307) );
  AND2_X1 U11350 ( .A1(n10310), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3297) );
  AND2_X1 U11351 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10310), .ZN(P2_U3298) );
  AND2_X1 U11352 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10310), .ZN(P2_U3299) );
  NOR2_X1 U11353 ( .A1(n10307), .A2(n10299), .ZN(P2_U3300) );
  AND2_X1 U11354 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10310), .ZN(P2_U3301) );
  AND2_X1 U11355 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10310), .ZN(P2_U3302) );
  AND2_X1 U11356 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10310), .ZN(P2_U3303) );
  AND2_X1 U11357 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10310), .ZN(P2_U3304) );
  AND2_X1 U11358 ( .A1(n10310), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3305) );
  AND2_X1 U11359 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10310), .ZN(P2_U3306) );
  NOR2_X1 U11360 ( .A1(n10307), .A2(n10300), .ZN(P2_U3307) );
  AND2_X1 U11361 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10310), .ZN(P2_U3308) );
  AND2_X1 U11362 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10310), .ZN(P2_U3309) );
  AND2_X1 U11363 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10310), .ZN(P2_U3310) );
  AND2_X1 U11364 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10310), .ZN(P2_U3311) );
  NOR2_X1 U11365 ( .A1(n10307), .A2(n10301), .ZN(P2_U3312) );
  NOR2_X1 U11366 ( .A1(n10307), .A2(n10302), .ZN(P2_U3313) );
  AND2_X1 U11367 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10310), .ZN(P2_U3314) );
  AND2_X1 U11368 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10310), .ZN(P2_U3315) );
  NOR2_X1 U11369 ( .A1(n10307), .A2(n10303), .ZN(P2_U3316) );
  AND2_X1 U11370 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10310), .ZN(P2_U3317) );
  NOR2_X1 U11371 ( .A1(n10307), .A2(n10304), .ZN(P2_U3318) );
  AND2_X1 U11372 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10310), .ZN(P2_U3319) );
  AND2_X1 U11373 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10310), .ZN(P2_U3320) );
  NOR2_X1 U11374 ( .A1(n10307), .A2(n10305), .ZN(P2_U3321) );
  AND2_X1 U11375 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10310), .ZN(P2_U3322) );
  AND2_X1 U11376 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10310), .ZN(P2_U3323) );
  NOR2_X1 U11377 ( .A1(n10307), .A2(n10306), .ZN(P2_U3324) );
  AND2_X1 U11378 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10310), .ZN(P2_U3325) );
  AND2_X1 U11379 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10310), .ZN(P2_U3326) );
  AOI22_X1 U11380 ( .A1(n10313), .A2(n10309), .B1(n10308), .B2(n10310), .ZN(
        P2_U3437) );
  AOI22_X1 U11381 ( .A1(n10313), .A2(n10312), .B1(n10311), .B2(n10310), .ZN(
        P2_U3438) );
  INV_X1 U11382 ( .A(n10314), .ZN(n10316) );
  OAI22_X1 U11383 ( .A1(n10316), .A2(n10364), .B1(n10315), .B2(n10362), .ZN(
        n10317) );
  AOI211_X1 U11384 ( .C1(n10368), .C2(n10319), .A(n10318), .B(n10317), .ZN(
        n10372) );
  INV_X1 U11385 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U11386 ( .A1(n10371), .A2(n10372), .B1(n10320), .B2(n10370), .ZN(
        P2_U3463) );
  INV_X1 U11387 ( .A(n10321), .ZN(n10323) );
  OAI21_X1 U11388 ( .B1(n10323), .B2(n10362), .A(n10322), .ZN(n10326) );
  INV_X1 U11389 ( .A(n10324), .ZN(n10325) );
  AOI211_X1 U11390 ( .C1(n10327), .C2(n10368), .A(n10326), .B(n10325), .ZN(
        n10373) );
  INV_X1 U11391 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10328) );
  AOI22_X1 U11392 ( .A1(n10371), .A2(n10373), .B1(n10328), .B2(n10370), .ZN(
        P2_U3469) );
  OAI211_X1 U11393 ( .C1(n10331), .C2(n10362), .A(n10330), .B(n10329), .ZN(
        n10332) );
  AOI21_X1 U11394 ( .B1(n10368), .B2(n10333), .A(n10332), .ZN(n10374) );
  INV_X1 U11395 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U11396 ( .A1(n10371), .A2(n10374), .B1(n10334), .B2(n10370), .ZN(
        P2_U3472) );
  INV_X1 U11397 ( .A(n10335), .ZN(n10353) );
  OAI22_X1 U11398 ( .A1(n10337), .A2(n10364), .B1(n10336), .B2(n10362), .ZN(
        n10339) );
  AOI211_X1 U11399 ( .C1(n10353), .C2(n10340), .A(n10339), .B(n10338), .ZN(
        n10375) );
  AOI22_X1 U11400 ( .A1(n10371), .A2(n10375), .B1(n5321), .B2(n10370), .ZN(
        P2_U3475) );
  OAI22_X1 U11401 ( .A1(n10342), .A2(n10364), .B1(n10341), .B2(n10362), .ZN(
        n10344) );
  AOI211_X1 U11402 ( .C1(n10353), .C2(n10345), .A(n10344), .B(n10343), .ZN(
        n10377) );
  INV_X1 U11403 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U11404 ( .A1(n10371), .A2(n10377), .B1(n10346), .B2(n10370), .ZN(
        P2_U3478) );
  INV_X1 U11405 ( .A(n10347), .ZN(n10352) );
  OAI22_X1 U11406 ( .A1(n10349), .A2(n10364), .B1(n10348), .B2(n10362), .ZN(
        n10351) );
  AOI211_X1 U11407 ( .C1(n10353), .C2(n10352), .A(n10351), .B(n10350), .ZN(
        n10378) );
  INV_X1 U11408 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10354) );
  AOI22_X1 U11409 ( .A1(n10371), .A2(n10378), .B1(n10354), .B2(n10370), .ZN(
        P2_U3481) );
  OAI21_X1 U11410 ( .B1(n10356), .B2(n10362), .A(n10355), .ZN(n10357) );
  AOI211_X1 U11411 ( .C1(n10359), .C2(n10368), .A(n10358), .B(n10357), .ZN(
        n10379) );
  INV_X1 U11412 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10360) );
  AOI22_X1 U11413 ( .A1(n10371), .A2(n10379), .B1(n10360), .B2(n10370), .ZN(
        P2_U3484) );
  INV_X1 U11414 ( .A(n10361), .ZN(n10369) );
  OAI22_X1 U11415 ( .A1(n10365), .A2(n10364), .B1(n10363), .B2(n10362), .ZN(
        n10366) );
  AOI211_X1 U11416 ( .C1(n10369), .C2(n10368), .A(n10367), .B(n10366), .ZN(
        n10381) );
  AOI22_X1 U11417 ( .A1(n10371), .A2(n10381), .B1(n5274), .B2(n10370), .ZN(
        P2_U3487) );
  AOI22_X1 U11418 ( .A1(n10382), .A2(n10372), .B1(n5384), .B2(n10380), .ZN(
        P2_U3524) );
  AOI22_X1 U11419 ( .A1(n10382), .A2(n10373), .B1(n7148), .B2(n10380), .ZN(
        P2_U3526) );
  AOI22_X1 U11420 ( .A1(n10382), .A2(n10374), .B1(n7173), .B2(n10380), .ZN(
        P2_U3527) );
  AOI22_X1 U11421 ( .A1(n10382), .A2(n10375), .B1(n7334), .B2(n10380), .ZN(
        P2_U3528) );
  AOI22_X1 U11422 ( .A1(n10382), .A2(n10377), .B1(n10376), .B2(n10380), .ZN(
        P2_U3529) );
  AOI22_X1 U11423 ( .A1(n10382), .A2(n10378), .B1(n7336), .B2(n10380), .ZN(
        P2_U3530) );
  AOI22_X1 U11424 ( .A1(n10382), .A2(n10379), .B1(n7763), .B2(n10380), .ZN(
        P2_U3531) );
  AOI22_X1 U11425 ( .A1(n10382), .A2(n10381), .B1(n7767), .B2(n10380), .ZN(
        P2_U3532) );
  NOR2_X1 U11426 ( .A1(n10384), .A2(n10383), .ZN(n10385) );
  XOR2_X1 U11427 ( .A(n10385), .B(P2_ADDR_REG_1__SCAN_IN), .Z(ADD_1071_U5) );
  XOR2_X1 U11428 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11429 ( .B1(n10388), .B2(n10387), .A(n10386), .ZN(ADD_1071_U56) );
  OAI21_X1 U11430 ( .B1(n10391), .B2(n10390), .A(n10389), .ZN(ADD_1071_U57) );
  OAI21_X1 U11431 ( .B1(n10394), .B2(n10393), .A(n10392), .ZN(ADD_1071_U58) );
  OAI21_X1 U11432 ( .B1(n10397), .B2(n10396), .A(n10395), .ZN(ADD_1071_U59) );
  OAI21_X1 U11433 ( .B1(n10400), .B2(n10399), .A(n10398), .ZN(ADD_1071_U60) );
  OAI21_X1 U11434 ( .B1(n10403), .B2(n10402), .A(n10401), .ZN(ADD_1071_U61) );
  AOI21_X1 U11435 ( .B1(n10406), .B2(n10405), .A(n10404), .ZN(ADD_1071_U62) );
  AOI21_X1 U11436 ( .B1(n10409), .B2(n10408), .A(n10407), .ZN(ADD_1071_U63) );
  XOR2_X1 U11437 ( .A(n10410), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  XOR2_X1 U11438 ( .A(n10412), .B(n10411), .Z(ADD_1071_U54) );
  NOR2_X1 U11439 ( .A1(n10414), .A2(n10413), .ZN(n10415) );
  XOR2_X1 U11440 ( .A(n10415), .B(P1_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  OAI21_X1 U11441 ( .B1(n10418), .B2(n10417), .A(n10416), .ZN(n10419) );
  XNOR2_X1 U11442 ( .A(n10419), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11443 ( .B1(n10422), .B2(n10421), .A(n10420), .ZN(ADD_1071_U47) );
  AOI21_X1 U11444 ( .B1(n10425), .B2(n10424), .A(n10423), .ZN(ADD_1071_U48) );
  XOR2_X1 U11445 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10426), .Z(ADD_1071_U49) );
  XOR2_X1 U11446 ( .A(n10428), .B(n10427), .Z(ADD_1071_U53) );
  XNOR2_X1 U11447 ( .A(n10430), .B(n10429), .ZN(ADD_1071_U52) );
  XNOR2_X1 U5019 ( .A(n5092), .B(n5091), .ZN(n8231) );
  INV_X1 U5052 ( .A(n7263), .ZN(n7511) );
  BUF_X2 U5050 ( .A(n5880), .Z(n4482) );
  NAND2_X2 U5040 ( .A1(n6672), .A2(n7263), .ZN(n8358) );
  CLKBUF_X2 U5048 ( .A(n6398), .Z(n8329) );
  CLKBUF_X2 U8056 ( .A(n5923), .Z(n6514) );
endmodule

