

module b14_C_SARLock_k_128_7 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2170, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938;

  CLKBUF_X2 U2413 ( .A(n2925), .Z(n3659) );
  INV_X1 U2414 ( .A(n2923), .ZN(n3665) );
  AND2_X1 U2415 ( .A1(n2653), .A2(n2722), .ZN(n4413) );
  CLKBUF_X2 U2416 ( .A(n2465), .Z(n3906) );
  NAND2_X1 U2417 ( .A1(n2818), .A2(n2430), .ZN(n2732) );
  INV_X1 U2418 ( .A(n2922), .ZN(n3145) );
  INV_X1 U2419 ( .A(n2925), .ZN(n3679) );
  INV_X1 U2420 ( .A(n4408), .ZN(n2435) );
  NOR2_X1 U2421 ( .A1(n3086), .A2(n3016), .ZN(n3109) );
  NAND2_X1 U2422 ( .A1(n2722), .A2(IR_REG_31__SCAN_IN), .ZN(n2223) );
  NAND4_X1 U2423 ( .A1(n2488), .A2(n2487), .A3(n2486), .A4(n2485), .ZN(n4010)
         );
  INV_X2 U2424 ( .A(n4245), .ZN(n4557) );
  OAI21_X2 U2425 ( .B1(n3774), .B2(n2229), .A(n2179), .ZN(n3699) );
  NAND2_X2 U2426 ( .A1(n3725), .A2(n3776), .ZN(n3774) );
  NOR2_X2 U2427 ( .A1(n3315), .A2(n3311), .ZN(n3363) );
  NAND3_X2 U2428 ( .A1(n2294), .A2(n2293), .A3(n2290), .ZN(n4408) );
  AOI21_X2 U2429 ( .B1(n4205), .B2(n2677), .A(n2676), .ZN(n4191) );
  NAND2_X2 U2430 ( .A1(n4329), .A2(n2669), .ZN(n4205) );
  NAND2_X1 U2431 ( .A1(n2916), .A2(n2915), .ZN(n2170) );
  OAI21_X2 U2432 ( .B1(n2732), .B2(n2431), .A(IR_REG_29__SCAN_IN), .ZN(n2358)
         );
  AND2_X4 U2433 ( .A1(n2936), .A2(n2730), .ZN(n4361) );
  AND2_X2 U2434 ( .A1(n2903), .A2(n2774), .ZN(n2936) );
  INV_X1 U2435 ( .A(n3676), .ZN(n2173) );
  INV_X1 U2436 ( .A(n4011), .ZN(n4539) );
  INV_X1 U2437 ( .A(n4012), .ZN(n2917) );
  NAND4_X1 U2438 ( .A1(n2464), .A2(n2463), .A3(n2462), .A4(n2461), .ZN(n4013)
         );
  AND4_X1 U2439 ( .A1(n2455), .A2(n2454), .A3(n2453), .A4(n2452), .ZN(n2950)
         );
  INV_X1 U2440 ( .A(n2443), .ZN(n2468) );
  AND2_X2 U2441 ( .A1(n2435), .A2(n2434), .ZN(n2460) );
  NAND2_X1 U2442 ( .A1(n3653), .A2(n3647), .ZN(n3766) );
  INV_X1 U2443 ( .A(n2322), .ZN(n4241) );
  OR2_X1 U2444 ( .A1(n2218), .A2(n2217), .ZN(n2215) );
  NAND2_X1 U2445 ( .A1(n2325), .A2(n2411), .ZN(n4249) );
  AOI22_X1 U2446 ( .A1(n3582), .A2(n2198), .B1(n2216), .B2(n2220), .ZN(n2214)
         );
  NAND2_X1 U2447 ( .A1(n3525), .A2(n2641), .ZN(n3550) );
  OAI21_X1 U2448 ( .B1(n2809), .B2(n3685), .A(n2808), .ZN(n4126) );
  AOI21_X1 U2449 ( .B1(n3380), .B2(n2607), .A(n2412), .ZN(n3419) );
  OAI21_X1 U2450 ( .B1(n3226), .B2(n3225), .A(n3224), .ZN(n3259) );
  NAND2_X1 U2451 ( .A1(n2578), .A2(n2577), .ZN(n3305) );
  OAI22_X1 U2452 ( .A1(n3197), .A2(n3196), .B1(n3195), .B2(n3194), .ZN(n3226)
         );
  AOI21_X1 U2453 ( .B1(n3159), .B2(n3158), .A(n3157), .ZN(n3160) );
  OAI21_X2 U2454 ( .B1(n3080), .B2(n3079), .A(n2233), .ZN(n3081) );
  NAND2_X1 U2455 ( .A1(n2235), .A2(n2404), .ZN(n2234) );
  NOR2_X1 U2456 ( .A1(n3127), .A2(n2402), .ZN(n2401) );
  AND2_X1 U2457 ( .A1(n3082), .A2(n2403), .ZN(n2402) );
  NOR2_X1 U2458 ( .A1(n2982), .A2(n3114), .ZN(n3020) );
  NAND2_X1 U2459 ( .A1(n2447), .A2(n2446), .ZN(n4012) );
  AND2_X1 U2460 ( .A1(n2494), .A2(n2493), .ZN(n3149) );
  CLKBUF_X3 U2461 ( .A(n2468), .Z(n2670) );
  INV_X2 U2462 ( .A(n2642), .ZN(n2484) );
  INV_X1 U2463 ( .A(n4413), .ZN(n4099) );
  CLKBUF_X2 U2464 ( .A(n2458), .Z(n2642) );
  NAND2_X1 U2465 ( .A1(n2435), .A2(n2844), .ZN(n2458) );
  MUX2_X1 U2466 ( .A(n2211), .B(n2249), .S(n2465), .Z(n3055) );
  NAND2_X1 U2469 ( .A1(n2650), .A2(IR_REG_31__SCAN_IN), .ZN(n2725) );
  XNOR2_X1 U2470 ( .A(n2781), .B(IR_REG_25__SCAN_IN), .ZN(n2848) );
  INV_X1 U2471 ( .A(n2628), .ZN(n2244) );
  NAND2_X1 U2472 ( .A1(n2777), .A2(IR_REG_31__SCAN_IN), .ZN(n2792) );
  XNOR2_X1 U2473 ( .A(n2448), .B(IR_REG_2__SCAN_IN), .ZN(n4420) );
  AND2_X1 U2474 ( .A1(n2367), .A2(n2194), .ZN(n2366) );
  AND2_X1 U2475 ( .A1(n2298), .A2(n2361), .ZN(n2176) );
  INV_X1 U2476 ( .A(n2213), .ZN(n2475) );
  AND2_X1 U2477 ( .A1(n2427), .A2(n2428), .ZN(n2367) );
  AND4_X1 U2478 ( .A1(n2248), .A2(n2247), .A3(n2246), .A4(n2245), .ZN(n2427)
         );
  AND3_X1 U2479 ( .A1(n2477), .A2(n2420), .A3(n2474), .ZN(n2421) );
  NOR2_X1 U2480 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2422)
         );
  NOR2_X1 U2481 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2423)
         );
  NOR2_X1 U2482 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2424)
         );
  NOR2_X1 U2483 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2425)
         );
  NOR2_X1 U2484 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2245)
         );
  NOR2_X1 U2485 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2246)
         );
  NOR2_X1 U2486 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2247)
         );
  NOR2_X1 U2487 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .ZN(n2248)
         );
  INV_X1 U2488 ( .A(IR_REG_23__SCAN_IN), .ZN(n2791) );
  INV_X1 U2489 ( .A(IR_REG_24__SCAN_IN), .ZN(n2778) );
  INV_X1 U2490 ( .A(IR_REG_25__SCAN_IN), .ZN(n4795) );
  OAI221_X1 U2491 ( .B1(n2469), .B2(keyinput122), .C1(n2211), .C2(keyinput48), 
        .A(n4901), .ZN(n4910) );
  INV_X2 U2492 ( .A(IR_REG_0__SCAN_IN), .ZN(n2211) );
  AOI21_X2 U2493 ( .B1(n3516), .B2(n2632), .A(n2631), .ZN(n3526) );
  NAND2_X1 U2494 ( .A1(n2917), .A2(n4552), .ZN(n2738) );
  INV_X2 U2495 ( .A(n2950), .ZN(n2456) );
  NOR2_X4 U2496 ( .A1(n4361), .A2(n2170), .ZN(n2925) );
  NAND2_X1 U2497 ( .A1(n2435), .A2(n2844), .ZN(n2172) );
  OAI22_X2 U2498 ( .A1(n3305), .A2(n2590), .B1(n3503), .B2(n3433), .ZN(n3359)
         );
  XNOR2_X2 U2499 ( .A(n2223), .B(n2723), .ZN(n2730) );
  OAI21_X2 U2500 ( .B1(n3359), .B2(n3925), .A(n2598), .ZN(n3380) );
  NAND2_X2 U2501 ( .A1(n2730), .A2(n2735), .ZN(n2916) );
  AND2_X4 U2502 ( .A1(n2434), .A2(n4408), .ZN(n2459) );
  AND2_X1 U2503 ( .A1(n2435), .A2(n2434), .ZN(n2174) );
  NAND2_X1 U2504 ( .A1(n2818), .A2(n2731), .ZN(n2438) );
  OAI21_X1 U2505 ( .B1(n2180), .B2(n2196), .A(n2356), .ZN(n2355) );
  NAND2_X1 U2506 ( .A1(n3612), .A2(n2221), .ZN(n2220) );
  INV_X1 U2507 ( .A(n2383), .ZN(n2221) );
  NAND2_X1 U2508 ( .A1(n2388), .A2(n3722), .ZN(n2387) );
  AND2_X1 U2509 ( .A1(n2698), .A2(REG3_REG_26__SCAN_IN), .ZN(n2704) );
  AND2_X1 U2510 ( .A1(n2704), .A2(REG3_REG_27__SCAN_IN), .ZN(n2712) );
  NOR2_X1 U2511 ( .A1(n2344), .A2(n2341), .ZN(n2340) );
  INV_X1 U2512 ( .A(n2351), .ZN(n2341) );
  INV_X1 U2513 ( .A(n2345), .ZN(n2344) );
  NAND2_X1 U2514 ( .A1(n3489), .A2(n3488), .ZN(n2240) );
  NAND2_X1 U2515 ( .A1(n2379), .A2(n2377), .ZN(n2376) );
  NAND2_X1 U2516 ( .A1(n2378), .A2(n2382), .ZN(n2377) );
  NAND2_X1 U2517 ( .A1(n2380), .A2(n2413), .ZN(n2379) );
  NAND2_X1 U2518 ( .A1(n2382), .A2(n3689), .ZN(n2380) );
  INV_X1 U2519 ( .A(n3054), .ZN(n3049) );
  INV_X1 U2520 ( .A(n2224), .ZN(n3653) );
  AOI21_X1 U2521 ( .B1(n3774), .B2(n2179), .A(n2225), .ZN(n2224) );
  NAND2_X1 U2522 ( .A1(n2226), .A2(n3651), .ZN(n2225) );
  NAND2_X1 U2523 ( .A1(n2321), .A2(n2320), .ZN(n2319) );
  INV_X1 U2524 ( .A(n2885), .ZN(n2320) );
  NAND2_X1 U2525 ( .A1(n4441), .A2(n4442), .ZN(n4440) );
  NAND2_X1 U2526 ( .A1(n4453), .A2(n4454), .ZN(n4452) );
  NOR2_X1 U2527 ( .A1(n4306), .A2(n4147), .ZN(n2710) );
  INV_X1 U2528 ( .A(n4001), .ZN(n3503) );
  AND2_X1 U2529 ( .A1(n2915), .A2(n4560), .ZN(n2951) );
  OAI21_X1 U2530 ( .B1(n2176), .B2(n2295), .A(n2292), .ZN(n2291) );
  NAND2_X1 U2531 ( .A1(n2553), .A2(IR_REG_30__SCAN_IN), .ZN(n2292) );
  NAND2_X1 U2532 ( .A1(n2268), .A2(n2267), .ZN(n2266) );
  INV_X1 U2533 ( .A(n2416), .ZN(n2268) );
  NOR2_X1 U2534 ( .A1(n4113), .A2(n4599), .ZN(n2267) );
  NAND2_X1 U2535 ( .A1(n2220), .A2(n3820), .ZN(n2217) );
  INV_X1 U2536 ( .A(n3743), .ZN(n2218) );
  NAND2_X1 U2537 ( .A1(n3612), .A2(n2384), .ZN(n2216) );
  NOR2_X1 U2538 ( .A1(n3930), .A2(n2346), .ZN(n2345) );
  INV_X1 U2539 ( .A(n2555), .ZN(n2346) );
  NOR2_X1 U2540 ( .A1(n2352), .A2(n2546), .ZN(n2351) );
  INV_X1 U2541 ( .A(n2531), .ZN(n2352) );
  NAND2_X1 U2542 ( .A1(n2299), .A2(n2187), .ZN(n2742) );
  INV_X1 U2543 ( .A(n2738), .ZN(n2288) );
  AND2_X1 U2544 ( .A1(n3844), .A2(n4543), .ZN(n2284) );
  NAND2_X1 U2545 ( .A1(n4539), .A2(n3042), .ZN(n3847) );
  NAND2_X1 U2546 ( .A1(n2296), .A2(IR_REG_31__SCAN_IN), .ZN(n2295) );
  AND2_X1 U2547 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .ZN(n2431)
         );
  NAND2_X1 U2548 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2430) );
  AND3_X1 U2549 ( .A1(n2624), .A2(n2623), .A3(n4853), .ZN(n2625) );
  INV_X1 U2550 ( .A(IR_REG_15__SCAN_IN), .ZN(n2623) );
  INV_X1 U2551 ( .A(IR_REG_11__SCAN_IN), .ZN(n4855) );
  NAND2_X1 U2552 ( .A1(n2388), .A2(n2228), .ZN(n2227) );
  AND2_X1 U2553 ( .A1(n2608), .A2(n2417), .ZN(n2619) );
  OAI21_X1 U2554 ( .B1(n2963), .B2(n3679), .A(n2919), .ZN(n2971) );
  NAND2_X1 U2555 ( .A1(n3391), .A2(n2399), .ZN(n2398) );
  INV_X1 U2556 ( .A(n3388), .ZN(n2399) );
  NOR2_X1 U2557 ( .A1(n2393), .A2(n2238), .ZN(n2237) );
  INV_X1 U2558 ( .A(n2394), .ZN(n2393) );
  INV_X1 U2559 ( .A(n2408), .ZN(n2238) );
  NOR2_X1 U2560 ( .A1(n2395), .A2(n3428), .ZN(n2394) );
  INV_X1 U2561 ( .A(n2397), .ZN(n2395) );
  OR2_X1 U2562 ( .A1(n2580), .A2(n2579), .ZN(n2591) );
  AOI21_X1 U2563 ( .B1(n2456), .B2(n3659), .A(n2926), .ZN(n2927) );
  AND2_X1 U2564 ( .A1(n3604), .A2(n3603), .ZN(n3796) );
  NAND2_X1 U2565 ( .A1(n3081), .A2(n2178), .ZN(n2232) );
  INV_X1 U2566 ( .A(n2401), .ZN(n2235) );
  OR2_X1 U2567 ( .A1(n2712), .A2(n2705), .ZN(n3691) );
  OR2_X1 U2568 ( .A1(n2704), .A2(n2699), .ZN(n3813) );
  AND2_X1 U2569 ( .A1(n2174), .A2(REG0_REG_2__SCAN_IN), .ZN(n2415) );
  NAND2_X1 U2570 ( .A1(n2212), .A2(n2211), .ZN(n2213) );
  INV_X1 U2571 ( .A(IR_REG_1__SCAN_IN), .ZN(n2212) );
  NOR2_X1 U2572 ( .A1(n4022), .A2(n2186), .ZN(n2882) );
  OAI21_X1 U2573 ( .B1(n4030), .B2(n2892), .A(n2894), .ZN(n2895) );
  NOR2_X1 U2574 ( .A1(n3026), .A2(n2261), .ZN(n2260) );
  NAND2_X1 U2575 ( .A1(n3024), .A2(n2258), .ZN(n2257) );
  INV_X1 U2576 ( .A(n3026), .ZN(n2258) );
  NOR2_X1 U2577 ( .A1(n2210), .A2(n3020), .ZN(n3443) );
  NAND2_X1 U2578 ( .A1(n4440), .A2(n3446), .ZN(n3447) );
  XNOR2_X1 U2579 ( .A(n3469), .B(n2265), .ZN(n4046) );
  NAND2_X1 U2580 ( .A1(n4452), .A2(n3449), .ZN(n3450) );
  NAND2_X1 U2581 ( .A1(n4465), .A2(REG2_REG_12__SCAN_IN), .ZN(n4463) );
  NAND2_X1 U2582 ( .A1(n3455), .A2(n3454), .ZN(n4058) );
  XNOR2_X1 U2583 ( .A(n2315), .B(n4066), .ZN(n4060) );
  NAND2_X1 U2584 ( .A1(n4058), .A2(n2316), .ZN(n2315) );
  NAND2_X1 U2585 ( .A1(n4414), .A2(REG1_REG_13__SCAN_IN), .ZN(n2316) );
  NAND2_X1 U2586 ( .A1(n4060), .A2(REG1_REG_14__SCAN_IN), .ZN(n4068) );
  NOR2_X1 U2587 ( .A1(n4473), .A2(n2208), .ZN(n4082) );
  NAND2_X1 U2588 ( .A1(n4478), .A2(n4070), .ZN(n4071) );
  NAND2_X1 U2589 ( .A1(n2244), .A2(n2243), .ZN(n2650) );
  AND2_X1 U2590 ( .A1(n2629), .A2(n2639), .ZN(n2243) );
  INV_X1 U2591 ( .A(IR_REG_18__SCAN_IN), .ZN(n2639) );
  NOR2_X1 U2592 ( .A1(n2697), .A2(n2686), .ZN(n2357) );
  NOR2_X1 U2593 ( .A1(n4316), .A2(n2696), .ZN(n2697) );
  OR2_X1 U2594 ( .A1(n4175), .A2(n4198), .ZN(n2685) );
  OAI21_X1 U2595 ( .B1(n4249), .B2(n2324), .A(n2323), .ZN(n2322) );
  AND2_X1 U2596 ( .A1(n4226), .A2(n4332), .ZN(n2324) );
  NAND2_X1 U2597 ( .A1(n4271), .A2(n4253), .ZN(n2323) );
  NOR2_X1 U2598 ( .A1(n2656), .A2(n4875), .ZN(n2657) );
  NAND2_X1 U2599 ( .A1(n2619), .A2(REG3_REG_17__SCAN_IN), .ZN(n2646) );
  AOI21_X1 U2600 ( .B1(n2276), .B2(n3925), .A(n2275), .ZN(n2274) );
  INV_X1 U2601 ( .A(n3879), .ZN(n2275) );
  NAND2_X1 U2602 ( .A1(n2278), .A2(n3883), .ZN(n3958) );
  NAND2_X1 U2603 ( .A1(n3292), .A2(n2746), .ZN(n2278) );
  AND2_X1 U2604 ( .A1(n3281), .A2(n3283), .ZN(n3930) );
  INV_X1 U2605 ( .A(n4008), .ZN(n3166) );
  INV_X1 U2606 ( .A(n4215), .ZN(n4548) );
  INV_X1 U2607 ( .A(n2735), .ZN(n2903) );
  NOR2_X2 U2608 ( .A1(n4143), .A2(n4127), .ZN(n2824) );
  OAI21_X1 U2609 ( .B1(n2465), .B2(n2450), .A(n2449), .ZN(n4552) );
  NAND2_X1 U2610 ( .A1(n2465), .A2(DATAI_2_), .ZN(n2449) );
  AND2_X1 U2611 ( .A1(n2785), .A2(n2789), .ZN(n2846) );
  INV_X1 U2612 ( .A(n2295), .ZN(n2289) );
  AND2_X1 U2613 ( .A1(n2190), .A2(n2428), .ZN(n2406) );
  NAND2_X1 U2614 ( .A1(n2242), .A2(n3490), .ZN(n2241) );
  NAND2_X1 U2615 ( .A1(n2240), .A2(n3491), .ZN(n2239) );
  NOR2_X1 U2616 ( .A1(n2374), .A2(n3834), .ZN(n2372) );
  AND2_X1 U2617 ( .A1(n2376), .A2(n2201), .ZN(n2374) );
  NAND2_X1 U2618 ( .A1(n2376), .A2(n2381), .ZN(n2375) );
  OR2_X1 U2619 ( .A1(n2382), .A2(n3689), .ZN(n2381) );
  OAI21_X2 U2620 ( .B1(n3736), .B2(n2195), .A(n2230), .ZN(n3690) );
  INV_X1 U2621 ( .A(n2231), .ZN(n2230) );
  OAI21_X1 U2622 ( .B1(n2195), .B2(n3734), .A(n3808), .ZN(n2231) );
  INV_X1 U2623 ( .A(n4213), .ZN(n4175) );
  AND2_X1 U2624 ( .A1(n2954), .A2(n4615), .ZN(n3824) );
  INV_X1 U2625 ( .A(n4319), .ZN(n4231) );
  INV_X1 U2626 ( .A(n3799), .ZN(n4356) );
  NAND4_X1 U2627 ( .A1(n2552), .A2(n2551), .A3(n2550), .A4(n2549), .ZN(n4004)
         );
  NAND2_X1 U2628 ( .A1(n4037), .A2(n2884), .ZN(n2321) );
  INV_X1 U2629 ( .A(n2319), .ZN(n2981) );
  NOR2_X1 U2630 ( .A1(n4502), .A2(n2209), .ZN(n4090) );
  INV_X1 U2631 ( .A(n4128), .ZN(n4306) );
  INV_X1 U2632 ( .A(n2333), .ZN(n2332) );
  INV_X2 U2633 ( .A(n4610), .ZN(n4612) );
  NAND2_X1 U2634 ( .A1(n2270), .A2(n2269), .ZN(n2416) );
  INV_X1 U2635 ( .A(n2822), .ZN(n2269) );
  INV_X1 U2636 ( .A(n4121), .ZN(n2270) );
  INV_X1 U2637 ( .A(n2433), .ZN(n2298) );
  INV_X1 U2638 ( .A(n3611), .ZN(n3612) );
  NAND2_X1 U2639 ( .A1(n2467), .A2(n4543), .ZN(n2362) );
  INV_X1 U2640 ( .A(IR_REG_14__SCAN_IN), .ZN(n2624) );
  OR2_X1 U2641 ( .A1(n2818), .A2(n2432), .ZN(n2439) );
  NAND2_X1 U2642 ( .A1(n2179), .A2(n2229), .ZN(n2226) );
  INV_X1 U2643 ( .A(IR_REG_17__SCAN_IN), .ZN(n2629) );
  INV_X1 U2644 ( .A(n3948), .ZN(n2356) );
  AND2_X1 U2645 ( .A1(n4209), .A2(n4207), .ZN(n3967) );
  OR2_X1 U2646 ( .A1(n3996), .A2(n4228), .ZN(n4209) );
  AND2_X1 U2647 ( .A1(n4208), .A2(n4207), .ZN(n4224) );
  AND2_X1 U2648 ( .A1(n4265), .A2(n2753), .ZN(n3960) );
  NOR2_X1 U2649 ( .A1(n2277), .A2(n2273), .ZN(n2272) );
  INV_X1 U2650 ( .A(n2746), .ZN(n2273) );
  INV_X1 U2651 ( .A(n3883), .ZN(n2276) );
  INV_X1 U2652 ( .A(n3207), .ZN(n3201) );
  AOI21_X1 U2653 ( .B1(n2304), .B2(n2302), .A(n2301), .ZN(n2300) );
  INV_X1 U2654 ( .A(n3863), .ZN(n2302) );
  INV_X1 U2655 ( .A(n3853), .ZN(n2301) );
  OR2_X1 U2656 ( .A1(n3012), .A2(n2303), .ZN(n2299) );
  INV_X1 U2657 ( .A(n2304), .ZN(n2303) );
  INV_X1 U2658 ( .A(IR_REG_16__SCAN_IN), .ZN(n4853) );
  NAND2_X1 U2659 ( .A1(n4117), .A2(n4127), .ZN(n2339) );
  OR2_X1 U2660 ( .A1(n3421), .A2(n4354), .ZN(n3420) );
  NAND2_X1 U2661 ( .A1(n2253), .A2(n2252), .ZN(n3136) );
  NOR2_X1 U2662 ( .A1(n3176), .A2(n3201), .ZN(n2253) );
  INV_X1 U2663 ( .A(IR_REG_27__SCAN_IN), .ZN(n2432) );
  INV_X1 U2664 ( .A(IR_REG_28__SCAN_IN), .ZN(n2731) );
  INV_X1 U2665 ( .A(IR_REG_26__SCAN_IN), .ZN(n2429) );
  NOR2_X1 U2666 ( .A1(n2426), .A2(IR_REG_13__SCAN_IN), .ZN(n2369) );
  INV_X1 U2667 ( .A(IR_REG_6__SCAN_IN), .ZN(n2516) );
  AND2_X1 U2668 ( .A1(n2465), .A2(DATAI_23_), .ZN(n3638) );
  INV_X1 U2669 ( .A(n2413), .ZN(n2378) );
  INV_X1 U2670 ( .A(n3682), .ZN(n2382) );
  AND2_X1 U2671 ( .A1(n3632), .A2(n3633), .ZN(n3722) );
  NAND2_X1 U2672 ( .A1(n3388), .A2(n3389), .ZN(n2397) );
  NOR2_X1 U2673 ( .A1(n2689), .A2(n4886), .ZN(n2698) );
  NOR2_X1 U2674 ( .A1(n3648), .A2(n3647), .ZN(n3649) );
  INV_X1 U2675 ( .A(n3619), .ZN(n3620) );
  INV_X1 U2676 ( .A(n3723), .ZN(n2389) );
  OR2_X1 U2677 ( .A1(n3728), .A2(n3722), .ZN(n2390) );
  INV_X1 U2678 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2556) );
  NOR2_X1 U2679 ( .A1(n2557), .A2(n2556), .ZN(n2568) );
  AND2_X1 U2680 ( .A1(n2386), .A2(n3753), .ZN(n2383) );
  NAND2_X1 U2681 ( .A1(n3591), .A2(n3754), .ZN(n2386) );
  AND2_X1 U2682 ( .A1(n3746), .A2(n3754), .ZN(n2384) );
  NAND2_X1 U2683 ( .A1(n3743), .A2(n3820), .ZN(n3590) );
  NOR2_X1 U2684 ( .A1(n2591), .A2(n4826), .ZN(n2608) );
  NAND2_X1 U2685 ( .A1(n2891), .A2(n2890), .ZN(n2893) );
  NAND2_X1 U2686 ( .A1(n2311), .A2(n2880), .ZN(n2883) );
  NAND2_X1 U2687 ( .A1(n2312), .A2(n4419), .ZN(n2311) );
  INV_X1 U2688 ( .A(n2882), .ZN(n2312) );
  NOR2_X1 U2689 ( .A1(n2495), .A2(IR_REG_5__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U2690 ( .A1(n4417), .A2(REG1_REG_5__SCAN_IN), .ZN(n2318) );
  NAND2_X1 U2691 ( .A1(n4436), .A2(n3445), .ZN(n4441) );
  NAND2_X1 U2692 ( .A1(n4443), .A2(n3468), .ZN(n3469) );
  NAND2_X1 U2693 ( .A1(n4042), .A2(n3448), .ZN(n4453) );
  NAND2_X1 U2694 ( .A1(n4469), .A2(n3451), .ZN(n3455) );
  NAND2_X1 U2695 ( .A1(n2263), .A2(n4052), .ZN(n4055) );
  INV_X1 U2696 ( .A(n4053), .ZN(n2264) );
  NOR2_X1 U2697 ( .A1(n4055), .A2(n4066), .ZN(n4079) );
  XNOR2_X1 U2698 ( .A(n4082), .B(n4563), .ZN(n4485) );
  NAND2_X1 U2699 ( .A1(n4485), .A2(n4922), .ZN(n4484) );
  AND2_X1 U2700 ( .A1(n2764), .A2(n2763), .ZN(n4139) );
  NOR2_X1 U2701 ( .A1(n3972), .A2(n2308), .ZN(n2306) );
  NAND2_X1 U2702 ( .A1(n2309), .A2(n2307), .ZN(n4172) );
  AND2_X1 U2703 ( .A1(n3912), .A2(n4171), .ZN(n4153) );
  NAND2_X1 U2704 ( .A1(n3996), .A2(n4234), .ZN(n2669) );
  NAND2_X1 U2705 ( .A1(n4272), .A2(n2661), .ZN(n2325) );
  NAND2_X1 U2706 ( .A1(n3729), .A2(n3942), .ZN(n2661) );
  INV_X1 U2707 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4875) );
  OR2_X1 U2708 ( .A1(n2646), .A2(n2418), .ZN(n2656) );
  INV_X1 U2709 ( .A(n3602), .ZN(n3800) );
  OR2_X1 U2710 ( .A1(n3377), .A2(n3921), .ZN(n3378) );
  NAND2_X1 U2711 ( .A1(n2343), .A2(n2342), .ZN(n3274) );
  AOI21_X1 U2712 ( .B1(n2345), .B2(n2349), .A(n2189), .ZN(n2342) );
  NAND2_X1 U2713 ( .A1(n2532), .A2(n2340), .ZN(n2343) );
  OAI21_X1 U2714 ( .B1(n2743), .B2(n2282), .A(n2280), .ZN(n2744) );
  INV_X1 U2715 ( .A(n2281), .ZN(n2280) );
  OAI21_X1 U2716 ( .B1(n2175), .B2(n2282), .A(n3870), .ZN(n2281) );
  NAND2_X1 U2717 ( .A1(n2279), .A2(n3857), .ZN(n3242) );
  NAND2_X1 U2718 ( .A1(n2743), .A2(n2175), .ZN(n2279) );
  INV_X1 U2719 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4829) );
  NOR2_X1 U2720 ( .A1(n2510), .A2(n2509), .ZN(n2521) );
  NAND2_X1 U2721 ( .A1(n2299), .A2(n2300), .ZN(n3060) );
  AND3_X1 U2722 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2502) );
  NAND2_X1 U2723 ( .A1(n2502), .A2(REG3_REG_6__SCAN_IN), .ZN(n2510) );
  AND2_X2 U2724 ( .A1(n3848), .A2(n3851), .ZN(n3924) );
  AND2_X1 U2725 ( .A1(n3847), .A2(n2286), .ZN(n2285) );
  NAND2_X1 U2726 ( .A1(n3844), .A2(n2288), .ZN(n2286) );
  NAND2_X1 U2727 ( .A1(n4533), .A2(n2738), .ZN(n3034) );
  INV_X1 U2728 ( .A(n4543), .ZN(n2364) );
  INV_X1 U2729 ( .A(n4542), .ZN(n2365) );
  NAND2_X1 U2730 ( .A1(n4534), .A2(n4543), .ZN(n4533) );
  INV_X1 U2731 ( .A(DATAI_1_), .ZN(n2250) );
  INV_X1 U2732 ( .A(DATAI_0_), .ZN(n2249) );
  AND2_X1 U2733 ( .A1(n3954), .A2(n2338), .ZN(n2336) );
  NAND2_X1 U2734 ( .A1(n3951), .A2(n2339), .ZN(n2337) );
  OAI21_X1 U2735 ( .B1(n3954), .B2(n2337), .A(n2334), .ZN(n2333) );
  NAND2_X1 U2736 ( .A1(n2335), .A2(n2338), .ZN(n2334) );
  INV_X1 U2737 ( .A(n2339), .ZN(n2335) );
  NOR2_X1 U2738 ( .A1(n4289), .A2(n4290), .ZN(n4288) );
  AND2_X1 U2739 ( .A1(n2465), .A2(DATAI_28_), .ZN(n4127) );
  INV_X1 U2740 ( .A(n4294), .ZN(n4147) );
  NAND2_X1 U2741 ( .A1(n4160), .A2(n4147), .ZN(n4143) );
  AND2_X1 U2742 ( .A1(n2465), .A2(DATAI_27_), .ZN(n4294) );
  NOR2_X1 U2743 ( .A1(n4193), .A2(n2251), .ZN(n4160) );
  NAND2_X1 U2744 ( .A1(n4181), .A2(n4162), .ZN(n2251) );
  INV_X1 U2745 ( .A(n4162), .ZN(n4303) );
  NOR2_X1 U2746 ( .A1(n4193), .A2(n2696), .ZN(n4179) );
  OR2_X1 U2747 ( .A1(n4217), .A2(n4315), .ZN(n4193) );
  NAND2_X1 U2748 ( .A1(n4235), .A2(n4218), .ZN(n4217) );
  NOR2_X1 U2749 ( .A1(n4234), .A2(n4252), .ZN(n4235) );
  NAND2_X1 U2750 ( .A1(n2255), .A2(n4253), .ZN(n4252) );
  AND2_X1 U2751 ( .A1(n3534), .A2(n3800), .ZN(n3559) );
  NAND2_X1 U2752 ( .A1(n3559), .A2(n3715), .ZN(n4278) );
  NOR2_X2 U2753 ( .A1(n3420), .A2(n3594), .ZN(n3534) );
  INV_X1 U2754 ( .A(n3756), .ZN(n3594) );
  INV_X1 U2755 ( .A(n3576), .ZN(n3823) );
  NAND2_X1 U2756 ( .A1(n3363), .A2(n2254), .ZN(n3421) );
  AND2_X1 U2757 ( .A1(n3504), .A2(n3823), .ZN(n2254) );
  INV_X1 U2758 ( .A(n4000), .ZN(n3822) );
  INV_X1 U2759 ( .A(n3495), .ZN(n3504) );
  AND2_X1 U2760 ( .A1(n3363), .A2(n3504), .ZN(n3381) );
  INV_X1 U2761 ( .A(n3311), .ZN(n3433) );
  OR2_X1 U2762 ( .A1(n3297), .A2(n3395), .ZN(n3315) );
  INV_X1 U2763 ( .A(n4003), .ZN(n3400) );
  INV_X1 U2764 ( .A(n3291), .ZN(n3329) );
  NAND2_X1 U2765 ( .A1(n3298), .A2(n3329), .ZN(n3297) );
  INV_X1 U2766 ( .A(n4355), .ZN(n4538) );
  AND2_X1 U2767 ( .A1(n2947), .A2(n2938), .ZN(n4355) );
  INV_X1 U2768 ( .A(n4229), .ZN(n4535) );
  INV_X1 U2769 ( .A(n4358), .ZN(n4536) );
  NAND2_X1 U2770 ( .A1(n3111), .A2(n3167), .ZN(n3176) );
  INV_X1 U2771 ( .A(n2253), .ZN(n3177) );
  AND2_X1 U2772 ( .A1(n3109), .A2(n3150), .ZN(n3111) );
  NAND2_X1 U2773 ( .A1(n3087), .A2(n3089), .ZN(n3086) );
  INV_X1 U2774 ( .A(n3126), .ZN(n3016) );
  AND2_X1 U2775 ( .A1(n4550), .A2(n3001), .ZN(n3087) );
  NAND2_X1 U2776 ( .A1(n3054), .A2(n3055), .ZN(n4551) );
  INV_X1 U2777 ( .A(n4592), .ZN(n4585) );
  NAND2_X1 U2778 ( .A1(n2360), .A2(n2361), .ZN(n2359) );
  INV_X1 U2779 ( .A(n2431), .ZN(n2360) );
  INV_X1 U2780 ( .A(IR_REG_20__SCAN_IN), .ZN(n2723) );
  AND2_X1 U2781 ( .A1(n2614), .A2(n2606), .ZN(n4081) );
  AND2_X1 U2782 ( .A1(n2574), .A2(n2567), .ZN(n3462) );
  INV_X1 U2783 ( .A(IR_REG_7__SCAN_IN), .ZN(n4843) );
  AOI21_X1 U2784 ( .B1(n3162), .B2(n3161), .A(n3160), .ZN(n3197) );
  INV_X1 U2785 ( .A(n3638), .ZN(n4218) );
  INV_X1 U2786 ( .A(n3608), .ZN(n3715) );
  NAND2_X1 U2787 ( .A1(n3774), .A2(n3775), .ZN(n3728) );
  NAND2_X1 U2788 ( .A1(n2396), .A2(n2397), .ZN(n3429) );
  NAND2_X1 U2789 ( .A1(n3390), .A2(n2398), .ZN(n2396) );
  NOR2_X1 U2790 ( .A1(n3124), .A2(n2410), .ZN(n3128) );
  OR2_X1 U2791 ( .A1(n3078), .A2(n3077), .ZN(n2233) );
  NOR2_X1 U2792 ( .A1(n3081), .A2(n3082), .ZN(n3124) );
  NAND2_X1 U2793 ( .A1(n2236), .A2(n2391), .ZN(n3489) );
  AOI21_X1 U2794 ( .B1(n2392), .B2(n2394), .A(n2206), .ZN(n2391) );
  INV_X1 U2795 ( .A(n2398), .ZN(n2392) );
  NAND2_X1 U2796 ( .A1(n2390), .A2(n3723), .ZN(n3787) );
  OR2_X1 U2797 ( .A1(n2953), .A2(n2949), .ZN(n3821) );
  NAND2_X1 U2798 ( .A1(n2405), .A2(n3735), .ZN(n3812) );
  NAND2_X1 U2799 ( .A1(n3736), .A2(n3734), .ZN(n2405) );
  OAI21_X1 U2800 ( .B1(n3691), .B2(n2443), .A(n2709), .ZN(n4128) );
  OAI21_X1 U2801 ( .B1(n3813), .B2(n2443), .A(n2703), .ZN(n4295) );
  NAND2_X1 U2802 ( .A1(n2684), .A2(n2683), .ZN(n4213) );
  OAI211_X1 U2803 ( .C1(n4254), .C2(n2443), .A(n2437), .B(n2436), .ZN(n4226)
         );
  NAND4_X1 U2804 ( .A1(n2585), .A2(n2584), .A3(n2583), .A4(n2582), .ZN(n4001)
         );
  NOR2_X1 U2805 ( .A1(n2415), .A2(n2414), .ZN(n2447) );
  OR2_X1 U2806 ( .A1(n2642), .A2(n2457), .ZN(n2464) );
  XNOR2_X1 U2807 ( .A(n2882), .B(n4419), .ZN(n2876) );
  NAND2_X1 U2808 ( .A1(n2876), .A2(REG1_REG_3__SCAN_IN), .ZN(n2880) );
  XNOR2_X1 U2809 ( .A(n2883), .B(n2310), .ZN(n4038) );
  INV_X1 U2810 ( .A(n4418), .ZN(n2310) );
  XNOR2_X1 U2811 ( .A(n2893), .B(n4418), .ZN(n4030) );
  XNOR2_X1 U2812 ( .A(n2317), .B(n3022), .ZN(n2982) );
  NAND2_X1 U2813 ( .A1(n2257), .A2(n2256), .ZN(n3463) );
  AND2_X1 U2814 ( .A1(n2262), .A2(n2259), .ZN(n3027) );
  NAND2_X1 U2815 ( .A1(n3025), .A2(REG2_REG_6__SCAN_IN), .ZN(n2259) );
  NAND2_X1 U2816 ( .A1(n4431), .A2(n3467), .ZN(n4444) );
  NAND2_X1 U2817 ( .A1(n4444), .A2(n4445), .ZN(n4443) );
  XNOR2_X1 U2818 ( .A(n3447), .B(n2265), .ZN(n4043) );
  NAND2_X1 U2819 ( .A1(n4043), .A2(REG1_REG_10__SCAN_IN), .ZN(n4042) );
  NAND2_X1 U2820 ( .A1(n4463), .A2(n3474), .ZN(n4054) );
  INV_X1 U2821 ( .A(n2315), .ZN(n4067) );
  NOR2_X1 U2822 ( .A1(n4475), .A2(n4474), .ZN(n4473) );
  OR2_X1 U2823 ( .A1(n4430), .A2(n4019), .ZN(n4492) );
  AOI21_X1 U2824 ( .B1(n4094), .B2(REG2_REG_18__SCAN_IN), .A(n4093), .ZN(n4096) );
  INV_X1 U2825 ( .A(n4492), .ZN(n4464) );
  INV_X1 U2826 ( .A(n4298), .ZN(n4117) );
  AOI21_X1 U2827 ( .B1(n2688), .B2(n2357), .A(n2180), .ZN(n4158) );
  NAND2_X1 U2828 ( .A1(n2309), .A2(n2761), .ZN(n4188) );
  AND2_X1 U2829 ( .A1(n2675), .A2(n2674), .ZN(n4319) );
  NAND2_X1 U2830 ( .A1(n3906), .A2(DATAI_24_), .ZN(n4198) );
  AND4_X1 U2831 ( .A1(n2636), .A2(n2635), .A3(n2634), .A4(n2633), .ZN(n3758)
         );
  AND2_X1 U2832 ( .A1(n2622), .A2(n2621), .ZN(n3799) );
  OR2_X1 U2833 ( .A1(n3536), .A2(n4579), .ZN(n4239) );
  NAND2_X1 U2834 ( .A1(n2347), .A2(n2555), .ZN(n3290) );
  NAND2_X1 U2835 ( .A1(n2350), .A2(n2348), .ZN(n2347) );
  NAND2_X1 U2836 ( .A1(n2350), .A2(n2353), .ZN(n3241) );
  NAND2_X1 U2837 ( .A1(n2743), .A2(n3855), .ZN(n3133) );
  NOR2_X1 U2838 ( .A1(n2409), .A2(n3927), .ZN(n2326) );
  INV_X1 U2839 ( .A(n4239), .ZN(n4618) );
  NAND2_X1 U2840 ( .A1(n4592), .A2(n2904), .ZN(n4615) );
  OR2_X1 U2841 ( .A1(n2827), .A2(n2902), .ZN(n4610) );
  NAND2_X1 U2842 ( .A1(n2847), .A2(n2951), .ZN(n4559) );
  INV_X1 U2843 ( .A(n2291), .ZN(n2290) );
  NAND2_X1 U2844 ( .A1(n2783), .A2(n2289), .ZN(n2294) );
  INV_X1 U2845 ( .A(n2947), .ZN(n4409) );
  NAND2_X1 U2846 ( .A1(n2794), .A2(IR_REG_31__SCAN_IN), .ZN(n2779) );
  INV_X1 U2847 ( .A(n2774), .ZN(n4411) );
  INV_X1 U2848 ( .A(n4075), .ZN(n4094) );
  INV_X1 U2849 ( .A(n4084), .ZN(n4562) );
  INV_X1 U2850 ( .A(n4448), .ZN(n4569) );
  INV_X1 U2851 ( .A(n3465), .ZN(n4571) );
  OR2_X1 U2852 ( .A1(n2475), .A2(n2553), .ZN(n2448) );
  NAND2_X1 U2853 ( .A1(n2375), .A2(n3777), .ZN(n2373) );
  INV_X1 U2854 ( .A(n2321), .ZN(n2886) );
  XNOR2_X1 U2855 ( .A(n4090), .B(n4089), .ZN(n2314) );
  OR2_X1 U2856 ( .A1(n4119), .A2(n4350), .ZN(n2825) );
  OR2_X1 U2857 ( .A1(n4126), .A2(n4350), .ZN(n2810) );
  OAI211_X1 U2858 ( .C1(n2331), .C2(n2416), .A(n2266), .B(n2181), .ZN(n2831)
         );
  NAND2_X1 U2859 ( .A1(n4601), .A2(n4365), .ZN(n2331) );
  AND2_X1 U2860 ( .A1(n3855), .A2(n2283), .ZN(n2175) );
  NOR2_X1 U2861 ( .A1(n4087), .A2(n4088), .ZN(n2177) );
  AND2_X1 U2862 ( .A1(n2404), .A2(n2403), .ZN(n2178) );
  INV_X1 U2863 ( .A(n2349), .ZN(n2348) );
  NAND2_X1 U2864 ( .A1(n2188), .A2(n2353), .ZN(n2349) );
  INV_X1 U2865 ( .A(n3227), .ZN(n2252) );
  AND2_X1 U2866 ( .A1(n2200), .A2(n2227), .ZN(n2179) );
  OAI211_X1 U2867 ( .C1(n4279), .C2(n2443), .A(n2660), .B(n2659), .ZN(n4333)
         );
  AND2_X1 U2868 ( .A1(n4316), .A2(n2696), .ZN(n2180) );
  INV_X1 U2869 ( .A(n2388), .ZN(n2229) );
  NOR2_X1 U2870 ( .A1(n3788), .A2(n2389), .ZN(n2388) );
  OR2_X1 U2871 ( .A1(n4601), .A2(REG0_REG_29__SCAN_IN), .ZN(n2181) );
  AND2_X1 U2872 ( .A1(n2327), .A2(n2328), .ZN(n2182) );
  NAND2_X1 U2873 ( .A1(n3582), .A2(n3581), .ZN(n3742) );
  AND2_X1 U2874 ( .A1(n2390), .A2(n2388), .ZN(n2183) );
  NAND2_X1 U2875 ( .A1(n4008), .A2(n3146), .ZN(n2184) );
  NAND2_X1 U2876 ( .A1(n2588), .A2(n2367), .ZN(n2777) );
  NOR2_X1 U2877 ( .A1(n4488), .A2(REG1_REG_16__SCAN_IN), .ZN(n2185) );
  NAND2_X1 U2878 ( .A1(n2688), .A2(n2687), .ZN(n4170) );
  NAND2_X1 U2879 ( .A1(n2385), .A2(n3592), .ZN(n3752) );
  NAND2_X1 U2880 ( .A1(n2219), .A2(n2383), .ZN(n3706) );
  INV_X1 U2881 ( .A(IR_REG_3__SCAN_IN), .ZN(n2477) );
  AND2_X1 U2882 ( .A1(n4420), .A2(REG1_REG_2__SCAN_IN), .ZN(n2186) );
  AND2_X1 U2883 ( .A1(n2300), .A2(n2741), .ZN(n2187) );
  INV_X1 U2884 ( .A(n4419), .ZN(n2881) );
  AND2_X1 U2885 ( .A1(n2489), .A2(n2479), .ZN(n4419) );
  OR2_X1 U2886 ( .A1(n4004), .A2(n3263), .ZN(n2188) );
  NAND2_X1 U2887 ( .A1(n3142), .A2(n3143), .ZN(n2404) );
  AND2_X1 U2888 ( .A1(n3400), .A2(n3329), .ZN(n2189) );
  INV_X1 U2889 ( .A(IR_REG_29__SCAN_IN), .ZN(n2361) );
  INV_X1 U2890 ( .A(IR_REG_31__SCAN_IN), .ZN(n2553) );
  INV_X1 U2891 ( .A(n3024), .ZN(n2262) );
  AND3_X1 U2892 ( .A1(n2791), .A2(n4795), .A3(n2778), .ZN(n2190) );
  INV_X1 U2893 ( .A(n2410), .ZN(n2403) );
  INV_X1 U2894 ( .A(n2868), .ZN(n4421) );
  OAI211_X1 U2895 ( .C1(IR_REG_1__SCAN_IN), .C2(IR_REG_31__SCAN_IN), .A(n2213), 
        .B(n2313), .ZN(n2868) );
  AND2_X1 U2896 ( .A1(n2500), .A2(n2184), .ZN(n2191) );
  AND2_X1 U2897 ( .A1(n3474), .A2(n2264), .ZN(n2192) );
  NAND2_X1 U2898 ( .A1(n2319), .A2(n2318), .ZN(n2317) );
  AND2_X1 U2899 ( .A1(n2176), .A2(IR_REG_30__SCAN_IN), .ZN(n2193) );
  AND2_X1 U2900 ( .A1(n2190), .A2(n2429), .ZN(n2194) );
  INV_X1 U2901 ( .A(IR_REG_2__SCAN_IN), .ZN(n2474) );
  NAND2_X2 U2902 ( .A1(n2844), .A2(n4408), .ZN(n2443) );
  INV_X1 U2903 ( .A(n4415), .ZN(n2265) );
  NAND2_X1 U2904 ( .A1(n2532), .A2(n2351), .ZN(n2350) );
  NAND2_X1 U2905 ( .A1(n3668), .A2(n3735), .ZN(n2195) );
  NAND2_X1 U2906 ( .A1(n2244), .A2(n2629), .ZN(n2638) );
  NAND2_X1 U2907 ( .A1(n3325), .A2(n2408), .ZN(n3390) );
  AND2_X1 U2908 ( .A1(n2241), .A2(n2239), .ZN(n3572) );
  INV_X1 U2909 ( .A(IR_REG_22__SCAN_IN), .ZN(n2428) );
  AND2_X1 U2910 ( .A1(n4295), .A2(n4303), .ZN(n2196) );
  INV_X1 U2911 ( .A(n3951), .ZN(n2338) );
  OR2_X1 U2912 ( .A1(n4128), .A2(n4294), .ZN(n2197) );
  INV_X1 U2913 ( .A(n2255), .ZN(n4342) );
  NOR2_X1 U2914 ( .A1(n4278), .A2(n4277), .ZN(n2255) );
  INV_X1 U2915 ( .A(n4316), .ZN(n4196) );
  NAND2_X1 U2916 ( .A1(n2695), .A2(n2694), .ZN(n4316) );
  AND2_X1 U2917 ( .A1(n2220), .A2(n3581), .ZN(n2198) );
  NOR2_X1 U2918 ( .A1(n3290), .A2(n3930), .ZN(n2199) );
  BUF_X1 U2919 ( .A(n2588), .Z(n2626) );
  INV_X1 U2920 ( .A(n2686), .ZN(n2687) );
  NOR2_X1 U2921 ( .A1(n4213), .A2(n4315), .ZN(n2686) );
  INV_X1 U2922 ( .A(n2308), .ZN(n2307) );
  OR2_X1 U2923 ( .A1(n3946), .A2(n3941), .ZN(n2308) );
  AND2_X1 U2924 ( .A1(n2387), .A2(n3643), .ZN(n2200) );
  OR2_X1 U2925 ( .A1(n3682), .A2(n2378), .ZN(n2201) );
  OR2_X1 U2926 ( .A1(n3464), .A2(n4814), .ZN(n2202) );
  AND2_X1 U2927 ( .A1(n4319), .A2(n3638), .ZN(n3946) );
  AND2_X1 U2928 ( .A1(n2356), .A2(n2357), .ZN(n2203) );
  INV_X1 U2929 ( .A(n3775), .ZN(n2228) );
  NAND2_X1 U2930 ( .A1(n2327), .A2(n2326), .ZN(n3067) );
  INV_X2 U2931 ( .A(n4599), .ZN(n4601) );
  AND2_X1 U2932 ( .A1(n3847), .A2(n3844), .ZN(n2204) );
  AND2_X1 U2933 ( .A1(n3906), .A2(DATAI_20_), .ZN(n4277) );
  INV_X1 U2934 ( .A(n4277), .ZN(n3942) );
  XNOR2_X1 U2935 ( .A(n2779), .B(n2778), .ZN(n2788) );
  INV_X1 U2936 ( .A(n3861), .ZN(n2305) );
  NAND2_X1 U2937 ( .A1(n2532), .A2(n2531), .ZN(n3135) );
  NAND2_X1 U2938 ( .A1(n2501), .A2(n2500), .ZN(n3102) );
  INV_X1 U2939 ( .A(n3857), .ZN(n2282) );
  AND2_X1 U2940 ( .A1(n2401), .A2(n2400), .ZN(n2205) );
  INV_X1 U2941 ( .A(n4253), .ZN(n4332) );
  NAND2_X1 U2942 ( .A1(n3906), .A2(DATAI_21_), .ZN(n4253) );
  AND2_X1 U2943 ( .A1(n3879), .A2(n3836), .ZN(n3925) );
  INV_X1 U2944 ( .A(n3925), .ZN(n2277) );
  AND2_X1 U2945 ( .A1(n3884), .A2(n3885), .ZN(n3931) );
  INV_X1 U2946 ( .A(n3874), .ZN(n2283) );
  OR2_X1 U2947 ( .A1(n4430), .A2(n2861), .ZN(n4103) );
  NAND2_X1 U2948 ( .A1(n4544), .A2(n4585), .ZN(n4594) );
  INV_X1 U2949 ( .A(n3834), .ZN(n3777) );
  AND2_X1 U2950 ( .A1(n3398), .A2(n3397), .ZN(n2206) );
  OR2_X1 U2951 ( .A1(n2783), .A2(n2433), .ZN(n2207) );
  AND2_X1 U2952 ( .A1(n4081), .A2(REG2_REG_15__SCAN_IN), .ZN(n2208) );
  INV_X1 U2953 ( .A(n2409), .ZN(n2328) );
  INV_X1 U2954 ( .A(IR_REG_21__SCAN_IN), .ZN(n2222) );
  INV_X1 U2955 ( .A(IR_REG_4__SCAN_IN), .ZN(n2420) );
  NAND2_X1 U2956 ( .A1(n2297), .A2(n2176), .ZN(n2837) );
  NOR2_X1 U2957 ( .A1(n4084), .A2(REG1_REG_17__SCAN_IN), .ZN(n2209) );
  INV_X1 U2958 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2261) );
  INV_X1 U2959 ( .A(IR_REG_30__SCAN_IN), .ZN(n2296) );
  NAND2_X1 U2960 ( .A1(n4437), .A2(REG1_REG_8__SCAN_IN), .ZN(n4436) );
  AND2_X1 U2961 ( .A1(n2317), .A2(n3022), .ZN(n2210) );
  XNOR2_X1 U2962 ( .A(n4071), .B(n4563), .ZN(n4488) );
  NAND2_X1 U2963 ( .A1(n4479), .A2(n4480), .ZN(n4478) );
  NAND2_X1 U2964 ( .A1(n2215), .A2(n2214), .ZN(n3621) );
  NAND3_X1 U2965 ( .A1(n3590), .A2(n3742), .A3(n2384), .ZN(n2219) );
  NAND2_X4 U2966 ( .A1(n2916), .A2(n2915), .ZN(n3676) );
  XNOR2_X2 U2967 ( .A(n2726), .B(n2222), .ZN(n2735) );
  XNOR2_X1 U2968 ( .A(n3690), .B(n3689), .ZN(n3696) );
  NAND2_X2 U2969 ( .A1(n2234), .A2(n2232), .ZN(n3159) );
  NAND2_X1 U2970 ( .A1(n3325), .A2(n2237), .ZN(n2236) );
  INV_X1 U2971 ( .A(n3489), .ZN(n2242) );
  INV_X1 U2972 ( .A(n3055), .ZN(n2973) );
  MUX2_X1 U2973 ( .A(n2868), .B(n2250), .S(n2465), .Z(n3054) );
  NOR2_X2 U2974 ( .A1(n3136), .A2(n3263), .ZN(n3298) );
  NAND2_X2 U2975 ( .A1(n2368), .A2(IR_REG_31__SCAN_IN), .ZN(n2818) );
  NAND2_X1 U2976 ( .A1(n3025), .A2(n2260), .ZN(n2256) );
  NAND3_X1 U2977 ( .A1(n2257), .A2(n2256), .A3(n2202), .ZN(n3466) );
  XNOR2_X1 U2978 ( .A(n3473), .B(n4567), .ZN(n4465) );
  NAND2_X1 U2979 ( .A1(n4463), .A2(n2192), .ZN(n2263) );
  NOR2_X1 U2980 ( .A1(n4810), .A2(n4057), .ZN(n4078) );
  OAI21_X1 U2981 ( .B1(n2314), .B2(n4103), .A(n2177), .ZN(U3258) );
  NAND2_X1 U2982 ( .A1(n3292), .A2(n2272), .ZN(n2271) );
  NAND2_X1 U2983 ( .A1(n2271), .A2(n2274), .ZN(n3377) );
  NAND2_X1 U2984 ( .A1(n4534), .A2(n2284), .ZN(n2287) );
  NAND2_X1 U2985 ( .A1(n2287), .A2(n2285), .ZN(n3088) );
  INV_X1 U2986 ( .A(n2783), .ZN(n2297) );
  NAND2_X1 U2987 ( .A1(n2297), .A2(n2193), .ZN(n2293) );
  OAI21_X1 U2988 ( .B1(n3012), .B2(n3010), .A(n3863), .ZN(n3103) );
  AOI21_X1 U2989 ( .B1(n3010), .B2(n3863), .A(n2305), .ZN(n2304) );
  NAND2_X1 U2990 ( .A1(n2760), .A2(n2759), .ZN(n2309) );
  NAND2_X1 U2991 ( .A1(n2309), .A2(n2306), .ZN(n2764) );
  NAND3_X1 U2992 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .A3(
        IR_REG_0__SCAN_IN), .ZN(n2313) );
  NAND2_X1 U2993 ( .A1(n2501), .A2(n2191), .ZN(n2327) );
  NAND2_X1 U2994 ( .A1(n2812), .A2(n2336), .ZN(n2329) );
  OR2_X1 U2995 ( .A1(n2812), .A2(n2337), .ZN(n2330) );
  AOI21_X1 U2996 ( .B1(n4113), .B2(n4594), .A(n2416), .ZN(n2828) );
  NAND3_X1 U2997 ( .A1(n2330), .A2(n2332), .A3(n2329), .ZN(n4113) );
  OR2_X1 U2998 ( .A1(n4005), .A2(n3227), .ZN(n2353) );
  NAND2_X1 U2999 ( .A1(n2688), .A2(n2203), .ZN(n2354) );
  NAND2_X1 U3000 ( .A1(n2354), .A2(n2355), .ZN(n4142) );
  INV_X2 U3001 ( .A(n2434), .ZN(n2844) );
  OAI21_X2 U3002 ( .B1(n2732), .B2(n2359), .A(n2358), .ZN(n2434) );
  NAND2_X1 U3003 ( .A1(n4542), .A2(n2467), .ZN(n2363) );
  NAND3_X1 U3004 ( .A1(n2363), .A2(n2480), .A3(n2362), .ZN(n2482) );
  NAND2_X1 U3005 ( .A1(n4540), .A2(n2467), .ZN(n3033) );
  NAND2_X1 U3006 ( .A1(n2365), .A2(n2364), .ZN(n4540) );
  NAND2_X1 U3007 ( .A1(n2588), .A2(n2366), .ZN(n2368) );
  AND2_X1 U3008 ( .A1(n2588), .A2(n2427), .ZN(n2407) );
  INV_X1 U3009 ( .A(n2407), .ZN(n2727) );
  NAND2_X1 U3010 ( .A1(n2962), .A2(n2960), .ZN(n2961) );
  XNOR2_X1 U3011 ( .A(n2929), .B(n2927), .ZN(n2960) );
  NOR2_X1 U3012 ( .A1(n2495), .A2(n2426), .ZN(n2586) );
  AND2_X2 U3013 ( .A1(n2370), .A2(n2369), .ZN(n2588) );
  INV_X1 U3014 ( .A(n2495), .ZN(n2370) );
  NAND2_X1 U3015 ( .A1(n3690), .A2(n2372), .ZN(n2371) );
  OAI211_X1 U3016 ( .C1(n3690), .C2(n2373), .A(n2371), .B(n3688), .ZN(U3217)
         );
  NAND3_X1 U3017 ( .A1(n3590), .A2(n3742), .A3(n3746), .ZN(n2385) );
  NAND2_X1 U3018 ( .A1(n3081), .A2(n2403), .ZN(n2400) );
  NAND2_X1 U3019 ( .A1(n2407), .A2(n2406), .ZN(n2783) );
  NAND2_X2 U3020 ( .A1(n2916), .A2(n2944), .ZN(n2923) );
  OAI22_X1 U3021 ( .A1(n2950), .A2(n2922), .B1(n3054), .B2(n3676), .ZN(n2924)
         );
  OAI22_X1 U3022 ( .A1(n2917), .A2(n2922), .B1(n3676), .B2(n2955), .ZN(n2918)
         );
  NAND2_X1 U3023 ( .A1(n2920), .A2(n3665), .ZN(n2921) );
  OR2_X1 U3024 ( .A1(n3324), .A2(n3323), .ZN(n2408) );
  AND2_X1 U3025 ( .A1(n3166), .A2(n3150), .ZN(n2409) );
  AND2_X1 U3026 ( .A1(n3123), .A2(n3122), .ZN(n2410) );
  OR2_X1 U3027 ( .A1(n3729), .A2(n3942), .ZN(n2411) );
  AND2_X1 U3028 ( .A1(n4359), .A2(n3823), .ZN(n2412) );
  OR2_X1 U3029 ( .A1(n3675), .A2(n3674), .ZN(n2413) );
  INV_X1 U3030 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2509) );
  AND2_X1 U3031 ( .A1(n2459), .A2(REG2_REG_2__SCAN_IN), .ZN(n2414) );
  INV_X1 U3032 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2533) );
  NAND2_X1 U3033 ( .A1(n3906), .A2(DATAI_25_), .ZN(n4181) );
  AOI21_X1 U3034 ( .B1(n3550), .B2(n2655), .A(n2654), .ZN(n4272) );
  NAND2_X1 U3035 ( .A1(n3906), .A2(DATAI_22_), .ZN(n4228) );
  INV_X1 U3036 ( .A(n4228), .ZN(n4234) );
  OAI21_X1 U3037 ( .B1(n3797), .B2(n3796), .A(n3711), .ZN(n3611) );
  OAI21_X1 U3038 ( .B1(n3618), .B2(n3617), .A(n3710), .ZN(n3619) );
  INV_X1 U3039 ( .A(n4181), .ZN(n2696) );
  INV_X1 U3040 ( .A(n3652), .ZN(n3647) );
  AND2_X1 U3041 ( .A1(n4298), .A2(n4127), .ZN(n3903) );
  INV_X1 U3042 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U3043 ( .A1(n2929), .A2(n2928), .ZN(n2930) );
  CLKBUF_X3 U3044 ( .A(n3145), .Z(n3662) );
  INV_X1 U3045 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4826) );
  AND2_X1 U3046 ( .A1(n4231), .A2(n3638), .ZN(n2676) );
  AND2_X1 U3047 ( .A1(n2735), .A2(n4411), .ZN(n2938) );
  NAND2_X1 U3048 ( .A1(n2950), .A2(n3049), .ZN(n3842) );
  OR3_X1 U3049 ( .A1(n2541), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2543) );
  INV_X1 U3050 ( .A(n3042), .ZN(n3001) );
  OR3_X1 U3051 ( .A1(n2678), .A2(n3701), .A3(n3769), .ZN(n2689) );
  NAND2_X1 U3052 ( .A1(n3699), .A2(n3649), .ZN(n3765) );
  AOI22_X1 U3053 ( .A1(n3145), .A2(n2973), .B1(IR_REG_0__SCAN_IN), .B2(n2914), 
        .ZN(n2919) );
  NAND2_X1 U3054 ( .A1(n2662), .A2(REG3_REG_22__SCAN_IN), .ZN(n2678) );
  INV_X1 U3055 ( .A(n3146), .ZN(n3150) );
  OR2_X1 U3056 ( .A1(n3683), .A2(n2443), .ZN(n2719) );
  NAND2_X1 U3057 ( .A1(n2883), .A2(n4418), .ZN(n2884) );
  INV_X1 U3058 ( .A(n3954), .ZN(n2721) );
  INV_X1 U3059 ( .A(n3996), .ZN(n4336) );
  INV_X1 U3060 ( .A(n3931), .ZN(n2617) );
  INV_X1 U3061 ( .A(n3999), .ZN(n4359) );
  OR2_X1 U3062 ( .A1(n2547), .A2(n4829), .ZN(n2557) );
  NAND2_X1 U3063 ( .A1(n2521), .A2(REG3_REG_8__SCAN_IN), .ZN(n2534) );
  INV_X1 U3064 ( .A(n4198), .ZN(n4315) );
  INV_X1 U3065 ( .A(n3163), .ZN(n3167) );
  AND2_X1 U3066 ( .A1(n2767), .A2(n2766), .ZN(n4215) );
  AND2_X1 U3067 ( .A1(n2988), .A2(n2951), .ZN(n2943) );
  NOR2_X1 U3068 ( .A1(n2543), .A2(IR_REG_9__SCAN_IN), .ZN(n2564) );
  AND2_X1 U3069 ( .A1(n2657), .A2(REG3_REG_21__SCAN_IN), .ZN(n2662) );
  OR2_X1 U3070 ( .A1(n2534), .A2(n2533), .ZN(n2547) );
  AND2_X1 U3071 ( .A1(n2991), .A2(STATE_REG_SCAN_IN), .ZN(n3831) );
  AND2_X1 U3072 ( .A1(n2719), .A2(n2718), .ZN(n4298) );
  NAND2_X1 U3073 ( .A1(n4038), .A2(REG1_REG_4__SCAN_IN), .ZN(n4037) );
  INV_X1 U3074 ( .A(n4103), .ZN(n4499) );
  AND2_X1 U3075 ( .A1(n4245), .A2(n4536), .ZN(n4256) );
  INV_X1 U3076 ( .A(n4621), .ZN(n4251) );
  INV_X1 U3077 ( .A(n4615), .ZN(n4549) );
  INV_X1 U3078 ( .A(n4127), .ZN(n3685) );
  AND2_X1 U3079 ( .A1(n2908), .A2(n2774), .ZN(n4592) );
  AND2_X1 U3080 ( .A1(n2856), .A2(n2854), .ZN(n4498) );
  INV_X1 U3081 ( .A(n3831), .ZN(n3786) );
  OR2_X1 U3082 ( .A1(n2953), .A2(n2941), .ZN(n3834) );
  OAI211_X1 U3083 ( .C1(n2642), .C2(n4348), .A(n2649), .B(n2648), .ZN(n4269)
         );
  OR2_X1 U3084 ( .A1(n4430), .A2(n4409), .ZN(n4505) );
  AND2_X1 U3085 ( .A1(n3304), .A2(n3068), .ZN(n4621) );
  NAND2_X1 U3086 ( .A1(n4612), .A2(n4361), .ZN(n4350) );
  OR2_X1 U3087 ( .A1(n4119), .A2(n4404), .ZN(n2830) );
  NAND2_X1 U3088 ( .A1(n4601), .A2(n4361), .ZN(n4404) );
  OR2_X1 U3089 ( .A1(n2827), .A2(n2935), .ZN(n4599) );
  INV_X1 U3090 ( .A(n4559), .ZN(n4558) );
  AND2_X1 U3091 ( .A1(n2987), .A2(STATE_REG_SCAN_IN), .ZN(n4560) );
  XNOR2_X1 U3092 ( .A(n2554), .B(IR_REG_10__SCAN_IN), .ZN(n4415) );
  AND2_X1 U3093 ( .A1(n2527), .A2(n2519), .ZN(n4416) );
  INV_X1 U3094 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2807) );
  NAND2_X1 U3095 ( .A1(n2568), .A2(REG3_REG_12__SCAN_IN), .ZN(n2580) );
  AND2_X1 U3096 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2417) );
  NAND2_X1 U3097 ( .A1(REG3_REG_19__SCAN_IN), .A2(REG3_REG_18__SCAN_IN), .ZN(
        n2418) );
  NOR2_X1 U3098 ( .A1(n2657), .A2(REG3_REG_21__SCAN_IN), .ZN(n2419) );
  OR2_X1 U3099 ( .A1(n2662), .A2(n2419), .ZN(n4254) );
  NAND2_X1 U3100 ( .A1(n2421), .A2(n2475), .ZN(n2495) );
  NAND4_X1 U3101 ( .A1(n2425), .A2(n2424), .A3(n2423), .A4(n2422), .ZN(n2426)
         );
  NAND3_X1 U3102 ( .A1(n2432), .A2(n2731), .A3(n2429), .ZN(n2433) );
  AOI22_X1 U3103 ( .A1(n2459), .A2(REG2_REG_21__SCAN_IN), .B1(n2460), .B2(
        REG0_REG_21__SCAN_IN), .ZN(n2437) );
  NAND2_X1 U3104 ( .A1(n2484), .A2(REG1_REG_21__SCAN_IN), .ZN(n2436) );
  INV_X1 U3105 ( .A(n4226), .ZN(n4271) );
  NAND2_X1 U3106 ( .A1(n2439), .A2(n2438), .ZN(n2441) );
  NAND2_X1 U3107 ( .A1(n2731), .A2(IR_REG_27__SCAN_IN), .ZN(n2440) );
  INV_X1 U3108 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2442) );
  OR2_X1 U3109 ( .A1(n2458), .A2(n2442), .ZN(n2445) );
  NAND2_X1 U3110 ( .A1(n2468), .A2(REG3_REG_2__SCAN_IN), .ZN(n2444) );
  AND2_X1 U3111 ( .A1(n2445), .A2(n2444), .ZN(n2446) );
  INV_X1 U3112 ( .A(n4420), .ZN(n2450) );
  INV_X1 U3113 ( .A(n4552), .ZN(n2955) );
  NAND2_X1 U3114 ( .A1(n4012), .A2(n2955), .ZN(n3845) );
  AND2_X2 U3115 ( .A1(n3845), .A2(n2738), .ZN(n4543) );
  NAND2_X1 U3116 ( .A1(n2459), .A2(REG2_REG_1__SCAN_IN), .ZN(n2455) );
  NAND2_X1 U3117 ( .A1(n2174), .A2(REG0_REG_1__SCAN_IN), .ZN(n2454) );
  INV_X1 U3118 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2451) );
  OR2_X1 U3119 ( .A1(n2172), .A2(n2451), .ZN(n2453) );
  NAND2_X1 U3120 ( .A1(n2468), .A2(REG3_REG_1__SCAN_IN), .ZN(n2452) );
  NAND2_X1 U3121 ( .A1(n2456), .A2(n3054), .ZN(n3840) );
  NAND2_X1 U3122 ( .A1(n3840), .A2(n3842), .ZN(n2736) );
  INV_X1 U3123 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2457) );
  NAND2_X1 U3124 ( .A1(n2468), .A2(REG3_REG_0__SCAN_IN), .ZN(n2463) );
  NAND2_X1 U3125 ( .A1(n2459), .A2(REG2_REG_0__SCAN_IN), .ZN(n2462) );
  NAND2_X1 U3126 ( .A1(n2460), .A2(REG0_REG_0__SCAN_IN), .ZN(n2461) );
  AND2_X1 U3127 ( .A1(n4013), .A2(n2973), .ZN(n3046) );
  NAND2_X1 U3128 ( .A1(n2736), .A2(n3046), .ZN(n3048) );
  NAND2_X1 U3129 ( .A1(n2456), .A2(n3049), .ZN(n2466) );
  NAND2_X1 U3130 ( .A1(n3048), .A2(n2466), .ZN(n4542) );
  NAND2_X1 U3131 ( .A1(n2917), .A2(n2955), .ZN(n2467) );
  INV_X1 U3132 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2469) );
  NAND2_X1 U3133 ( .A1(n2670), .A2(n2469), .ZN(n2473) );
  NAND2_X1 U3134 ( .A1(n2484), .A2(REG1_REG_3__SCAN_IN), .ZN(n2472) );
  NAND2_X1 U3135 ( .A1(n2460), .A2(REG0_REG_3__SCAN_IN), .ZN(n2471) );
  NAND2_X1 U3136 ( .A1(n2459), .A2(REG2_REG_3__SCAN_IN), .ZN(n2470) );
  NAND4_X1 U3137 ( .A1(n2473), .A2(n2472), .A3(n2471), .A4(n2470), .ZN(n4011)
         );
  NAND2_X1 U3138 ( .A1(n2475), .A2(n2474), .ZN(n2476) );
  NAND2_X1 U3139 ( .A1(n2476), .A2(IR_REG_31__SCAN_IN), .ZN(n2478) );
  NAND2_X1 U3140 ( .A1(n2478), .A2(n2477), .ZN(n2489) );
  OR2_X1 U3141 ( .A1(n2478), .A2(n2477), .ZN(n2479) );
  MUX2_X1 U3142 ( .A(n4419), .B(DATAI_3_), .S(n2465), .Z(n3042) );
  NAND2_X1 U3143 ( .A1(n4011), .A2(n3042), .ZN(n2480) );
  NAND2_X1 U3144 ( .A1(n4539), .A2(n3001), .ZN(n2481) );
  NAND2_X1 U3145 ( .A1(n2482), .A2(n2481), .ZN(n3090) );
  INV_X1 U3146 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2483) );
  XNOR2_X1 U3147 ( .A(n2483), .B(REG3_REG_3__SCAN_IN), .ZN(n3098) );
  NAND2_X1 U31480 ( .A1(n2670), .A2(n3098), .ZN(n2488) );
  NAND2_X1 U31490 ( .A1(n2484), .A2(REG1_REG_4__SCAN_IN), .ZN(n2487) );
  NAND2_X1 U3150 ( .A1(n2459), .A2(REG2_REG_4__SCAN_IN), .ZN(n2486) );
  NAND2_X1 U3151 ( .A1(n2460), .A2(REG0_REG_4__SCAN_IN), .ZN(n2485) );
  INV_X1 U3152 ( .A(n4010), .ZN(n3004) );
  NAND2_X1 U3153 ( .A1(n2489), .A2(IR_REG_31__SCAN_IN), .ZN(n2490) );
  XNOR2_X1 U3154 ( .A(n2490), .B(IR_REG_4__SCAN_IN), .ZN(n4418) );
  MUX2_X1 U3155 ( .A(n4418), .B(DATAI_4_), .S(n3906), .Z(n3073) );
  NAND2_X1 U3156 ( .A1(n3004), .A2(n3073), .ZN(n3848) );
  INV_X1 U3157 ( .A(n3073), .ZN(n3089) );
  NAND2_X1 U3158 ( .A1(n4010), .A2(n3089), .ZN(n3851) );
  NAND2_X1 U3159 ( .A1(n4010), .A2(n3073), .ZN(n2491) );
  OAI21_X2 U3160 ( .B1(n3090), .B2(n3924), .A(n2491), .ZN(n3011) );
  AOI22_X1 U3161 ( .A1(n2484), .A2(REG1_REG_5__SCAN_IN), .B1(n2460), .B2(
        REG0_REG_5__SCAN_IN), .ZN(n2494) );
  AOI21_X1 U3162 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2492) );
  NOR2_X1 U3163 ( .A1(n2492), .A2(n2502), .ZN(n4614) );
  AOI22_X1 U3164 ( .A1(n2670), .A2(n4614), .B1(n2459), .B2(REG2_REG_5__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U3165 ( .A1(n2495), .A2(IR_REG_31__SCAN_IN), .ZN(n2496) );
  MUX2_X1 U3166 ( .A(IR_REG_31__SCAN_IN), .B(n2496), .S(IR_REG_5__SCAN_IN), 
        .Z(n2498) );
  INV_X1 U3167 ( .A(n2517), .ZN(n2497) );
  NAND2_X1 U3168 ( .A1(n2498), .A2(n2497), .ZN(n2976) );
  INV_X1 U3169 ( .A(DATAI_5_), .ZN(n4755) );
  MUX2_X1 U3170 ( .A(n2976), .B(n4755), .S(n2465), .Z(n3126) );
  NAND2_X1 U3171 ( .A1(n3149), .A2(n3126), .ZN(n2499) );
  NAND2_X1 U3172 ( .A1(n3011), .A2(n2499), .ZN(n2501) );
  INV_X1 U3173 ( .A(n3149), .ZN(n4009) );
  NAND2_X1 U3174 ( .A1(n4009), .A2(n3016), .ZN(n2500) );
  OAI21_X1 U3175 ( .B1(n2502), .B2(REG3_REG_6__SCAN_IN), .A(n2510), .ZN(n4520)
         );
  INV_X1 U3176 ( .A(n4520), .ZN(n2503) );
  NAND2_X1 U3177 ( .A1(n2670), .A2(n2503), .ZN(n2507) );
  NAND2_X1 U3178 ( .A1(n2484), .A2(REG1_REG_6__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U3179 ( .A1(n2459), .A2(REG2_REG_6__SCAN_IN), .ZN(n2505) );
  NAND2_X1 U3180 ( .A1(n2460), .A2(REG0_REG_6__SCAN_IN), .ZN(n2504) );
  NAND4_X1 U3181 ( .A1(n2507), .A2(n2506), .A3(n2505), .A4(n2504), .ZN(n4008)
         );
  OR2_X1 U3182 ( .A1(n2517), .A2(n2553), .ZN(n2508) );
  XNOR2_X1 U3183 ( .A(n2508), .B(IR_REG_6__SCAN_IN), .ZN(n3022) );
  MUX2_X1 U3184 ( .A(n3022), .B(DATAI_6_), .S(n2465), .Z(n3146) );
  AND2_X1 U3185 ( .A1(n2510), .A2(n2509), .ZN(n2511) );
  NOR2_X1 U3186 ( .A1(n2521), .A2(n2511), .ZN(n3172) );
  NAND2_X1 U3187 ( .A1(n2670), .A2(n3172), .ZN(n2515) );
  NAND2_X1 U3188 ( .A1(n2484), .A2(REG1_REG_7__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U3189 ( .A1(n2459), .A2(REG2_REG_7__SCAN_IN), .ZN(n2513) );
  NAND2_X1 U3190 ( .A1(n2460), .A2(REG0_REG_7__SCAN_IN), .ZN(n2512) );
  NAND4_X1 U3191 ( .A1(n2515), .A2(n2514), .A3(n2513), .A4(n2512), .ZN(n4007)
         );
  INV_X1 U3192 ( .A(n4007), .ZN(n3206) );
  NAND2_X1 U3193 ( .A1(n2517), .A2(n2516), .ZN(n2541) );
  NAND2_X1 U3194 ( .A1(n2541), .A2(IR_REG_31__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U3195 ( .A1(n2518), .A2(n4843), .ZN(n2527) );
  OR2_X1 U3196 ( .A1(n2518), .A2(n4843), .ZN(n2519) );
  MUX2_X1 U3197 ( .A(n4416), .B(DATAI_7_), .S(n2465), .Z(n3163) );
  NAND2_X1 U3198 ( .A1(n3206), .A2(n3163), .ZN(n2741) );
  NAND2_X1 U3199 ( .A1(n4007), .A2(n3167), .ZN(n3856) );
  NAND2_X1 U3200 ( .A1(n2741), .A2(n3856), .ZN(n3066) );
  NAND2_X1 U3201 ( .A1(n4007), .A2(n3163), .ZN(n2520) );
  NAND2_X1 U3202 ( .A1(n3067), .A2(n2520), .ZN(n3179) );
  OR2_X1 U3203 ( .A1(n2521), .A2(REG3_REG_8__SCAN_IN), .ZN(n2522) );
  AND2_X1 U3204 ( .A1(n2534), .A2(n2522), .ZN(n4513) );
  NAND2_X1 U3205 ( .A1(n2670), .A2(n4513), .ZN(n2526) );
  NAND2_X1 U3206 ( .A1(n2484), .A2(REG1_REG_8__SCAN_IN), .ZN(n2525) );
  NAND2_X1 U3207 ( .A1(n2459), .A2(REG2_REG_8__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U3208 ( .A1(n2460), .A2(REG0_REG_8__SCAN_IN), .ZN(n2523) );
  NAND4_X1 U3209 ( .A1(n2526), .A2(n2525), .A3(n2524), .A4(n2523), .ZN(n4006)
         );
  INV_X1 U32100 ( .A(n4006), .ZN(n3232) );
  NAND2_X1 U32110 ( .A1(n2527), .A2(IR_REG_31__SCAN_IN), .ZN(n2528) );
  XNOR2_X1 U32120 ( .A(n2528), .B(IR_REG_8__SCAN_IN), .ZN(n3465) );
  INV_X1 U32130 ( .A(DATAI_8_), .ZN(n2529) );
  MUX2_X1 U32140 ( .A(n4571), .B(n2529), .S(n2465), .Z(n3207) );
  NAND2_X1 U32150 ( .A1(n3232), .A2(n3207), .ZN(n2530) );
  NAND2_X1 U32160 ( .A1(n3179), .A2(n2530), .ZN(n2532) );
  NAND2_X1 U32170 ( .A1(n4006), .A2(n3201), .ZN(n2531) );
  NAND2_X1 U32180 ( .A1(n2534), .A2(n2533), .ZN(n2535) );
  NAND2_X1 U32190 ( .A1(n2547), .A2(n2535), .ZN(n3238) );
  INV_X1 U32200 ( .A(n3238), .ZN(n2536) );
  NAND2_X1 U32210 ( .A1(n2670), .A2(n2536), .ZN(n2540) );
  NAND2_X1 U32220 ( .A1(n2484), .A2(REG1_REG_9__SCAN_IN), .ZN(n2539) );
  NAND2_X1 U32230 ( .A1(n2460), .A2(REG0_REG_9__SCAN_IN), .ZN(n2538) );
  NAND2_X1 U32240 ( .A1(n2459), .A2(REG2_REG_9__SCAN_IN), .ZN(n2537) );
  NAND4_X1 U32250 ( .A1(n2540), .A2(n2539), .A3(n2538), .A4(n2537), .ZN(n4005)
         );
  NAND2_X1 U32260 ( .A1(n2543), .A2(IR_REG_31__SCAN_IN), .ZN(n2542) );
  MUX2_X1 U32270 ( .A(IR_REG_31__SCAN_IN), .B(n2542), .S(IR_REG_9__SCAN_IN), 
        .Z(n2545) );
  INV_X1 U32280 ( .A(n2564), .ZN(n2544) );
  NAND2_X1 U32290 ( .A1(n2545), .A2(n2544), .ZN(n4448) );
  MUX2_X1 U32300 ( .A(n4569), .B(DATAI_9_), .S(n2465), .Z(n3227) );
  AND2_X1 U32310 ( .A1(n4005), .A2(n3227), .ZN(n2546) );
  NAND2_X1 U32320 ( .A1(n2547), .A2(n4829), .ZN(n2548) );
  AND2_X1 U32330 ( .A1(n2557), .A2(n2548), .ZN(n4506) );
  NAND2_X1 U32340 ( .A1(n2670), .A2(n4506), .ZN(n2552) );
  NAND2_X1 U32350 ( .A1(n2484), .A2(REG1_REG_10__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U32360 ( .A1(n2459), .A2(REG2_REG_10__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U32370 ( .A1(n2460), .A2(REG0_REG_10__SCAN_IN), .ZN(n2549) );
  OR2_X1 U32380 ( .A1(n2564), .A2(n2553), .ZN(n2554) );
  MUX2_X1 U32390 ( .A(n4415), .B(DATAI_10_), .S(n3906), .Z(n3263) );
  NAND2_X1 U32400 ( .A1(n4004), .A2(n3263), .ZN(n2555) );
  NAND2_X1 U32410 ( .A1(n2484), .A2(REG1_REG_11__SCAN_IN), .ZN(n2562) );
  AND2_X1 U32420 ( .A1(n2557), .A2(n2556), .ZN(n2558) );
  NOR2_X1 U32430 ( .A1(n2568), .A2(n2558), .ZN(n3333) );
  NAND2_X1 U32440 ( .A1(n2670), .A2(n3333), .ZN(n2561) );
  NAND2_X1 U32450 ( .A1(n2460), .A2(REG0_REG_11__SCAN_IN), .ZN(n2560) );
  NAND2_X1 U32460 ( .A1(n2459), .A2(REG2_REG_11__SCAN_IN), .ZN(n2559) );
  NAND4_X1 U32470 ( .A1(n2562), .A2(n2561), .A3(n2560), .A4(n2559), .ZN(n4003)
         );
  INV_X1 U32480 ( .A(IR_REG_10__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U32490 ( .A1(n2564), .A2(n2563), .ZN(n2565) );
  NAND2_X1 U32500 ( .A1(n2565), .A2(IR_REG_31__SCAN_IN), .ZN(n2566) );
  NAND2_X1 U32510 ( .A1(n2566), .A2(n4855), .ZN(n2574) );
  OR2_X1 U32520 ( .A1(n2566), .A2(n4855), .ZN(n2567) );
  MUX2_X1 U32530 ( .A(n3462), .B(DATAI_11_), .S(n3906), .Z(n3291) );
  NAND2_X1 U32540 ( .A1(n3400), .A2(n3291), .ZN(n3281) );
  NAND2_X1 U32550 ( .A1(n4003), .A2(n3329), .ZN(n3283) );
  OR2_X1 U32560 ( .A1(n2568), .A2(REG3_REG_12__SCAN_IN), .ZN(n2569) );
  AND2_X1 U32570 ( .A1(n2569), .A2(n2580), .ZN(n3404) );
  NAND2_X1 U32580 ( .A1(n2670), .A2(n3404), .ZN(n2573) );
  NAND2_X1 U32590 ( .A1(n2484), .A2(REG1_REG_12__SCAN_IN), .ZN(n2572) );
  NAND2_X1 U32600 ( .A1(n2459), .A2(REG2_REG_12__SCAN_IN), .ZN(n2571) );
  NAND2_X1 U32610 ( .A1(n2460), .A2(REG0_REG_12__SCAN_IN), .ZN(n2570) );
  NAND4_X1 U32620 ( .A1(n2573), .A2(n2572), .A3(n2571), .A4(n2570), .ZN(n4002)
         );
  NAND2_X1 U32630 ( .A1(n2574), .A2(IR_REG_31__SCAN_IN), .ZN(n2575) );
  XNOR2_X1 U32640 ( .A(n2575), .B(IR_REG_12__SCAN_IN), .ZN(n3472) );
  MUX2_X1 U32650 ( .A(n3472), .B(DATAI_12_), .S(n2465), .Z(n3395) );
  NAND2_X1 U32660 ( .A1(n4002), .A2(n3395), .ZN(n2576) );
  NAND2_X1 U32670 ( .A1(n3274), .A2(n2576), .ZN(n2578) );
  INV_X1 U32680 ( .A(n4002), .ZN(n3432) );
  INV_X1 U32690 ( .A(n3395), .ZN(n3401) );
  NAND2_X1 U32700 ( .A1(n3432), .A2(n3401), .ZN(n2577) );
  NAND2_X1 U32710 ( .A1(n2580), .A2(n2579), .ZN(n2581) );
  AND2_X1 U32720 ( .A1(n2591), .A2(n2581), .ZN(n3437) );
  NAND2_X1 U32730 ( .A1(n2670), .A2(n3437), .ZN(n2585) );
  NAND2_X1 U32740 ( .A1(n2484), .A2(REG1_REG_13__SCAN_IN), .ZN(n2584) );
  NAND2_X1 U32750 ( .A1(n2459), .A2(REG2_REG_13__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U32760 ( .A1(n2460), .A2(REG0_REG_13__SCAN_IN), .ZN(n2582) );
  NOR2_X1 U32770 ( .A1(n2586), .A2(n2553), .ZN(n2587) );
  MUX2_X1 U32780 ( .A(n2553), .B(n2587), .S(IR_REG_13__SCAN_IN), .Z(n2589) );
  OR2_X1 U32790 ( .A1(n2589), .A2(n2626), .ZN(n3459) );
  INV_X1 U32800 ( .A(n3459), .ZN(n4414) );
  MUX2_X1 U32810 ( .A(n4414), .B(DATAI_13_), .S(n2465), .Z(n3311) );
  NOR2_X1 U32820 ( .A1(n4001), .A2(n3311), .ZN(n2590) );
  NAND2_X1 U32830 ( .A1(n2484), .A2(REG1_REG_14__SCAN_IN), .ZN(n2596) );
  AND2_X1 U32840 ( .A1(n2591), .A2(n4826), .ZN(n2592) );
  NOR2_X1 U32850 ( .A1(n2608), .A2(n2592), .ZN(n3508) );
  NAND2_X1 U32860 ( .A1(n2670), .A2(n3508), .ZN(n2595) );
  NAND2_X1 U32870 ( .A1(n2460), .A2(REG0_REG_14__SCAN_IN), .ZN(n2594) );
  NAND2_X1 U32880 ( .A1(n2459), .A2(REG2_REG_14__SCAN_IN), .ZN(n2593) );
  NAND4_X1 U32890 ( .A1(n2596), .A2(n2595), .A3(n2594), .A4(n2593), .ZN(n4000)
         );
  OR2_X1 U32900 ( .A1(n2626), .A2(n2553), .ZN(n2597) );
  XNOR2_X1 U32910 ( .A(n2597), .B(IR_REG_14__SCAN_IN), .ZN(n4059) );
  MUX2_X1 U32920 ( .A(n4059), .B(DATAI_14_), .S(n2465), .Z(n3495) );
  NAND2_X1 U32930 ( .A1(n3822), .A2(n3495), .ZN(n3879) );
  NAND2_X1 U32940 ( .A1(n4000), .A2(n3504), .ZN(n3836) );
  NAND2_X1 U32950 ( .A1(n3822), .A2(n3504), .ZN(n2598) );
  INV_X1 U32960 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2599) );
  XNOR2_X1 U32970 ( .A(n2608), .B(n2599), .ZN(n3830) );
  NAND2_X1 U32980 ( .A1(n2670), .A2(n3830), .ZN(n2603) );
  NAND2_X1 U32990 ( .A1(n2484), .A2(REG1_REG_15__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U33000 ( .A1(n2459), .A2(REG2_REG_15__SCAN_IN), .ZN(n2601) );
  NAND2_X1 U33010 ( .A1(n2460), .A2(REG0_REG_15__SCAN_IN), .ZN(n2600) );
  NAND4_X1 U33020 ( .A1(n2603), .A2(n2602), .A3(n2601), .A4(n2600), .ZN(n3999)
         );
  NAND2_X1 U33030 ( .A1(n2626), .A2(n2624), .ZN(n2604) );
  NAND2_X1 U33040 ( .A1(n2604), .A2(IR_REG_31__SCAN_IN), .ZN(n2605) );
  NAND2_X1 U33050 ( .A1(n2605), .A2(n2623), .ZN(n2614) );
  OR2_X1 U33060 ( .A1(n2605), .A2(n2623), .ZN(n2606) );
  MUX2_X1 U33070 ( .A(n4081), .B(DATAI_15_), .S(n2465), .Z(n3576) );
  NAND2_X1 U33080 ( .A1(n3999), .A2(n3576), .ZN(n2607) );
  AOI21_X1 U33090 ( .B1(n2608), .B2(REG3_REG_15__SCAN_IN), .A(
        REG3_REG_16__SCAN_IN), .ZN(n2609) );
  NOR2_X1 U33100 ( .A1(n2619), .A2(n2609), .ZN(n3749) );
  NAND2_X1 U33110 ( .A1(n2670), .A2(n3749), .ZN(n2613) );
  NAND2_X1 U33120 ( .A1(n2484), .A2(REG1_REG_16__SCAN_IN), .ZN(n2612) );
  NAND2_X1 U33130 ( .A1(n2459), .A2(REG2_REG_16__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U33140 ( .A1(n2460), .A2(REG0_REG_16__SCAN_IN), .ZN(n2610) );
  NAND4_X1 U33150 ( .A1(n2613), .A2(n2612), .A3(n2611), .A4(n2610), .ZN(n3998)
         );
  INV_X1 U33160 ( .A(n3998), .ZN(n3826) );
  NAND2_X1 U33170 ( .A1(n2614), .A2(IR_REG_31__SCAN_IN), .ZN(n2615) );
  XNOR2_X1 U33180 ( .A(n2615), .B(IR_REG_16__SCAN_IN), .ZN(n4563) );
  MUX2_X1 U33190 ( .A(n4563), .B(DATAI_16_), .S(n3906), .Z(n4354) );
  NAND2_X1 U33200 ( .A1(n3826), .A2(n4354), .ZN(n3884) );
  INV_X1 U33210 ( .A(n4354), .ZN(n2616) );
  NAND2_X1 U33220 ( .A1(n3998), .A2(n2616), .ZN(n3885) );
  NAND2_X1 U33230 ( .A1(n3419), .A2(n2617), .ZN(n3418) );
  NAND2_X1 U33240 ( .A1(n3998), .A2(n4354), .ZN(n2618) );
  NAND2_X1 U33250 ( .A1(n3418), .A2(n2618), .ZN(n3516) );
  AOI22_X1 U33260 ( .A1(n2484), .A2(REG1_REG_17__SCAN_IN), .B1(n2460), .B2(
        REG0_REG_17__SCAN_IN), .ZN(n2622) );
  OR2_X1 U33270 ( .A1(n2619), .A2(REG3_REG_17__SCAN_IN), .ZN(n2620) );
  AND2_X1 U33280 ( .A1(n2646), .A2(n2620), .ZN(n3761) );
  AOI22_X1 U33290 ( .A1(n2670), .A2(n3761), .B1(n2459), .B2(
        REG2_REG_17__SCAN_IN), .ZN(n2621) );
  NAND2_X1 U33300 ( .A1(n2626), .A2(n2625), .ZN(n2628) );
  NAND2_X1 U33310 ( .A1(n2628), .A2(IR_REG_31__SCAN_IN), .ZN(n2627) );
  MUX2_X1 U33320 ( .A(IR_REG_31__SCAN_IN), .B(n2627), .S(IR_REG_17__SCAN_IN), 
        .Z(n2630) );
  AND2_X1 U33330 ( .A1(n2630), .A2(n2638), .ZN(n4084) );
  INV_X1 U33340 ( .A(DATAI_17_), .ZN(n4561) );
  MUX2_X1 U33350 ( .A(n4562), .B(n4561), .S(n2465), .Z(n3756) );
  NAND2_X1 U33360 ( .A1(n3799), .A2(n3756), .ZN(n2632) );
  AND2_X1 U33370 ( .A1(n4356), .A2(n3594), .ZN(n2631) );
  XNOR2_X1 U33380 ( .A(n2646), .B(REG3_REG_18__SCAN_IN), .ZN(n3804) );
  NAND2_X1 U33390 ( .A1(n3804), .A2(n2670), .ZN(n2636) );
  NAND2_X1 U33400 ( .A1(n2484), .A2(REG1_REG_18__SCAN_IN), .ZN(n2635) );
  NAND2_X1 U33410 ( .A1(n2460), .A2(REG0_REG_18__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U33420 ( .A1(n2459), .A2(REG2_REG_18__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U33430 ( .A1(n2638), .A2(IR_REG_31__SCAN_IN), .ZN(n2637) );
  MUX2_X1 U33440 ( .A(IR_REG_31__SCAN_IN), .B(n2637), .S(IR_REG_18__SCAN_IN), 
        .Z(n2640) );
  NAND2_X1 U33450 ( .A1(n2640), .A2(n2650), .ZN(n4075) );
  MUX2_X1 U33460 ( .A(n4094), .B(DATAI_18_), .S(n2465), .Z(n3602) );
  NAND2_X1 U33470 ( .A1(n3758), .A2(n3602), .ZN(n3551) );
  INV_X1 U33480 ( .A(n3758), .ZN(n3997) );
  NAND2_X1 U33490 ( .A1(n3997), .A2(n3800), .ZN(n3552) );
  NAND2_X1 U33500 ( .A1(n3551), .A2(n3552), .ZN(n3529) );
  NAND2_X1 U33510 ( .A1(n3526), .A2(n3529), .ZN(n3525) );
  NAND2_X1 U33520 ( .A1(n3758), .A2(n3800), .ZN(n2641) );
  INV_X1 U3353 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4348) );
  NAND2_X1 U33540 ( .A1(n2459), .A2(REG2_REG_19__SCAN_IN), .ZN(n2644) );
  NAND2_X1 U3355 ( .A1(n2460), .A2(REG0_REG_19__SCAN_IN), .ZN(n2643) );
  AND2_X1 U3356 ( .A1(n2644), .A2(n2643), .ZN(n2649) );
  INV_X1 U3357 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2645) );
  INV_X1 U3358 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4709) );
  OAI21_X1 U3359 ( .B1(n2646), .B2(n2645), .A(n4709), .ZN(n2647) );
  NAND2_X1 U3360 ( .A1(n2647), .A2(n2656), .ZN(n3721) );
  OR2_X1 U3361 ( .A1(n3721), .A2(n2443), .ZN(n2648) );
  INV_X1 U3362 ( .A(n2725), .ZN(n2651) );
  NAND2_X1 U3363 ( .A1(n2651), .A2(IR_REG_19__SCAN_IN), .ZN(n2653) );
  INV_X1 U3364 ( .A(IR_REG_19__SCAN_IN), .ZN(n2652) );
  NAND2_X1 U3365 ( .A1(n2725), .A2(n2652), .ZN(n2722) );
  MUX2_X1 U3366 ( .A(n4413), .B(DATAI_19_), .S(n3906), .Z(n3608) );
  NAND2_X1 U3367 ( .A1(n4269), .A2(n3608), .ZN(n2655) );
  NOR2_X1 U3368 ( .A1(n4269), .A2(n3608), .ZN(n2654) );
  AND2_X1 U3369 ( .A1(n2656), .A2(n4875), .ZN(n2658) );
  OR2_X1 U3370 ( .A1(n2658), .A2(n2657), .ZN(n4279) );
  AOI22_X1 U3371 ( .A1(n2459), .A2(REG2_REG_20__SCAN_IN), .B1(n2460), .B2(
        REG0_REG_20__SCAN_IN), .ZN(n2660) );
  NAND2_X1 U3372 ( .A1(n2484), .A2(REG1_REG_20__SCAN_IN), .ZN(n2659) );
  INV_X1 U3373 ( .A(n4333), .ZN(n3729) );
  OR2_X1 U3374 ( .A1(n2662), .A2(REG3_REG_22__SCAN_IN), .ZN(n2663) );
  AND2_X1 U3375 ( .A1(n2678), .A2(n2663), .ZN(n4237) );
  NAND2_X1 U3376 ( .A1(n4237), .A2(n2670), .ZN(n2668) );
  INV_X1 U3377 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4717) );
  NAND2_X1 U3378 ( .A1(n2460), .A2(REG0_REG_22__SCAN_IN), .ZN(n2665) );
  NAND2_X1 U3379 ( .A1(n2459), .A2(REG2_REG_22__SCAN_IN), .ZN(n2664) );
  OAI211_X1 U3380 ( .C1(n2642), .C2(n4717), .A(n2665), .B(n2664), .ZN(n2666)
         );
  INV_X1 U3381 ( .A(n2666), .ZN(n2667) );
  NAND2_X1 U3382 ( .A1(n2668), .A2(n2667), .ZN(n3996) );
  NAND2_X1 U3383 ( .A1(n3996), .A2(n4228), .ZN(n2757) );
  NAND2_X1 U3384 ( .A1(n4209), .A2(n2757), .ZN(n4240) );
  NAND2_X1 U3385 ( .A1(n4241), .A2(n4240), .ZN(n4329) );
  XNOR2_X1 U3386 ( .A(n2678), .B(REG3_REG_23__SCAN_IN), .ZN(n4219) );
  NAND2_X1 U3387 ( .A1(n4219), .A2(n2670), .ZN(n2675) );
  INV_X1 U3388 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4325) );
  NAND2_X1 U3389 ( .A1(n2460), .A2(REG0_REG_23__SCAN_IN), .ZN(n2672) );
  NAND2_X1 U3390 ( .A1(n2459), .A2(REG2_REG_23__SCAN_IN), .ZN(n2671) );
  OAI211_X1 U3391 ( .C1(n2642), .C2(n4325), .A(n2672), .B(n2671), .ZN(n2673)
         );
  INV_X1 U3392 ( .A(n2673), .ZN(n2674) );
  NAND2_X1 U3393 ( .A1(n4319), .A2(n4218), .ZN(n2677) );
  INV_X1 U3394 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3701) );
  INV_X1 U3395 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3769) );
  OAI21_X1 U3396 ( .B1(n2678), .B2(n3701), .A(n3769), .ZN(n2679) );
  AND2_X1 U3397 ( .A1(n2679), .A2(n2689), .ZN(n4194) );
  NAND2_X1 U3398 ( .A1(n4194), .A2(n2670), .ZN(n2684) );
  INV_X1 U3399 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4724) );
  NAND2_X1 U3400 ( .A1(n2460), .A2(REG0_REG_24__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U3401 ( .A1(n2459), .A2(REG2_REG_24__SCAN_IN), .ZN(n2680) );
  OAI211_X1 U3402 ( .C1(n2458), .C2(n4724), .A(n2681), .B(n2680), .ZN(n2682)
         );
  INV_X1 U3403 ( .A(n2682), .ZN(n2683) );
  NAND2_X1 U3404 ( .A1(n4191), .A2(n2685), .ZN(n2688) );
  INV_X1 U3405 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4886) );
  AND2_X1 U3406 ( .A1(n2689), .A2(n4886), .ZN(n2690) );
  NOR2_X1 U3407 ( .A1(n2698), .A2(n2690), .ZN(n4183) );
  NAND2_X1 U3408 ( .A1(n4183), .A2(n2670), .ZN(n2695) );
  INV_X1 U3409 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4313) );
  NAND2_X1 U3410 ( .A1(n2460), .A2(REG0_REG_25__SCAN_IN), .ZN(n2692) );
  NAND2_X1 U3411 ( .A1(n2459), .A2(REG2_REG_25__SCAN_IN), .ZN(n2691) );
  OAI211_X1 U3412 ( .C1(n4313), .C2(n2642), .A(n2692), .B(n2691), .ZN(n2693)
         );
  INV_X1 U3413 ( .A(n2693), .ZN(n2694) );
  NOR2_X1 U3414 ( .A1(n2698), .A2(REG3_REG_26__SCAN_IN), .ZN(n2699) );
  INV_X1 U3415 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4309) );
  NAND2_X1 U3416 ( .A1(n2460), .A2(REG0_REG_26__SCAN_IN), .ZN(n2701) );
  NAND2_X1 U3417 ( .A1(n2459), .A2(REG2_REG_26__SCAN_IN), .ZN(n2700) );
  OAI211_X1 U3418 ( .C1(n2642), .C2(n4309), .A(n2701), .B(n2700), .ZN(n2702)
         );
  INV_X1 U3419 ( .A(n2702), .ZN(n2703) );
  NAND2_X1 U3420 ( .A1(n3906), .A2(DATAI_26_), .ZN(n4162) );
  NOR2_X1 U3421 ( .A1(n4295), .A2(n4303), .ZN(n3948) );
  NOR2_X1 U3422 ( .A1(n2704), .A2(REG3_REG_27__SCAN_IN), .ZN(n2705) );
  INV_X1 U3423 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4301) );
  NAND2_X1 U3424 ( .A1(n2460), .A2(REG0_REG_27__SCAN_IN), .ZN(n2707) );
  NAND2_X1 U3425 ( .A1(n2459), .A2(REG2_REG_27__SCAN_IN), .ZN(n2706) );
  OAI211_X1 U3426 ( .C1(n2172), .C2(n4301), .A(n2707), .B(n2706), .ZN(n2708)
         );
  INV_X1 U3427 ( .A(n2708), .ZN(n2709) );
  AOI21_X1 U3428 ( .B1(n4142), .B2(n2197), .A(n2710), .ZN(n2711) );
  INV_X1 U3429 ( .A(n2711), .ZN(n2812) );
  NAND2_X1 U3430 ( .A1(n2712), .A2(REG3_REG_28__SCAN_IN), .ZN(n4118) );
  INV_X1 U3431 ( .A(n2712), .ZN(n2713) );
  INV_X1 U3432 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3684) );
  NAND2_X1 U3433 ( .A1(n2713), .A2(n3684), .ZN(n2714) );
  NAND2_X1 U3434 ( .A1(n4118), .A2(n2714), .ZN(n3683) );
  NAND2_X1 U3435 ( .A1(n2460), .A2(REG0_REG_28__SCAN_IN), .ZN(n2716) );
  NAND2_X1 U3436 ( .A1(n2459), .A2(REG2_REG_28__SCAN_IN), .ZN(n2715) );
  OAI211_X1 U3437 ( .C1(n2458), .C2(n2807), .A(n2716), .B(n2715), .ZN(n2717)
         );
  INV_X1 U3438 ( .A(n2717), .ZN(n2718) );
  INV_X1 U3439 ( .A(n3903), .ZN(n2720) );
  NAND2_X1 U3440 ( .A1(n4117), .A2(n3685), .ZN(n3897) );
  NAND2_X1 U3441 ( .A1(n2720), .A2(n3897), .ZN(n3954) );
  XNOR2_X1 U3442 ( .A(n2812), .B(n2721), .ZN(n4125) );
  OAI21_X1 U3443 ( .B1(IR_REG_19__SCAN_IN), .B2(IR_REG_20__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2724) );
  NAND2_X1 U3444 ( .A1(n2725), .A2(n2724), .ZN(n2726) );
  NAND2_X1 U3445 ( .A1(n2727), .A2(IR_REG_31__SCAN_IN), .ZN(n2728) );
  XNOR2_X1 U3446 ( .A(n2728), .B(n2428), .ZN(n2774) );
  XNOR2_X1 U3447 ( .A(n2916), .B(n4411), .ZN(n2729) );
  NAND2_X1 U3448 ( .A1(n2729), .A2(n4099), .ZN(n4544) );
  AND2_X1 U3449 ( .A1(n2730), .A2(n4413), .ZN(n2908) );
  MUX2_X1 U3450 ( .A(n2732), .B(n2553), .S(n2731), .Z(n2733) );
  INV_X1 U3451 ( .A(n2733), .ZN(n2734) );
  NAND2_X1 U3452 ( .A1(n2734), .A2(n2207), .ZN(n2947) );
  NAND2_X1 U3453 ( .A1(n4409), .A2(n2938), .ZN(n4358) );
  INV_X1 U3454 ( .A(n4013), .ZN(n2963) );
  NAND2_X1 U3455 ( .A1(n2963), .A2(n2973), .ZN(n3838) );
  OR2_X1 U3456 ( .A1(n2736), .A2(n3838), .ZN(n2737) );
  NAND2_X1 U3457 ( .A1(n2737), .A2(n3842), .ZN(n4534) );
  NAND2_X1 U34580 ( .A1(n4011), .A2(n3001), .ZN(n3844) );
  INV_X1 U34590 ( .A(n3848), .ZN(n2739) );
  OR2_X1 U3460 ( .A1(n3088), .A2(n2739), .ZN(n2740) );
  NAND2_X1 U3461 ( .A1(n2740), .A2(n3851), .ZN(n3012) );
  AND2_X1 U3462 ( .A1(n4009), .A2(n3126), .ZN(n3010) );
  NAND2_X1 U3463 ( .A1(n3149), .A2(n3016), .ZN(n3863) );
  NAND2_X1 U3464 ( .A1(n4008), .A2(n3150), .ZN(n3861) );
  NAND2_X1 U3465 ( .A1(n3166), .A2(n3146), .ZN(n3853) );
  NAND2_X1 U3466 ( .A1(n2742), .A2(n3856), .ZN(n3181) );
  NAND2_X1 U34670 ( .A1(n3232), .A2(n3201), .ZN(n3858) );
  NAND2_X1 U3468 ( .A1(n3181), .A2(n3858), .ZN(n2743) );
  NAND2_X1 U34690 ( .A1(n4006), .A2(n3207), .ZN(n3855) );
  AND2_X1 U3470 ( .A1(n4005), .A2(n2252), .ZN(n3874) );
  INV_X1 U34710 ( .A(n4005), .ZN(n3267) );
  NAND2_X1 U3472 ( .A1(n3267), .A2(n3227), .ZN(n3857) );
  INV_X1 U34730 ( .A(n3263), .ZN(n3268) );
  NAND2_X1 U3474 ( .A1(n4004), .A2(n3268), .ZN(n3870) );
  INV_X1 U34750 ( .A(n4004), .ZN(n3328) );
  NAND2_X1 U3476 ( .A1(n3328), .A2(n3263), .ZN(n3873) );
  NAND2_X1 U34770 ( .A1(n2744), .A2(n3873), .ZN(n3292) );
  NAND2_X1 U3478 ( .A1(n4002), .A2(n3401), .ZN(n3306) );
  NAND2_X1 U34790 ( .A1(n4001), .A2(n3433), .ZN(n2745) );
  NAND2_X1 U3480 ( .A1(n3306), .A2(n2745), .ZN(n2747) );
  INV_X1 U34810 ( .A(n3283), .ZN(n3871) );
  NOR2_X1 U3482 ( .A1(n2747), .A2(n3871), .ZN(n2746) );
  NAND2_X1 U34830 ( .A1(n3432), .A2(n3395), .ZN(n3308) );
  NAND2_X1 U3484 ( .A1(n3281), .A2(n3308), .ZN(n2749) );
  INV_X1 U34850 ( .A(n2747), .ZN(n3876) );
  NOR2_X1 U3486 ( .A1(n4001), .A2(n3433), .ZN(n2748) );
  AOI21_X1 U34870 ( .B1(n2749), .B2(n3876), .A(n2748), .ZN(n3883) );
  NAND2_X1 U3488 ( .A1(n4359), .A2(n3576), .ZN(n3878) );
  NAND2_X1 U34890 ( .A1(n3999), .A2(n3823), .ZN(n3837) );
  NAND2_X1 U3490 ( .A1(n3878), .A2(n3837), .ZN(n3921) );
  NAND2_X1 U34910 ( .A1(n3378), .A2(n3837), .ZN(n3424) );
  NAND2_X1 U3492 ( .A1(n3424), .A2(n3931), .ZN(n3512) );
  NAND2_X1 U34930 ( .A1(n4356), .A2(n3756), .ZN(n3887) );
  AND2_X1 U3494 ( .A1(n3885), .A2(n3887), .ZN(n3959) );
  NAND2_X1 U34950 ( .A1(n3512), .A2(n3959), .ZN(n4267) );
  NAND2_X1 U3496 ( .A1(n3799), .A2(n3594), .ZN(n3528) );
  NAND2_X1 U34970 ( .A1(n3551), .A2(n3528), .ZN(n2752) );
  NAND2_X1 U3498 ( .A1(n4269), .A2(n3715), .ZN(n2750) );
  AND2_X1 U34990 ( .A1(n2750), .A2(n3552), .ZN(n2754) );
  NOR2_X1 U3500 ( .A1(n4269), .A2(n3715), .ZN(n2751) );
  AOI21_X1 U35010 ( .B1(n2752), .B2(n2754), .A(n2751), .ZN(n4265) );
  OR2_X1 U3502 ( .A1(n4333), .A2(n3942), .ZN(n2753) );
  NAND2_X1 U35030 ( .A1(n4267), .A2(n3960), .ZN(n2756) );
  INV_X1 U3504 ( .A(n2754), .ZN(n4266) );
  AND2_X1 U35050 ( .A1(n4333), .A2(n3942), .ZN(n2755) );
  AOI21_X1 U35060 ( .B1(n3960), .B2(n4266), .A(n2755), .ZN(n3963) );
  NAND2_X1 U35070 ( .A1(n2756), .A2(n3963), .ZN(n4247) );
  OR2_X1 U35080 ( .A1(n4226), .A2(n4253), .ZN(n4207) );
  NAND2_X1 U35090 ( .A1(n4247), .A2(n3967), .ZN(n2760) );
  OR2_X1 U35100 ( .A1(n4319), .A2(n3638), .ZN(n3945) );
  AND2_X1 U35110 ( .A1(n3945), .A2(n2757), .ZN(n3895) );
  AND2_X1 U35120 ( .A1(n4226), .A2(n4253), .ZN(n4206) );
  NAND2_X1 U35130 ( .A1(n4209), .A2(n4206), .ZN(n2758) );
  NAND2_X1 U35140 ( .A1(n3895), .A2(n2758), .ZN(n3968) );
  INV_X1 U35150 ( .A(n3968), .ZN(n2759) );
  INV_X1 U35160 ( .A(n3946), .ZN(n2761) );
  NOR2_X1 U35170 ( .A1(n4213), .A2(n4198), .ZN(n3941) );
  OR2_X1 U35180 ( .A1(n4295), .A2(n4162), .ZN(n2762) );
  OR2_X1 U35190 ( .A1(n4316), .A2(n4181), .ZN(n4154) );
  NAND2_X1 U35200 ( .A1(n2762), .A2(n4154), .ZN(n3972) );
  NAND2_X1 U35210 ( .A1(n4316), .A2(n4181), .ZN(n3912) );
  NAND2_X1 U35220 ( .A1(n4213), .A2(n4198), .ZN(n4171) );
  NAND2_X1 U35230 ( .A1(n4295), .A2(n4162), .ZN(n3973) );
  OAI21_X1 U35240 ( .B1(n3972), .B2(n4153), .A(n3973), .ZN(n3899) );
  INV_X1 U35250 ( .A(n3899), .ZN(n2763) );
  XNOR2_X1 U35260 ( .A(n4128), .B(n4294), .ZN(n4141) );
  NAND2_X1 U35270 ( .A1(n4139), .A2(n4141), .ZN(n4138) );
  NOR2_X1 U35280 ( .A1(n4128), .A2(n4147), .ZN(n3902) );
  INV_X1 U35290 ( .A(n3902), .ZN(n2765) );
  NAND2_X1 U35300 ( .A1(n4138), .A2(n2765), .ZN(n2813) );
  XNOR2_X1 U35310 ( .A(n2813), .B(n2721), .ZN(n2768) );
  INV_X1 U35320 ( .A(n2730), .ZN(n4412) );
  NAND2_X1 U35330 ( .A1(n4412), .A2(n2735), .ZN(n2767) );
  NAND2_X1 U35340 ( .A1(n4413), .A2(n4411), .ZN(n2766) );
  NAND2_X1 U35350 ( .A1(n2768), .A2(n4548), .ZN(n4137) );
  OR2_X1 U35360 ( .A1(n4118), .A2(n2443), .ZN(n2773) );
  INV_X1 U35370 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2823) );
  NAND2_X1 U35380 ( .A1(n2459), .A2(REG2_REG_29__SCAN_IN), .ZN(n2770) );
  NAND2_X1 U35390 ( .A1(n2460), .A2(REG0_REG_29__SCAN_IN), .ZN(n2769) );
  OAI211_X1 U35400 ( .C1(n2458), .C2(n2823), .A(n2770), .B(n2769), .ZN(n2771)
         );
  INV_X1 U35410 ( .A(n2771), .ZN(n2772) );
  NAND2_X1 U35420 ( .A1(n2773), .A2(n2772), .ZN(n3908) );
  NAND2_X1 U35430 ( .A1(n2936), .A2(n4412), .ZN(n4229) );
  AOI22_X1 U35440 ( .A1(n3908), .A2(n4355), .B1(n4535), .B2(n4127), .ZN(n2775)
         );
  OAI211_X1 U35450 ( .C1(n4306), .C2(n4358), .A(n4137), .B(n2775), .ZN(n2776)
         );
  AOI21_X1 U35460 ( .B1(n4125), .B2(n4594), .A(n2776), .ZN(n3565) );
  NAND2_X1 U35470 ( .A1(n2792), .A2(n2791), .ZN(n2794) );
  OAI21_X1 U35480 ( .B1(IR_REG_23__SCAN_IN), .B2(IR_REG_24__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2780) );
  NAND2_X1 U35490 ( .A1(n2792), .A2(n2780), .ZN(n2781) );
  NAND2_X1 U35500 ( .A1(n2788), .A2(n2848), .ZN(n2782) );
  MUX2_X1 U35510 ( .A(n2788), .B(n2782), .S(B_REG_SCAN_IN), .Z(n2785) );
  NAND2_X1 U35520 ( .A1(n2783), .A2(IR_REG_31__SCAN_IN), .ZN(n2784) );
  XNOR2_X1 U35530 ( .A(n2784), .B(IR_REG_26__SCAN_IN), .ZN(n2789) );
  INV_X1 U35540 ( .A(D_REG_1__SCAN_IN), .ZN(n2850) );
  NAND2_X1 U35550 ( .A1(n2846), .A2(n2850), .ZN(n2787) );
  INV_X1 U35560 ( .A(n2789), .ZN(n3568) );
  NAND2_X1 U35570 ( .A1(n3568), .A2(n2848), .ZN(n2786) );
  NAND2_X1 U35580 ( .A1(n2787), .A2(n2786), .ZN(n2901) );
  NAND2_X1 U35590 ( .A1(n2730), .A2(n4099), .ZN(n2937) );
  NAND2_X1 U35600 ( .A1(n2937), .A2(n2938), .ZN(n2988) );
  INV_X1 U35610 ( .A(n2788), .ZN(n2790) );
  INV_X1 U35620 ( .A(n2848), .ZN(n4410) );
  NAND3_X1 U35630 ( .A1(n2790), .A2(n4410), .A3(n2789), .ZN(n2915) );
  OR2_X1 U35640 ( .A1(n2792), .A2(n2791), .ZN(n2793) );
  NAND2_X1 U35650 ( .A1(n2794), .A2(n2793), .ZN(n2987) );
  NOR4_X1 U35660 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_31__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2803) );
  NOR4_X1 U35670 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n2802) );
  INV_X1 U35680 ( .A(D_REG_16__SCAN_IN), .ZN(n4747) );
  INV_X1 U35690 ( .A(D_REG_14__SCAN_IN), .ZN(n4749) );
  INV_X1 U35700 ( .A(D_REG_10__SCAN_IN), .ZN(n4753) );
  INV_X1 U35710 ( .A(D_REG_22__SCAN_IN), .ZN(n4752) );
  NAND4_X1 U35720 ( .A1(n4747), .A2(n4749), .A3(n4753), .A4(n4752), .ZN(n2800)
         );
  NOR4_X1 U35730 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2798) );
  NOR4_X1 U35740 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2797) );
  NOR4_X1 U35750 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2796) );
  NOR4_X1 U35760 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2795) );
  NAND4_X1 U35770 ( .A1(n2798), .A2(n2797), .A3(n2796), .A4(n2795), .ZN(n2799)
         );
  NOR4_X1 U35780 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(n2800), 
        .A4(n2799), .ZN(n2801) );
  NAND3_X1 U35790 ( .A1(n2803), .A2(n2802), .A3(n2801), .ZN(n2804) );
  NAND2_X1 U35800 ( .A1(n2846), .A2(n2804), .ZN(n2933) );
  NAND2_X1 U35810 ( .A1(n4592), .A2(n2903), .ZN(n2942) );
  NAND4_X1 U3582 ( .A1(n2901), .A2(n2943), .A3(n2933), .A4(n2942), .ZN(n2827)
         );
  INV_X1 U3583 ( .A(D_REG_0__SCAN_IN), .ZN(n3570) );
  NAND2_X1 U3584 ( .A1(n2846), .A2(n3570), .ZN(n2806) );
  NAND2_X1 U3585 ( .A1(n2788), .A2(n3568), .ZN(n2805) );
  NAND2_X1 U3586 ( .A1(n2806), .A2(n2805), .ZN(n2902) );
  MUX2_X1 U3587 ( .A(n2807), .B(n3565), .S(n4612), .Z(n2811) );
  NOR2_X1 U3588 ( .A1(n4551), .A2(n4552), .ZN(n4550) );
  INV_X1 U3589 ( .A(n4143), .ZN(n2809) );
  INV_X1 U3590 ( .A(n2824), .ZN(n2808) );
  NAND2_X1 U3591 ( .A1(n2811), .A2(n2810), .ZN(U3546) );
  NAND2_X1 U3592 ( .A1(n3906), .A2(DATAI_29_), .ZN(n4115) );
  XNOR2_X1 U3593 ( .A(n3908), .B(n4115), .ZN(n3951) );
  AOI21_X1 U3594 ( .B1(n2813), .B2(n3897), .A(n3903), .ZN(n2814) );
  XOR2_X1 U3595 ( .A(n3951), .B(n2814), .Z(n2821) );
  INV_X1 U3596 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2817) );
  NAND2_X1 U3597 ( .A1(n2459), .A2(REG2_REG_30__SCAN_IN), .ZN(n2816) );
  NAND2_X1 U3598 ( .A1(n2460), .A2(REG0_REG_30__SCAN_IN), .ZN(n2815) );
  OAI211_X1 U3599 ( .C1(n2172), .C2(n2817), .A(n2816), .B(n2815), .ZN(n3995)
         );
  INV_X1 U3600 ( .A(n3995), .ZN(n2820) );
  XNOR2_X1 U3601 ( .A(n2818), .B(IR_REG_27__SCAN_IN), .ZN(n2861) );
  NAND2_X1 U3602 ( .A1(n2861), .A2(B_REG_SCAN_IN), .ZN(n2819) );
  NAND2_X1 U3603 ( .A1(n4355), .A2(n2819), .ZN(n4105) );
  OAI22_X1 U3604 ( .A1(n2821), .A2(n4215), .B1(n2820), .B2(n4105), .ZN(n4121)
         );
  OAI22_X1 U3605 ( .A1(n4298), .A2(n4358), .B1(n4115), .B2(n4229), .ZN(n2822)
         );
  MUX2_X1 U3606 ( .A(n2823), .B(n2828), .S(n4612), .Z(n2826) );
  NAND2_X1 U3607 ( .A1(n2824), .A2(n4115), .ZN(n4289) );
  OAI21_X1 U3608 ( .B1(n2824), .B2(n4115), .A(n4289), .ZN(n4119) );
  NAND2_X1 U3609 ( .A1(n2826), .A2(n2825), .ZN(U3547) );
  INV_X1 U3610 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2829) );
  INV_X1 U3611 ( .A(n2902), .ZN(n2935) );
  NAND2_X1 U3612 ( .A1(n2831), .A2(n2830), .ZN(U3515) );
  INV_X1 U3613 ( .A(n4560), .ZN(n2832) );
  NOR2_X2 U3614 ( .A1(n2915), .A2(n2832), .ZN(U4043) );
  INV_X2 U3615 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3616 ( .A(DATAI_14_), .ZN(n2834) );
  NAND2_X1 U3617 ( .A1(n4059), .A2(STATE_REG_SCAN_IN), .ZN(n2833) );
  OAI21_X1 U3618 ( .B1(STATE_REG_SCAN_IN), .B2(n2834), .A(n2833), .ZN(U3338)
         );
  INV_X1 U3619 ( .A(n3022), .ZN(n2980) );
  INV_X1 U3620 ( .A(DATAI_6_), .ZN(n2835) );
  MUX2_X1 U3621 ( .A(n2980), .B(n2835), .S(U3149), .Z(n2836) );
  INV_X1 U3622 ( .A(n2836), .ZN(U3346) );
  NAND3_X1 U3623 ( .A1(n2296), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n2838) );
  INV_X1 U3624 ( .A(DATAI_31_), .ZN(n4921) );
  OAI22_X1 U3625 ( .A1(n2837), .A2(n2838), .B1(STATE_REG_SCAN_IN), .B2(n4921), 
        .ZN(U3321) );
  INV_X1 U3626 ( .A(DATAI_18_), .ZN(n4918) );
  NAND2_X1 U3627 ( .A1(n4094), .A2(STATE_REG_SCAN_IN), .ZN(n2839) );
  OAI21_X1 U3628 ( .B1(STATE_REG_SCAN_IN), .B2(n4918), .A(n2839), .ZN(U3334)
         );
  INV_X1 U3629 ( .A(DATAI_24_), .ZN(n2840) );
  MUX2_X1 U3630 ( .A(n2840), .B(n2788), .S(STATE_REG_SCAN_IN), .Z(n2841) );
  INV_X1 U3631 ( .A(n2841), .ZN(U3328) );
  INV_X1 U3632 ( .A(DATAI_27_), .ZN(n2843) );
  NAND2_X1 U3633 ( .A1(n2861), .A2(STATE_REG_SCAN_IN), .ZN(n2842) );
  OAI21_X1 U3634 ( .B1(STATE_REG_SCAN_IN), .B2(n2843), .A(n2842), .ZN(U3325)
         );
  INV_X1 U3635 ( .A(DATAI_29_), .ZN(n4777) );
  NAND2_X1 U3636 ( .A1(n2844), .A2(STATE_REG_SCAN_IN), .ZN(n2845) );
  OAI21_X1 U3637 ( .B1(STATE_REG_SCAN_IN), .B2(n4777), .A(n2845), .ZN(U3323)
         );
  INV_X1 U3638 ( .A(n2846), .ZN(n2847) );
  AND2_X1 U3639 ( .A1(n2848), .A2(n4560), .ZN(n2849) );
  AOI22_X1 U3640 ( .A1(n4559), .A2(n2850), .B1(n2849), .B2(n3568), .ZN(U3459)
         );
  INV_X1 U3641 ( .A(n2951), .ZN(n2852) );
  INV_X1 U3642 ( .A(n2987), .ZN(n2851) );
  NAND2_X1 U3643 ( .A1(n2851), .A2(STATE_REG_SCAN_IN), .ZN(n3993) );
  NAND2_X1 U3644 ( .A1(n2852), .A2(n3993), .ZN(n2856) );
  NAND2_X1 U3645 ( .A1(n2938), .A2(n2987), .ZN(n2853) );
  AND2_X1 U3646 ( .A1(n2853), .A2(n2465), .ZN(n2855) );
  INV_X1 U3647 ( .A(n2855), .ZN(n2854) );
  NOR2_X1 U3648 ( .A1(n4498), .A2(U4043), .ZN(U3148) );
  NAND2_X1 U3649 ( .A1(n2856), .A2(n2855), .ZN(n4430) );
  NAND2_X1 U3650 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4018) );
  INV_X1 U3651 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2857) );
  MUX2_X1 U3652 ( .A(REG2_REG_1__SCAN_IN), .B(n2857), .S(n2868), .Z(n2860) );
  NAND2_X1 U3653 ( .A1(n4421), .A2(REG2_REG_1__SCAN_IN), .ZN(n2869) );
  AOI21_X1 U3654 ( .B1(n2868), .B2(n2857), .A(n4018), .ZN(n2858) );
  NAND2_X1 U3655 ( .A1(n2869), .A2(n2858), .ZN(n2870) );
  INV_X1 U3656 ( .A(n2870), .ZN(n2859) );
  INV_X1 U3657 ( .A(n2861), .ZN(n4426) );
  NOR2_X1 U3658 ( .A1(n2947), .A2(n4426), .ZN(n3989) );
  INV_X1 U3659 ( .A(n3989), .ZN(n4019) );
  AOI211_X1 U3660 ( .C1(n4018), .C2(n2860), .A(n2859), .B(n4492), .ZN(n2865)
         );
  NAND2_X1 U3661 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2863) );
  XNOR2_X1 U3662 ( .A(n4421), .B(REG1_REG_1__SCAN_IN), .ZN(n2862) );
  NOR2_X1 U3663 ( .A1(n2862), .A2(n2863), .ZN(n2875) );
  AOI211_X1 U3664 ( .C1(n2863), .C2(n2862), .A(n2875), .B(n4103), .ZN(n2864)
         );
  NOR2_X1 U3665 ( .A1(n2865), .A2(n2864), .ZN(n2867) );
  AOI22_X1 U3666 ( .A1(n4498), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n2866) );
  OAI211_X1 U3667 ( .C1(n2868), .C2(n4505), .A(n2867), .B(n2866), .ZN(U3241)
         );
  NAND2_X1 U3668 ( .A1(n2870), .A2(n2869), .ZN(n4020) );
  INV_X1 U3669 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2871) );
  XNOR2_X1 U3670 ( .A(n4420), .B(n2871), .ZN(n4021) );
  NAND2_X1 U3671 ( .A1(n4020), .A2(n4021), .ZN(n2873) );
  NAND2_X1 U3672 ( .A1(n4420), .A2(REG2_REG_2__SCAN_IN), .ZN(n2872) );
  NAND2_X1 U3673 ( .A1(n2873), .A2(n2872), .ZN(n2889) );
  XNOR2_X1 U3674 ( .A(n2889), .B(n2881), .ZN(n2888) );
  XNOR2_X1 U3675 ( .A(n2888), .B(REG2_REG_3__SCAN_IN), .ZN(n2879) );
  NOR2_X1 U3676 ( .A1(STATE_REG_SCAN_IN), .A2(n2469), .ZN(n3002) );
  NOR2_X1 U3677 ( .A1(n4505), .A2(n2881), .ZN(n2874) );
  AOI211_X1 U3678 ( .C1(n4498), .C2(ADDR_REG_3__SCAN_IN), .A(n3002), .B(n2874), 
        .ZN(n2878) );
  AOI21_X1 U3679 ( .B1(REG1_REG_1__SCAN_IN), .B2(n4421), .A(n2875), .ZN(n4024)
         );
  MUX2_X1 U3680 ( .A(n2442), .B(REG1_REG_2__SCAN_IN), .S(n4420), .Z(n4023) );
  NOR2_X1 U3681 ( .A1(n4024), .A2(n4023), .ZN(n4022) );
  OAI211_X1 U3682 ( .C1(REG1_REG_3__SCAN_IN), .C2(n2876), .A(n4499), .B(n2880), 
        .ZN(n2877) );
  OAI211_X1 U3683 ( .C1(n2879), .C2(n4492), .A(n2878), .B(n2877), .ZN(U3243)
         );
  XOR2_X1 U3684 ( .A(REG1_REG_5__SCAN_IN), .B(n2976), .Z(n2885) );
  AOI211_X1 U3685 ( .C1(n2886), .C2(n2885), .A(n4103), .B(n2981), .ZN(n2900)
         );
  INV_X1 U3686 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2887) );
  MUX2_X1 U3687 ( .A(n2887), .B(REG2_REG_5__SCAN_IN), .S(n2976), .Z(n2896) );
  NAND2_X1 U3688 ( .A1(n2888), .A2(REG2_REG_3__SCAN_IN), .ZN(n2891) );
  NAND2_X1 U3689 ( .A1(n2889), .A2(n4419), .ZN(n2890) );
  INV_X1 U3690 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2892) );
  NAND2_X1 U3691 ( .A1(n2893), .A2(n4418), .ZN(n2894) );
  NAND2_X1 U3692 ( .A1(n2895), .A2(n2896), .ZN(n2978) );
  OAI211_X1 U3693 ( .C1(n2896), .C2(n2895), .A(n4464), .B(n2978), .ZN(n2898)
         );
  INV_X1 U3694 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4770) );
  NOR2_X1 U3695 ( .A1(STATE_REG_SCAN_IN), .A2(n4770), .ZN(n3118) );
  AOI21_X1 U3696 ( .B1(n4498), .B2(ADDR_REG_5__SCAN_IN), .A(n3118), .ZN(n2897)
         );
  OAI211_X1 U3697 ( .C1(n4505), .C2(n2976), .A(n2898), .B(n2897), .ZN(n2899)
         );
  OR2_X1 U3698 ( .A1(n2900), .A2(n2899), .ZN(U3245) );
  NAND2_X1 U3699 ( .A1(n4013), .A2(n3055), .ZN(n3839) );
  AND2_X1 U3700 ( .A1(n3838), .A2(n3839), .ZN(n4575) );
  INV_X1 U3701 ( .A(n2901), .ZN(n2934) );
  NAND4_X1 U3702 ( .A1(n2934), .A2(n2943), .A3(n2902), .A4(n2933), .ZN(n2905)
         );
  AND2_X1 U3703 ( .A1(n2903), .A2(n2951), .ZN(n2904) );
  NAND2_X2 U3704 ( .A1(n2905), .A2(n4615), .ZN(n4245) );
  NOR2_X1 U3705 ( .A1(n2916), .A2(n4099), .ZN(n2906) );
  NAND2_X1 U3706 ( .A1(n4245), .A2(n2906), .ZN(n3304) );
  NAND2_X1 U3707 ( .A1(n2973), .A2(n2936), .ZN(n4573) );
  AOI21_X1 U3708 ( .B1(n4215), .B2(n4544), .A(n4575), .ZN(n2907) );
  AOI21_X1 U3709 ( .B1(n4355), .B2(n2456), .A(n2907), .ZN(n4574) );
  OAI21_X1 U3710 ( .B1(n2908), .B2(n4573), .A(n4574), .ZN(n2912) );
  INV_X1 U3711 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2910) );
  INV_X1 U3712 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2909) );
  OAI22_X1 U3713 ( .A1(n4245), .A2(n2910), .B1(n2909), .B2(n4615), .ZN(n2911)
         );
  AOI21_X1 U3714 ( .B1(n2912), .B2(n4245), .A(n2911), .ZN(n2913) );
  OAI21_X1 U3715 ( .B1(n4575), .B2(n3304), .A(n2913), .ZN(U3290) );
  INV_X1 U3716 ( .A(n2915), .ZN(n2914) );
  OR2_X2 U3717 ( .A1(n2914), .A2(n2916), .ZN(n2922) );
  NAND2_X1 U3718 ( .A1(n4099), .A2(n4411), .ZN(n2944) );
  XNOR2_X1 U3719 ( .A(n2918), .B(n2923), .ZN(n2993) );
  INV_X2 U3720 ( .A(n3145), .ZN(n3678) );
  OAI22_X1 U3721 ( .A1(n2917), .A2(n3679), .B1(n3678), .B2(n2955), .ZN(n2992)
         );
  XNOR2_X1 U3722 ( .A(n2993), .B(n2992), .ZN(n2932) );
  AOI22_X1 U3723 ( .A1(n4013), .A2(n3145), .B1(n2173), .B2(n2973), .ZN(n2920)
         );
  OAI21_X1 U3724 ( .B1(n2457), .B2(n2915), .A(n2920), .ZN(n2970) );
  NAND2_X1 U3725 ( .A1(n2970), .A2(n2971), .ZN(n2969) );
  NAND2_X1 U3726 ( .A1(n2969), .A2(n2921), .ZN(n2962) );
  XNOR2_X1 U3727 ( .A(n2924), .B(n2923), .ZN(n2929) );
  AND2_X1 U3728 ( .A1(n3049), .A2(n3145), .ZN(n2926) );
  INV_X1 U3729 ( .A(n2927), .ZN(n2928) );
  NAND2_X1 U3730 ( .A1(n2961), .A2(n2930), .ZN(n2931) );
  NOR2_X1 U3731 ( .A1(n2931), .A2(n2932), .ZN(n2994) );
  AOI21_X1 U3732 ( .B1(n2932), .B2(n2931), .A(n2994), .ZN(n2959) );
  NAND3_X1 U3733 ( .A1(n2935), .A2(n2934), .A3(n2933), .ZN(n2953) );
  NAND2_X1 U3734 ( .A1(n2937), .A2(n2936), .ZN(n2940) );
  INV_X1 U3735 ( .A(n2938), .ZN(n2939) );
  NAND3_X1 U3736 ( .A1(n2951), .A2(n2940), .A3(n2939), .ZN(n2941) );
  NAND2_X1 U3737 ( .A1(n2953), .A2(n2942), .ZN(n2990) );
  NAND2_X1 U3738 ( .A1(n2990), .A2(n2943), .ZN(n2972) );
  INV_X1 U3739 ( .A(n2944), .ZN(n2945) );
  NAND2_X1 U3740 ( .A1(n2945), .A2(n4560), .ZN(n2946) );
  NOR2_X1 U3741 ( .A1(n2922), .A2(n2946), .ZN(n3990) );
  NAND2_X1 U3742 ( .A1(n3990), .A2(n2947), .ZN(n2948) );
  OR2_X2 U3743 ( .A1(n2953), .A2(n2948), .ZN(n3827) );
  NAND2_X1 U3744 ( .A1(n3990), .A2(n4409), .ZN(n2949) );
  OAI22_X1 U3745 ( .A1(n4539), .A2(n3827), .B1(n3821), .B2(n2950), .ZN(n2957)
         );
  NAND2_X1 U3746 ( .A1(n4535), .A2(n2951), .ZN(n2952) );
  OR2_X1 U3747 ( .A1(n2953), .A2(n2952), .ZN(n2954) );
  NOR2_X1 U3748 ( .A1(n3824), .A2(n2955), .ZN(n2956) );
  AOI211_X1 U3749 ( .C1(REG3_REG_2__SCAN_IN), .C2(n2972), .A(n2957), .B(n2956), 
        .ZN(n2958) );
  OAI21_X1 U3750 ( .B1(n2959), .B2(n3834), .A(n2958), .ZN(U3234) );
  INV_X1 U3751 ( .A(n2972), .ZN(n2968) );
  INV_X1 U3752 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2967) );
  OAI211_X1 U3753 ( .C1(n2960), .C2(n2962), .A(n2961), .B(n3777), .ZN(n2966)
         );
  INV_X1 U3754 ( .A(n3824), .ZN(n3790) );
  OAI22_X1 U3755 ( .A1(n2963), .A2(n3821), .B1(n3827), .B2(n2917), .ZN(n2964)
         );
  AOI21_X1 U3756 ( .B1(n3049), .B2(n3790), .A(n2964), .ZN(n2965) );
  OAI211_X1 U3757 ( .C1(n2968), .C2(n2967), .A(n2966), .B(n2965), .ZN(U3219)
         );
  OAI21_X1 U3758 ( .B1(n2971), .B2(n2970), .A(n2969), .ZN(n4014) );
  AOI22_X1 U3759 ( .A1(n3790), .A2(n2973), .B1(REG3_REG_0__SCAN_IN), .B2(n2972), .ZN(n2975) );
  INV_X1 U3760 ( .A(n3827), .ZN(n3780) );
  NAND2_X1 U3761 ( .A1(n3780), .A2(n2456), .ZN(n2974) );
  OAI211_X1 U3762 ( .C1(n4014), .C2(n3834), .A(n2975), .B(n2974), .ZN(U3229)
         );
  INV_X1 U3763 ( .A(n2976), .ZN(n4417) );
  NAND2_X1 U3764 ( .A1(n4417), .A2(REG2_REG_5__SCAN_IN), .ZN(n2977) );
  NAND2_X1 U3765 ( .A1(n2978), .A2(n2977), .ZN(n3023) );
  XNOR2_X1 U3766 ( .A(n3023), .B(n2980), .ZN(n3025) );
  XOR2_X1 U3767 ( .A(REG2_REG_6__SCAN_IN), .B(n3025), .Z(n2985) );
  INV_X1 U3768 ( .A(REG3_REG_6__SCAN_IN), .ZN(n4750) );
  NOR2_X1 U3769 ( .A1(STATE_REG_SCAN_IN), .A2(n4750), .ZN(n3151) );
  AOI21_X1 U3770 ( .B1(n4498), .B2(ADDR_REG_6__SCAN_IN), .A(n3151), .ZN(n2979)
         );
  OAI21_X1 U3771 ( .B1(n4505), .B2(n2980), .A(n2979), .ZN(n2984) );
  INV_X1 U3772 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3114) );
  AOI211_X1 U3773 ( .C1(n3114), .C2(n2982), .A(n4103), .B(n3020), .ZN(n2983)
         );
  AOI211_X1 U3774 ( .C1(n4464), .C2(n2985), .A(n2984), .B(n2983), .ZN(n2986)
         );
  INV_X1 U3775 ( .A(n2986), .ZN(U3246) );
  AND3_X1 U3776 ( .A1(n2988), .A2(n2987), .A3(n2915), .ZN(n2989) );
  NAND2_X1 U3777 ( .A1(n2990), .A2(n2989), .ZN(n2991) );
  INV_X1 U3778 ( .A(n2992), .ZN(n2996) );
  INV_X1 U3779 ( .A(n2993), .ZN(n2995) );
  AOI21_X1 U3780 ( .B1(n2996), .B2(n2995), .A(n2994), .ZN(n3080) );
  NAND2_X1 U3781 ( .A1(n4011), .A2(n3662), .ZN(n2998) );
  NAND2_X1 U3782 ( .A1(n3042), .A2(n2173), .ZN(n2997) );
  NAND2_X1 U3783 ( .A1(n2998), .A2(n2997), .ZN(n2999) );
  XNOR2_X1 U3784 ( .A(n2999), .B(n2923), .ZN(n3078) );
  OAI22_X1 U3785 ( .A1(n4539), .A2(n3679), .B1(n3001), .B2(n3678), .ZN(n3077)
         );
  XNOR2_X1 U3786 ( .A(n3078), .B(n3077), .ZN(n3079) );
  XNOR2_X1 U3787 ( .A(n3080), .B(n3079), .ZN(n3000) );
  NAND2_X1 U3788 ( .A1(n3000), .A2(n3777), .ZN(n3008) );
  OAI22_X1 U3789 ( .A1(n3001), .A2(n3824), .B1(n2917), .B2(n3821), .ZN(n3006)
         );
  INV_X1 U3790 ( .A(n3002), .ZN(n3003) );
  OAI21_X1 U3791 ( .B1(n3827), .B2(n3004), .A(n3003), .ZN(n3005) );
  NOR2_X1 U3792 ( .A1(n3006), .A2(n3005), .ZN(n3007) );
  OAI211_X1 U3793 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3786), .A(n3008), .B(n3007), 
        .ZN(U3215) );
  INV_X1 U3794 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n4884) );
  NAND2_X1 U3795 ( .A1(n3908), .A2(U4043), .ZN(n3009) );
  OAI21_X1 U3796 ( .B1(U4043), .B2(n4884), .A(n3009), .ZN(U3579) );
  INV_X1 U3797 ( .A(n3010), .ZN(n3850) );
  AND2_X1 U3798 ( .A1(n3850), .A2(n3863), .ZN(n3926) );
  XNOR2_X1 U3799 ( .A(n3011), .B(n3926), .ZN(n4613) );
  XNOR2_X1 U3800 ( .A(n3012), .B(n3926), .ZN(n3015) );
  OAI22_X1 U3801 ( .A1(n3166), .A2(n4538), .B1(n4229), .B2(n3126), .ZN(n3013)
         );
  AOI21_X1 U3802 ( .B1(n4536), .B2(n4010), .A(n3013), .ZN(n3014) );
  OAI21_X1 U3803 ( .B1(n3015), .B2(n4215), .A(n3014), .ZN(n4624) );
  AOI21_X1 U3804 ( .B1(n4613), .B2(n4594), .A(n4624), .ZN(n3019) );
  AOI21_X1 U3805 ( .B1(n3016), .B2(n3086), .A(n3109), .ZN(n4619) );
  INV_X1 U3806 ( .A(n4350), .ZN(n4605) );
  AOI22_X1 U3807 ( .A1(n4619), .A2(n4605), .B1(REG1_REG_5__SCAN_IN), .B2(n4610), .ZN(n3017) );
  OAI21_X1 U3808 ( .B1(n3019), .B2(n4610), .A(n3017), .ZN(U3523) );
  INV_X1 U3809 ( .A(n4404), .ZN(n4587) );
  AOI22_X1 U3810 ( .A1(n4619), .A2(n4587), .B1(REG0_REG_5__SCAN_IN), .B2(n4599), .ZN(n3018) );
  OAI21_X1 U3811 ( .B1(n3019), .B2(n4599), .A(n3018), .ZN(U3477) );
  INV_X1 U3812 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4831) );
  MUX2_X1 U3813 ( .A(REG1_REG_7__SCAN_IN), .B(n4831), .S(n4416), .Z(n3021) );
  XNOR2_X1 U3814 ( .A(n3443), .B(n3021), .ZN(n3031) );
  AND2_X1 U3815 ( .A1(n3023), .A2(n3022), .ZN(n3024) );
  INV_X1 U3816 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4814) );
  MUX2_X1 U3817 ( .A(n4814), .B(REG2_REG_7__SCAN_IN), .S(n4416), .Z(n3026) );
  AOI211_X1 U3818 ( .C1(n3027), .C2(n3026), .A(n4492), .B(n3463), .ZN(n3030)
         );
  INV_X1 U3819 ( .A(n4416), .ZN(n3464) );
  NOR2_X1 U3820 ( .A1(STATE_REG_SCAN_IN), .A2(n2509), .ZN(n3168) );
  AOI21_X1 U3821 ( .B1(n4498), .B2(ADDR_REG_7__SCAN_IN), .A(n3168), .ZN(n3028)
         );
  OAI21_X1 U3822 ( .B1(n4505), .B2(n3464), .A(n3028), .ZN(n3029) );
  AOI211_X1 U3823 ( .C1(n3031), .C2(n4499), .A(n3030), .B(n3029), .ZN(n3032)
         );
  INV_X1 U3824 ( .A(n3032), .ZN(U3247) );
  XNOR2_X1 U3825 ( .A(n3033), .B(n2204), .ZN(n3036) );
  INV_X1 U3826 ( .A(n3036), .ZN(n4529) );
  XNOR2_X1 U3827 ( .A(n3034), .B(n2204), .ZN(n3039) );
  AOI22_X1 U3828 ( .A1(n4010), .A2(n4355), .B1(n4535), .B2(n3042), .ZN(n3035)
         );
  OAI21_X1 U3829 ( .B1(n2917), .B2(n4358), .A(n3035), .ZN(n3038) );
  NOR2_X1 U3830 ( .A1(n3036), .A2(n4544), .ZN(n3037) );
  AOI211_X1 U3831 ( .C1(n3039), .C2(n4548), .A(n3038), .B(n3037), .ZN(n4532)
         );
  INV_X1 U3832 ( .A(n4532), .ZN(n3040) );
  AOI21_X1 U3833 ( .B1(n4592), .B2(n4529), .A(n3040), .ZN(n3045) );
  INV_X1 U3834 ( .A(n4550), .ZN(n3041) );
  AOI21_X1 U3835 ( .B1(n3042), .B2(n3041), .A(n3087), .ZN(n4528) );
  AOI22_X1 U3836 ( .A1(n4528), .A2(n4587), .B1(REG0_REG_3__SCAN_IN), .B2(n4599), .ZN(n3043) );
  OAI21_X1 U3837 ( .B1(n3045), .B2(n4599), .A(n3043), .ZN(U3473) );
  AOI22_X1 U3838 ( .A1(n4528), .A2(n4605), .B1(REG1_REG_3__SCAN_IN), .B2(n4610), .ZN(n3044) );
  OAI21_X1 U3839 ( .B1(n3045), .B2(n4610), .A(n3044), .ZN(U3521) );
  XNOR2_X1 U3840 ( .A(n2736), .B(n3838), .ZN(n3053) );
  OR2_X1 U3841 ( .A1(n2736), .A2(n3046), .ZN(n3047) );
  NAND2_X1 U3842 ( .A1(n3048), .A2(n3047), .ZN(n4580) );
  AOI22_X1 U3843 ( .A1(n4012), .A2(n4355), .B1(n4535), .B2(n3049), .ZN(n3051)
         );
  NAND2_X1 U3844 ( .A1(n4013), .A2(n4536), .ZN(n3050) );
  OAI211_X1 U3845 ( .C1(n4580), .C2(n4544), .A(n3051), .B(n3050), .ZN(n3052)
         );
  AOI21_X1 U3846 ( .B1(n4548), .B2(n3053), .A(n3052), .ZN(n4577) );
  NAND2_X1 U3847 ( .A1(n4245), .A2(n4099), .ZN(n3536) );
  INV_X1 U3848 ( .A(n4361), .ZN(n4579) );
  OAI21_X1 U3849 ( .B1(n3055), .B2(n3054), .A(n4551), .ZN(n4578) );
  INV_X1 U3850 ( .A(n4578), .ZN(n3058) );
  AOI22_X1 U3851 ( .A1(n4557), .A2(REG2_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4549), .ZN(n3056) );
  OAI21_X1 U3852 ( .B1(n4580), .B2(n3304), .A(n3056), .ZN(n3057) );
  AOI21_X1 U3853 ( .B1(n4618), .B2(n3058), .A(n3057), .ZN(n3059) );
  OAI21_X1 U3854 ( .B1(n4577), .B2(n4557), .A(n3059), .ZN(U3289) );
  INV_X1 U3855 ( .A(n3066), .ZN(n3927) );
  XNOR2_X1 U3856 ( .A(n3060), .B(n3927), .ZN(n3063) );
  AOI22_X1 U3857 ( .A1(n4006), .A2(n4355), .B1(n3163), .B2(n4535), .ZN(n3061)
         );
  OAI21_X1 U3858 ( .B1(n3166), .B2(n4358), .A(n3061), .ZN(n3062) );
  AOI21_X1 U3859 ( .B1(n3063), .B2(n4548), .A(n3062), .ZN(n4597) );
  NOR2_X1 U3860 ( .A1(n4245), .A2(n4814), .ZN(n3065) );
  OAI211_X1 U3861 ( .C1(n3111), .C2(n3167), .A(n4361), .B(n3176), .ZN(n4596)
         );
  NOR2_X1 U3862 ( .A1(n4596), .A2(n3536), .ZN(n3064) );
  AOI211_X1 U3863 ( .C1(n4549), .C2(n3172), .A(n3065), .B(n3064), .ZN(n3070)
         );
  OR2_X1 U3864 ( .A1(n2182), .A2(n3066), .ZN(n4595) );
  INV_X1 U3865 ( .A(n4544), .ZN(n3247) );
  NAND2_X1 U3866 ( .A1(n4245), .A2(n3247), .ZN(n3068) );
  NAND3_X1 U3867 ( .A1(n4595), .A2(n3067), .A3(n4251), .ZN(n3069) );
  OAI211_X1 U3868 ( .C1(n4597), .C2(n4557), .A(n3070), .B(n3069), .ZN(U3283)
         );
  INV_X1 U3869 ( .A(n3821), .ZN(n3789) );
  AOI22_X1 U3870 ( .A1(n3790), .A2(n3073), .B1(n3789), .B2(n4011), .ZN(n3071)
         );
  NAND2_X1 U3871 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n4031) );
  OAI211_X1 U3872 ( .C1(n3149), .C2(n3827), .A(n3071), .B(n4031), .ZN(n3084)
         );
  AND2_X1 U3873 ( .A1(n3073), .A2(n3662), .ZN(n3072) );
  AOI21_X1 U3874 ( .B1(n4010), .B2(n3659), .A(n3072), .ZN(n3121) );
  NAND2_X1 U3875 ( .A1(n4010), .A2(n3145), .ZN(n3075) );
  NAND2_X1 U3876 ( .A1(n3073), .A2(n2173), .ZN(n3074) );
  NAND2_X1 U3877 ( .A1(n3075), .A2(n3074), .ZN(n3076) );
  XNOR2_X1 U3878 ( .A(n3076), .B(n2923), .ZN(n3123) );
  XOR2_X1 U3879 ( .A(n3121), .B(n3123), .Z(n3082) );
  AOI211_X1 U3880 ( .C1(n3082), .C2(n3081), .A(n3834), .B(n3124), .ZN(n3083)
         );
  AOI211_X1 U3881 ( .C1(n3831), .C2(n3098), .A(n3084), .B(n3083), .ZN(n3085)
         );
  INV_X1 U3882 ( .A(n3085), .ZN(U3227) );
  OAI211_X1 U3883 ( .C1(n3087), .C2(n3089), .A(n4361), .B(n3086), .ZN(n4589)
         );
  NOR2_X1 U3884 ( .A1(n4589), .A2(n4413), .ZN(n3097) );
  XOR2_X1 U3885 ( .A(n3924), .B(n3088), .Z(n3096) );
  OAI22_X1 U3886 ( .A1(n4539), .A2(n4358), .B1(n3089), .B2(n4229), .ZN(n3094)
         );
  OR2_X1 U3887 ( .A1(n3090), .A2(n3924), .ZN(n3092) );
  NAND2_X1 U3888 ( .A1(n3090), .A2(n3924), .ZN(n3091) );
  NAND2_X1 U3889 ( .A1(n3092), .A2(n3091), .ZN(n3099) );
  NOR2_X1 U3890 ( .A1(n3099), .A2(n4544), .ZN(n3093) );
  AOI211_X1 U3891 ( .C1(n4355), .C2(n4009), .A(n3094), .B(n3093), .ZN(n3095)
         );
  OAI21_X1 U3892 ( .B1(n4215), .B2(n3096), .A(n3095), .ZN(n4590) );
  AOI211_X1 U3893 ( .C1(n4549), .C2(n3098), .A(n3097), .B(n4590), .ZN(n3101)
         );
  INV_X1 U3894 ( .A(n3099), .ZN(n4593) );
  INV_X1 U3895 ( .A(n3304), .ZN(n4553) );
  AOI22_X1 U3896 ( .A1(n4593), .A2(n4553), .B1(REG2_REG_4__SCAN_IN), .B2(n4557), .ZN(n3100) );
  OAI21_X1 U3897 ( .B1(n3101), .B2(n4557), .A(n3100), .ZN(U3286) );
  NAND2_X1 U3898 ( .A1(n3853), .A2(n3861), .ZN(n3933) );
  XOR2_X1 U3899 ( .A(n3102), .B(n3933), .Z(n4524) );
  INV_X1 U3900 ( .A(n4524), .ZN(n3108) );
  XNOR2_X1 U3901 ( .A(n3103), .B(n3933), .ZN(n3106) );
  OAI22_X1 U3902 ( .A1(n3149), .A2(n4358), .B1(n3150), .B2(n4229), .ZN(n3104)
         );
  AOI21_X1 U3903 ( .B1(n4355), .B2(n4007), .A(n3104), .ZN(n3105) );
  OAI21_X1 U3904 ( .B1(n3106), .B2(n4215), .A(n3105), .ZN(n3107) );
  AOI21_X1 U3905 ( .B1(n4524), .B2(n3247), .A(n3107), .ZN(n4527) );
  OAI21_X1 U3906 ( .B1(n4585), .B2(n3108), .A(n4527), .ZN(n3116) );
  NOR2_X1 U3907 ( .A1(n3109), .A2(n3150), .ZN(n3110) );
  OR2_X1 U3908 ( .A1(n3111), .A2(n3110), .ZN(n4522) );
  INV_X1 U3909 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4736) );
  OAI22_X1 U3910 ( .A1(n4522), .A2(n4404), .B1(n4601), .B2(n4736), .ZN(n3112)
         );
  AOI21_X1 U3911 ( .B1(n3116), .B2(n4601), .A(n3112), .ZN(n3113) );
  INV_X1 U3912 ( .A(n3113), .ZN(U3479) );
  OAI22_X1 U3913 ( .A1(n4522), .A2(n4350), .B1(n4612), .B2(n3114), .ZN(n3115)
         );
  AOI21_X1 U3914 ( .B1(n3116), .B2(n4612), .A(n3115), .ZN(n3117) );
  INV_X1 U3915 ( .A(n3117), .ZN(U3524) );
  AOI21_X1 U3916 ( .B1(n3780), .B2(n4008), .A(n3118), .ZN(n3120) );
  NAND2_X1 U3917 ( .A1(n3789), .A2(n4010), .ZN(n3119) );
  OAI211_X1 U3918 ( .C1(n3824), .C2(n3126), .A(n3120), .B(n3119), .ZN(n3130)
         );
  INV_X1 U3919 ( .A(n3121), .ZN(n3122) );
  OAI22_X1 U3920 ( .A1(n3149), .A2(n3678), .B1(n3676), .B2(n3126), .ZN(n3125)
         );
  XNOR2_X1 U3921 ( .A(n3125), .B(n2923), .ZN(n3142) );
  OAI22_X1 U3922 ( .A1(n3149), .A2(n3679), .B1(n3678), .B2(n3126), .ZN(n3143)
         );
  XNOR2_X1 U3923 ( .A(n3142), .B(n3143), .ZN(n3127) );
  AOI211_X1 U3924 ( .C1(n3128), .C2(n3127), .A(n3834), .B(n2205), .ZN(n3129)
         );
  AOI211_X1 U3925 ( .C1(n3831), .C2(n4614), .A(n3130), .B(n3129), .ZN(n3131)
         );
  INV_X1 U3926 ( .A(n3131), .ZN(U3224) );
  AND2_X1 U3927 ( .A1(n2283), .A2(n3857), .ZN(n3917) );
  INV_X1 U3928 ( .A(n3917), .ZN(n3132) );
  XNOR2_X1 U3929 ( .A(n3133), .B(n3132), .ZN(n3134) );
  NAND2_X1 U3930 ( .A1(n3134), .A2(n4548), .ZN(n3215) );
  XNOR2_X1 U3931 ( .A(n3135), .B(n3917), .ZN(n3213) );
  NAND2_X1 U3932 ( .A1(n3213), .A2(n4251), .ZN(n3141) );
  INV_X1 U3933 ( .A(n3136), .ZN(n3240) );
  AOI21_X1 U3934 ( .B1(n3227), .B2(n3177), .A(n3240), .ZN(n3222) );
  NAND2_X1 U3935 ( .A1(n4245), .A2(n4535), .ZN(n4197) );
  NAND2_X1 U3936 ( .A1(n4245), .A2(n4355), .ZN(n4260) );
  INV_X1 U3937 ( .A(n4260), .ZN(n3301) );
  AOI22_X1 U3938 ( .A1(n3301), .A2(n4004), .B1(n4256), .B2(n4006), .ZN(n3137)
         );
  OAI21_X1 U3939 ( .B1(n2252), .B2(n4197), .A(n3137), .ZN(n3139) );
  INV_X1 U3940 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4813) );
  OAI22_X1 U3941 ( .A1(n3238), .A2(n4615), .B1(n4813), .B2(n4245), .ZN(n3138)
         );
  AOI211_X1 U3942 ( .C1(n3222), .C2(n4618), .A(n3139), .B(n3138), .ZN(n3140)
         );
  OAI211_X1 U3943 ( .C1(n4557), .C2(n3215), .A(n3141), .B(n3140), .ZN(U3281)
         );
  OAI22_X1 U3944 ( .A1(n3166), .A2(n3678), .B1(n3676), .B2(n3150), .ZN(n3144)
         );
  XOR2_X1 U3945 ( .A(n2923), .B(n3144), .Z(n3157) );
  AOI22_X1 U3946 ( .A1(n4008), .A2(n3659), .B1(n3662), .B2(n3146), .ZN(n3158)
         );
  INV_X1 U3947 ( .A(n3158), .ZN(n3162) );
  XNOR2_X1 U3948 ( .A(n3157), .B(n3162), .ZN(n3147) );
  XNOR2_X1 U3949 ( .A(n3159), .B(n3147), .ZN(n3148) );
  NAND2_X1 U3950 ( .A1(n3148), .A2(n3777), .ZN(n3156) );
  OAI22_X1 U3951 ( .A1(n3824), .A2(n3150), .B1(n3149), .B2(n3821), .ZN(n3154)
         );
  INV_X1 U3952 ( .A(n3151), .ZN(n3152) );
  OAI21_X1 U3953 ( .B1(n3827), .B2(n3206), .A(n3152), .ZN(n3153) );
  NOR2_X1 U3954 ( .A1(n3154), .A2(n3153), .ZN(n3155) );
  OAI211_X1 U3955 ( .C1(n3786), .C2(n4520), .A(n3156), .B(n3155), .ZN(U3236)
         );
  INV_X1 U3956 ( .A(n3159), .ZN(n3161) );
  AND2_X1 U3957 ( .A1(n3163), .A2(n3662), .ZN(n3164) );
  AOI21_X1 U3958 ( .B1(n4007), .B2(n3659), .A(n3164), .ZN(n3195) );
  OAI22_X1 U3959 ( .A1(n3206), .A2(n3678), .B1(n3676), .B2(n3167), .ZN(n3165)
         );
  XNOR2_X1 U3960 ( .A(n3165), .B(n2923), .ZN(n3193) );
  XOR2_X1 U3961 ( .A(n3195), .B(n3193), .Z(n3196) );
  XNOR2_X1 U3962 ( .A(n3197), .B(n3196), .ZN(n3175) );
  OAI22_X1 U3963 ( .A1(n3824), .A2(n3167), .B1(n3166), .B2(n3821), .ZN(n3171)
         );
  INV_X1 U3964 ( .A(n3168), .ZN(n3169) );
  OAI21_X1 U3965 ( .B1(n3827), .B2(n3232), .A(n3169), .ZN(n3170) );
  NOR2_X1 U3966 ( .A1(n3171), .A2(n3170), .ZN(n3174) );
  NAND2_X1 U3967 ( .A1(n3831), .A2(n3172), .ZN(n3173) );
  OAI211_X1 U3968 ( .C1(n3175), .C2(n3834), .A(n3174), .B(n3173), .ZN(U3210)
         );
  INV_X1 U3969 ( .A(n3176), .ZN(n3178) );
  OAI21_X1 U3970 ( .B1(n3178), .B2(n3207), .A(n3177), .ZN(n4514) );
  AND2_X1 U3971 ( .A1(n3858), .A2(n3855), .ZN(n3914) );
  XNOR2_X1 U3972 ( .A(n3179), .B(n3914), .ZN(n4516) );
  NAND2_X1 U3973 ( .A1(n4516), .A2(n3247), .ZN(n3187) );
  INV_X1 U3974 ( .A(n3914), .ZN(n3180) );
  XNOR2_X1 U3975 ( .A(n3181), .B(n3180), .ZN(n3185) );
  NAND2_X1 U3976 ( .A1(n4005), .A2(n4355), .ZN(n3183) );
  NAND2_X1 U3977 ( .A1(n4007), .A2(n4536), .ZN(n3182) );
  OAI211_X1 U3978 ( .C1(n4229), .C2(n3207), .A(n3183), .B(n3182), .ZN(n3184)
         );
  AOI21_X1 U3979 ( .B1(n3185), .B2(n4548), .A(n3184), .ZN(n3186) );
  AND2_X1 U3980 ( .A1(n3187), .A2(n3186), .ZN(n4519) );
  NAND2_X1 U3981 ( .A1(n4516), .A2(n4592), .ZN(n3188) );
  AND2_X1 U3982 ( .A1(n4519), .A2(n3188), .ZN(n3191) );
  INV_X1 U3983 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4839) );
  MUX2_X1 U3984 ( .A(n3191), .B(n4839), .S(n4610), .Z(n3189) );
  OAI21_X1 U3985 ( .B1(n4514), .B2(n4350), .A(n3189), .ZN(U3526) );
  INV_X1 U3986 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3190) );
  MUX2_X1 U3987 ( .A(n3191), .B(n3190), .S(n4599), .Z(n3192) );
  OAI21_X1 U3988 ( .B1(n4514), .B2(n4404), .A(n3192), .ZN(U3483) );
  INV_X1 U3989 ( .A(n3193), .ZN(n3194) );
  NAND2_X1 U3990 ( .A1(n4006), .A2(n3662), .ZN(n3199) );
  NAND2_X1 U3991 ( .A1(n3201), .A2(n2173), .ZN(n3198) );
  NAND2_X1 U3992 ( .A1(n3199), .A2(n3198), .ZN(n3200) );
  XNOR2_X1 U3993 ( .A(n3200), .B(n3665), .ZN(n3203) );
  AOI22_X1 U3994 ( .A1(n4006), .A2(n3659), .B1(n3201), .B2(n3662), .ZN(n3202)
         );
  NOR2_X1 U3995 ( .A1(n3203), .A2(n3202), .ZN(n3225) );
  NAND2_X1 U3996 ( .A1(n3203), .A2(n3202), .ZN(n3224) );
  INV_X1 U3997 ( .A(n3224), .ZN(n3204) );
  NOR2_X1 U3998 ( .A1(n3225), .A2(n3204), .ZN(n3205) );
  XNOR2_X1 U3999 ( .A(n3226), .B(n3205), .ZN(n3212) );
  OAI22_X1 U4000 ( .A1(n3824), .A2(n3207), .B1(n3206), .B2(n3821), .ZN(n3209)
         );
  NAND2_X1 U4001 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4434) );
  OAI21_X1 U4002 ( .B1(n3827), .B2(n3267), .A(n4434), .ZN(n3208) );
  NOR2_X1 U4003 ( .A1(n3209), .A2(n3208), .ZN(n3211) );
  NAND2_X1 U4004 ( .A1(n3831), .A2(n4513), .ZN(n3210) );
  OAI211_X1 U4005 ( .C1(n3212), .C2(n3834), .A(n3211), .B(n3210), .ZN(U3218)
         );
  NAND2_X1 U4006 ( .A1(n3213), .A2(n4594), .ZN(n3217) );
  AOI22_X1 U4007 ( .A1(n4004), .A2(n4355), .B1(n4535), .B2(n3227), .ZN(n3216)
         );
  NAND2_X1 U4008 ( .A1(n4006), .A2(n4536), .ZN(n3214) );
  NAND4_X1 U4009 ( .A1(n3217), .A2(n3216), .A3(n3215), .A4(n3214), .ZN(n3220)
         );
  MUX2_X1 U4010 ( .A(n3220), .B(REG1_REG_9__SCAN_IN), .S(n4610), .Z(n3218) );
  AOI21_X1 U4011 ( .B1(n4605), .B2(n3222), .A(n3218), .ZN(n3219) );
  INV_X1 U4012 ( .A(n3219), .ZN(U3527) );
  MUX2_X1 U4013 ( .A(n3220), .B(REG0_REG_9__SCAN_IN), .S(n4599), .Z(n3221) );
  AOI21_X1 U4014 ( .B1(n3222), .B2(n4587), .A(n3221), .ZN(n3223) );
  INV_X1 U4015 ( .A(n3223), .ZN(U3485) );
  OAI22_X1 U4016 ( .A1(n3267), .A2(n3679), .B1(n2252), .B2(n3678), .ZN(n3255)
         );
  NAND2_X1 U4017 ( .A1(n4005), .A2(n3662), .ZN(n3229) );
  NAND2_X1 U4018 ( .A1(n3227), .A2(n2173), .ZN(n3228) );
  NAND2_X1 U4019 ( .A1(n3229), .A2(n3228), .ZN(n3230) );
  XNOR2_X1 U4020 ( .A(n3230), .B(n2923), .ZN(n3254) );
  XOR2_X1 U4021 ( .A(n3255), .B(n3254), .Z(n3258) );
  XNOR2_X1 U4022 ( .A(n3259), .B(n3258), .ZN(n3231) );
  NAND2_X1 U4023 ( .A1(n3231), .A2(n3777), .ZN(n3237) );
  OAI22_X1 U4024 ( .A1(n3824), .A2(n2252), .B1(n3232), .B2(n3821), .ZN(n3235)
         );
  NOR2_X1 U4025 ( .A1(STATE_REG_SCAN_IN), .A2(n2533), .ZN(n4450) );
  INV_X1 U4026 ( .A(n4450), .ZN(n3233) );
  OAI21_X1 U4027 ( .B1(n3827), .B2(n3328), .A(n3233), .ZN(n3234) );
  NOR2_X1 U4028 ( .A1(n3235), .A2(n3234), .ZN(n3236) );
  OAI211_X1 U4029 ( .C1(n3786), .C2(n3238), .A(n3237), .B(n3236), .ZN(U3228)
         );
  INV_X1 U4030 ( .A(n3298), .ZN(n3239) );
  OAI21_X1 U4031 ( .B1(n3240), .B2(n3268), .A(n3239), .ZN(n4507) );
  INV_X1 U4032 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3249) );
  NAND2_X1 U4033 ( .A1(n3873), .A2(n3870), .ZN(n3934) );
  XNOR2_X1 U4034 ( .A(n3241), .B(n3934), .ZN(n4509) );
  XNOR2_X1 U4035 ( .A(n3242), .B(n3934), .ZN(n3245) );
  OAI22_X1 U4036 ( .A1(n3267), .A2(n4358), .B1(n3268), .B2(n4229), .ZN(n3243)
         );
  AOI21_X1 U4037 ( .B1(n4355), .B2(n4003), .A(n3243), .ZN(n3244) );
  OAI21_X1 U4038 ( .B1(n3245), .B2(n4215), .A(n3244), .ZN(n3246) );
  AOI21_X1 U4039 ( .B1(n4509), .B2(n3247), .A(n3246), .ZN(n4512) );
  INV_X1 U4040 ( .A(n4512), .ZN(n3248) );
  AOI21_X1 U4041 ( .B1(n4592), .B2(n4509), .A(n3248), .ZN(n3251) );
  MUX2_X1 U4042 ( .A(n3249), .B(n3251), .S(n4601), .Z(n3250) );
  OAI21_X1 U40430 ( .B1(n4507), .B2(n4404), .A(n3250), .ZN(U3487) );
  INV_X1 U4044 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3252) );
  MUX2_X1 U4045 ( .A(n3252), .B(n3251), .S(n4612), .Z(n3253) );
  OAI21_X1 U4046 ( .B1(n4507), .B2(n4350), .A(n3253), .ZN(U3528) );
  INV_X1 U4047 ( .A(n4506), .ZN(n3273) );
  INV_X1 U4048 ( .A(n3254), .ZN(n3257) );
  INV_X1 U4049 ( .A(n3255), .ZN(n3256) );
  AOI22_X1 U4050 ( .A1(n3259), .A2(n3258), .B1(n3257), .B2(n3256), .ZN(n3266)
         );
  NAND2_X1 U4051 ( .A1(n4004), .A2(n3662), .ZN(n3261) );
  NAND2_X1 U4052 ( .A1(n3263), .A2(n2173), .ZN(n3260) );
  NAND2_X1 U4053 ( .A1(n3261), .A2(n3260), .ZN(n3262) );
  XNOR2_X1 U4054 ( .A(n3262), .B(n2923), .ZN(n3322) );
  AND2_X1 U4055 ( .A1(n3263), .A2(n3662), .ZN(n3264) );
  AOI21_X1 U4056 ( .B1(n4004), .B2(n3659), .A(n3264), .ZN(n3323) );
  XNOR2_X1 U4057 ( .A(n3322), .B(n3323), .ZN(n3265) );
  NAND2_X1 U4058 ( .A1(n3266), .A2(n3265), .ZN(n3325) );
  OAI211_X1 U4059 ( .C1(n3266), .C2(n3265), .A(n3325), .B(n3777), .ZN(n3272)
         );
  NAND2_X1 U4060 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4048) );
  INV_X1 U4061 ( .A(n4048), .ZN(n3270) );
  OAI22_X1 U4062 ( .A1(n3824), .A2(n3268), .B1(n3267), .B2(n3821), .ZN(n3269)
         );
  AOI211_X1 U4063 ( .C1(n3780), .C2(n4003), .A(n3270), .B(n3269), .ZN(n3271)
         );
  OAI211_X1 U4064 ( .C1(n3786), .C2(n3273), .A(n3272), .B(n3271), .ZN(U3214)
         );
  AND2_X1 U4065 ( .A1(n3308), .A2(n3306), .ZN(n3915) );
  INV_X1 U4066 ( .A(n3915), .ZN(n3285) );
  XNOR2_X1 U4067 ( .A(n3274), .B(n3285), .ZN(n3346) );
  NAND2_X1 U4068 ( .A1(n3297), .A2(n3395), .ZN(n3275) );
  NAND2_X1 U4069 ( .A1(n3315), .A2(n3275), .ZN(n3357) );
  INV_X1 U4070 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3277) );
  INV_X1 U4071 ( .A(n3404), .ZN(n3276) );
  OAI22_X1 U4072 ( .A1(n4245), .A2(n3277), .B1(n3276), .B2(n4615), .ZN(n3278)
         );
  AOI21_X1 U4073 ( .B1(n3301), .B2(n4001), .A(n3278), .ZN(n3280) );
  INV_X1 U4074 ( .A(n4197), .ZN(n4257) );
  AOI22_X1 U4075 ( .A1(n4257), .A2(n3395), .B1(n4256), .B2(n4003), .ZN(n3279)
         );
  OAI211_X1 U4076 ( .C1(n3357), .C2(n4239), .A(n3280), .B(n3279), .ZN(n3288)
         );
  INV_X1 U4077 ( .A(n3281), .ZN(n3282) );
  OR2_X1 U4078 ( .A1(n3292), .A2(n3282), .ZN(n3284) );
  NAND2_X1 U4079 ( .A1(n3284), .A2(n3283), .ZN(n3309) );
  XNOR2_X1 U4080 ( .A(n3309), .B(n3285), .ZN(n3286) );
  NAND2_X1 U4081 ( .A1(n3286), .A2(n4548), .ZN(n3348) );
  NOR2_X1 U4082 ( .A1(n3348), .A2(n4557), .ZN(n3287) );
  AOI211_X1 U4083 ( .C1(n4251), .C2(n3346), .A(n3288), .B(n3287), .ZN(n3289)
         );
  INV_X1 U4084 ( .A(n3289), .ZN(U3278) );
  AOI21_X1 U4085 ( .B1(n3930), .B2(n3290), .A(n2199), .ZN(n3337) );
  AOI22_X1 U4086 ( .A1(n4004), .A2(n4536), .B1(n3291), .B2(n4535), .ZN(n3295)
         );
  XNOR2_X1 U4087 ( .A(n3292), .B(n3930), .ZN(n3293) );
  NAND2_X1 U4088 ( .A1(n3293), .A2(n4548), .ZN(n3294) );
  OAI211_X1 U4089 ( .C1(n3337), .C2(n4544), .A(n3295), .B(n3294), .ZN(n3339)
         );
  NAND2_X1 U4090 ( .A1(n3339), .A2(n4245), .ZN(n3303) );
  INV_X1 U4091 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3461) );
  INV_X1 U4092 ( .A(n3333), .ZN(n3296) );
  OAI22_X1 U4093 ( .A1(n4245), .A2(n3461), .B1(n3296), .B2(n4615), .ZN(n3300)
         );
  OAI21_X1 U4094 ( .B1(n3298), .B2(n3329), .A(n3297), .ZN(n3345) );
  NOR2_X1 U4095 ( .A1(n3345), .A2(n4239), .ZN(n3299) );
  AOI211_X1 U4096 ( .C1(n3301), .C2(n4002), .A(n3300), .B(n3299), .ZN(n3302)
         );
  OAI211_X1 U4097 ( .C1(n3337), .C2(n3304), .A(n3303), .B(n3302), .ZN(U3279)
         );
  XNOR2_X1 U4098 ( .A(n4001), .B(n3433), .ZN(n3943) );
  XNOR2_X1 U4099 ( .A(n3305), .B(n3943), .ZN(n3371) );
  INV_X1 U4100 ( .A(n3371), .ZN(n3321) );
  INV_X1 U4101 ( .A(n3306), .ZN(n3307) );
  AOI21_X1 U4102 ( .B1(n3309), .B2(n3308), .A(n3307), .ZN(n3310) );
  XNOR2_X1 U4103 ( .A(n3310), .B(n3943), .ZN(n3314) );
  AOI22_X1 U4104 ( .A1(n4000), .A2(n4355), .B1(n4535), .B2(n3311), .ZN(n3313)
         );
  NAND2_X1 U4105 ( .A1(n4002), .A2(n4536), .ZN(n3312) );
  OAI211_X1 U4106 ( .C1(n3314), .C2(n4215), .A(n3313), .B(n3312), .ZN(n3370)
         );
  INV_X1 U4107 ( .A(n3315), .ZN(n3317) );
  INV_X1 U4108 ( .A(n3363), .ZN(n3316) );
  OAI21_X1 U4109 ( .B1(n3317), .B2(n3433), .A(n3316), .ZN(n3376) );
  AOI22_X1 U4110 ( .A1(n4557), .A2(REG2_REG_13__SCAN_IN), .B1(n3437), .B2(
        n4549), .ZN(n3318) );
  OAI21_X1 U4111 ( .B1(n3376), .B2(n4239), .A(n3318), .ZN(n3319) );
  AOI21_X1 U4112 ( .B1(n3370), .B2(n4245), .A(n3319), .ZN(n3320) );
  OAI21_X1 U4113 ( .B1(n4621), .B2(n3321), .A(n3320), .ZN(U3277) );
  INV_X1 U4114 ( .A(n3322), .ZN(n3324) );
  OAI22_X1 U4115 ( .A1(n3400), .A2(n3678), .B1(n3676), .B2(n3329), .ZN(n3326)
         );
  XNOR2_X1 U4116 ( .A(n3326), .B(n2923), .ZN(n3388) );
  OAI22_X1 U4117 ( .A1(n3400), .A2(n3679), .B1(n3678), .B2(n3329), .ZN(n3389)
         );
  INV_X1 U4118 ( .A(n3389), .ZN(n3391) );
  XNOR2_X1 U4119 ( .A(n3388), .B(n3391), .ZN(n3327) );
  XNOR2_X1 U4120 ( .A(n3390), .B(n3327), .ZN(n3336) );
  OAI22_X1 U4121 ( .A1(n3824), .A2(n3329), .B1(n3328), .B2(n3821), .ZN(n3332)
         );
  AND2_X1 U4122 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4461) );
  INV_X1 U4123 ( .A(n4461), .ZN(n3330) );
  OAI21_X1 U4124 ( .B1(n3827), .B2(n3432), .A(n3330), .ZN(n3331) );
  NOR2_X1 U4125 ( .A1(n3332), .A2(n3331), .ZN(n3335) );
  NAND2_X1 U4126 ( .A1(n3831), .A2(n3333), .ZN(n3334) );
  OAI211_X1 U4127 ( .C1(n3336), .C2(n3834), .A(n3335), .B(n3334), .ZN(U3233)
         );
  INV_X1 U4128 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3340) );
  OAI22_X1 U4129 ( .A1(n3337), .A2(n4585), .B1(n3432), .B2(n4538), .ZN(n3338)
         );
  NOR2_X1 U4130 ( .A1(n3339), .A2(n3338), .ZN(n3342) );
  MUX2_X1 U4131 ( .A(n3340), .B(n3342), .S(n4601), .Z(n3341) );
  OAI21_X1 U4132 ( .B1(n3345), .B2(n4404), .A(n3341), .ZN(U3489) );
  INV_X1 U4133 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3343) );
  MUX2_X1 U4134 ( .A(n3343), .B(n3342), .S(n4612), .Z(n3344) );
  OAI21_X1 U4135 ( .B1(n4350), .B2(n3345), .A(n3344), .ZN(U3529) );
  NAND2_X1 U4136 ( .A1(n3346), .A2(n4594), .ZN(n3351) );
  AOI22_X1 U4137 ( .A1(n4001), .A2(n4355), .B1(n4535), .B2(n3395), .ZN(n3347)
         );
  OAI211_X1 U4138 ( .C1(n3400), .C2(n4358), .A(n3348), .B(n3347), .ZN(n3349)
         );
  INV_X1 U4139 ( .A(n3349), .ZN(n3350) );
  NAND2_X1 U4140 ( .A1(n3351), .A2(n3350), .ZN(n3354) );
  MUX2_X1 U4141 ( .A(n3354), .B(REG0_REG_12__SCAN_IN), .S(n4599), .Z(n3352) );
  INV_X1 U4142 ( .A(n3352), .ZN(n3353) );
  OAI21_X1 U4143 ( .B1(n3357), .B2(n4404), .A(n3353), .ZN(U3491) );
  MUX2_X1 U4144 ( .A(n3354), .B(REG1_REG_12__SCAN_IN), .S(n4610), .Z(n3355) );
  INV_X1 U4145 ( .A(n3355), .ZN(n3356) );
  OAI21_X1 U4146 ( .B1(n4350), .B2(n3357), .A(n3356), .ZN(U3530) );
  XNOR2_X1 U4147 ( .A(n3958), .B(n3925), .ZN(n3358) );
  NAND2_X1 U4148 ( .A1(n3358), .A2(n4548), .ZN(n3409) );
  INV_X1 U4149 ( .A(n3359), .ZN(n3361) );
  OR2_X1 U4150 ( .A1(n3359), .A2(n3925), .ZN(n3360) );
  OAI21_X1 U4151 ( .B1(n3361), .B2(n2277), .A(n3360), .ZN(n3411) );
  NAND2_X1 U4152 ( .A1(n3411), .A2(n4251), .ZN(n3369) );
  INV_X1 U4153 ( .A(n3381), .ZN(n3362) );
  OAI21_X1 U4154 ( .B1(n3363), .B2(n3504), .A(n3362), .ZN(n3417) );
  INV_X1 U4155 ( .A(n3417), .ZN(n3367) );
  AOI22_X1 U4156 ( .A1(n4257), .A2(n3495), .B1(n4256), .B2(n4001), .ZN(n3365)
         );
  AOI22_X1 U4157 ( .A1(n4557), .A2(REG2_REG_14__SCAN_IN), .B1(n3508), .B2(
        n4549), .ZN(n3364) );
  OAI211_X1 U4158 ( .C1(n4359), .C2(n4260), .A(n3365), .B(n3364), .ZN(n3366)
         );
  AOI21_X1 U4159 ( .B1(n3367), .B2(n4618), .A(n3366), .ZN(n3368) );
  OAI211_X1 U4160 ( .C1(n4557), .C2(n3409), .A(n3369), .B(n3368), .ZN(U3276)
         );
  INV_X1 U4161 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3452) );
  AOI21_X1 U4162 ( .B1(n4594), .B2(n3371), .A(n3370), .ZN(n3373) );
  MUX2_X1 U4163 ( .A(n3452), .B(n3373), .S(n4612), .Z(n3372) );
  OAI21_X1 U4164 ( .B1(n4350), .B2(n3376), .A(n3372), .ZN(U3531) );
  INV_X1 U4165 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3374) );
  MUX2_X1 U4166 ( .A(n3374), .B(n3373), .S(n4601), .Z(n3375) );
  OAI21_X1 U4167 ( .B1(n3376), .B2(n4404), .A(n3375), .ZN(U3493) );
  AOI21_X1 U4168 ( .B1(n3377), .B2(n3921), .A(n4215), .ZN(n3379) );
  NAND2_X1 U4169 ( .A1(n3379), .A2(n3378), .ZN(n3480) );
  XNOR2_X1 U4170 ( .A(n3380), .B(n3921), .ZN(n3482) );
  NAND2_X1 U4171 ( .A1(n3482), .A2(n4251), .ZN(n3387) );
  OAI21_X1 U4172 ( .B1(n3381), .B2(n3823), .A(n3421), .ZN(n3487) );
  INV_X1 U4173 ( .A(n3487), .ZN(n3385) );
  AOI22_X1 U4174 ( .A1(n4257), .A2(n3576), .B1(n4256), .B2(n4000), .ZN(n3383)
         );
  AOI22_X1 U4175 ( .A1(n4557), .A2(REG2_REG_15__SCAN_IN), .B1(n3830), .B2(
        n4549), .ZN(n3382) );
  OAI211_X1 U4176 ( .C1(n3826), .C2(n4260), .A(n3383), .B(n3382), .ZN(n3384)
         );
  AOI21_X1 U4177 ( .B1(n3385), .B2(n4618), .A(n3384), .ZN(n3386) );
  OAI211_X1 U4178 ( .C1(n4557), .C2(n3480), .A(n3387), .B(n3386), .ZN(U3275)
         );
  NAND2_X1 U4179 ( .A1(n4002), .A2(n3662), .ZN(n3393) );
  NAND2_X1 U4180 ( .A1(n3395), .A2(n2173), .ZN(n3392) );
  NAND2_X1 U4181 ( .A1(n3393), .A2(n3392), .ZN(n3394) );
  XNOR2_X1 U4182 ( .A(n3394), .B(n3665), .ZN(n3398) );
  AND2_X1 U4183 ( .A1(n3395), .A2(n3662), .ZN(n3396) );
  AOI21_X1 U4184 ( .B1(n4002), .B2(n3659), .A(n3396), .ZN(n3397) );
  NOR2_X1 U4185 ( .A1(n3398), .A2(n3397), .ZN(n3428) );
  NOR2_X1 U4186 ( .A1(n3428), .A2(n2206), .ZN(n3399) );
  XNOR2_X1 U4187 ( .A(n3429), .B(n3399), .ZN(n3407) );
  OAI22_X1 U4188 ( .A1(n3824), .A2(n3401), .B1(n3400), .B2(n3821), .ZN(n3403)
         );
  NAND2_X1 U4189 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4466) );
  OAI21_X1 U4190 ( .B1(n3827), .B2(n3503), .A(n4466), .ZN(n3402) );
  NOR2_X1 U4191 ( .A1(n3403), .A2(n3402), .ZN(n3406) );
  NAND2_X1 U4192 ( .A1(n3831), .A2(n3404), .ZN(n3405) );
  OAI211_X1 U4193 ( .C1(n3407), .C2(n3834), .A(n3406), .B(n3405), .ZN(U3221)
         );
  INV_X1 U4194 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3412) );
  AOI22_X1 U4195 ( .A1(n3999), .A2(n4355), .B1(n3495), .B2(n4535), .ZN(n3408)
         );
  OAI211_X1 U4196 ( .C1(n3503), .C2(n4358), .A(n3409), .B(n3408), .ZN(n3410)
         );
  AOI21_X1 U4197 ( .B1(n3411), .B2(n4594), .A(n3410), .ZN(n3414) );
  MUX2_X1 U4198 ( .A(n3412), .B(n3414), .S(n4612), .Z(n3413) );
  OAI21_X1 U4199 ( .B1(n4350), .B2(n3417), .A(n3413), .ZN(U3532) );
  INV_X1 U4200 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3415) );
  MUX2_X1 U4201 ( .A(n3415), .B(n3414), .S(n4601), .Z(n3416) );
  OAI21_X1 U4202 ( .B1(n3417), .B2(n4404), .A(n3416), .ZN(U3495) );
  OAI21_X1 U4203 ( .B1(n3419), .B2(n2617), .A(n3418), .ZN(n4366) );
  INV_X1 U4204 ( .A(n3420), .ZN(n3518) );
  AOI21_X1 U4205 ( .B1(n4354), .B2(n3421), .A(n3518), .ZN(n4362) );
  AOI22_X1 U4206 ( .A1(n4257), .A2(n4354), .B1(n4256), .B2(n3999), .ZN(n3423)
         );
  AOI22_X1 U4207 ( .A1(n4557), .A2(REG2_REG_16__SCAN_IN), .B1(n3749), .B2(
        n4549), .ZN(n3422) );
  OAI211_X1 U4208 ( .C1(n3799), .C2(n4260), .A(n3423), .B(n3422), .ZN(n3426)
         );
  OAI211_X1 U4209 ( .C1(n3424), .C2(n3931), .A(n3512), .B(n4548), .ZN(n4363)
         );
  NOR2_X1 U4210 ( .A1(n4363), .A2(n4557), .ZN(n3425) );
  AOI211_X1 U4211 ( .C1(n4362), .C2(n4618), .A(n3426), .B(n3425), .ZN(n3427)
         );
  OAI21_X1 U4212 ( .B1(n4366), .B2(n4621), .A(n3427), .ZN(U3274) );
  OAI22_X1 U4213 ( .A1(n3503), .A2(n3678), .B1(n3676), .B2(n3433), .ZN(n3430)
         );
  XOR2_X1 U4214 ( .A(n2923), .B(n3430), .Z(n3488) );
  INV_X1 U4215 ( .A(n3488), .ZN(n3490) );
  OAI22_X1 U4216 ( .A1(n3503), .A2(n3679), .B1(n2922), .B2(n3433), .ZN(n3491)
         );
  XNOR2_X1 U4217 ( .A(n3490), .B(n3491), .ZN(n3431) );
  XNOR2_X1 U4218 ( .A(n3489), .B(n3431), .ZN(n3440) );
  OAI22_X1 U4219 ( .A1(n3824), .A2(n3433), .B1(n3432), .B2(n3821), .ZN(n3436)
         );
  AND2_X1 U4220 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n3456) );
  INV_X1 U4221 ( .A(n3456), .ZN(n3434) );
  OAI21_X1 U4222 ( .B1(n3827), .B2(n3822), .A(n3434), .ZN(n3435) );
  NOR2_X1 U4223 ( .A1(n3436), .A2(n3435), .ZN(n3439) );
  NAND2_X1 U4224 ( .A1(n3831), .A2(n3437), .ZN(n3438) );
  OAI211_X1 U4225 ( .C1(n3440), .C2(n3834), .A(n3439), .B(n3438), .ZN(U3231)
         );
  NAND2_X1 U4226 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3462), .ZN(n3449) );
  INV_X1 U4227 ( .A(n3462), .ZN(n4568) );
  AOI22_X1 U4228 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3462), .B1(n4568), .B2(
        n3343), .ZN(n4454) );
  INV_X1 U4229 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3441) );
  AOI22_X1 U4230 ( .A1(n4569), .A2(REG1_REG_9__SCAN_IN), .B1(n3441), .B2(n4448), .ZN(n4442) );
  NOR2_X1 U4231 ( .A1(n4416), .A2(REG1_REG_7__SCAN_IN), .ZN(n3442) );
  OAI22_X1 U4232 ( .A1(n3443), .A2(n3442), .B1(n4831), .B2(n3464), .ZN(n3444)
         );
  NAND2_X1 U4233 ( .A1(n3444), .A2(n3465), .ZN(n3445) );
  XNOR2_X1 U4234 ( .A(n3444), .B(n4571), .ZN(n4437) );
  NAND2_X1 U4235 ( .A1(n4569), .A2(REG1_REG_9__SCAN_IN), .ZN(n3446) );
  NAND2_X1 U4236 ( .A1(n3447), .A2(n4415), .ZN(n3448) );
  NAND2_X1 U4237 ( .A1(n3472), .A2(n3450), .ZN(n3451) );
  INV_X1 U4238 ( .A(n3472), .ZN(n4567) );
  XNOR2_X1 U4239 ( .A(n3450), .B(n4567), .ZN(n4470) );
  NAND2_X1 U4240 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4470), .ZN(n4469) );
  NOR2_X1 U4241 ( .A1(n3459), .A2(n3452), .ZN(n3453) );
  AOI21_X1 U4242 ( .B1(n3452), .B2(n3459), .A(n3453), .ZN(n3454) );
  OAI211_X1 U4243 ( .C1(n3455), .C2(n3454), .A(n4058), .B(n4499), .ZN(n3458)
         );
  AOI21_X1 U4244 ( .B1(n4498), .B2(ADDR_REG_13__SCAN_IN), .A(n3456), .ZN(n3457) );
  OAI211_X1 U4245 ( .C1(n4505), .C2(n3459), .A(n3458), .B(n3457), .ZN(n3478)
         );
  INV_X1 U4246 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4816) );
  NOR2_X1 U4247 ( .A1(n3459), .A2(n4816), .ZN(n4053) );
  NAND2_X1 U4248 ( .A1(n3459), .A2(n4816), .ZN(n4052) );
  INV_X1 U4249 ( .A(n4052), .ZN(n3460) );
  NOR2_X1 U4250 ( .A1(n4053), .A2(n3460), .ZN(n3476) );
  NAND2_X1 U4251 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3462), .ZN(n3471) );
  AOI22_X1 U4252 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3462), .B1(n4568), .B2(
        n3461), .ZN(n4457) );
  NAND2_X1 U4253 ( .A1(n4569), .A2(REG2_REG_9__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4254 ( .A1(n4569), .A2(REG2_REG_9__SCAN_IN), .B1(n4813), .B2(n4448), .ZN(n4445) );
  NAND2_X1 U4255 ( .A1(n3465), .A2(n3466), .ZN(n3467) );
  XNOR2_X1 U4256 ( .A(n3466), .B(n4571), .ZN(n4432) );
  NAND2_X1 U4257 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4432), .ZN(n4431) );
  NAND2_X1 U4258 ( .A1(n3469), .A2(n4415), .ZN(n3470) );
  NAND2_X1 U4259 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4046), .ZN(n4045) );
  NAND2_X1 U4260 ( .A1(n3470), .A2(n4045), .ZN(n4456) );
  NAND2_X1 U4261 ( .A1(n4457), .A2(n4456), .ZN(n4455) );
  NAND2_X1 U4262 ( .A1(n3471), .A2(n4455), .ZN(n3473) );
  NAND2_X1 U4263 ( .A1(n3472), .A2(n3473), .ZN(n3474) );
  OAI21_X1 U4264 ( .B1(n3476), .B2(n4054), .A(n4464), .ZN(n3475) );
  AOI21_X1 U4265 ( .B1(n3476), .B2(n4054), .A(n3475), .ZN(n3477) );
  OR2_X1 U4266 ( .A1(n3478), .A2(n3477), .ZN(U3253) );
  INV_X1 U4267 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4268 ( .A1(n3998), .A2(n4355), .B1(n4535), .B2(n3576), .ZN(n3479)
         );
  OAI211_X1 U4269 ( .C1(n3822), .C2(n4358), .A(n3480), .B(n3479), .ZN(n3481)
         );
  AOI21_X1 U4270 ( .B1(n3482), .B2(n4594), .A(n3481), .ZN(n3485) );
  MUX2_X1 U4271 ( .A(n3483), .B(n3485), .S(n4601), .Z(n3484) );
  OAI21_X1 U4272 ( .B1(n3487), .B2(n4404), .A(n3484), .ZN(U3497) );
  MUX2_X1 U4273 ( .A(n4833), .B(n3485), .S(n4612), .Z(n3486) );
  OAI21_X1 U4274 ( .B1(n4350), .B2(n3487), .A(n3486), .ZN(U3533) );
  NAND2_X1 U4275 ( .A1(n4000), .A2(n3662), .ZN(n3493) );
  NAND2_X1 U4276 ( .A1(n3495), .A2(n2173), .ZN(n3492) );
  NAND2_X1 U4277 ( .A1(n3493), .A2(n3492), .ZN(n3494) );
  XNOR2_X1 U4278 ( .A(n3494), .B(n2923), .ZN(n3501) );
  INV_X1 U4279 ( .A(n3501), .ZN(n3499) );
  NAND2_X1 U4280 ( .A1(n4000), .A2(n2925), .ZN(n3497) );
  NAND2_X1 U4281 ( .A1(n3495), .A2(n3662), .ZN(n3496) );
  NAND2_X1 U4282 ( .A1(n3497), .A2(n3496), .ZN(n3500) );
  INV_X1 U4283 ( .A(n3500), .ZN(n3498) );
  NAND2_X1 U4284 ( .A1(n3499), .A2(n3498), .ZN(n3573) );
  NAND2_X1 U4285 ( .A1(n3501), .A2(n3500), .ZN(n3571) );
  NAND2_X1 U4286 ( .A1(n3573), .A2(n3571), .ZN(n3502) );
  XNOR2_X1 U4287 ( .A(n3572), .B(n3502), .ZN(n3511) );
  OAI22_X1 U4288 ( .A1(n3824), .A2(n3504), .B1(n3503), .B2(n3821), .ZN(n3507)
         );
  NOR2_X1 U4289 ( .A1(n4826), .A2(STATE_REG_SCAN_IN), .ZN(n4061) );
  INV_X1 U4290 ( .A(n4061), .ZN(n3505) );
  OAI21_X1 U4291 ( .B1(n3827), .B2(n4359), .A(n3505), .ZN(n3506) );
  NOR2_X1 U4292 ( .A1(n3507), .A2(n3506), .ZN(n3510) );
  NAND2_X1 U4293 ( .A1(n3831), .A2(n3508), .ZN(n3509) );
  OAI211_X1 U4294 ( .C1(n3511), .C2(n3834), .A(n3510), .B(n3509), .ZN(U3212)
         );
  NAND2_X1 U4295 ( .A1(n3512), .A2(n3885), .ZN(n3514) );
  AND2_X1 U4296 ( .A1(n3528), .A2(n3887), .ZN(n3916) );
  INV_X1 U4297 ( .A(n3916), .ZN(n3513) );
  XNOR2_X1 U4298 ( .A(n3514), .B(n3513), .ZN(n3515) );
  NAND2_X1 U4299 ( .A1(n3515), .A2(n4548), .ZN(n3541) );
  XNOR2_X1 U4300 ( .A(n3516), .B(n3916), .ZN(n3543) );
  NAND2_X1 U4301 ( .A1(n3543), .A2(n4251), .ZN(n3524) );
  INV_X1 U4302 ( .A(n3534), .ZN(n3517) );
  OAI21_X1 U4303 ( .B1(n3518), .B2(n3756), .A(n3517), .ZN(n3549) );
  INV_X1 U4304 ( .A(n3549), .ZN(n3522) );
  AOI22_X1 U4305 ( .A1(n4257), .A2(n3594), .B1(n4256), .B2(n3998), .ZN(n3520)
         );
  AOI22_X1 U4306 ( .A1(n4557), .A2(REG2_REG_17__SCAN_IN), .B1(n3761), .B2(
        n4549), .ZN(n3519) );
  OAI211_X1 U4307 ( .C1(n3758), .C2(n4260), .A(n3520), .B(n3519), .ZN(n3521)
         );
  AOI21_X1 U4308 ( .B1(n3522), .B2(n4618), .A(n3521), .ZN(n3523) );
  OAI211_X1 U4309 ( .C1(n4557), .C2(n3541), .A(n3524), .B(n3523), .ZN(U3273)
         );
  OAI21_X1 U4310 ( .B1(n3526), .B2(n3529), .A(n3525), .ZN(n3527) );
  INV_X1 U4311 ( .A(n3527), .ZN(n4353) );
  NAND2_X1 U4312 ( .A1(n4267), .A2(n3528), .ZN(n3554) );
  INV_X1 U4313 ( .A(n3529), .ZN(n3932) );
  XNOR2_X1 U4314 ( .A(n3554), .B(n3932), .ZN(n3532) );
  AOI22_X1 U4315 ( .A1(n4269), .A2(n4355), .B1(n3602), .B2(n4535), .ZN(n3530)
         );
  OAI21_X1 U4316 ( .B1(n3799), .B2(n4358), .A(n3530), .ZN(n3531) );
  AOI21_X1 U4317 ( .B1(n3532), .B2(n4548), .A(n3531), .ZN(n4352) );
  INV_X1 U4318 ( .A(n4352), .ZN(n3538) );
  INV_X1 U4319 ( .A(n3559), .ZN(n3533) );
  OAI211_X1 U4320 ( .C1(n3534), .C2(n3800), .A(n3533), .B(n4361), .ZN(n4351)
         );
  AOI22_X1 U4321 ( .A1(n4557), .A2(REG2_REG_18__SCAN_IN), .B1(n3804), .B2(
        n4549), .ZN(n3535) );
  OAI21_X1 U4322 ( .B1(n4351), .B2(n3536), .A(n3535), .ZN(n3537) );
  AOI21_X1 U4323 ( .B1(n3538), .B2(n4245), .A(n3537), .ZN(n3539) );
  OAI21_X1 U4324 ( .B1(n4353), .B2(n4621), .A(n3539), .ZN(U3272) );
  AOI22_X1 U4325 ( .A1(n3998), .A2(n4536), .B1(n3594), .B2(n4535), .ZN(n3540)
         );
  OAI211_X1 U4326 ( .C1(n3758), .C2(n4538), .A(n3541), .B(n3540), .ZN(n3542)
         );
  AOI21_X1 U4327 ( .B1(n3543), .B2(n4594), .A(n3542), .ZN(n3547) );
  INV_X1 U4328 ( .A(REG0_REG_17__SCAN_IN), .ZN(n3544) );
  MUX2_X1 U4329 ( .A(n3547), .B(n3544), .S(n4599), .Z(n3545) );
  OAI21_X1 U4330 ( .B1(n3549), .B2(n4404), .A(n3545), .ZN(U3501) );
  INV_X1 U4331 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3546) );
  MUX2_X1 U4332 ( .A(n3547), .B(n3546), .S(n4610), .Z(n3548) );
  OAI21_X1 U4333 ( .B1(n4350), .B2(n3549), .A(n3548), .ZN(U3535) );
  XNOR2_X1 U4334 ( .A(n4269), .B(n3715), .ZN(n3944) );
  XNOR2_X1 U4335 ( .A(n3550), .B(n3944), .ZN(n4347) );
  INV_X1 U4336 ( .A(n4347), .ZN(n3564) );
  INV_X1 U4337 ( .A(n3551), .ZN(n3553) );
  OAI21_X1 U4338 ( .B1(n3554), .B2(n3553), .A(n3552), .ZN(n3555) );
  XOR2_X1 U4339 ( .A(n3944), .B(n3555), .Z(n3558) );
  OAI22_X1 U4340 ( .A1(n3729), .A2(n4538), .B1(n4229), .B2(n3715), .ZN(n3556)
         );
  AOI21_X1 U4341 ( .B1(n4536), .B2(n3997), .A(n3556), .ZN(n3557) );
  OAI21_X1 U4342 ( .B1(n3558), .B2(n4215), .A(n3557), .ZN(n4346) );
  OAI21_X1 U4343 ( .B1(n3559), .B2(n3715), .A(n4278), .ZN(n4405) );
  NOR2_X1 U4344 ( .A1(n4405), .A2(n4239), .ZN(n3562) );
  INV_X1 U4345 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3560) );
  OAI22_X1 U4346 ( .A1(n4245), .A2(n3560), .B1(n3721), .B2(n4615), .ZN(n3561)
         );
  AOI211_X1 U4347 ( .C1(n4346), .C2(n4245), .A(n3562), .B(n3561), .ZN(n3563)
         );
  OAI21_X1 U4348 ( .B1(n3564), .B2(n4621), .A(n3563), .ZN(U3271) );
  INV_X1 U4349 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3566) );
  MUX2_X1 U4350 ( .A(n3566), .B(n3565), .S(n4601), .Z(n3567) );
  OAI21_X1 U4351 ( .B1(n4126), .B2(n4404), .A(n3567), .ZN(U3514) );
  AND2_X1 U4352 ( .A1(n3568), .A2(n4560), .ZN(n3569) );
  AOI22_X1 U4353 ( .A1(n4559), .A2(n3570), .B1(n3569), .B2(n2788), .ZN(U3458)
         );
  NAND2_X1 U4354 ( .A1(n3572), .A2(n3571), .ZN(n3574) );
  NAND2_X1 U4355 ( .A1(n3574), .A2(n3573), .ZN(n3579) );
  OAI22_X1 U4356 ( .A1(n4359), .A2(n3678), .B1(n3676), .B2(n3823), .ZN(n3575)
         );
  XOR2_X1 U4357 ( .A(n2923), .B(n3575), .Z(n3580) );
  NAND2_X1 U4358 ( .A1(n3579), .A2(n3580), .ZN(n3743) );
  NAND2_X1 U4359 ( .A1(n3999), .A2(n2925), .ZN(n3578) );
  NAND2_X1 U4360 ( .A1(n3576), .A2(n3662), .ZN(n3577) );
  NAND2_X1 U4361 ( .A1(n3578), .A2(n3577), .ZN(n3820) );
  INV_X1 U4362 ( .A(n3579), .ZN(n3582) );
  INV_X1 U4363 ( .A(n3580), .ZN(n3581) );
  NAND2_X1 U4364 ( .A1(n3998), .A2(n3662), .ZN(n3584) );
  NAND2_X1 U4365 ( .A1(n4354), .A2(n2173), .ZN(n3583) );
  NAND2_X1 U4366 ( .A1(n3584), .A2(n3583), .ZN(n3585) );
  XNOR2_X1 U4367 ( .A(n3585), .B(n2923), .ZN(n3589) );
  NAND2_X1 U4368 ( .A1(n3998), .A2(n3659), .ZN(n3587) );
  NAND2_X1 U4369 ( .A1(n4354), .A2(n3662), .ZN(n3586) );
  NAND2_X1 U4370 ( .A1(n3587), .A2(n3586), .ZN(n3588) );
  NOR2_X1 U4371 ( .A1(n3589), .A2(n3588), .ZN(n3591) );
  AOI21_X1 U4372 ( .B1(n3589), .B2(n3588), .A(n3591), .ZN(n3746) );
  INV_X1 U4373 ( .A(n3591), .ZN(n3592) );
  OAI22_X1 U4374 ( .A1(n3799), .A2(n3678), .B1(n3676), .B2(n3756), .ZN(n3593)
         );
  XNOR2_X1 U4375 ( .A(n3593), .B(n2923), .ZN(n3597) );
  OR2_X1 U4376 ( .A1(n3799), .A2(n3679), .ZN(n3596) );
  NAND2_X1 U4377 ( .A1(n3594), .A2(n3662), .ZN(n3595) );
  NAND2_X1 U4378 ( .A1(n3596), .A2(n3595), .ZN(n3598) );
  NAND2_X1 U4379 ( .A1(n3597), .A2(n3598), .ZN(n3754) );
  INV_X1 U4380 ( .A(n3597), .ZN(n3600) );
  INV_X1 U4381 ( .A(n3598), .ZN(n3599) );
  NAND2_X1 U4382 ( .A1(n3600), .A2(n3599), .ZN(n3753) );
  OAI22_X1 U4383 ( .A1(n3758), .A2(n3678), .B1(n3676), .B2(n3800), .ZN(n3601)
         );
  XNOR2_X1 U4384 ( .A(n3601), .B(n3665), .ZN(n3797) );
  OR2_X1 U4385 ( .A1(n3758), .A2(n3679), .ZN(n3604) );
  NAND2_X1 U4386 ( .A1(n3602), .A2(n3662), .ZN(n3603) );
  NAND2_X1 U4387 ( .A1(n4269), .A2(n3662), .ZN(n3606) );
  NAND2_X1 U4388 ( .A1(n3608), .A2(n2173), .ZN(n3605) );
  NAND2_X1 U4389 ( .A1(n3606), .A2(n3605), .ZN(n3607) );
  XNOR2_X1 U4390 ( .A(n3607), .B(n2923), .ZN(n3613) );
  NAND2_X1 U4391 ( .A1(n4269), .A2(n3659), .ZN(n3610) );
  NAND2_X1 U4392 ( .A1(n3608), .A2(n3662), .ZN(n3609) );
  NAND2_X1 U4393 ( .A1(n3610), .A2(n3609), .ZN(n3614) );
  NAND2_X1 U4394 ( .A1(n3613), .A2(n3614), .ZN(n3711) );
  INV_X1 U4395 ( .A(n3711), .ZN(n3618) );
  NAND2_X1 U4396 ( .A1(n3797), .A2(n3796), .ZN(n3617) );
  INV_X1 U4397 ( .A(n3613), .ZN(n3616) );
  INV_X1 U4398 ( .A(n3614), .ZN(n3615) );
  NAND2_X1 U4399 ( .A1(n3616), .A2(n3615), .ZN(n3710) );
  NAND2_X1 U4400 ( .A1(n3621), .A2(n3620), .ZN(n3725) );
  NAND2_X1 U4401 ( .A1(n4333), .A2(n3662), .ZN(n3623) );
  NAND2_X1 U4402 ( .A1(n2173), .A2(n4277), .ZN(n3622) );
  NAND2_X1 U4403 ( .A1(n3623), .A2(n3622), .ZN(n3624) );
  XNOR2_X1 U4404 ( .A(n3624), .B(n3665), .ZN(n3627) );
  NOR2_X1 U4405 ( .A1(n3942), .A2(n2922), .ZN(n3625) );
  AOI21_X1 U4406 ( .B1(n4333), .B2(n2925), .A(n3625), .ZN(n3626) );
  OR2_X1 U4407 ( .A1(n3627), .A2(n3626), .ZN(n3776) );
  NAND2_X1 U4408 ( .A1(n3627), .A2(n3626), .ZN(n3775) );
  NAND2_X1 U4409 ( .A1(n4226), .A2(n3662), .ZN(n3629) );
  NAND2_X1 U4410 ( .A1(n4332), .A2(n2173), .ZN(n3628) );
  NAND2_X1 U4411 ( .A1(n3629), .A2(n3628), .ZN(n3630) );
  XNOR2_X1 U4412 ( .A(n3630), .B(n3665), .ZN(n3632) );
  NOR2_X1 U4413 ( .A1(n2922), .A2(n4253), .ZN(n3631) );
  AOI21_X1 U4414 ( .B1(n4226), .B2(n3659), .A(n3631), .ZN(n3633) );
  INV_X1 U4415 ( .A(n3632), .ZN(n3635) );
  INV_X1 U4416 ( .A(n3633), .ZN(n3634) );
  NAND2_X1 U4417 ( .A1(n3635), .A2(n3634), .ZN(n3723) );
  OAI22_X1 U4418 ( .A1(n4336), .A2(n3678), .B1(n4228), .B2(n3676), .ZN(n3636)
         );
  XNOR2_X1 U4419 ( .A(n3636), .B(n2923), .ZN(n3642) );
  OAI22_X1 U4420 ( .A1(n4336), .A2(n3679), .B1(n4228), .B2(n3678), .ZN(n3641)
         );
  XNOR2_X1 U4421 ( .A(n3642), .B(n3641), .ZN(n3788) );
  OAI22_X1 U4422 ( .A1(n4319), .A2(n3678), .B1(n3676), .B2(n4218), .ZN(n3637)
         );
  XNOR2_X1 U4423 ( .A(n3637), .B(n2923), .ZN(n3645) );
  OR2_X1 U4424 ( .A1(n4319), .A2(n3679), .ZN(n3640) );
  NAND2_X1 U4425 ( .A1(n3662), .A2(n3638), .ZN(n3639) );
  NAND2_X1 U4426 ( .A1(n3640), .A2(n3639), .ZN(n3644) );
  XNOR2_X1 U4427 ( .A(n3645), .B(n3644), .ZN(n3697) );
  NOR2_X1 U4428 ( .A1(n3642), .A2(n3641), .ZN(n3698) );
  NOR2_X1 U4429 ( .A1(n3697), .A2(n3698), .ZN(n3643) );
  NAND2_X1 U4430 ( .A1(n3645), .A2(n3644), .ZN(n3651) );
  INV_X1 U4431 ( .A(n3651), .ZN(n3648) );
  NOR2_X1 U4432 ( .A1(n2922), .A2(n4198), .ZN(n3646) );
  AOI21_X1 U4433 ( .B1(n4213), .B2(n2925), .A(n3646), .ZN(n3652) );
  OAI22_X1 U4434 ( .A1(n4175), .A2(n3678), .B1(n3676), .B2(n4198), .ZN(n3650)
         );
  XNOR2_X1 U4435 ( .A(n3650), .B(n2923), .ZN(n3768) );
  NAND2_X1 U4436 ( .A1(n3765), .A2(n3768), .ZN(n3654) );
  NAND2_X1 U4437 ( .A1(n3654), .A2(n3766), .ZN(n3736) );
  NAND2_X1 U4438 ( .A1(n4316), .A2(n3662), .ZN(n3656) );
  NAND2_X1 U4439 ( .A1(n2696), .A2(n2173), .ZN(n3655) );
  NAND2_X1 U4440 ( .A1(n3656), .A2(n3655), .ZN(n3657) );
  XNOR2_X1 U4441 ( .A(n3657), .B(n3665), .ZN(n3661) );
  NOR2_X1 U4442 ( .A1(n2922), .A2(n4181), .ZN(n3658) );
  AOI21_X1 U4443 ( .B1(n4316), .B2(n3659), .A(n3658), .ZN(n3660) );
  NAND2_X1 U4444 ( .A1(n3661), .A2(n3660), .ZN(n3734) );
  OR2_X1 U4445 ( .A1(n3661), .A2(n3660), .ZN(n3735) );
  NAND2_X1 U4446 ( .A1(n4295), .A2(n3662), .ZN(n3664) );
  NAND2_X1 U4447 ( .A1(n4303), .A2(n2173), .ZN(n3663) );
  NAND2_X1 U4448 ( .A1(n3664), .A2(n3663), .ZN(n3666) );
  XNOR2_X1 U4449 ( .A(n3666), .B(n3665), .ZN(n3670) );
  NOR2_X1 U4450 ( .A1(n2922), .A2(n4162), .ZN(n3667) );
  AOI21_X1 U4451 ( .B1(n4295), .B2(n2925), .A(n3667), .ZN(n3669) );
  NOR2_X1 U4452 ( .A1(n3670), .A2(n3669), .ZN(n3810) );
  INV_X1 U4453 ( .A(n3810), .ZN(n3668) );
  NAND2_X1 U4454 ( .A1(n3670), .A2(n3669), .ZN(n3808) );
  OAI22_X1 U4455 ( .A1(n4306), .A2(n3678), .B1(n3676), .B2(n4147), .ZN(n3671)
         );
  XNOR2_X1 U4456 ( .A(n3671), .B(n2923), .ZN(n3672) );
  OAI22_X1 U4457 ( .A1(n4306), .A2(n3679), .B1(n3678), .B2(n4147), .ZN(n3673)
         );
  XNOR2_X1 U4458 ( .A(n3672), .B(n3673), .ZN(n3689) );
  INV_X1 U4459 ( .A(n3672), .ZN(n3675) );
  INV_X1 U4460 ( .A(n3673), .ZN(n3674) );
  OAI22_X1 U4461 ( .A1(n4298), .A2(n3678), .B1(n3685), .B2(n3676), .ZN(n3677)
         );
  XNOR2_X1 U4462 ( .A(n3677), .B(n2923), .ZN(n3681) );
  OAI22_X1 U4463 ( .A1(n4298), .A2(n3679), .B1(n3685), .B2(n3678), .ZN(n3680)
         );
  XNOR2_X1 U4464 ( .A(n3681), .B(n3680), .ZN(n3682) );
  INV_X1 U4465 ( .A(n3683), .ZN(n4129) );
  INV_X1 U4466 ( .A(n3908), .ZN(n4132) );
  OAI22_X1 U4467 ( .A1(n4132), .A2(n3827), .B1(STATE_REG_SCAN_IN), .B2(n3684), 
        .ZN(n3687) );
  OAI22_X1 U4468 ( .A1(n4306), .A2(n3821), .B1(n3824), .B2(n3685), .ZN(n3686)
         );
  AOI211_X1 U4469 ( .C1(n4129), .C2(n3831), .A(n3687), .B(n3686), .ZN(n3688)
         );
  INV_X1 U4470 ( .A(n3691), .ZN(n4144) );
  AOI22_X1 U4471 ( .A1(n4295), .A2(n3789), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3693) );
  NAND2_X1 U4472 ( .A1(n3790), .A2(n4294), .ZN(n3692) );
  OAI211_X1 U4473 ( .C1(n4298), .C2(n3827), .A(n3693), .B(n3692), .ZN(n3694)
         );
  AOI21_X1 U4474 ( .B1(n4144), .B2(n3831), .A(n3694), .ZN(n3695) );
  OAI21_X1 U4475 ( .B1(n3696), .B2(n3834), .A(n3695), .ZN(U3211) );
  OAI21_X1 U4476 ( .B1(n2183), .B2(n3698), .A(n3697), .ZN(n3700) );
  NAND3_X1 U4477 ( .A1(n3700), .A2(n3777), .A3(n3699), .ZN(n3705) );
  OAI22_X1 U4478 ( .A1(n4336), .A2(n3821), .B1(n3824), .B2(n4218), .ZN(n3703)
         );
  OAI22_X1 U4479 ( .A1(n4175), .A2(n3827), .B1(STATE_REG_SCAN_IN), .B2(n3701), 
        .ZN(n3702) );
  AOI211_X1 U4480 ( .C1(n4219), .C2(n3831), .A(n3703), .B(n3702), .ZN(n3704)
         );
  NAND2_X1 U4481 ( .A1(n3705), .A2(n3704), .ZN(U3213) );
  INV_X1 U4482 ( .A(n3706), .ZN(n3708) );
  INV_X1 U4483 ( .A(n3796), .ZN(n3707) );
  NOR2_X1 U4484 ( .A1(n3708), .A2(n3707), .ZN(n3709) );
  OAI22_X1 U4485 ( .A1(n3709), .A2(n3797), .B1(n3796), .B2(n3706), .ZN(n3713)
         );
  NAND2_X1 U4486 ( .A1(n3711), .A2(n3710), .ZN(n3712) );
  XNOR2_X1 U4487 ( .A(n3713), .B(n3712), .ZN(n3714) );
  NAND2_X1 U4488 ( .A1(n3714), .A2(n3777), .ZN(n3720) );
  OAI22_X1 U4489 ( .A1(n3824), .A2(n3715), .B1(n3758), .B2(n3821), .ZN(n3718)
         );
  NAND2_X1 U4490 ( .A1(n3780), .A2(n4333), .ZN(n3716) );
  NAND2_X1 U4491 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4098) );
  NAND2_X1 U4492 ( .A1(n3716), .A2(n4098), .ZN(n3717) );
  NOR2_X1 U4493 ( .A1(n3718), .A2(n3717), .ZN(n3719) );
  OAI211_X1 U4494 ( .C1(n3786), .C2(n3721), .A(n3720), .B(n3719), .ZN(U3216)
         );
  INV_X1 U4495 ( .A(n3722), .ZN(n3724) );
  NAND2_X1 U4496 ( .A1(n3724), .A2(n3723), .ZN(n3727) );
  OAI211_X1 U4497 ( .C1(n3725), .C2(n2228), .A(n3776), .B(n3727), .ZN(n3726)
         );
  OAI211_X1 U4498 ( .C1(n3728), .C2(n3727), .A(n3777), .B(n3726), .ZN(n3733)
         );
  OAI22_X1 U4499 ( .A1(n3824), .A2(n4253), .B1(n3729), .B2(n3821), .ZN(n3731)
         );
  NOR2_X1 U4500 ( .A1(n4336), .A2(n3827), .ZN(n3730) );
  AOI211_X1 U4501 ( .C1(REG3_REG_21__SCAN_IN), .C2(U3149), .A(n3731), .B(n3730), .ZN(n3732) );
  OAI211_X1 U4502 ( .C1(n3786), .C2(n4254), .A(n3733), .B(n3732), .ZN(U3220)
         );
  NAND2_X1 U4503 ( .A1(n3735), .A2(n3734), .ZN(n3737) );
  XOR2_X1 U4504 ( .A(n3737), .B(n3736), .Z(n3741) );
  OAI22_X1 U4505 ( .A1(n4175), .A2(n3821), .B1(n3824), .B2(n4181), .ZN(n3739)
         );
  INV_X1 U4506 ( .A(n4295), .ZN(n4146) );
  OAI22_X1 U4507 ( .A1(n4146), .A2(n3827), .B1(STATE_REG_SCAN_IN), .B2(n4886), 
        .ZN(n3738) );
  AOI211_X1 U4508 ( .C1(n4183), .C2(n3831), .A(n3739), .B(n3738), .ZN(n3740)
         );
  OAI21_X1 U4509 ( .B1(n3741), .B2(n3834), .A(n3740), .ZN(U3222) );
  INV_X1 U4510 ( .A(n3742), .ZN(n3744) );
  OAI21_X1 U4511 ( .B1(n3744), .B2(n3820), .A(n3743), .ZN(n3745) );
  XOR2_X1 U4512 ( .A(n3746), .B(n3745), .Z(n3751) );
  AOI22_X1 U4513 ( .A1(n3790), .A2(n4354), .B1(n3789), .B2(n3999), .ZN(n3747)
         );
  NAND2_X1 U4514 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4483) );
  OAI211_X1 U4515 ( .C1(n3799), .C2(n3827), .A(n3747), .B(n4483), .ZN(n3748)
         );
  AOI21_X1 U4516 ( .B1(n3749), .B2(n3831), .A(n3748), .ZN(n3750) );
  OAI21_X1 U4517 ( .B1(n3751), .B2(n3834), .A(n3750), .ZN(U3223) );
  NAND2_X1 U4518 ( .A1(n3754), .A2(n3753), .ZN(n3755) );
  XNOR2_X1 U4519 ( .A(n3752), .B(n3755), .ZN(n3764) );
  OAI22_X1 U4520 ( .A1(n3824), .A2(n3756), .B1(n3826), .B2(n3821), .ZN(n3760)
         );
  INV_X1 U4521 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4703) );
  NOR2_X1 U4522 ( .A1(STATE_REG_SCAN_IN), .A2(n4703), .ZN(n4497) );
  INV_X1 U4523 ( .A(n4497), .ZN(n3757) );
  OAI21_X1 U4524 ( .B1(n3827), .B2(n3758), .A(n3757), .ZN(n3759) );
  NOR2_X1 U4525 ( .A1(n3760), .A2(n3759), .ZN(n3763) );
  NAND2_X1 U4526 ( .A1(n3831), .A2(n3761), .ZN(n3762) );
  OAI211_X1 U4527 ( .C1(n3764), .C2(n3834), .A(n3763), .B(n3762), .ZN(U3225)
         );
  NAND2_X1 U4528 ( .A1(n3766), .A2(n3765), .ZN(n3767) );
  XOR2_X1 U4529 ( .A(n3768), .B(n3767), .Z(n3773) );
  OAI22_X1 U4530 ( .A1(n4319), .A2(n3821), .B1(n3824), .B2(n4198), .ZN(n3771)
         );
  OAI22_X1 U4531 ( .A1(n4196), .A2(n3827), .B1(STATE_REG_SCAN_IN), .B2(n3769), 
        .ZN(n3770) );
  AOI211_X1 U4532 ( .C1(n4194), .C2(n3831), .A(n3771), .B(n3770), .ZN(n3772)
         );
  OAI21_X1 U4533 ( .B1(n3773), .B2(n3834), .A(n3772), .ZN(U3226) );
  NOR2_X1 U4534 ( .A1(n3774), .A2(n2228), .ZN(n3779) );
  AOI21_X1 U4535 ( .B1(n3776), .B2(n3775), .A(n3725), .ZN(n3778) );
  OAI21_X1 U4536 ( .B1(n3779), .B2(n3778), .A(n3777), .ZN(n3785) );
  NAND2_X1 U4537 ( .A1(n4226), .A2(n3780), .ZN(n3781) );
  OAI21_X1 U4538 ( .B1(STATE_REG_SCAN_IN), .B2(n4875), .A(n3781), .ZN(n3783)
         );
  INV_X1 U4539 ( .A(n4269), .ZN(n3801) );
  OAI22_X1 U4540 ( .A1(n3824), .A2(n3942), .B1(n3801), .B2(n3821), .ZN(n3782)
         );
  NOR2_X1 U4541 ( .A1(n3783), .A2(n3782), .ZN(n3784) );
  OAI211_X1 U4542 ( .C1(n3786), .C2(n4279), .A(n3785), .B(n3784), .ZN(U3230)
         );
  AOI21_X1 U4543 ( .B1(n3788), .B2(n3787), .A(n2183), .ZN(n3795) );
  AOI22_X1 U4544 ( .A1(n3790), .A2(n4234), .B1(n4226), .B2(n3789), .ZN(n3792)
         );
  NAND2_X1 U4545 ( .A1(U3149), .A2(REG3_REG_22__SCAN_IN), .ZN(n3791) );
  OAI211_X1 U4546 ( .C1(n4319), .C2(n3827), .A(n3792), .B(n3791), .ZN(n3793)
         );
  AOI21_X1 U4547 ( .B1(n4237), .B2(n3831), .A(n3793), .ZN(n3794) );
  OAI21_X1 U4548 ( .B1(n3795), .B2(n3834), .A(n3794), .ZN(U3232) );
  XNOR2_X1 U4549 ( .A(n3797), .B(n3796), .ZN(n3798) );
  XNOR2_X1 U4550 ( .A(n3706), .B(n3798), .ZN(n3807) );
  OAI22_X1 U4551 ( .A1(n3824), .A2(n3800), .B1(n3799), .B2(n3821), .ZN(n3803)
         );
  NAND2_X1 U4552 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4074) );
  OAI21_X1 U4553 ( .B1(n3827), .B2(n3801), .A(n4074), .ZN(n3802) );
  NOR2_X1 U4554 ( .A1(n3803), .A2(n3802), .ZN(n3806) );
  NAND2_X1 U4555 ( .A1(n3831), .A2(n3804), .ZN(n3805) );
  OAI211_X1 U4556 ( .C1(n3807), .C2(n3834), .A(n3806), .B(n3805), .ZN(U3235)
         );
  INV_X1 U4557 ( .A(n3808), .ZN(n3809) );
  NOR2_X1 U4558 ( .A1(n3810), .A2(n3809), .ZN(n3811) );
  XNOR2_X1 U4559 ( .A(n3812), .B(n3811), .ZN(n3818) );
  INV_X1 U4560 ( .A(n3813), .ZN(n4163) );
  INV_X1 U4561 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3814) );
  OAI22_X1 U4562 ( .A1(n4196), .A2(n3821), .B1(STATE_REG_SCAN_IN), .B2(n3814), 
        .ZN(n3816) );
  OAI22_X1 U4563 ( .A1(n4306), .A2(n3827), .B1(n3824), .B2(n4162), .ZN(n3815)
         );
  AOI211_X1 U4564 ( .C1(n4163), .C2(n3831), .A(n3816), .B(n3815), .ZN(n3817)
         );
  OAI21_X1 U4565 ( .B1(n3818), .B2(n3834), .A(n3817), .ZN(U3237) );
  NAND2_X1 U4566 ( .A1(n3742), .A2(n3743), .ZN(n3819) );
  XOR2_X1 U4567 ( .A(n3820), .B(n3819), .Z(n3835) );
  OAI22_X1 U4568 ( .A1(n3824), .A2(n3823), .B1(n3822), .B2(n3821), .ZN(n3829)
         );
  NOR2_X1 U4569 ( .A1(STATE_REG_SCAN_IN), .A2(n2599), .ZN(n4477) );
  INV_X1 U4570 ( .A(n4477), .ZN(n3825) );
  OAI21_X1 U4571 ( .B1(n3827), .B2(n3826), .A(n3825), .ZN(n3828) );
  NOR2_X1 U4572 ( .A1(n3829), .A2(n3828), .ZN(n3833) );
  NAND2_X1 U4573 ( .A1(n3831), .A2(n3830), .ZN(n3832) );
  OAI211_X1 U4574 ( .C1(n3835), .C2(n3834), .A(n3833), .B(n3832), .ZN(U3238)
         );
  NOR2_X1 U4575 ( .A1(n4306), .A2(n4294), .ZN(n3901) );
  NAND2_X1 U4576 ( .A1(n3837), .A2(n3836), .ZN(n3868) );
  AND2_X1 U4577 ( .A1(n3868), .A2(n3878), .ZN(n3882) );
  INV_X1 U4578 ( .A(n3838), .ZN(n3841) );
  OAI211_X1 U4579 ( .C1(n3841), .C2(n2735), .A(n3840), .B(n3839), .ZN(n3843)
         );
  NAND3_X1 U4580 ( .A1(n3843), .A2(n2738), .A3(n3842), .ZN(n3846) );
  NAND3_X1 U4581 ( .A1(n3846), .A2(n3845), .A3(n3844), .ZN(n3849) );
  NAND3_X1 U4582 ( .A1(n3849), .A2(n3848), .A3(n3847), .ZN(n3852) );
  NAND4_X1 U4583 ( .A1(n3852), .A2(n3851), .A3(n3850), .A4(n3861), .ZN(n3854)
         );
  NAND3_X1 U4584 ( .A1(n3854), .A2(n3927), .A3(n3853), .ZN(n3860) );
  AND2_X1 U4585 ( .A1(n3856), .A2(n3855), .ZN(n3862) );
  INV_X1 U4586 ( .A(n3858), .ZN(n3859) );
  AOI211_X1 U4587 ( .C1(n3860), .C2(n3862), .A(n2282), .B(n3859), .ZN(n3869)
         );
  INV_X1 U4588 ( .A(n3862), .ZN(n3864) );
  NOR3_X1 U4589 ( .A1(n2305), .A2(n3864), .A3(n3863), .ZN(n3866) );
  INV_X1 U4590 ( .A(n3873), .ZN(n3865) );
  INV_X1 U4591 ( .A(n3882), .ZN(n3957) );
  OAI21_X1 U4592 ( .B1(n3866), .B2(n3865), .A(n3957), .ZN(n3867) );
  OAI21_X1 U4593 ( .B1(n3869), .B2(n3868), .A(n3867), .ZN(n3877) );
  INV_X1 U4594 ( .A(n3870), .ZN(n3872) );
  AOI211_X1 U4595 ( .C1(n3874), .C2(n3873), .A(n3872), .B(n3871), .ZN(n3875)
         );
  NAND3_X1 U4596 ( .A1(n3877), .A2(n3876), .A3(n3875), .ZN(n3881) );
  AOI21_X1 U4597 ( .B1(n3879), .B2(n3878), .A(n3882), .ZN(n3955) );
  INV_X1 U4598 ( .A(n3955), .ZN(n3880) );
  OAI211_X1 U4599 ( .C1(n3883), .C2(n3882), .A(n3881), .B(n3880), .ZN(n3886)
         );
  INV_X1 U4600 ( .A(n3884), .ZN(n3956) );
  AOI21_X1 U4601 ( .B1(n3886), .B2(n3885), .A(n3956), .ZN(n3889) );
  INV_X1 U4602 ( .A(n3887), .ZN(n3888) );
  OAI21_X1 U4603 ( .B1(n3889), .B2(n3888), .A(n3960), .ZN(n3891) );
  INV_X1 U4604 ( .A(n4206), .ZN(n3890) );
  NAND3_X1 U4605 ( .A1(n3891), .A2(n3963), .A3(n3890), .ZN(n3892) );
  NAND2_X1 U4606 ( .A1(n3967), .A2(n3892), .ZN(n3894) );
  NOR2_X1 U4607 ( .A1(n3941), .A2(n3946), .ZN(n3965) );
  INV_X1 U4608 ( .A(n3965), .ZN(n3893) );
  AOI211_X1 U4609 ( .C1(n3895), .C2(n3894), .A(n3972), .B(n3893), .ZN(n3900)
         );
  NAND2_X1 U4610 ( .A1(n3908), .A2(n4115), .ZN(n3896) );
  AND2_X1 U4611 ( .A1(n3897), .A2(n3896), .ZN(n3974) );
  INV_X1 U4612 ( .A(n3974), .ZN(n3898) );
  OR4_X1 U4613 ( .A1(n3901), .A2(n3900), .A3(n3899), .A4(n3898), .ZN(n3911) );
  OR2_X1 U4614 ( .A1(n3903), .A2(n3902), .ZN(n3970) );
  AND2_X1 U4615 ( .A1(n3906), .A2(DATAI_30_), .ZN(n4290) );
  INV_X1 U4616 ( .A(n4290), .ZN(n3909) );
  INV_X1 U4617 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4285) );
  NAND2_X1 U4618 ( .A1(n2459), .A2(REG2_REG_31__SCAN_IN), .ZN(n3905) );
  NAND2_X1 U4619 ( .A1(n2460), .A2(REG0_REG_31__SCAN_IN), .ZN(n3904) );
  OAI211_X1 U4620 ( .C1(n2172), .C2(n4285), .A(n3905), .B(n3904), .ZN(n4107)
         );
  NAND2_X1 U4621 ( .A1(n3906), .A2(DATAI_31_), .ZN(n4108) );
  NAND2_X1 U4622 ( .A1(n4107), .A2(n4108), .ZN(n3910) );
  OAI21_X1 U4623 ( .B1(n3995), .B2(n3909), .A(n3910), .ZN(n3918) );
  INV_X1 U4624 ( .A(n3918), .ZN(n3907) );
  OAI21_X1 U4625 ( .B1(n3908), .B2(n4115), .A(n3907), .ZN(n3969) );
  AOI21_X1 U4626 ( .B1(n3974), .B2(n3970), .A(n3969), .ZN(n3976) );
  NAND2_X1 U4627 ( .A1(n3995), .A2(n3909), .ZN(n3981) );
  OAI21_X1 U4628 ( .B1(n4107), .B2(n4108), .A(n3981), .ZN(n3919) );
  AOI22_X1 U4629 ( .A1(n3911), .A2(n3976), .B1(n3919), .B2(n3910), .ZN(n3987)
         );
  INV_X1 U4630 ( .A(n4141), .ZN(n3953) );
  NAND2_X1 U4631 ( .A1(n4154), .A2(n3912), .ZN(n4174) );
  INV_X1 U4632 ( .A(n4174), .ZN(n3939) );
  INV_X1 U4633 ( .A(n4207), .ZN(n3913) );
  OR2_X1 U4634 ( .A1(n3913), .A2(n4206), .ZN(n4250) );
  NAND4_X1 U4635 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n3914), .ZN(n3920)
         );
  NOR4_X1 U4636 ( .A1(n4250), .A2(n3920), .A3(n3919), .A4(n3918), .ZN(n3938)
         );
  INV_X1 U4637 ( .A(n2736), .ZN(n3923) );
  INV_X1 U4638 ( .A(n3921), .ZN(n3922) );
  NAND4_X1 U4639 ( .A1(n3923), .A2(n3922), .A3(n4543), .A4(n2204), .ZN(n3929)
         );
  NAND4_X1 U4640 ( .A1(n3927), .A2(n3926), .A3(n3925), .A4(n3924), .ZN(n3928)
         );
  NOR2_X1 U4641 ( .A1(n3929), .A2(n3928), .ZN(n3937) );
  NAND4_X1 U4642 ( .A1(n3932), .A2(n3931), .A3(n3930), .A4(n4575), .ZN(n3935)
         );
  NOR4_X1 U4643 ( .A1(n4240), .A2(n3935), .A3(n3934), .A4(n3933), .ZN(n3936)
         );
  AND4_X1 U4644 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(n3950)
         );
  INV_X1 U4645 ( .A(n4171), .ZN(n3940) );
  OR2_X1 U4646 ( .A1(n3941), .A2(n3940), .ZN(n4190) );
  XNOR2_X1 U4647 ( .A(n4333), .B(n3942), .ZN(n4273) );
  NOR4_X1 U4648 ( .A1(n4190), .A2(n4273), .A3(n3944), .A4(n3943), .ZN(n3949)
         );
  INV_X1 U4649 ( .A(n3945), .ZN(n3947) );
  NOR2_X1 U4650 ( .A1(n3947), .A2(n3946), .ZN(n4211) );
  OR2_X1 U4651 ( .A1(n3948), .A2(n2196), .ZN(n4159) );
  NAND4_X1 U4652 ( .A1(n3950), .A2(n3949), .A3(n4211), .A4(n4159), .ZN(n3952)
         );
  NOR4_X1 U4653 ( .A1(n3954), .A2(n3953), .A3(n3952), .A4(n3951), .ZN(n3985)
         );
  INV_X1 U4654 ( .A(n4107), .ZN(n3980) );
  AOI211_X1 U4655 ( .C1(n3958), .C2(n3957), .A(n3956), .B(n3955), .ZN(n3962)
         );
  INV_X1 U4656 ( .A(n3959), .ZN(n3961) );
  OAI21_X1 U4657 ( .B1(n3962), .B2(n3961), .A(n3960), .ZN(n3964) );
  NAND2_X1 U4658 ( .A1(n3964), .A2(n3963), .ZN(n3966) );
  OAI221_X1 U4659 ( .B1(n3968), .B2(n3967), .C1(n3968), .C2(n3966), .A(n3965), 
        .ZN(n3971) );
  AOI211_X1 U4660 ( .C1(n4153), .C2(n3971), .A(n3970), .B(n3969), .ZN(n3978)
         );
  INV_X1 U4661 ( .A(n3972), .ZN(n3977) );
  NAND3_X1 U4662 ( .A1(n4141), .A2(n3974), .A3(n3973), .ZN(n3975) );
  AOI22_X1 U4663 ( .A1(n3978), .A2(n3977), .B1(n3976), .B2(n3975), .ZN(n3979)
         );
  AOI21_X1 U4664 ( .B1(n4290), .B2(n3980), .A(n3979), .ZN(n3983) );
  AOI21_X1 U4665 ( .B1(n3981), .B2(n4107), .A(n4108), .ZN(n3982) );
  NOR2_X1 U4666 ( .A1(n3983), .A2(n3982), .ZN(n3984) );
  MUX2_X1 U4667 ( .A(n3985), .B(n3984), .S(n2735), .Z(n3986) );
  MUX2_X1 U4668 ( .A(n3987), .B(n3986), .S(n4412), .Z(n3988) );
  XNOR2_X1 U4669 ( .A(n3988), .B(n4413), .ZN(n3994) );
  NAND2_X1 U4670 ( .A1(n3990), .A2(n3989), .ZN(n3991) );
  OAI211_X1 U4671 ( .C1(n4411), .C2(n3993), .A(n3991), .B(B_REG_SCAN_IN), .ZN(
        n3992) );
  OAI21_X1 U4672 ( .B1(n3994), .B2(n3993), .A(n3992), .ZN(U3239) );
  INV_X2 U4673 ( .A(U4043), .ZN(n4015) );
  MUX2_X1 U4674 ( .A(n4107), .B(DATAO_REG_31__SCAN_IN), .S(n4015), .Z(U3581)
         );
  MUX2_X1 U4675 ( .A(n3995), .B(DATAO_REG_30__SCAN_IN), .S(n4015), .Z(U3580)
         );
  MUX2_X1 U4676 ( .A(DATAO_REG_28__SCAN_IN), .B(n4117), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4677 ( .A(DATAO_REG_27__SCAN_IN), .B(n4128), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4678 ( .A(DATAO_REG_26__SCAN_IN), .B(n4295), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4679 ( .A(DATAO_REG_25__SCAN_IN), .B(n4316), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4680 ( .A(n4213), .B(DATAO_REG_24__SCAN_IN), .S(n4015), .Z(U3574)
         );
  MUX2_X1 U4681 ( .A(DATAO_REG_23__SCAN_IN), .B(n4231), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4682 ( .A(DATAO_REG_22__SCAN_IN), .B(n3996), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4683 ( .A(n4226), .B(DATAO_REG_21__SCAN_IN), .S(n4015), .Z(U3571)
         );
  MUX2_X1 U4684 ( .A(DATAO_REG_20__SCAN_IN), .B(n4333), .S(U4043), .Z(U3570)
         );
  MUX2_X1 U4685 ( .A(n4269), .B(DATAO_REG_19__SCAN_IN), .S(n4015), .Z(U3569)
         );
  MUX2_X1 U4686 ( .A(DATAO_REG_18__SCAN_IN), .B(n3997), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4687 ( .A(DATAO_REG_17__SCAN_IN), .B(n4356), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4688 ( .A(n3998), .B(DATAO_REG_16__SCAN_IN), .S(n4015), .Z(U3566)
         );
  MUX2_X1 U4689 ( .A(n3999), .B(DATAO_REG_15__SCAN_IN), .S(n4015), .Z(U3565)
         );
  MUX2_X1 U4690 ( .A(n4000), .B(DATAO_REG_14__SCAN_IN), .S(n4015), .Z(U3564)
         );
  MUX2_X1 U4691 ( .A(n4001), .B(DATAO_REG_13__SCAN_IN), .S(n4015), .Z(U3563)
         );
  MUX2_X1 U4692 ( .A(n4002), .B(DATAO_REG_12__SCAN_IN), .S(n4015), .Z(U3562)
         );
  MUX2_X1 U4693 ( .A(n4003), .B(DATAO_REG_11__SCAN_IN), .S(n4015), .Z(U3561)
         );
  MUX2_X1 U4694 ( .A(n4004), .B(DATAO_REG_10__SCAN_IN), .S(n4015), .Z(U3560)
         );
  MUX2_X1 U4695 ( .A(n4005), .B(DATAO_REG_9__SCAN_IN), .S(n4015), .Z(U3559) );
  MUX2_X1 U4696 ( .A(n4006), .B(DATAO_REG_8__SCAN_IN), .S(n4015), .Z(U3558) );
  MUX2_X1 U4697 ( .A(n4007), .B(DATAO_REG_7__SCAN_IN), .S(n4015), .Z(U3557) );
  MUX2_X1 U4698 ( .A(n4008), .B(DATAO_REG_6__SCAN_IN), .S(n4015), .Z(U3556) );
  MUX2_X1 U4699 ( .A(DATAO_REG_5__SCAN_IN), .B(n4009), .S(U4043), .Z(U3555) );
  MUX2_X1 U4700 ( .A(n4010), .B(DATAO_REG_4__SCAN_IN), .S(n4015), .Z(U3554) );
  MUX2_X1 U4701 ( .A(n4011), .B(DATAO_REG_3__SCAN_IN), .S(n4015), .Z(U3553) );
  MUX2_X1 U4702 ( .A(n4012), .B(DATAO_REG_2__SCAN_IN), .S(n4015), .Z(U3552) );
  MUX2_X1 U4703 ( .A(n2456), .B(DATAO_REG_1__SCAN_IN), .S(n4015), .Z(U3551) );
  MUX2_X1 U4704 ( .A(n4013), .B(DATAO_REG_0__SCAN_IN), .S(n4015), .Z(U3550) );
  NAND3_X1 U4705 ( .A1(n4014), .A2(n4409), .A3(n4426), .ZN(n4017) );
  OAI21_X1 U4706 ( .B1(REG2_REG_0__SCAN_IN), .B2(n4426), .A(n4409), .ZN(n4425)
         );
  AOI21_X1 U4707 ( .B1(n4425), .B2(n2211), .A(n4015), .ZN(n4016) );
  OAI211_X1 U4708 ( .C1(n4019), .C2(n4018), .A(n4017), .B(n4016), .ZN(n4041)
         );
  AOI22_X1 U4709 ( .A1(n4498), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4029) );
  XOR2_X1 U4710 ( .A(n4021), .B(n4020), .Z(n4026) );
  AOI211_X1 U4711 ( .C1(n4024), .C2(n4023), .A(n4022), .B(n4103), .ZN(n4025)
         );
  AOI21_X1 U4712 ( .B1(n4464), .B2(n4026), .A(n4025), .ZN(n4028) );
  INV_X1 U4713 ( .A(n4505), .ZN(n4044) );
  NAND2_X1 U4714 ( .A1(n4044), .A2(n4420), .ZN(n4027) );
  NAND4_X1 U4715 ( .A1(n4041), .A2(n4029), .A3(n4028), .A4(n4027), .ZN(U3242)
         );
  XNOR2_X1 U4716 ( .A(n4030), .B(REG2_REG_4__SCAN_IN), .ZN(n4036) );
  INV_X1 U4717 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4034) );
  INV_X1 U4718 ( .A(n4498), .ZN(n4033) );
  NAND2_X1 U4719 ( .A1(n4044), .A2(n4418), .ZN(n4032) );
  OAI211_X1 U4720 ( .C1(n4034), .C2(n4033), .A(n4032), .B(n4031), .ZN(n4035)
         );
  AOI21_X1 U4721 ( .B1(n4464), .B2(n4036), .A(n4035), .ZN(n4040) );
  OAI211_X1 U4722 ( .C1(n4038), .C2(REG1_REG_4__SCAN_IN), .A(n4037), .B(n4499), 
        .ZN(n4039) );
  NAND3_X1 U4723 ( .A1(n4041), .A2(n4040), .A3(n4039), .ZN(U3244) );
  OAI211_X1 U4724 ( .C1(n4043), .C2(REG1_REG_10__SCAN_IN), .A(n4499), .B(n4042), .ZN(n4051) );
  AOI22_X1 U4725 ( .A1(n4044), .A2(n4415), .B1(n4498), .B2(
        ADDR_REG_10__SCAN_IN), .ZN(n4050) );
  OAI211_X1 U4726 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4046), .A(n4464), .B(n4045), .ZN(n4047) );
  AND2_X1 U4727 ( .A1(n4048), .A2(n4047), .ZN(n4049) );
  NAND3_X1 U4728 ( .A1(n4051), .A2(n4050), .A3(n4049), .ZN(U3250) );
  INV_X1 U4729 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4810) );
  INV_X1 U4730 ( .A(n4059), .ZN(n4066) );
  AOI21_X1 U4731 ( .B1(n4066), .B2(n4055), .A(n4079), .ZN(n4056) );
  INV_X1 U4732 ( .A(n4056), .ZN(n4057) );
  AOI211_X1 U4733 ( .C1(n4810), .C2(n4057), .A(n4078), .B(n4492), .ZN(n4065)
         );
  OAI211_X1 U4734 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4060), .A(n4499), .B(n4068), .ZN(n4063) );
  AOI21_X1 U4735 ( .B1(n4498), .B2(ADDR_REG_14__SCAN_IN), .A(n4061), .ZN(n4062) );
  OAI211_X1 U4736 ( .C1(n4505), .C2(n4066), .A(n4063), .B(n4062), .ZN(n4064)
         );
  OR2_X1 U4737 ( .A1(n4065), .A2(n4064), .ZN(U3254) );
  XNOR2_X1 U4738 ( .A(n4075), .B(REG1_REG_18__SCAN_IN), .ZN(n4089) );
  NAND2_X1 U4739 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4081), .ZN(n4070) );
  INV_X1 U4740 ( .A(n4081), .ZN(n4565) );
  INV_X1 U4741 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4833) );
  AOI22_X1 U4742 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4081), .B1(n4565), .B2(
        n4833), .ZN(n4480) );
  OR2_X1 U4743 ( .A1(n4067), .A2(n4066), .ZN(n4069) );
  NAND2_X1 U4744 ( .A1(n4069), .A2(n4068), .ZN(n4479) );
  NOR2_X1 U4745 ( .A1(n4563), .A2(n4071), .ZN(n4072) );
  INV_X1 U4746 ( .A(n4563), .ZN(n4491) );
  NOR2_X1 U4747 ( .A1(n4072), .A2(n2185), .ZN(n4501) );
  AOI22_X1 U4748 ( .A1(n4084), .A2(n3546), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4562), .ZN(n4500) );
  NOR2_X1 U4749 ( .A1(n4501), .A2(n4500), .ZN(n4502) );
  NAND2_X1 U4750 ( .A1(n4498), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4073) );
  OAI211_X1 U4751 ( .C1(n4505), .C2(n4075), .A(n4074), .B(n4073), .ZN(n4088)
         );
  INV_X1 U4752 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4893) );
  NOR2_X1 U4753 ( .A1(n4094), .A2(n4893), .ZN(n4076) );
  AOI21_X1 U4754 ( .B1(n4094), .B2(n4893), .A(n4076), .ZN(n4086) );
  NOR2_X1 U4755 ( .A1(n4084), .A2(REG2_REG_17__SCAN_IN), .ZN(n4077) );
  AOI21_X1 U4756 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4084), .A(n4077), .ZN(n4495) );
  NOR2_X1 U4757 ( .A1(n4079), .A2(n4078), .ZN(n4475) );
  NAND2_X1 U4758 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4081), .ZN(n4080) );
  OAI21_X1 U4759 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4081), .A(n4080), .ZN(n4474) );
  NAND2_X1 U4760 ( .A1(n4082), .A2(n4491), .ZN(n4083) );
  INV_X1 U4761 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4922) );
  NAND2_X1 U4762 ( .A1(n4083), .A2(n4484), .ZN(n4493) );
  NAND2_X1 U4763 ( .A1(n4495), .A2(n4493), .ZN(n4494) );
  OAI21_X1 U4764 ( .B1(n4084), .B2(REG2_REG_17__SCAN_IN), .A(n4494), .ZN(n4085) );
  NOR2_X1 U4765 ( .A1(n4085), .A2(n4086), .ZN(n4093) );
  AOI211_X1 U4766 ( .C1(n4086), .C2(n4085), .A(n4093), .B(n4492), .ZN(n4087)
         );
  AOI22_X1 U4767 ( .A1(n4090), .A2(n4089), .B1(REG1_REG_18__SCAN_IN), .B2(
        n4094), .ZN(n4092) );
  MUX2_X1 U4768 ( .A(n4348), .B(REG1_REG_19__SCAN_IN), .S(n4413), .Z(n4091) );
  XNOR2_X1 U4769 ( .A(n4092), .B(n4091), .ZN(n4104) );
  MUX2_X1 U4770 ( .A(REG2_REG_19__SCAN_IN), .B(n3560), .S(n4413), .Z(n4095) );
  XNOR2_X1 U4771 ( .A(n4096), .B(n4095), .ZN(n4101) );
  NAND2_X1 U4772 ( .A1(n4498), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4097) );
  OAI211_X1 U4773 ( .C1(n4505), .C2(n4099), .A(n4098), .B(n4097), .ZN(n4100)
         );
  AOI21_X1 U4774 ( .B1(n4101), .B2(n4464), .A(n4100), .ZN(n4102) );
  OAI21_X1 U4775 ( .B1(n4104), .B2(n4103), .A(n4102), .ZN(U3259) );
  XNOR2_X1 U4776 ( .A(n4288), .B(n4108), .ZN(n4370) );
  INV_X1 U4777 ( .A(n4105), .ZN(n4106) );
  NAND2_X1 U4778 ( .A1(n4107), .A2(n4106), .ZN(n4292) );
  INV_X1 U4779 ( .A(n4108), .ZN(n4109) );
  NAND2_X1 U4780 ( .A1(n4109), .A2(n4535), .ZN(n4110) );
  NAND2_X1 U4781 ( .A1(n4292), .A2(n4110), .ZN(n4367) );
  NAND2_X1 U4782 ( .A1(n4245), .A2(n4367), .ZN(n4112) );
  NAND2_X1 U4783 ( .A1(n4557), .A2(REG2_REG_31__SCAN_IN), .ZN(n4111) );
  OAI211_X1 U4784 ( .C1(n4370), .C2(n4239), .A(n4112), .B(n4111), .ZN(U3260)
         );
  INV_X1 U4785 ( .A(n4113), .ZN(n4124) );
  INV_X1 U4786 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4114) );
  OAI22_X1 U4787 ( .A1(n4197), .A2(n4115), .B1(n4114), .B2(n4245), .ZN(n4116)
         );
  AOI21_X1 U4788 ( .B1(n4117), .B2(n4256), .A(n4116), .ZN(n4123) );
  OAI22_X1 U4789 ( .A1(n4119), .A2(n4239), .B1(n4118), .B2(n4615), .ZN(n4120)
         );
  OAI21_X1 U4790 ( .B1(n4121), .B2(n4120), .A(n4245), .ZN(n4122) );
  OAI211_X1 U4791 ( .C1(n4124), .C2(n4621), .A(n4123), .B(n4122), .ZN(U3354)
         );
  NAND2_X1 U4792 ( .A1(n4125), .A2(n4251), .ZN(n4136) );
  INV_X1 U4793 ( .A(n4126), .ZN(n4134) );
  AOI22_X1 U4794 ( .A1(n4128), .A2(n4256), .B1(n4127), .B2(n4257), .ZN(n4131)
         );
  AOI22_X1 U4795 ( .A1(n4129), .A2(n4549), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4557), .ZN(n4130) );
  OAI211_X1 U4796 ( .C1(n4132), .C2(n4260), .A(n4131), .B(n4130), .ZN(n4133)
         );
  AOI21_X1 U4797 ( .B1(n4134), .B2(n4618), .A(n4133), .ZN(n4135) );
  OAI211_X1 U4798 ( .C1(n4557), .C2(n4137), .A(n4136), .B(n4135), .ZN(U3262)
         );
  OAI21_X1 U4799 ( .B1(n4141), .B2(n4139), .A(n4138), .ZN(n4140) );
  NAND2_X1 U4800 ( .A1(n4140), .A2(n4548), .ZN(n4297) );
  XNOR2_X1 U4801 ( .A(n4142), .B(n4141), .ZN(n4300) );
  NAND2_X1 U4802 ( .A1(n4300), .A2(n4251), .ZN(n4152) );
  OAI21_X1 U4803 ( .B1(n4160), .B2(n4147), .A(n4143), .ZN(n4377) );
  INV_X1 U4804 ( .A(n4377), .ZN(n4150) );
  INV_X1 U4805 ( .A(n4256), .ZN(n4199) );
  AOI22_X1 U4806 ( .A1(n4144), .A2(n4549), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4557), .ZN(n4145) );
  OAI21_X1 U4807 ( .B1(n4146), .B2(n4199), .A(n4145), .ZN(n4149) );
  OAI22_X1 U4808 ( .A1(n4298), .A2(n4260), .B1(n4197), .B2(n4147), .ZN(n4148)
         );
  AOI211_X1 U4809 ( .C1(n4150), .C2(n4618), .A(n4149), .B(n4148), .ZN(n4151)
         );
  OAI211_X1 U4810 ( .C1(n4557), .C2(n4297), .A(n4152), .B(n4151), .ZN(U3263)
         );
  NAND2_X1 U4811 ( .A1(n4172), .A2(n4153), .ZN(n4155) );
  NAND2_X1 U4812 ( .A1(n4155), .A2(n4154), .ZN(n4156) );
  XNOR2_X1 U4813 ( .A(n4156), .B(n4159), .ZN(n4157) );
  NAND2_X1 U4814 ( .A1(n4157), .A2(n4548), .ZN(n4305) );
  XOR2_X1 U4815 ( .A(n4159), .B(n4158), .Z(n4308) );
  NAND2_X1 U4816 ( .A1(n4308), .A2(n4251), .ZN(n4169) );
  INV_X1 U4817 ( .A(n4160), .ZN(n4161) );
  OAI21_X1 U4818 ( .B1(n4179), .B2(n4162), .A(n4161), .ZN(n4381) );
  INV_X1 U4819 ( .A(n4381), .ZN(n4167) );
  AOI22_X1 U4820 ( .A1(n4163), .A2(n4549), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4557), .ZN(n4165) );
  AOI22_X1 U4821 ( .A1(n4316), .A2(n4256), .B1(n4303), .B2(n4257), .ZN(n4164)
         );
  OAI211_X1 U4822 ( .C1(n4306), .C2(n4260), .A(n4165), .B(n4164), .ZN(n4166)
         );
  AOI21_X1 U4823 ( .B1(n4167), .B2(n4618), .A(n4166), .ZN(n4168) );
  OAI211_X1 U4824 ( .C1(n4557), .C2(n4305), .A(n4169), .B(n4168), .ZN(U3264)
         );
  XNOR2_X1 U4825 ( .A(n4170), .B(n4174), .ZN(n4312) );
  INV_X1 U4826 ( .A(n4312), .ZN(n4187) );
  NAND2_X1 U4827 ( .A1(n4172), .A2(n4171), .ZN(n4173) );
  XOR2_X1 U4828 ( .A(n4174), .B(n4173), .Z(n4178) );
  OAI22_X1 U4829 ( .A1(n4175), .A2(n4358), .B1(n4181), .B2(n4229), .ZN(n4176)
         );
  AOI21_X1 U4830 ( .B1(n4295), .B2(n4355), .A(n4176), .ZN(n4177) );
  OAI21_X1 U4831 ( .B1(n4178), .B2(n4215), .A(n4177), .ZN(n4311) );
  INV_X1 U4832 ( .A(n4193), .ZN(n4182) );
  INV_X1 U4833 ( .A(n4179), .ZN(n4180) );
  OAI21_X1 U4834 ( .B1(n4182), .B2(n4181), .A(n4180), .ZN(n4385) );
  AOI22_X1 U4835 ( .A1(n4183), .A2(n4549), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4557), .ZN(n4184) );
  OAI21_X1 U4836 ( .B1(n4385), .B2(n4239), .A(n4184), .ZN(n4185) );
  AOI21_X1 U4837 ( .B1(n4311), .B2(n4245), .A(n4185), .ZN(n4186) );
  OAI21_X1 U4838 ( .B1(n4187), .B2(n4621), .A(n4186), .ZN(U3265) );
  XOR2_X1 U4839 ( .A(n4190), .B(n4188), .Z(n4189) );
  NAND2_X1 U4840 ( .A1(n4189), .A2(n4548), .ZN(n4318) );
  XNOR2_X1 U4841 ( .A(n4191), .B(n4190), .ZN(n4321) );
  NAND2_X1 U4842 ( .A1(n4321), .A2(n4251), .ZN(n4204) );
  NAND2_X1 U4843 ( .A1(n4217), .A2(n4315), .ZN(n4192) );
  NAND2_X1 U4844 ( .A1(n4193), .A2(n4192), .ZN(n4388) );
  INV_X1 U4845 ( .A(n4388), .ZN(n4202) );
  AOI22_X1 U4846 ( .A1(n4194), .A2(n4549), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4557), .ZN(n4195) );
  OAI21_X1 U4847 ( .B1(n4196), .B2(n4260), .A(n4195), .ZN(n4201) );
  OAI22_X1 U4848 ( .A1(n4319), .A2(n4199), .B1(n4198), .B2(n4197), .ZN(n4200)
         );
  AOI211_X1 U4849 ( .C1(n4202), .C2(n4618), .A(n4201), .B(n4200), .ZN(n4203)
         );
  OAI211_X1 U4850 ( .C1(n4557), .C2(n4318), .A(n4204), .B(n4203), .ZN(U3266)
         );
  XNOR2_X1 U4851 ( .A(n4205), .B(n4211), .ZN(n4324) );
  INV_X1 U4852 ( .A(n4324), .ZN(n4223) );
  OR2_X1 U4853 ( .A1(n4247), .A2(n4206), .ZN(n4208) );
  OAI21_X1 U4854 ( .B1(n4224), .B2(n4240), .A(n4209), .ZN(n4210) );
  XOR2_X1 U4855 ( .A(n4211), .B(n4210), .Z(n4216) );
  OAI22_X1 U4856 ( .A1(n4336), .A2(n4358), .B1(n4229), .B2(n4218), .ZN(n4212)
         );
  AOI21_X1 U4857 ( .B1(n4355), .B2(n4213), .A(n4212), .ZN(n4214) );
  OAI21_X1 U4858 ( .B1(n4216), .B2(n4215), .A(n4214), .ZN(n4323) );
  OAI21_X1 U4859 ( .B1(n4235), .B2(n4218), .A(n4217), .ZN(n4392) );
  AOI22_X1 U4860 ( .A1(n4219), .A2(n4549), .B1(n4557), .B2(
        REG2_REG_23__SCAN_IN), .ZN(n4220) );
  OAI21_X1 U4861 ( .B1(n4392), .B2(n4239), .A(n4220), .ZN(n4221) );
  AOI21_X1 U4862 ( .B1(n4323), .B2(n4245), .A(n4221), .ZN(n4222) );
  OAI21_X1 U4863 ( .B1(n4223), .B2(n4621), .A(n4222), .ZN(U3267) );
  XNOR2_X1 U4864 ( .A(n4224), .B(n4240), .ZN(n4225) );
  NAND2_X1 U4865 ( .A1(n4225), .A2(n4548), .ZN(n4233) );
  NAND2_X1 U4866 ( .A1(n4226), .A2(n4536), .ZN(n4227) );
  OAI21_X1 U4867 ( .B1(n4229), .B2(n4228), .A(n4227), .ZN(n4230) );
  AOI21_X1 U4868 ( .B1(n4231), .B2(n4355), .A(n4230), .ZN(n4232) );
  NAND2_X1 U4869 ( .A1(n4233), .A2(n4232), .ZN(n4328) );
  AND2_X1 U4870 ( .A1(n4252), .A2(n4234), .ZN(n4236) );
  OR2_X1 U4871 ( .A1(n4236), .A2(n4235), .ZN(n4395) );
  AOI22_X1 U4872 ( .A1(n4237), .A2(n4549), .B1(n4557), .B2(
        REG2_REG_22__SCAN_IN), .ZN(n4238) );
  OAI21_X1 U4873 ( .B1(n4395), .B2(n4239), .A(n4238), .ZN(n4244) );
  NOR2_X1 U4874 ( .A1(n4241), .A2(n4240), .ZN(n4327) );
  INV_X1 U4875 ( .A(n4329), .ZN(n4242) );
  NOR3_X1 U4876 ( .A1(n4327), .A2(n4242), .A3(n4621), .ZN(n4243) );
  AOI211_X1 U4877 ( .C1(n4245), .C2(n4328), .A(n4244), .B(n4243), .ZN(n4246)
         );
  INV_X1 U4878 ( .A(n4246), .ZN(U3268) );
  XNOR2_X1 U4879 ( .A(n4247), .B(n4250), .ZN(n4248) );
  NAND2_X1 U4880 ( .A1(n4248), .A2(n4548), .ZN(n4335) );
  XOR2_X1 U4881 ( .A(n4250), .B(n4249), .Z(n4338) );
  NAND2_X1 U4882 ( .A1(n4338), .A2(n4251), .ZN(n4264) );
  OAI21_X1 U4883 ( .B1(n2255), .B2(n4253), .A(n4252), .ZN(n4399) );
  INV_X1 U4884 ( .A(n4399), .ZN(n4262) );
  INV_X1 U4885 ( .A(n4254), .ZN(n4255) );
  AOI22_X1 U4886 ( .A1(n4557), .A2(REG2_REG_21__SCAN_IN), .B1(n4255), .B2(
        n4549), .ZN(n4259) );
  AOI22_X1 U4887 ( .A1(n4257), .A2(n4332), .B1(n4256), .B2(n4333), .ZN(n4258)
         );
  OAI211_X1 U4888 ( .C1(n4336), .C2(n4260), .A(n4259), .B(n4258), .ZN(n4261)
         );
  AOI21_X1 U4889 ( .B1(n4262), .B2(n4618), .A(n4261), .ZN(n4263) );
  OAI211_X1 U4890 ( .C1(n4557), .C2(n4335), .A(n4264), .B(n4263), .ZN(U3269)
         );
  OAI21_X1 U4891 ( .B1(n4267), .B2(n4266), .A(n4265), .ZN(n4268) );
  XOR2_X1 U4892 ( .A(n4273), .B(n4268), .Z(n4276) );
  AOI22_X1 U4893 ( .A1(n4269), .A2(n4536), .B1(n4277), .B2(n4535), .ZN(n4270)
         );
  OAI21_X1 U4894 ( .B1(n4271), .B2(n4538), .A(n4270), .ZN(n4275) );
  XNOR2_X1 U4895 ( .A(n4272), .B(n4273), .ZN(n4345) );
  NOR2_X1 U4896 ( .A1(n4345), .A2(n4544), .ZN(n4274) );
  AOI211_X1 U4897 ( .C1(n4276), .C2(n4548), .A(n4275), .B(n4274), .ZN(n4344)
         );
  INV_X1 U4898 ( .A(n4345), .ZN(n4283) );
  NAND2_X1 U4899 ( .A1(n4278), .A2(n4277), .ZN(n4341) );
  AND3_X1 U4900 ( .A1(n4342), .A2(n4618), .A3(n4341), .ZN(n4282) );
  INV_X1 U4901 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4280) );
  OAI22_X1 U4902 ( .A1(n4245), .A2(n4280), .B1(n4279), .B2(n4615), .ZN(n4281)
         );
  AOI211_X1 U4903 ( .C1(n4283), .C2(n4553), .A(n4282), .B(n4281), .ZN(n4284)
         );
  OAI21_X1 U4904 ( .B1(n4344), .B2(n4557), .A(n4284), .ZN(U3270) );
  NOR2_X1 U4905 ( .A1(n4612), .A2(n4285), .ZN(n4286) );
  AOI21_X1 U4906 ( .B1(n4612), .B2(n4367), .A(n4286), .ZN(n4287) );
  OAI21_X1 U4907 ( .B1(n4370), .B2(n4350), .A(n4287), .ZN(U3549) );
  AOI21_X1 U4908 ( .B1(n4290), .B2(n4289), .A(n4288), .ZN(n4422) );
  INV_X1 U4909 ( .A(n4422), .ZN(n4373) );
  NAND2_X1 U4910 ( .A1(n4535), .A2(n4290), .ZN(n4291) );
  AND2_X1 U4911 ( .A1(n4292), .A2(n4291), .ZN(n4424) );
  MUX2_X1 U4912 ( .A(n4424), .B(n2817), .S(n4610), .Z(n4293) );
  OAI21_X1 U4913 ( .B1(n4373), .B2(n4350), .A(n4293), .ZN(U3548) );
  AOI22_X1 U4914 ( .A1(n4295), .A2(n4536), .B1(n4294), .B2(n4535), .ZN(n4296)
         );
  OAI211_X1 U4915 ( .C1(n4298), .C2(n4538), .A(n4297), .B(n4296), .ZN(n4299)
         );
  AOI21_X1 U4916 ( .B1(n4300), .B2(n4594), .A(n4299), .ZN(n4374) );
  MUX2_X1 U4917 ( .A(n4301), .B(n4374), .S(n4612), .Z(n4302) );
  OAI21_X1 U4918 ( .B1(n4350), .B2(n4377), .A(n4302), .ZN(U3545) );
  AOI22_X1 U4919 ( .A1(n4316), .A2(n4536), .B1(n4303), .B2(n4535), .ZN(n4304)
         );
  OAI211_X1 U4920 ( .C1(n4306), .C2(n4538), .A(n4305), .B(n4304), .ZN(n4307)
         );
  AOI21_X1 U4921 ( .B1(n4308), .B2(n4594), .A(n4307), .ZN(n4378) );
  MUX2_X1 U4922 ( .A(n4309), .B(n4378), .S(n4612), .Z(n4310) );
  OAI21_X1 U4923 ( .B1(n4350), .B2(n4381), .A(n4310), .ZN(U3544) );
  AOI21_X1 U4924 ( .B1(n4312), .B2(n4594), .A(n4311), .ZN(n4382) );
  MUX2_X1 U4925 ( .A(n4313), .B(n4382), .S(n4612), .Z(n4314) );
  OAI21_X1 U4926 ( .B1(n4350), .B2(n4385), .A(n4314), .ZN(U3543) );
  AOI22_X1 U4927 ( .A1(n4316), .A2(n4355), .B1(n4535), .B2(n4315), .ZN(n4317)
         );
  OAI211_X1 U4928 ( .C1(n4319), .C2(n4358), .A(n4318), .B(n4317), .ZN(n4320)
         );
  AOI21_X1 U4929 ( .B1(n4321), .B2(n4594), .A(n4320), .ZN(n4386) );
  MUX2_X1 U4930 ( .A(n4724), .B(n4386), .S(n4612), .Z(n4322) );
  OAI21_X1 U4931 ( .B1(n4350), .B2(n4388), .A(n4322), .ZN(U3542) );
  AOI21_X1 U4932 ( .B1(n4324), .B2(n4594), .A(n4323), .ZN(n4389) );
  MUX2_X1 U4933 ( .A(n4325), .B(n4389), .S(n4612), .Z(n4326) );
  OAI21_X1 U4934 ( .B1(n4350), .B2(n4392), .A(n4326), .ZN(U3541) );
  INV_X1 U4935 ( .A(n4594), .ZN(n4365) );
  NOR2_X1 U4936 ( .A1(n4327), .A2(n4365), .ZN(n4330) );
  AOI21_X1 U4937 ( .B1(n4330), .B2(n4329), .A(n4328), .ZN(n4393) );
  MUX2_X1 U4938 ( .A(n4717), .B(n4393), .S(n4612), .Z(n4331) );
  OAI21_X1 U4939 ( .B1(n4350), .B2(n4395), .A(n4331), .ZN(U3540) );
  INV_X1 U4940 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4339) );
  AOI22_X1 U4941 ( .A1(n4333), .A2(n4536), .B1(n4332), .B2(n4535), .ZN(n4334)
         );
  OAI211_X1 U4942 ( .C1(n4336), .C2(n4538), .A(n4335), .B(n4334), .ZN(n4337)
         );
  AOI21_X1 U4943 ( .B1(n4338), .B2(n4594), .A(n4337), .ZN(n4396) );
  MUX2_X1 U4944 ( .A(n4339), .B(n4396), .S(n4612), .Z(n4340) );
  OAI21_X1 U4945 ( .B1(n4350), .B2(n4399), .A(n4340), .ZN(U3539) );
  NAND3_X1 U4946 ( .A1(n4342), .A2(n4361), .A3(n4341), .ZN(n4343) );
  OAI211_X1 U4947 ( .C1(n4345), .C2(n4585), .A(n4344), .B(n4343), .ZN(n4400)
         );
  MUX2_X1 U4948 ( .A(REG1_REG_20__SCAN_IN), .B(n4400), .S(n4612), .Z(U3538) );
  AOI21_X1 U4949 ( .B1(n4347), .B2(n4594), .A(n4346), .ZN(n4401) );
  MUX2_X1 U4950 ( .A(n4348), .B(n4401), .S(n4612), .Z(n4349) );
  OAI21_X1 U4951 ( .B1(n4350), .B2(n4405), .A(n4349), .ZN(U3537) );
  OAI211_X1 U4952 ( .C1(n4353), .C2(n4365), .A(n4352), .B(n4351), .ZN(n4406)
         );
  MUX2_X1 U4953 ( .A(REG1_REG_18__SCAN_IN), .B(n4406), .S(n4612), .Z(U3536) );
  AOI22_X1 U4954 ( .A1(n4356), .A2(n4355), .B1(n4354), .B2(n4535), .ZN(n4357)
         );
  OAI21_X1 U4955 ( .B1(n4359), .B2(n4358), .A(n4357), .ZN(n4360) );
  AOI21_X1 U4956 ( .B1(n4362), .B2(n4361), .A(n4360), .ZN(n4364) );
  OAI211_X1 U4957 ( .C1(n4366), .C2(n4365), .A(n4364), .B(n4363), .ZN(n4407)
         );
  MUX2_X1 U4958 ( .A(REG1_REG_16__SCAN_IN), .B(n4407), .S(n4612), .Z(U3534) );
  NAND2_X1 U4959 ( .A1(n4601), .A2(n4367), .ZN(n4369) );
  NAND2_X1 U4960 ( .A1(n4599), .A2(REG0_REG_31__SCAN_IN), .ZN(n4368) );
  OAI211_X1 U4961 ( .C1(n4370), .C2(n4404), .A(n4369), .B(n4368), .ZN(U3517)
         );
  INV_X1 U4962 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4371) );
  MUX2_X1 U4963 ( .A(n4424), .B(n4371), .S(n4599), .Z(n4372) );
  OAI21_X1 U4964 ( .B1(n4373), .B2(n4404), .A(n4372), .ZN(U3516) );
  INV_X1 U4965 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4375) );
  MUX2_X1 U4966 ( .A(n4375), .B(n4374), .S(n4601), .Z(n4376) );
  OAI21_X1 U4967 ( .B1(n4377), .B2(n4404), .A(n4376), .ZN(U3513) );
  INV_X1 U4968 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4379) );
  MUX2_X1 U4969 ( .A(n4379), .B(n4378), .S(n4601), .Z(n4380) );
  OAI21_X1 U4970 ( .B1(n4381), .B2(n4404), .A(n4380), .ZN(U3512) );
  INV_X1 U4971 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4383) );
  MUX2_X1 U4972 ( .A(n4383), .B(n4382), .S(n4601), .Z(n4384) );
  OAI21_X1 U4973 ( .B1(n4385), .B2(n4404), .A(n4384), .ZN(U3511) );
  INV_X1 U4974 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4725) );
  MUX2_X1 U4975 ( .A(n4725), .B(n4386), .S(n4601), .Z(n4387) );
  OAI21_X1 U4976 ( .B1(n4388), .B2(n4404), .A(n4387), .ZN(U3510) );
  INV_X1 U4977 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4390) );
  MUX2_X1 U4978 ( .A(n4390), .B(n4389), .S(n4601), .Z(n4391) );
  OAI21_X1 U4979 ( .B1(n4392), .B2(n4404), .A(n4391), .ZN(U3509) );
  INV_X1 U4980 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4718) );
  MUX2_X1 U4981 ( .A(n4718), .B(n4393), .S(n4601), .Z(n4394) );
  OAI21_X1 U4982 ( .B1(n4395), .B2(n4404), .A(n4394), .ZN(U3508) );
  INV_X1 U4983 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4397) );
  MUX2_X1 U4984 ( .A(n4397), .B(n4396), .S(n4601), .Z(n4398) );
  OAI21_X1 U4985 ( .B1(n4399), .B2(n4404), .A(n4398), .ZN(U3507) );
  MUX2_X1 U4986 ( .A(REG0_REG_20__SCAN_IN), .B(n4400), .S(n4601), .Z(U3506) );
  INV_X1 U4987 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4402) );
  MUX2_X1 U4988 ( .A(n4402), .B(n4401), .S(n4601), .Z(n4403) );
  OAI21_X1 U4989 ( .B1(n4405), .B2(n4404), .A(n4403), .ZN(U3505) );
  MUX2_X1 U4990 ( .A(REG0_REG_18__SCAN_IN), .B(n4406), .S(n4601), .Z(U3503) );
  MUX2_X1 U4991 ( .A(REG0_REG_16__SCAN_IN), .B(n4407), .S(n4601), .Z(U3499) );
  MUX2_X1 U4992 ( .A(n4408), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U4993 ( .A(n4409), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U4994 ( .A(n2789), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4995 ( .A(DATAI_25_), .B(n4410), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U4996 ( .A(DATAI_22_), .B(n4411), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4997 ( .A(n2735), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4998 ( .A(DATAI_20_), .B(n4412), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4999 ( .A(n4413), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5000 ( .A(n4414), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5001 ( .A(n4415), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5002 ( .A(n4416), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5003 ( .A(n4417), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5004 ( .A(DATAI_4_), .B(n4418), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5005 ( .A(n4419), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5006 ( .A(n4420), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5007 ( .A(n4421), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U5008 ( .A1(n4422), .A2(n4618), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4557), .ZN(n4423) );
  OAI21_X1 U5009 ( .B1(n4557), .B2(n4424), .A(n4423), .ZN(U3261) );
  AOI21_X1 U5010 ( .B1(n2457), .B2(n4426), .A(n4425), .ZN(n4427) );
  XOR2_X1 U5011 ( .A(n4427), .B(n2211), .Z(n4429) );
  AOI22_X1 U5012 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4498), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4428) );
  OAI21_X1 U5013 ( .B1(n4430), .B2(n4429), .A(n4428), .ZN(U3240) );
  OAI211_X1 U5014 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4432), .A(n4464), .B(n4431), 
        .ZN(n4433) );
  NAND2_X1 U5015 ( .A1(n4434), .A2(n4433), .ZN(n4435) );
  AOI21_X1 U5016 ( .B1(n4498), .B2(ADDR_REG_8__SCAN_IN), .A(n4435), .ZN(n4439)
         );
  OAI211_X1 U5017 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4437), .A(n4499), .B(n4436), 
        .ZN(n4438) );
  OAI211_X1 U5018 ( .C1(n4505), .C2(n4571), .A(n4439), .B(n4438), .ZN(U3248)
         );
  OAI211_X1 U5019 ( .C1(n4442), .C2(n4441), .A(n4499), .B(n4440), .ZN(n4447)
         );
  OAI211_X1 U5020 ( .C1(n4445), .C2(n4444), .A(n4464), .B(n4443), .ZN(n4446)
         );
  OAI211_X1 U5021 ( .C1(n4505), .C2(n4448), .A(n4447), .B(n4446), .ZN(n4449)
         );
  AOI211_X1 U5022 ( .C1(n4498), .C2(ADDR_REG_9__SCAN_IN), .A(n4450), .B(n4449), 
        .ZN(n4451) );
  INV_X1 U5023 ( .A(n4451), .ZN(U3249) );
  OAI211_X1 U5024 ( .C1(n4454), .C2(n4453), .A(n4499), .B(n4452), .ZN(n4459)
         );
  OAI211_X1 U5025 ( .C1(n4457), .C2(n4456), .A(n4464), .B(n4455), .ZN(n4458)
         );
  OAI211_X1 U5026 ( .C1(n4505), .C2(n4568), .A(n4459), .B(n4458), .ZN(n4460)
         );
  AOI211_X1 U5027 ( .C1(n4498), .C2(ADDR_REG_11__SCAN_IN), .A(n4461), .B(n4460), .ZN(n4462) );
  INV_X1 U5028 ( .A(n4462), .ZN(U3251) );
  OAI211_X1 U5029 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4465), .A(n4464), .B(n4463), .ZN(n4467) );
  NAND2_X1 U5030 ( .A1(n4467), .A2(n4466), .ZN(n4468) );
  AOI21_X1 U5031 ( .B1(n4498), .B2(ADDR_REG_12__SCAN_IN), .A(n4468), .ZN(n4472) );
  OAI211_X1 U5032 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4470), .A(n4499), .B(n4469), .ZN(n4471) );
  OAI211_X1 U5033 ( .C1(n4505), .C2(n4567), .A(n4472), .B(n4471), .ZN(U3252)
         );
  AOI211_X1 U5034 ( .C1(n4475), .C2(n4474), .A(n4473), .B(n4492), .ZN(n4476)
         );
  AOI211_X1 U5035 ( .C1(n4498), .C2(ADDR_REG_15__SCAN_IN), .A(n4477), .B(n4476), .ZN(n4482) );
  OAI211_X1 U5036 ( .C1(n4480), .C2(n4479), .A(n4499), .B(n4478), .ZN(n4481)
         );
  OAI211_X1 U5037 ( .C1(n4505), .C2(n4565), .A(n4482), .B(n4481), .ZN(U3255)
         );
  INV_X1 U5038 ( .A(n4483), .ZN(n4487) );
  AOI221_X1 U5039 ( .B1(n4485), .B2(n4484), .C1(n4922), .C2(n4484), .A(n4492), 
        .ZN(n4486) );
  AOI211_X1 U5040 ( .C1(n4498), .C2(ADDR_REG_16__SCAN_IN), .A(n4487), .B(n4486), .ZN(n4490) );
  OAI221_X1 U5041 ( .B1(n2185), .B2(REG1_REG_16__SCAN_IN), .C1(n2185), .C2(
        n4488), .A(n4499), .ZN(n4489) );
  OAI211_X1 U5042 ( .C1(n4505), .C2(n4491), .A(n4490), .B(n4489), .ZN(U3256)
         );
  AOI221_X1 U5043 ( .B1(n4495), .B2(n4494), .C1(n4493), .C2(n4494), .A(n4492), 
        .ZN(n4496) );
  AOI211_X1 U5044 ( .C1(n4498), .C2(ADDR_REG_17__SCAN_IN), .A(n4497), .B(n4496), .ZN(n4504) );
  OAI221_X1 U5045 ( .B1(n4502), .B2(n4501), .C1(n4502), .C2(n4500), .A(n4499), 
        .ZN(n4503) );
  OAI211_X1 U5046 ( .C1(n4505), .C2(n4562), .A(n4504), .B(n4503), .ZN(U3257)
         );
  AOI22_X1 U5047 ( .A1(n4506), .A2(n4549), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4557), .ZN(n4511) );
  INV_X1 U5048 ( .A(n4507), .ZN(n4508) );
  AOI22_X1 U5049 ( .A1(n4509), .A2(n4553), .B1(n4618), .B2(n4508), .ZN(n4510)
         );
  OAI211_X1 U5050 ( .C1(n4557), .C2(n4512), .A(n4511), .B(n4510), .ZN(U3280)
         );
  AOI22_X1 U5051 ( .A1(n4513), .A2(n4549), .B1(REG2_REG_8__SCAN_IN), .B2(n4557), .ZN(n4518) );
  INV_X1 U5052 ( .A(n4514), .ZN(n4515) );
  AOI22_X1 U5053 ( .A1(n4516), .A2(n4553), .B1(n4618), .B2(n4515), .ZN(n4517)
         );
  OAI211_X1 U5054 ( .C1(n4557), .C2(n4519), .A(n4518), .B(n4517), .ZN(U3282)
         );
  OAI22_X1 U5055 ( .A1(n4245), .A2(n2261), .B1(n4520), .B2(n4615), .ZN(n4521)
         );
  INV_X1 U5056 ( .A(n4521), .ZN(n4526) );
  INV_X1 U5057 ( .A(n4522), .ZN(n4523) );
  AOI22_X1 U5058 ( .A1(n4524), .A2(n4553), .B1(n4618), .B2(n4523), .ZN(n4525)
         );
  OAI211_X1 U5059 ( .C1(n4557), .C2(n4527), .A(n4526), .B(n4525), .ZN(U3284)
         );
  AOI22_X1 U5060 ( .A1(n4557), .A2(REG2_REG_3__SCAN_IN), .B1(n4549), .B2(n2469), .ZN(n4531) );
  AOI22_X1 U5061 ( .A1(n4529), .A2(n4553), .B1(n4618), .B2(n4528), .ZN(n4530)
         );
  OAI211_X1 U5062 ( .C1(n4557), .C2(n4532), .A(n4531), .B(n4530), .ZN(U3287)
         );
  OAI21_X1 U5063 ( .B1(n4543), .B2(n4534), .A(n4533), .ZN(n4547) );
  AOI22_X1 U5064 ( .A1(n2456), .A2(n4536), .B1(n4552), .B2(n4535), .ZN(n4537)
         );
  OAI21_X1 U5065 ( .B1(n4539), .B2(n4538), .A(n4537), .ZN(n4546) );
  INV_X1 U5066 ( .A(n4540), .ZN(n4541) );
  AOI21_X1 U5067 ( .B1(n4543), .B2(n4542), .A(n4541), .ZN(n4586) );
  NOR2_X1 U5068 ( .A1(n4586), .A2(n4544), .ZN(n4545) );
  AOI211_X1 U5069 ( .C1(n4548), .C2(n4547), .A(n4546), .B(n4545), .ZN(n4584)
         );
  AOI22_X1 U5070 ( .A1(REG3_REG_2__SCAN_IN), .A2(n4549), .B1(
        REG2_REG_2__SCAN_IN), .B2(n4557), .ZN(n4556) );
  INV_X1 U5071 ( .A(n4586), .ZN(n4554) );
  AOI21_X1 U5072 ( .B1(n4552), .B2(n4551), .A(n4550), .ZN(n4604) );
  AOI22_X1 U5073 ( .A1(n4554), .A2(n4553), .B1(n4618), .B2(n4604), .ZN(n4555)
         );
  OAI211_X1 U5074 ( .C1(n4557), .C2(n4584), .A(n4556), .B(n4555), .ZN(U3288)
         );
  INV_X1 U5075 ( .A(D_REG_31__SCAN_IN), .ZN(n4771) );
  NOR2_X1 U5076 ( .A1(n4558), .A2(n4771), .ZN(U3291) );
  AND2_X1 U5077 ( .A1(D_REG_30__SCAN_IN), .A2(n4559), .ZN(U3292) );
  INV_X1 U5078 ( .A(D_REG_29__SCAN_IN), .ZN(n4800) );
  NOR2_X1 U5079 ( .A1(n4558), .A2(n4800), .ZN(U3293) );
  AND2_X1 U5080 ( .A1(D_REG_28__SCAN_IN), .A2(n4559), .ZN(U3294) );
  AND2_X1 U5081 ( .A1(D_REG_27__SCAN_IN), .A2(n4559), .ZN(U3295) );
  INV_X1 U5082 ( .A(D_REG_26__SCAN_IN), .ZN(n4779) );
  NOR2_X1 U5083 ( .A1(n4558), .A2(n4779), .ZN(U3296) );
  AND2_X1 U5084 ( .A1(D_REG_25__SCAN_IN), .A2(n4559), .ZN(U3297) );
  AND2_X1 U5085 ( .A1(D_REG_24__SCAN_IN), .A2(n4559), .ZN(U3298) );
  AND2_X1 U5086 ( .A1(D_REG_23__SCAN_IN), .A2(n4559), .ZN(U3299) );
  NOR2_X1 U5087 ( .A1(n4558), .A2(n4752), .ZN(U3300) );
  AND2_X1 U5088 ( .A1(D_REG_21__SCAN_IN), .A2(n4559), .ZN(U3301) );
  INV_X1 U5089 ( .A(D_REG_20__SCAN_IN), .ZN(n4782) );
  NOR2_X1 U5090 ( .A1(n4558), .A2(n4782), .ZN(U3302) );
  INV_X1 U5091 ( .A(D_REG_19__SCAN_IN), .ZN(n4756) );
  NOR2_X1 U5092 ( .A1(n4558), .A2(n4756), .ZN(U3303) );
  AND2_X1 U5093 ( .A1(D_REG_18__SCAN_IN), .A2(n4559), .ZN(U3304) );
  AND2_X1 U5094 ( .A1(D_REG_17__SCAN_IN), .A2(n4559), .ZN(U3305) );
  NOR2_X1 U5095 ( .A1(n4558), .A2(n4747), .ZN(U3306) );
  AND2_X1 U5096 ( .A1(D_REG_15__SCAN_IN), .A2(n4559), .ZN(U3307) );
  NOR2_X1 U5097 ( .A1(n4558), .A2(n4749), .ZN(U3308) );
  INV_X1 U5098 ( .A(D_REG_13__SCAN_IN), .ZN(n4769) );
  NOR2_X1 U5099 ( .A1(n4558), .A2(n4769), .ZN(U3309) );
  AND2_X1 U5100 ( .A1(D_REG_12__SCAN_IN), .A2(n4559), .ZN(U3310) );
  AND2_X1 U5101 ( .A1(D_REG_11__SCAN_IN), .A2(n4559), .ZN(U3311) );
  NOR2_X1 U5102 ( .A1(n4558), .A2(n4753), .ZN(U3312) );
  AND2_X1 U5103 ( .A1(D_REG_9__SCAN_IN), .A2(n4559), .ZN(U3313) );
  AND2_X1 U5104 ( .A1(D_REG_8__SCAN_IN), .A2(n4559), .ZN(U3314) );
  INV_X1 U5105 ( .A(D_REG_7__SCAN_IN), .ZN(n4791) );
  NOR2_X1 U5106 ( .A1(n4558), .A2(n4791), .ZN(U3315) );
  INV_X1 U5107 ( .A(D_REG_6__SCAN_IN), .ZN(n4801) );
  NOR2_X1 U5108 ( .A1(n4558), .A2(n4801), .ZN(U3316) );
  AND2_X1 U5109 ( .A1(D_REG_5__SCAN_IN), .A2(n4559), .ZN(U3317) );
  INV_X1 U5110 ( .A(D_REG_4__SCAN_IN), .ZN(n4780) );
  NOR2_X1 U5111 ( .A1(n4558), .A2(n4780), .ZN(U3318) );
  AND2_X1 U5112 ( .A1(D_REG_3__SCAN_IN), .A2(n4559), .ZN(U3319) );
  AND2_X1 U5113 ( .A1(D_REG_2__SCAN_IN), .A2(n4559), .ZN(U3320) );
  INV_X1 U5114 ( .A(DATAI_23_), .ZN(n4919) );
  AOI21_X1 U5115 ( .B1(U3149), .B2(n4919), .A(n4560), .ZN(U3329) );
  AOI22_X1 U5116 ( .A1(STATE_REG_SCAN_IN), .A2(n4562), .B1(n4561), .B2(U3149), 
        .ZN(U3335) );
  OAI22_X1 U5117 ( .A1(U3149), .A2(n4563), .B1(DATAI_16_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4564) );
  INV_X1 U5118 ( .A(n4564), .ZN(U3336) );
  INV_X1 U5119 ( .A(DATAI_15_), .ZN(n4811) );
  AOI22_X1 U5120 ( .A1(STATE_REG_SCAN_IN), .A2(n4565), .B1(n4811), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5121 ( .A(DATAI_12_), .ZN(n4566) );
  AOI22_X1 U5122 ( .A1(STATE_REG_SCAN_IN), .A2(n4567), .B1(n4566), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5123 ( .A(DATAI_11_), .ZN(n4692) );
  AOI22_X1 U5124 ( .A1(STATE_REG_SCAN_IN), .A2(n4568), .B1(n4692), .B2(U3149), 
        .ZN(U3341) );
  OAI22_X1 U5125 ( .A1(U3149), .A2(n4569), .B1(DATAI_9_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4570) );
  INV_X1 U5126 ( .A(n4570), .ZN(U3343) );
  AOI22_X1 U5127 ( .A1(STATE_REG_SCAN_IN), .A2(n4571), .B1(n2529), .B2(U3149), 
        .ZN(U3344) );
  OAI22_X1 U5128 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4572) );
  INV_X1 U5129 ( .A(n4572), .ZN(U3352) );
  OAI211_X1 U5130 ( .C1(n4575), .C2(n4585), .A(n4574), .B(n4573), .ZN(n4576)
         );
  INV_X1 U5131 ( .A(n4576), .ZN(n4602) );
  INV_X1 U5132 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4776) );
  AOI22_X1 U5133 ( .A1(n4601), .A2(n4602), .B1(n4776), .B2(n4599), .ZN(U3467)
         );
  INV_X1 U5134 ( .A(n4577), .ZN(n4582) );
  OAI22_X1 U5135 ( .A1(n4580), .A2(n4585), .B1(n4579), .B2(n4578), .ZN(n4581)
         );
  NOR2_X1 U5136 ( .A1(n4582), .A2(n4581), .ZN(n4603) );
  INV_X1 U5137 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4583) );
  AOI22_X1 U5138 ( .A1(n4601), .A2(n4603), .B1(n4583), .B2(n4599), .ZN(U3469)
         );
  INV_X1 U5139 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4783) );
  OAI21_X1 U5140 ( .B1(n4586), .B2(n4585), .A(n4584), .ZN(n4606) );
  AOI22_X1 U5141 ( .A1(n4606), .A2(n4601), .B1(n4587), .B2(n4604), .ZN(n4588)
         );
  OAI21_X1 U5142 ( .B1(n4601), .B2(n4783), .A(n4588), .ZN(U3471) );
  INV_X1 U5143 ( .A(n4589), .ZN(n4591) );
  AOI211_X1 U5144 ( .C1(n4593), .C2(n4592), .A(n4591), .B(n4590), .ZN(n4609)
         );
  INV_X1 U5145 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4763) );
  AOI22_X1 U5146 ( .A1(n4601), .A2(n4609), .B1(n4763), .B2(n4599), .ZN(U3475)
         );
  NAND3_X1 U5147 ( .A1(n4595), .A2(n4594), .A3(n3067), .ZN(n4598) );
  AND3_X1 U5148 ( .A1(n4598), .A2(n4597), .A3(n4596), .ZN(n4611) );
  INV_X1 U5149 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4600) );
  AOI22_X1 U5150 ( .A1(n4601), .A2(n4611), .B1(n4600), .B2(n4599), .ZN(U3481)
         );
  AOI22_X1 U5151 ( .A1(n4612), .A2(n4602), .B1(n2457), .B2(n4610), .ZN(U3518)
         );
  AOI22_X1 U5152 ( .A1(n4612), .A2(n4603), .B1(n2451), .B2(n4610), .ZN(U3519)
         );
  AOI22_X1 U5153 ( .A1(n4606), .A2(n4612), .B1(n4605), .B2(n4604), .ZN(n4607)
         );
  OAI21_X1 U5154 ( .B1(n4612), .B2(n2442), .A(n4607), .ZN(U3520) );
  INV_X1 U5155 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4608) );
  AOI22_X1 U5156 ( .A1(n4612), .A2(n4609), .B1(n4608), .B2(n4610), .ZN(U3522)
         );
  AOI22_X1 U5157 ( .A1(n4612), .A2(n4611), .B1(n4831), .B2(n4610), .ZN(U3525)
         );
  INV_X1 U5158 ( .A(n4613), .ZN(n4622) );
  INV_X1 U5159 ( .A(n4614), .ZN(n4616) );
  OAI22_X1 U5160 ( .A1(n4245), .A2(n2887), .B1(n4616), .B2(n4615), .ZN(n4617)
         );
  AOI21_X1 U5161 ( .B1(n4619), .B2(n4618), .A(n4617), .ZN(n4620) );
  OAI21_X1 U5162 ( .B1(n4622), .B2(n4621), .A(n4620), .ZN(n4623) );
  AOI21_X1 U5163 ( .B1(n4245), .B2(n4624), .A(n4623), .ZN(n4938) );
  NAND2_X1 U5164 ( .A1(keyinput67), .A2(keyinput80), .ZN(n4625) );
  NOR3_X1 U5165 ( .A1(keyinput35), .A2(keyinput103), .A3(n4625), .ZN(n4626) );
  NAND3_X1 U5166 ( .A1(keyinput98), .A2(keyinput99), .A3(n4626), .ZN(n4639) );
  NOR4_X1 U5167 ( .A1(keyinput22), .A2(keyinput94), .A3(keyinput24), .A4(
        keyinput110), .ZN(n4637) );
  NAND2_X1 U5168 ( .A1(keyinput44), .A2(keyinput77), .ZN(n4627) );
  NOR3_X1 U5169 ( .A1(keyinput72), .A2(keyinput64), .A3(n4627), .ZN(n4636) );
  NOR2_X1 U5170 ( .A1(keyinput73), .A2(keyinput111), .ZN(n4628) );
  NAND3_X1 U5171 ( .A1(keyinput63), .A2(keyinput100), .A3(n4628), .ZN(n4634)
         );
  INV_X1 U5172 ( .A(keyinput86), .ZN(n4629) );
  NAND4_X1 U5173 ( .A1(keyinput84), .A2(keyinput93), .A3(keyinput105), .A4(
        n4629), .ZN(n4633) );
  NAND4_X1 U5174 ( .A1(keyinput46), .A2(keyinput116), .A3(keyinput3), .A4(
        keyinput6), .ZN(n4632) );
  NOR3_X1 U5175 ( .A1(keyinput30), .A2(keyinput9), .A3(keyinput104), .ZN(n4630) );
  NAND2_X1 U5176 ( .A1(keyinput65), .A2(n4630), .ZN(n4631) );
  NOR4_X1 U5177 ( .A1(n4634), .A2(n4633), .A3(n4632), .A4(n4631), .ZN(n4635)
         );
  NAND3_X1 U5178 ( .A1(n4637), .A2(n4636), .A3(n4635), .ZN(n4638) );
  NOR4_X1 U5179 ( .A1(keyinput79), .A2(keyinput8), .A3(n4639), .A4(n4638), 
        .ZN(n4688) );
  NOR2_X1 U5180 ( .A1(keyinput82), .A2(keyinput91), .ZN(n4640) );
  NAND3_X1 U5181 ( .A1(keyinput87), .A2(keyinput95), .A3(n4640), .ZN(n4686) );
  INV_X1 U5182 ( .A(keyinput66), .ZN(n4641) );
  NAND4_X1 U5183 ( .A1(keyinput59), .A2(keyinput71), .A3(keyinput78), .A4(
        n4641), .ZN(n4685) );
  INV_X1 U5184 ( .A(keyinput47), .ZN(n4642) );
  NOR4_X1 U5185 ( .A1(keyinput27), .A2(keyinput43), .A3(keyinput54), .A4(n4642), .ZN(n4653) );
  NAND2_X1 U5186 ( .A1(keyinput23), .A2(keyinput10), .ZN(n4643) );
  NOR3_X1 U5187 ( .A1(keyinput18), .A2(keyinput26), .A3(n4643), .ZN(n4652) );
  NOR2_X1 U5188 ( .A1(keyinput13), .A2(keyinput49), .ZN(n4644) );
  NAND3_X1 U5189 ( .A1(keyinput53), .A2(keyinput12), .A3(n4644), .ZN(n4650) );
  NAND4_X1 U5190 ( .A1(keyinput97), .A2(keyinput113), .A3(keyinput125), .A4(
        keyinput69), .ZN(n4649) );
  NOR2_X1 U5191 ( .A1(keyinput36), .A2(keyinput40), .ZN(n4645) );
  NAND3_X1 U5192 ( .A1(keyinput28), .A2(keyinput52), .A3(n4645), .ZN(n4648) );
  INV_X1 U5193 ( .A(keyinput88), .ZN(n4646) );
  NAND4_X1 U5194 ( .A1(keyinput96), .A2(keyinput124), .A3(keyinput92), .A4(
        n4646), .ZN(n4647) );
  NOR4_X1 U5195 ( .A1(n4650), .A2(n4649), .A3(n4648), .A4(n4647), .ZN(n4651)
         );
  NAND3_X1 U5196 ( .A1(n4653), .A2(n4652), .A3(n4651), .ZN(n4684) );
  INV_X1 U5197 ( .A(keyinput39), .ZN(n4656) );
  INV_X1 U5198 ( .A(keyinput38), .ZN(n4654) );
  NAND4_X1 U5199 ( .A1(keyinput107), .A2(keyinput16), .A3(keyinput68), .A4(
        n4654), .ZN(n4655) );
  NOR4_X1 U5200 ( .A1(keyinput60), .A2(keyinput5), .A3(n4656), .A4(n4655), 
        .ZN(n4682) );
  NOR4_X1 U5201 ( .A1(keyinput51), .A2(keyinput42), .A3(keyinput55), .A4(
        keyinput127), .ZN(n4657) );
  NAND3_X1 U5202 ( .A1(keyinput2), .A2(keyinput102), .A3(n4657), .ZN(n4664) );
  NAND2_X1 U5203 ( .A1(keyinput112), .A2(keyinput85), .ZN(n4658) );
  NOR3_X1 U5204 ( .A1(keyinput41), .A2(keyinput14), .A3(n4658), .ZN(n4662) );
  NOR4_X1 U5205 ( .A1(keyinput114), .A2(keyinput123), .A3(keyinput7), .A4(
        keyinput31), .ZN(n4661) );
  NOR4_X1 U5206 ( .A1(keyinput89), .A2(keyinput90), .A3(keyinput11), .A4(
        keyinput119), .ZN(n4660) );
  AND4_X1 U5207 ( .A1(keyinput76), .A2(keyinput122), .A3(keyinput48), .A4(
        keyinput62), .ZN(n4659) );
  NAND4_X1 U5208 ( .A1(n4662), .A2(n4661), .A3(n4660), .A4(n4659), .ZN(n4663)
         );
  NOR4_X1 U5209 ( .A1(keyinput25), .A2(keyinput1), .A3(n4664), .A4(n4663), 
        .ZN(n4681) );
  NAND4_X1 U5210 ( .A1(keyinput126), .A2(keyinput108), .A3(keyinput120), .A4(
        keyinput117), .ZN(n4671) );
  NOR2_X1 U5211 ( .A1(keyinput34), .A2(keyinput56), .ZN(n4665) );
  NAND3_X1 U5212 ( .A1(keyinput70), .A2(keyinput57), .A3(n4665), .ZN(n4670) );
  INV_X1 U5213 ( .A(keyinput81), .ZN(n4666) );
  NAND4_X1 U5214 ( .A1(keyinput17), .A2(keyinput32), .A3(keyinput33), .A4(
        n4666), .ZN(n4669) );
  NOR2_X1 U5215 ( .A1(keyinput58), .A2(keyinput118), .ZN(n4667) );
  NAND3_X1 U5216 ( .A1(keyinput106), .A2(keyinput83), .A3(n4667), .ZN(n4668)
         );
  NOR4_X1 U5217 ( .A1(n4671), .A2(n4670), .A3(n4669), .A4(n4668), .ZN(n4680)
         );
  INV_X1 U5218 ( .A(keyinput20), .ZN(n4672) );
  NAND4_X1 U5219 ( .A1(keyinput0), .A2(keyinput37), .A3(keyinput4), .A4(n4672), 
        .ZN(n4678) );
  OR4_X1 U5220 ( .A1(keyinput115), .A2(keyinput21), .A3(keyinput61), .A4(
        keyinput109), .ZN(n4677) );
  NOR2_X1 U5221 ( .A1(keyinput19), .A2(keyinput101), .ZN(n4673) );
  NAND3_X1 U5222 ( .A1(keyinput75), .A2(keyinput45), .A3(n4673), .ZN(n4676) );
  NOR2_X1 U5223 ( .A1(keyinput50), .A2(keyinput15), .ZN(n4674) );
  NAND3_X1 U5224 ( .A1(keyinput74), .A2(keyinput29), .A3(n4674), .ZN(n4675) );
  NOR4_X1 U5225 ( .A1(n4678), .A2(n4677), .A3(n4676), .A4(n4675), .ZN(n4679)
         );
  NAND4_X1 U5226 ( .A1(n4682), .A2(n4681), .A3(n4680), .A4(n4679), .ZN(n4683)
         );
  NOR4_X1 U5227 ( .A1(n4686), .A2(n4685), .A3(n4684), .A4(n4683), .ZN(n4687)
         );
  AOI21_X1 U5228 ( .B1(n4688), .B2(n4687), .A(keyinput121), .ZN(n4936) );
  INV_X1 U5229 ( .A(IR_REG_8__SCAN_IN), .ZN(n4690) );
  AOI22_X1 U5230 ( .A1(n2529), .A2(keyinput21), .B1(n4690), .B2(keyinput61), 
        .ZN(n4689) );
  OAI221_X1 U5231 ( .B1(n2529), .B2(keyinput21), .C1(n4690), .C2(keyinput61), 
        .A(n4689), .ZN(n4701) );
  AOI22_X1 U5232 ( .A1(n2533), .A2(keyinput109), .B1(keyinput37), .B2(n4692), 
        .ZN(n4691) );
  OAI221_X1 U5233 ( .B1(n2533), .B2(keyinput109), .C1(n4692), .C2(keyinput37), 
        .A(n4691), .ZN(n4700) );
  INV_X1 U5234 ( .A(keyinput4), .ZN(n4694) );
  AOI22_X1 U5235 ( .A1(n3340), .A2(keyinput0), .B1(DATAO_REG_16__SCAN_IN), 
        .B2(n4694), .ZN(n4693) );
  OAI221_X1 U5236 ( .B1(n3340), .B2(keyinput0), .C1(n4694), .C2(
        DATAO_REG_16__SCAN_IN), .A(n4693), .ZN(n4699) );
  INV_X1 U5237 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4697) );
  INV_X1 U5238 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4696) );
  AOI22_X1 U5239 ( .A1(n4697), .A2(keyinput20), .B1(n4696), .B2(keyinput50), 
        .ZN(n4695) );
  OAI221_X1 U5240 ( .B1(n4697), .B2(keyinput20), .C1(n4696), .C2(keyinput50), 
        .A(n4695), .ZN(n4698) );
  NOR4_X1 U5241 ( .A1(n4701), .A2(n4700), .A3(n4699), .A4(n4698), .ZN(n4744)
         );
  AOI22_X1 U5242 ( .A1(n3544), .A2(keyinput74), .B1(n4703), .B2(keyinput29), 
        .ZN(n4702) );
  OAI221_X1 U5243 ( .B1(n3544), .B2(keyinput74), .C1(n4703), .C2(keyinput29), 
        .A(n4702), .ZN(n4715) );
  INV_X1 U5244 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4706) );
  INV_X1 U5245 ( .A(keyinput15), .ZN(n4705) );
  AOI22_X1 U5246 ( .A1(n4706), .A2(keyinput19), .B1(DATAO_REG_18__SCAN_IN), 
        .B2(n4705), .ZN(n4704) );
  OAI221_X1 U5247 ( .B1(n4706), .B2(keyinput19), .C1(n4705), .C2(
        DATAO_REG_18__SCAN_IN), .A(n4704), .ZN(n4714) );
  INV_X1 U5248 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4708) );
  AOI22_X1 U5249 ( .A1(n4709), .A2(keyinput75), .B1(keyinput101), .B2(n4708), 
        .ZN(n4707) );
  OAI221_X1 U5250 ( .B1(n4709), .B2(keyinput75), .C1(n4708), .C2(keyinput101), 
        .A(n4707), .ZN(n4713) );
  INV_X1 U5251 ( .A(keyinput34), .ZN(n4711) );
  AOI22_X1 U5252 ( .A1(n4339), .A2(keyinput45), .B1(DATAO_REG_22__SCAN_IN), 
        .B2(n4711), .ZN(n4710) );
  OAI221_X1 U5253 ( .B1(n4339), .B2(keyinput45), .C1(n4711), .C2(
        DATAO_REG_22__SCAN_IN), .A(n4710), .ZN(n4712) );
  NOR4_X1 U5254 ( .A1(n4715), .A2(n4714), .A3(n4713), .A4(n4712), .ZN(n4743)
         );
  AOI22_X1 U5255 ( .A1(n4718), .A2(keyinput70), .B1(n4717), .B2(keyinput57), 
        .ZN(n4716) );
  OAI221_X1 U5256 ( .B1(n4718), .B2(keyinput70), .C1(n4717), .C2(keyinput57), 
        .A(n4716), .ZN(n4729) );
  INV_X1 U5257 ( .A(keyinput56), .ZN(n4720) );
  AOI22_X1 U5258 ( .A1(n4390), .A2(keyinput126), .B1(DATAO_REG_23__SCAN_IN), 
        .B2(n4720), .ZN(n4719) );
  OAI221_X1 U5259 ( .B1(n4390), .B2(keyinput126), .C1(n4720), .C2(
        DATAO_REG_23__SCAN_IN), .A(n4719), .ZN(n4728) );
  INV_X1 U5260 ( .A(keyinput120), .ZN(n4722) );
  AOI22_X1 U5261 ( .A1(n4325), .A2(keyinput108), .B1(DATAO_REG_24__SCAN_IN), 
        .B2(n4722), .ZN(n4721) );
  OAI221_X1 U5262 ( .B1(n4325), .B2(keyinput108), .C1(n4722), .C2(
        DATAO_REG_24__SCAN_IN), .A(n4721), .ZN(n4727) );
  AOI22_X1 U5263 ( .A1(n4725), .A2(keyinput117), .B1(n4724), .B2(keyinput106), 
        .ZN(n4723) );
  OAI221_X1 U5264 ( .B1(n4725), .B2(keyinput117), .C1(n4724), .C2(keyinput106), 
        .A(n4723), .ZN(n4726) );
  NOR4_X1 U5265 ( .A1(n4729), .A2(n4728), .A3(n4727), .A4(n4726), .ZN(n4742)
         );
  INV_X1 U5266 ( .A(keyinput58), .ZN(n4731) );
  AOI22_X1 U5267 ( .A1(n4383), .A2(keyinput118), .B1(DATAO_REG_26__SCAN_IN), 
        .B2(n4731), .ZN(n4730) );
  OAI221_X1 U5268 ( .B1(n4383), .B2(keyinput118), .C1(n4731), .C2(
        DATAO_REG_26__SCAN_IN), .A(n4730), .ZN(n4740) );
  INV_X1 U5269 ( .A(keyinput17), .ZN(n4733) );
  AOI22_X1 U5270 ( .A1(n4375), .A2(keyinput83), .B1(DATAO_REG_28__SCAN_IN), 
        .B2(n4733), .ZN(n4732) );
  OAI221_X1 U5271 ( .B1(n4375), .B2(keyinput83), .C1(n4733), .C2(
        DATAO_REG_28__SCAN_IN), .A(n4732), .ZN(n4739) );
  AOI22_X1 U5272 ( .A1(n2829), .A2(keyinput81), .B1(n2823), .B2(keyinput32), 
        .ZN(n4734) );
  OAI221_X1 U5273 ( .B1(n2829), .B2(keyinput81), .C1(n2823), .C2(keyinput32), 
        .A(n4734), .ZN(n4738) );
  AOI22_X1 U5274 ( .A1(n4285), .A2(keyinput33), .B1(n4736), .B2(keyinput10), 
        .ZN(n4735) );
  OAI221_X1 U5275 ( .B1(n4285), .B2(keyinput33), .C1(n4736), .C2(keyinput10), 
        .A(n4735), .ZN(n4737) );
  NOR4_X1 U5276 ( .A1(n4740), .A2(n4739), .A3(n4738), .A4(n4737), .ZN(n4741)
         );
  NAND4_X1 U5277 ( .A1(n4744), .A2(n4743), .A3(n4742), .A4(n4741), .ZN(n4934)
         );
  INV_X1 U5278 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4746) );
  AOI22_X1 U5279 ( .A1(n4747), .A2(keyinput18), .B1(keyinput23), .B2(n4746), 
        .ZN(n4745) );
  OAI221_X1 U5280 ( .B1(n4747), .B2(keyinput18), .C1(n4746), .C2(keyinput23), 
        .A(n4745), .ZN(n4760) );
  AOI22_X1 U5281 ( .A1(n4750), .A2(keyinput26), .B1(n4749), .B2(keyinput27), 
        .ZN(n4748) );
  OAI221_X1 U5282 ( .B1(n4750), .B2(keyinput26), .C1(n4749), .C2(keyinput27), 
        .A(n4748), .ZN(n4759) );
  AOI22_X1 U5283 ( .A1(n4753), .A2(keyinput43), .B1(keyinput47), .B2(n4752), 
        .ZN(n4751) );
  OAI221_X1 U5284 ( .B1(n4753), .B2(keyinput43), .C1(n4752), .C2(keyinput47), 
        .A(n4751), .ZN(n4758) );
  AOI22_X1 U5285 ( .A1(n4756), .A2(keyinput54), .B1(keyinput59), .B2(n4755), 
        .ZN(n4754) );
  OAI221_X1 U5286 ( .B1(n4756), .B2(keyinput54), .C1(n4755), .C2(keyinput59), 
        .A(n4754), .ZN(n4757) );
  NOR4_X1 U5287 ( .A1(n4760), .A2(n4759), .A3(n4758), .A4(n4757), .ZN(n4808)
         );
  XOR2_X1 U5288 ( .A(DATAI_13_), .B(keyinput95), .Z(n4767) );
  XNOR2_X1 U5289 ( .A(IR_REG_30__SCAN_IN), .B(keyinput78), .ZN(n4762) );
  XNOR2_X1 U5290 ( .A(DATAI_3_), .B(keyinput66), .ZN(n4761) );
  NAND2_X1 U5291 ( .A1(n4762), .A2(n4761), .ZN(n4766) );
  XNOR2_X1 U5292 ( .A(n2420), .B(keyinput97), .ZN(n4765) );
  XNOR2_X1 U5293 ( .A(keyinput71), .B(n4763), .ZN(n4764) );
  OR4_X1 U5294 ( .A1(n4767), .A2(n4766), .A3(n4765), .A4(n4764), .ZN(n4774) );
  AOI22_X1 U5295 ( .A1(n4770), .A2(keyinput87), .B1(n4769), .B2(keyinput91), 
        .ZN(n4768) );
  OAI221_X1 U5296 ( .B1(n4770), .B2(keyinput87), .C1(n4769), .C2(keyinput91), 
        .A(n4768), .ZN(n4773) );
  XNOR2_X1 U5297 ( .A(n4771), .B(keyinput82), .ZN(n4772) );
  NOR3_X1 U5298 ( .A1(n4774), .A2(n4773), .A3(n4772), .ZN(n4807) );
  AOI22_X1 U5299 ( .A1(n4777), .A2(keyinput69), .B1(keyinput13), .B2(n4776), 
        .ZN(n4775) );
  OAI221_X1 U5300 ( .B1(n4777), .B2(keyinput69), .C1(n4776), .C2(keyinput13), 
        .A(n4775), .ZN(n4789) );
  AOI22_X1 U5301 ( .A1(n4780), .A2(keyinput113), .B1(keyinput125), .B2(n4779), 
        .ZN(n4778) );
  OAI221_X1 U5302 ( .B1(n4780), .B2(keyinput113), .C1(n4779), .C2(keyinput125), 
        .A(n4778), .ZN(n4788) );
  AOI22_X1 U5303 ( .A1(n4783), .A2(keyinput53), .B1(n4782), .B2(keyinput49), 
        .ZN(n4781) );
  OAI221_X1 U5304 ( .B1(n4783), .B2(keyinput53), .C1(n4782), .C2(keyinput49), 
        .A(n4781), .ZN(n4787) );
  XNOR2_X1 U5305 ( .A(IR_REG_28__SCAN_IN), .B(keyinput124), .ZN(n4785) );
  XNOR2_X1 U5306 ( .A(IR_REG_6__SCAN_IN), .B(keyinput12), .ZN(n4784) );
  NAND2_X1 U5307 ( .A1(n4785), .A2(n4784), .ZN(n4786) );
  NOR4_X1 U5308 ( .A1(n4789), .A2(n4788), .A3(n4787), .A4(n4786), .ZN(n4806)
         );
  INV_X1 U5309 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4792) );
  AOI22_X1 U5310 ( .A1(n4792), .A2(keyinput92), .B1(n4791), .B2(keyinput28), 
        .ZN(n4790) );
  OAI221_X1 U5311 ( .B1(n4792), .B2(keyinput92), .C1(n4791), .C2(keyinput28), 
        .A(n4790), .ZN(n4799) );
  INV_X1 U5312 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4794) );
  AOI22_X1 U5313 ( .A1(n2222), .A2(keyinput60), .B1(keyinput40), .B2(n4794), 
        .ZN(n4793) );
  OAI221_X1 U5314 ( .B1(n2222), .B2(keyinput60), .C1(n4794), .C2(keyinput40), 
        .A(n4793), .ZN(n4798) );
  XNOR2_X1 U5315 ( .A(n4795), .B(keyinput96), .ZN(n4797) );
  XNOR2_X1 U5316 ( .A(n2477), .B(keyinput52), .ZN(n4796) );
  OR4_X1 U5317 ( .A1(n4799), .A2(n4798), .A3(n4797), .A4(n4796), .ZN(n4804) );
  XNOR2_X1 U5318 ( .A(n4800), .B(keyinput88), .ZN(n4803) );
  XNOR2_X1 U5319 ( .A(n4801), .B(keyinput36), .ZN(n4802) );
  NOR3_X1 U5320 ( .A1(n4804), .A2(n4803), .A3(n4802), .ZN(n4805) );
  NAND4_X1 U5321 ( .A1(n4808), .A2(n4807), .A3(n4806), .A4(n4805), .ZN(n4933)
         );
  AOI22_X1 U5322 ( .A1(n4811), .A2(keyinput110), .B1(keyinput86), .B2(n4810), 
        .ZN(n4809) );
  OAI221_X1 U5323 ( .B1(n4811), .B2(keyinput110), .C1(n4810), .C2(keyinput86), 
        .A(n4809), .ZN(n4823) );
  AOI22_X1 U5324 ( .A1(n4814), .A2(keyinput94), .B1(n4813), .B2(keyinput24), 
        .ZN(n4812) );
  OAI221_X1 U5325 ( .B1(n4814), .B2(keyinput94), .C1(n4813), .C2(keyinput24), 
        .A(n4812), .ZN(n4822) );
  INV_X1 U5326 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4817) );
  AOI22_X1 U5327 ( .A1(n4817), .A2(keyinput77), .B1(keyinput64), .B2(n4816), 
        .ZN(n4815) );
  OAI221_X1 U5328 ( .B1(n4817), .B2(keyinput77), .C1(n4816), .C2(keyinput64), 
        .A(n4815), .ZN(n4821) );
  XNOR2_X1 U5329 ( .A(REG2_REG_2__SCAN_IN), .B(keyinput22), .ZN(n4819) );
  XNOR2_X1 U5330 ( .A(REG2_REG_0__SCAN_IN), .B(keyinput44), .ZN(n4818) );
  NAND2_X1 U5331 ( .A1(n4819), .A2(n4818), .ZN(n4820) );
  NOR4_X1 U5332 ( .A1(n4823), .A2(n4822), .A3(n4821), .A4(n4820), .ZN(n4866)
         );
  INV_X1 U5333 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4825) );
  AOI22_X1 U5334 ( .A1(n4826), .A2(keyinput99), .B1(keyinput103), .B2(n4825), 
        .ZN(n4824) );
  OAI221_X1 U5335 ( .B1(n4826), .B2(keyinput99), .C1(n4825), .C2(keyinput103), 
        .A(n4824), .ZN(n4837) );
  INV_X1 U5336 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4828) );
  AOI22_X1 U5337 ( .A1(n4829), .A2(keyinput80), .B1(n4828), .B2(keyinput98), 
        .ZN(n4827) );
  OAI221_X1 U5338 ( .B1(n4829), .B2(keyinput80), .C1(n4828), .C2(keyinput98), 
        .A(n4827), .ZN(n4836) );
  AOI22_X1 U5339 ( .A1(n3343), .A2(keyinput8), .B1(keyinput72), .B2(n4831), 
        .ZN(n4830) );
  OAI221_X1 U5340 ( .B1(n3343), .B2(keyinput8), .C1(n4831), .C2(keyinput72), 
        .A(n4830), .ZN(n4835) );
  AOI22_X1 U5341 ( .A1(n4833), .A2(keyinput67), .B1(keyinput79), .B2(n3452), 
        .ZN(n4832) );
  OAI221_X1 U5342 ( .B1(n4833), .B2(keyinput67), .C1(n3452), .C2(keyinput79), 
        .A(n4832), .ZN(n4834) );
  NOR4_X1 U5343 ( .A1(n4837), .A2(n4836), .A3(n4835), .A4(n4834), .ZN(n4865)
         );
  AOI22_X1 U5344 ( .A1(n2509), .A2(keyinput9), .B1(keyinput115), .B2(n4839), 
        .ZN(n4838) );
  OAI221_X1 U5345 ( .B1(n2509), .B2(keyinput9), .C1(n4839), .C2(keyinput115), 
        .A(n4838), .ZN(n4850) );
  INV_X1 U5346 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4841) );
  AOI22_X1 U5347 ( .A1(n4841), .A2(keyinput104), .B1(n3374), .B2(keyinput46), 
        .ZN(n4840) );
  OAI221_X1 U5348 ( .B1(n4841), .B2(keyinput104), .C1(n3374), .C2(keyinput46), 
        .A(n4840), .ZN(n4849) );
  INV_X1 U5349 ( .A(DATAI_7_), .ZN(n4844) );
  AOI22_X1 U5350 ( .A1(n4844), .A2(keyinput6), .B1(n4843), .B2(keyinput65), 
        .ZN(n4842) );
  OAI221_X1 U5351 ( .B1(n4844), .B2(keyinput6), .C1(n4843), .C2(keyinput65), 
        .A(n4842), .ZN(n4848) );
  XNOR2_X1 U5352 ( .A(IR_REG_13__SCAN_IN), .B(keyinput116), .ZN(n4846) );
  XNOR2_X1 U5353 ( .A(IR_REG_10__SCAN_IN), .B(keyinput3), .ZN(n4845) );
  NAND2_X1 U5354 ( .A1(n4846), .A2(n4845), .ZN(n4847) );
  NOR4_X1 U5355 ( .A1(n4850), .A2(n4849), .A3(n4848), .A4(n4847), .ZN(n4864)
         );
  AOI22_X1 U5356 ( .A1(n2850), .A2(keyinput105), .B1(keyinput73), .B2(n2599), 
        .ZN(n4851) );
  OAI221_X1 U5357 ( .B1(n2850), .B2(keyinput105), .C1(n2599), .C2(keyinput73), 
        .A(n4851), .ZN(n4862) );
  AOI22_X1 U5358 ( .A1(n4853), .A2(keyinput84), .B1(n3570), .B2(keyinput93), 
        .ZN(n4852) );
  OAI221_X1 U5359 ( .B1(n4853), .B2(keyinput84), .C1(n3570), .C2(keyinput93), 
        .A(n4852), .ZN(n4861) );
  INV_X1 U5360 ( .A(IR_REG_12__SCAN_IN), .ZN(n4856) );
  AOI22_X1 U5361 ( .A1(n4856), .A2(keyinput111), .B1(keyinput30), .B2(n4855), 
        .ZN(n4854) );
  OAI221_X1 U5362 ( .B1(n4856), .B2(keyinput111), .C1(n4855), .C2(keyinput30), 
        .A(n4854), .ZN(n4860) );
  XNOR2_X1 U5363 ( .A(REG1_REG_14__SCAN_IN), .B(keyinput63), .ZN(n4858) );
  XNOR2_X1 U5364 ( .A(IR_REG_14__SCAN_IN), .B(keyinput100), .ZN(n4857) );
  NAND2_X1 U5365 ( .A1(n4858), .A2(n4857), .ZN(n4859) );
  NOR4_X1 U5366 ( .A1(n4862), .A2(n4861), .A3(n4860), .A4(n4859), .ZN(n4863)
         );
  NAND4_X1 U5367 ( .A1(n4866), .A2(n4865), .A3(n4864), .A4(n4863), .ZN(n4932)
         );
  INV_X1 U5368 ( .A(keyinput42), .ZN(n4869) );
  INV_X1 U5369 ( .A(keyinput2), .ZN(n4868) );
  AOI22_X1 U5370 ( .A1(n4869), .A2(DATAO_REG_13__SCAN_IN), .B1(
        DATAO_REG_9__SCAN_IN), .B2(n4868), .ZN(n4867) );
  OAI221_X1 U5371 ( .B1(n4869), .B2(DATAO_REG_13__SCAN_IN), .C1(n4868), .C2(
        DATAO_REG_9__SCAN_IN), .A(n4867), .ZN(n4882) );
  INV_X1 U5372 ( .A(keyinput1), .ZN(n4872) );
  INV_X1 U5373 ( .A(keyinput51), .ZN(n4871) );
  AOI22_X1 U5374 ( .A1(n4872), .A2(DATAO_REG_12__SCAN_IN), .B1(
        DATAO_REG_1__SCAN_IN), .B2(n4871), .ZN(n4870) );
  OAI221_X1 U5375 ( .B1(n4872), .B2(DATAO_REG_12__SCAN_IN), .C1(n4871), .C2(
        DATAO_REG_1__SCAN_IN), .A(n4870), .ZN(n4881) );
  INV_X1 U5376 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4874) );
  AOI22_X1 U5377 ( .A1(n4875), .A2(keyinput127), .B1(n4874), .B2(keyinput114), 
        .ZN(n4873) );
  OAI221_X1 U5378 ( .B1(n4875), .B2(keyinput127), .C1(n4874), .C2(keyinput114), 
        .A(n4873), .ZN(n4880) );
  INV_X1 U5379 ( .A(keyinput102), .ZN(n4878) );
  INV_X1 U5380 ( .A(keyinput55), .ZN(n4877) );
  AOI22_X1 U5381 ( .A1(n4878), .A2(DATAO_REG_15__SCAN_IN), .B1(
        DATAO_REG_7__SCAN_IN), .B2(n4877), .ZN(n4876) );
  OAI221_X1 U5382 ( .B1(n4878), .B2(DATAO_REG_15__SCAN_IN), .C1(n4877), .C2(
        DATAO_REG_7__SCAN_IN), .A(n4876), .ZN(n4879) );
  NOR4_X1 U5383 ( .A1(n4882), .A2(n4881), .A3(n4880), .A4(n4879), .ZN(n4930)
         );
  XNOR2_X1 U5384 ( .A(keyinput16), .B(ADDR_REG_19__SCAN_IN), .ZN(n4883) );
  OAI21_X1 U5385 ( .B1(keyinput121), .B2(n4884), .A(n4883), .ZN(n4897) );
  INV_X1 U5386 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4887) );
  AOI22_X1 U5387 ( .A1(n4887), .A2(keyinput39), .B1(n4886), .B2(keyinput5), 
        .ZN(n4885) );
  OAI221_X1 U5388 ( .B1(n4887), .B2(keyinput39), .C1(n4886), .C2(keyinput5), 
        .A(n4885), .ZN(n4896) );
  INV_X1 U5389 ( .A(REG2_REG_3__SCAN_IN), .ZN(n4890) );
  INV_X1 U5390 ( .A(keyinput25), .ZN(n4889) );
  AOI22_X1 U5391 ( .A1(n4890), .A2(keyinput68), .B1(DATAO_REG_0__SCAN_IN), 
        .B2(n4889), .ZN(n4888) );
  OAI221_X1 U5392 ( .B1(n4890), .B2(keyinput68), .C1(n4889), .C2(
        DATAO_REG_0__SCAN_IN), .A(n4888), .ZN(n4895) );
  INV_X1 U5393 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4892) );
  AOI22_X1 U5394 ( .A1(n4893), .A2(keyinput107), .B1(n4892), .B2(keyinput38), 
        .ZN(n4891) );
  OAI221_X1 U5395 ( .B1(n4893), .B2(keyinput107), .C1(n4892), .C2(keyinput38), 
        .A(n4891), .ZN(n4894) );
  NOR4_X1 U5396 ( .A1(n4897), .A2(n4896), .A3(n4895), .A4(n4894), .ZN(n4929)
         );
  INV_X1 U5397 ( .A(keyinput62), .ZN(n4900) );
  INV_X1 U5398 ( .A(keyinput89), .ZN(n4899) );
  AOI22_X1 U5399 ( .A1(n4900), .A2(ADDR_REG_4__SCAN_IN), .B1(
        ADDR_REG_8__SCAN_IN), .B2(n4899), .ZN(n4898) );
  OAI221_X1 U5400 ( .B1(n4900), .B2(ADDR_REG_4__SCAN_IN), .C1(n4899), .C2(
        ADDR_REG_8__SCAN_IN), .A(n4898), .ZN(n4911) );
  AOI22_X1 U5401 ( .A1(n2469), .A2(keyinput122), .B1(n2211), .B2(keyinput48), 
        .ZN(n4901) );
  INV_X1 U5402 ( .A(REG2_REG_10__SCAN_IN), .ZN(n4904) );
  INV_X1 U5403 ( .A(keyinput35), .ZN(n4903) );
  AOI22_X1 U5404 ( .A1(n4904), .A2(keyinput119), .B1(ADDR_REG_10__SCAN_IN), 
        .B2(n4903), .ZN(n4902) );
  OAI221_X1 U5405 ( .B1(n4904), .B2(keyinput119), .C1(n4903), .C2(
        ADDR_REG_10__SCAN_IN), .A(n4902), .ZN(n4909) );
  INV_X1 U5406 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4907) );
  INV_X1 U5407 ( .A(keyinput11), .ZN(n4906) );
  AOI22_X1 U5408 ( .A1(n4907), .A2(keyinput90), .B1(ADDR_REG_9__SCAN_IN), .B2(
        n4906), .ZN(n4905) );
  OAI221_X1 U5409 ( .B1(n4907), .B2(keyinput90), .C1(n4906), .C2(
        ADDR_REG_9__SCAN_IN), .A(n4905), .ZN(n4908) );
  NOR4_X1 U5410 ( .A1(n4911), .A2(n4910), .A3(n4909), .A4(n4908), .ZN(n4928)
         );
  INV_X1 U5411 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4913) );
  AOI22_X1 U5412 ( .A1(n4913), .A2(keyinput41), .B1(n4280), .B2(keyinput7), 
        .ZN(n4912) );
  OAI221_X1 U5413 ( .B1(n4913), .B2(keyinput41), .C1(n4280), .C2(keyinput7), 
        .A(n4912), .ZN(n4926) );
  INV_X1 U5414 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4916) );
  INV_X1 U5415 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4915) );
  AOI22_X1 U5416 ( .A1(n4916), .A2(keyinput123), .B1(n4915), .B2(keyinput85), 
        .ZN(n4914) );
  OAI221_X1 U5417 ( .B1(n4916), .B2(keyinput123), .C1(n4915), .C2(keyinput85), 
        .A(n4914), .ZN(n4925) );
  AOI22_X1 U5418 ( .A1(n4919), .A2(keyinput14), .B1(keyinput76), .B2(n4918), 
        .ZN(n4917) );
  OAI221_X1 U5419 ( .B1(n4919), .B2(keyinput14), .C1(n4918), .C2(keyinput76), 
        .A(n4917), .ZN(n4924) );
  AOI22_X1 U5420 ( .A1(n4922), .A2(keyinput31), .B1(keyinput112), .B2(n4921), 
        .ZN(n4920) );
  OAI221_X1 U5421 ( .B1(n4922), .B2(keyinput31), .C1(n4921), .C2(keyinput112), 
        .A(n4920), .ZN(n4923) );
  NOR4_X1 U5422 ( .A1(n4926), .A2(n4925), .A3(n4924), .A4(n4923), .ZN(n4927)
         );
  NAND4_X1 U5423 ( .A1(n4930), .A2(n4929), .A3(n4928), .A4(n4927), .ZN(n4931)
         );
  NOR4_X1 U5424 ( .A1(n4934), .A2(n4933), .A3(n4932), .A4(n4931), .ZN(n4935)
         );
  OAI21_X1 U5425 ( .B1(DATAO_REG_29__SCAN_IN), .B2(n4936), .A(n4935), .ZN(
        n4937) );
  XOR2_X1 U5426 ( .A(n4938), .B(n4937), .Z(U3285) );
  NAND2_X4 U2468 ( .A1(n2441), .A2(n2440), .ZN(n2465) );
endmodule

