

module b20_C_SARLock_k_64_1 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137;

  XNOR2_X1 U4829 ( .A(n8494), .B(n9764), .ZN(n9773) );
  AND2_X1 U4830 ( .A1(n6669), .A2(n6908), .ZN(n6670) );
  INV_X1 U4831 ( .A(n7826), .ZN(n7847) );
  AND2_X1 U4832 ( .A1(n4700), .A2(n9705), .ZN(n6589) );
  INV_X1 U4833 ( .A(n6081), .ZN(n5786) );
  INV_X1 U4834 ( .A(n6565), .ZN(n8588) );
  AND2_X1 U4835 ( .A1(n6152), .A2(n8163), .ZN(n6514) );
  CLKBUF_X2 U4836 ( .A(n5713), .Z(n4332) );
  BUF_X1 U4837 ( .A(n5807), .Z(n4329) );
  INV_X1 U4838 ( .A(n5081), .ZN(n8948) );
  NAND2_X1 U4839 ( .A1(n4814), .A2(n5106), .ZN(n5171) );
  AND2_X1 U4840 ( .A1(n5025), .A2(n5201), .ZN(n5235) );
  NOR2_X1 U4841 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5025) );
  INV_X1 U4842 ( .A(n5727), .ZN(n6081) );
  OR2_X1 U4843 ( .A1(n5446), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5453) );
  INV_X1 U4844 ( .A(n7681), .ZN(n6872) );
  NAND2_X1 U4845 ( .A1(n6859), .A2(n8228), .ZN(n7682) );
  INV_X1 U4846 ( .A(n7622), .ZN(n5409) );
  INV_X2 U4847 ( .A(n5135), .ZN(n5516) );
  NAND2_X1 U4848 ( .A1(n7863), .A2(n5514), .ZN(n5117) );
  OR2_X1 U4849 ( .A1(n7192), .A2(n7191), .ZN(n4477) );
  INV_X2 U4850 ( .A(n6210), .ZN(n8110) );
  INV_X1 U4851 ( .A(n5117), .ZN(n6293) );
  AOI21_X1 U4852 ( .B1(n6928), .B2(n4858), .A(n4856), .ZN(n7047) );
  NAND2_X1 U4853 ( .A1(n5319), .A2(n5318), .ZN(n8286) );
  INV_X1 U4855 ( .A(n5703), .ZN(n7899) );
  CLKBUF_X3 U4856 ( .A(n4986), .Z(n4325) );
  INV_X1 U4857 ( .A(n9056), .ZN(n4495) );
  INV_X2 U4858 ( .A(n6098), .ZN(n6066) );
  INV_X1 U4859 ( .A(n5080), .ZN(n5079) );
  INV_X1 U4860 ( .A(n7626), .ZN(n4322) );
  BUF_X1 U4862 ( .A(n6177), .Z(n4324) );
  OAI21_X2 U4863 ( .B1(n5705), .B2(n5704), .A(n5718), .ZN(n6358) );
  XNOR2_X2 U4864 ( .A(n5625), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6152) );
  XNOR2_X2 U4865 ( .A(n5665), .B(n4533), .ZN(n6360) );
  NAND2_X4 U4866 ( .A1(n4838), .A2(n4837), .ZN(n6784) );
  OAI21_X2 U4867 ( .B1(n6588), .B2(n4354), .A(n4697), .ZN(n9705) );
  XNOR2_X2 U4868 ( .A(n8501), .B(n9830), .ZN(n9839) );
  AOI21_X1 U4869 ( .B1(n6276), .B2(n9352), .A(n6275), .ZN(n7594) );
  MUX2_X1 U4870 ( .A(n8225), .B(n8224), .S(n9901), .Z(n8227) );
  AOI21_X1 U4871 ( .B1(n4421), .B2(n6992), .A(n4420), .ZN(n4419) );
  NAND2_X1 U4872 ( .A1(n6271), .A2(n8191), .ZN(n9177) );
  NAND2_X1 U4873 ( .A1(n9054), .A2(n5987), .ZN(n4462) );
  OR2_X1 U4874 ( .A1(n8728), .A2(n8727), .ZN(n8730) );
  AOI21_X1 U4875 ( .B1(n4521), .B2(n4520), .A(n4519), .ZN(n7542) );
  AND2_X1 U4876 ( .A1(n5917), .A2(n4391), .ZN(n4491) );
  NAND2_X1 U4877 ( .A1(n6025), .A2(n6024), .ZN(n9464) );
  OAI21_X1 U4878 ( .B1(n5389), .B2(n5388), .A(n4985), .ZN(n5404) );
  OR2_X1 U4879 ( .A1(n6795), .A2(n6794), .ZN(n6928) );
  OR2_X1 U4880 ( .A1(n4353), .A2(n4483), .ZN(n4482) );
  OR2_X1 U4881 ( .A1(n5377), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5394) );
  OAI21_X1 U4882 ( .B1(n7696), .B2(n8837), .A(n7695), .ZN(n4424) );
  XNOR2_X1 U4883 ( .A(n5234), .B(n5233), .ZN(n6336) );
  NAND2_X1 U4884 ( .A1(n8121), .A2(n7990), .ZN(n7944) );
  INV_X2 U4885 ( .A(n9365), .ZN(n9358) );
  XNOR2_X1 U4886 ( .A(n5557), .B(n5556), .ZN(n7535) );
  INV_X1 U4887 ( .A(n6555), .ZN(n9107) );
  NAND2_X1 U4888 ( .A1(n5555), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5557) );
  CLKBUF_X3 U4889 ( .A(n5109), .Z(n5364) );
  NAND2_X1 U4890 ( .A1(n5554), .A2(n5555), .ZN(n7913) );
  AND4_X1 U4891 ( .A1(n5737), .A2(n5736), .A3(n5735), .A4(n5734), .ZN(n6555)
         );
  BUF_X2 U4892 ( .A(n5687), .Z(n5930) );
  CLKBUF_X1 U4893 ( .A(n6210), .Z(n7888) );
  OR2_X1 U4894 ( .A1(n5553), .A2(n5552), .ZN(n5554) );
  NAND2_X1 U4895 ( .A1(n9660), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9694) );
  OAI21_X1 U4896 ( .B1(n6250), .B2(n6514), .A(n6249), .ZN(n5659) );
  BUF_X2 U4897 ( .A(n5713), .Z(n4333) );
  AND2_X1 U4898 ( .A1(n9203), .A2(n8163), .ZN(n6250) );
  XNOR2_X1 U4899 ( .A(n5509), .B(n4836), .ZN(n7681) );
  NAND2_X1 U4900 ( .A1(n6151), .A2(n9203), .ZN(n6249) );
  NAND2_X1 U4901 ( .A1(n7310), .A2(n4331), .ZN(n8167) );
  INV_X1 U4902 ( .A(n5645), .ZN(n9491) );
  INV_X2 U4903 ( .A(n5724), .ZN(n6322) );
  NAND2_X1 U4904 ( .A1(n8939), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5076) );
  NAND2_X1 U4905 ( .A1(n5630), .A2(n5629), .ZN(n8163) );
  OR2_X1 U4906 ( .A1(n6132), .A2(n5624), .ZN(n5679) );
  XNOR2_X1 U4907 ( .A(n5639), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5645) );
  AND2_X1 U4908 ( .A1(n5502), .A2(n5501), .ZN(n5510) );
  XNOR2_X1 U4909 ( .A(n5607), .B(n5606), .ZN(n6177) );
  NAND2_X1 U4910 ( .A1(n5605), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U4911 ( .A1(n5633), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5620) );
  OR2_X2 U4912 ( .A1(n4616), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8947) );
  INV_X2 U4913 ( .A(n4907), .ZN(n4986) );
  OR2_X1 U4914 ( .A1(n4516), .A2(n4517), .ZN(n5604) );
  NOR2_X2 U4915 ( .A1(n4517), .A2(n4514), .ZN(n4809) );
  NAND2_X1 U4916 ( .A1(n5603), .A2(n5622), .ZN(n4514) );
  AND2_X2 U4917 ( .A1(n4904), .A2(n4903), .ZN(n4907) );
  AND3_X1 U4918 ( .A1(n4716), .A2(n5617), .A3(n5618), .ZN(n5603) );
  AND4_X1 U4919 ( .A1(n5752), .A2(n5704), .A3(n5592), .A4(n5897), .ZN(n5599)
         );
  AND4_X1 U4920 ( .A1(n5665), .A2(n5674), .A3(n5597), .A4(n5596), .ZN(n5598)
         );
  AND3_X1 U4921 ( .A1(n5892), .A2(n5801), .A3(n5595), .ZN(n5898) );
  INV_X1 U4922 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5892) );
  INV_X1 U4923 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5897) );
  INV_X1 U4924 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5075) );
  INV_X4 U4925 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4926 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5674) );
  INV_X4 U4927 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U4928 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5801) );
  INV_X1 U4929 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5704) );
  NOR2_X1 U4930 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n5631) );
  AND2_X4 U4931 ( .A1(n5640), .A2(n9491), .ZN(n5699) );
  NAND2_X1 U4932 ( .A1(n6354), .A2(n4323), .ZN(n4326) );
  NAND2_X1 U4933 ( .A1(n6354), .A2(n4324), .ZN(n4327) );
  AOI21_X2 U4934 ( .B1(n8529), .B2(P2_REG2_REG_10__SCAN_IN), .A(n9756), .ZN(
        n8494) );
  AND2_X4 U4935 ( .A1(n5641), .A2(n9491), .ZN(n5696) );
  BUF_X2 U4936 ( .A(n5807), .Z(n4328) );
  AND2_X1 U4937 ( .A1(n5641), .A2(n5645), .ZN(n5807) );
  NAND2_X1 U4938 ( .A1(n5724), .A2(n4907), .ZN(n4330) );
  XNOR2_X1 U4939 ( .A(n5654), .B(P1_IR_REG_19__SCAN_IN), .ZN(n5988) );
  OAI222_X1 U4940 ( .A1(n9493), .A2(n7583), .B1(P1_U3086), .B2(n6354), .C1(
        n7582), .C2(n9490), .ZN(P1_U3328) );
  AOI21_X2 U4941 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8525), .A(n9788), .ZN(
        n8497) );
  XNOR2_X2 U4942 ( .A(n9109), .B(n8110), .ZN(n6254) );
  AND2_X1 U4943 ( .A1(n5640), .A2(n5645), .ZN(n5713) );
  OAI211_X1 U4944 ( .C1(n8069), .C2(n8068), .A(n6270), .B(n8067), .ZN(n8073)
         );
  AOI21_X1 U4945 ( .B1(n4952), .B2(n4453), .A(n4390), .ZN(n4452) );
  NAND2_X1 U4946 ( .A1(n5243), .A2(n4453), .ZN(n4451) );
  OR2_X1 U4947 ( .A1(n8619), .A2(n8460), .ZN(n7846) );
  INV_X1 U4948 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5032) );
  NOR2_X1 U4949 ( .A1(n4892), .A2(n4364), .ZN(n4883) );
  INV_X1 U4950 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U4951 ( .A1(n4653), .A2(n4650), .ZN(n5370) );
  INV_X1 U4952 ( .A(n4651), .ZN(n4650) );
  OAI21_X1 U4953 ( .B1(n4971), .B2(n4652), .A(n4970), .ZN(n4651) );
  AOI21_X1 U4954 ( .B1(n4362), .B2(P2_D_REG_0__SCAN_IN), .A(n4344), .ZN(n4837)
         );
  AOI21_X1 U4955 ( .B1(n7865), .B2(n8592), .A(n5513), .ZN(n8679) );
  NAND2_X1 U4956 ( .A1(n5042), .A2(n5562), .ZN(n5565) );
  NAND2_X1 U4957 ( .A1(n4479), .A2(n5667), .ZN(n4478) );
  NAND2_X1 U4958 ( .A1(n5727), .A2(n7888), .ZN(n4479) );
  NAND2_X1 U4959 ( .A1(n8117), .A2(n8115), .ZN(n6257) );
  AND3_X1 U4960 ( .A1(n5679), .A2(P1_STATE_REG_SCAN_IN), .A3(n6323), .ZN(n6320) );
  NAND2_X1 U4961 ( .A1(n5638), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5639) );
  INV_X1 U4962 ( .A(n5633), .ZN(n5637) );
  NAND2_X1 U4963 ( .A1(n7821), .A2(n4378), .ZN(n4427) );
  NAND2_X1 U4964 ( .A1(n4562), .A2(n8167), .ZN(n4560) );
  OR2_X1 U4965 ( .A1(n9215), .A2(n9225), .ZN(n8083) );
  OR2_X1 U4966 ( .A1(n4987), .A2(n5401), .ZN(n4669) );
  INV_X1 U4967 ( .A(SI_9_), .ZN(n4943) );
  NAND2_X1 U4968 ( .A1(n5079), .A2(n5081), .ZN(n5109) );
  NAND2_X1 U4969 ( .A1(n4361), .A2(n5441), .ZN(n4597) );
  INV_X1 U4970 ( .A(n4737), .ZN(n4736) );
  OR2_X1 U4971 ( .A1(n8899), .A2(n8700), .ZN(n7805) );
  OR2_X1 U4972 ( .A1(n8909), .A2(n8699), .ZN(n7794) );
  NAND2_X1 U4973 ( .A1(n4358), .A2(n5327), .ZN(n4439) );
  INV_X1 U4974 ( .A(n7258), .ZN(n4614) );
  AOI21_X1 U4975 ( .B1(n4874), .B2(n4877), .A(n4387), .ZN(n4870) );
  INV_X1 U4976 ( .A(n4874), .ZN(n4871) );
  INV_X1 U4977 ( .A(n9039), .ZN(n4872) );
  NAND2_X1 U4978 ( .A1(n4449), .A2(n8962), .ZN(n4470) );
  OR2_X1 U4979 ( .A1(n6314), .A2(n6147), .ZN(n6247) );
  OR2_X1 U4980 ( .A1(n8098), .A2(n7896), .ZN(n4672) );
  NOR2_X1 U4981 ( .A1(n8098), .A2(n5703), .ZN(n4673) );
  OR2_X1 U4982 ( .A1(n8097), .A2(n7934), .ZN(n8099) );
  AND2_X1 U4983 ( .A1(n9282), .A2(n7971), .ZN(n4722) );
  NAND2_X1 U4984 ( .A1(n9047), .A2(n7391), .ZN(n4800) );
  OR2_X1 U4985 ( .A1(n8216), .A2(n7929), .ZN(n8093) );
  NOR2_X1 U4986 ( .A1(n6243), .A2(n4805), .ZN(n4804) );
  INV_X1 U4987 ( .A(n4806), .ZN(n4805) );
  AND2_X1 U4988 ( .A1(n4812), .A2(n4503), .ZN(n4502) );
  AND2_X1 U4989 ( .A1(n4368), .A2(n7975), .ZN(n4812) );
  NAND2_X1 U4990 ( .A1(n4811), .A2(n4504), .ZN(n4503) );
  XNOR2_X1 U4991 ( .A(n7607), .B(n7606), .ZN(n7610) );
  AOI21_X1 U4992 ( .B1(n4647), .B2(n4649), .A(n4645), .ZN(n4644) );
  INV_X1 U4993 ( .A(n5017), .ZN(n4645) );
  AND2_X1 U4994 ( .A1(n5012), .A2(n5011), .ZN(n5463) );
  AND2_X1 U4995 ( .A1(n5001), .A2(n5000), .ZN(n5442) );
  OAI21_X1 U4996 ( .B1(n5404), .B2(n4661), .A(n4404), .ZN(n5433) );
  INV_X1 U4997 ( .A(n4665), .ZN(n4661) );
  NOR2_X1 U4998 ( .A1(n5430), .A2(n4663), .ZN(n4662) );
  NAND2_X1 U4999 ( .A1(n5404), .A2(n4669), .ZN(n4668) );
  OAI21_X1 U5000 ( .B1(n5358), .B2(n4980), .A(n4979), .ZN(n5389) );
  AND2_X1 U5001 ( .A1(SI_14_), .A2(n5292), .ZN(n4960) );
  NAND2_X1 U5002 ( .A1(n4451), .A2(n4369), .ZN(n5291) );
  INV_X1 U5003 ( .A(n5254), .ZN(n4450) );
  NOR2_X1 U5004 ( .A1(n4941), .A2(n4639), .ZN(n4638) );
  INV_X1 U5005 ( .A(n4933), .ZN(n4639) );
  NAND2_X1 U5006 ( .A1(n7340), .A2(n4902), .ZN(n4903) );
  INV_X1 U5007 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4901) );
  NAND2_X1 U5008 ( .A1(n4847), .A2(n4846), .ZN(n4845) );
  NAND2_X1 U5009 ( .A1(n4848), .A2(n4849), .ZN(n4847) );
  OAI21_X1 U5010 ( .B1(n8327), .B2(n8325), .A(n4851), .ZN(n4846) );
  INV_X1 U5011 ( .A(n8327), .ZN(n4848) );
  NAND2_X1 U5012 ( .A1(n6928), .A2(n4860), .ZN(n7005) );
  AND2_X1 U5013 ( .A1(n5036), .A2(n5559), .ZN(n5037) );
  OAI21_X1 U5014 ( .B1(n7852), .B2(n8867), .A(n7842), .ZN(n4425) );
  AND4_X1 U5015 ( .A1(n5399), .A2(n5398), .A3(n5397), .A4(n5396), .ZN(n8426)
         );
  OR2_X1 U5016 ( .A1(n5477), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U5017 ( .A1(n5117), .A2(n4907), .ZN(n5221) );
  AND2_X1 U5018 ( .A1(n8646), .A2(n8791), .ZN(n4443) );
  AOI21_X1 U5019 ( .B1(n8667), .B2(n5461), .A(n5460), .ZN(n8654) );
  INV_X1 U5020 ( .A(n8462), .ZN(n8680) );
  OAI21_X1 U5021 ( .B1(n8730), .B2(n4600), .A(n4598), .ZN(n5429) );
  INV_X1 U5022 ( .A(n4599), .ZN(n4598) );
  OR2_X1 U5023 ( .A1(n8810), .A2(n8417), .ZN(n7800) );
  NAND2_X1 U5024 ( .A1(n5117), .A2(n4325), .ZN(n7636) );
  INV_X1 U5025 ( .A(n5221), .ZN(n7635) );
  INV_X1 U5026 ( .A(n7636), .ZN(n5491) );
  NAND2_X1 U5027 ( .A1(n5568), .A2(n5567), .ZN(n6431) );
  INV_X1 U5028 ( .A(n7541), .ZN(n5567) );
  NAND2_X1 U5029 ( .A1(n5558), .A2(n7535), .ZN(n5568) );
  INV_X1 U5030 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5503) );
  INV_X1 U5031 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5501) );
  XNOR2_X1 U5032 ( .A(n5390), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U5033 ( .A1(n5040), .A2(n5173), .ZN(n5041) );
  NAND2_X1 U5034 ( .A1(n4882), .A2(n4376), .ZN(n4488) );
  INV_X1 U5035 ( .A(n4864), .ZN(n4468) );
  AOI22_X1 U5036 ( .A1(n9108), .A2(n5695), .B1(n6215), .B2(n5727), .ZN(n5728)
         );
  NAND2_X1 U5037 ( .A1(n9458), .A2(n9238), .ZN(n8066) );
  NAND2_X1 U5038 ( .A1(n6056), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6075) );
  AND3_X1 U5039 ( .A1(n5928), .A2(n5927), .A3(n5926), .ZN(n9348) );
  NAND2_X1 U5040 ( .A1(n6225), .A2(n4893), .ZN(n7568) );
  OR2_X1 U5041 ( .A1(n7558), .A2(n9096), .ZN(n6224) );
  NAND2_X1 U5042 ( .A1(n4702), .A2(n4340), .ZN(n4701) );
  NOR2_X1 U5043 ( .A1(n6263), .A2(n7988), .ZN(n4705) );
  AND2_X1 U5044 ( .A1(n9354), .A2(n4331), .ZN(n6244) );
  NAND2_X1 U5045 ( .A1(n7943), .A2(n6977), .ZN(n4540) );
  XNOR2_X1 U5046 ( .A(n7610), .B(SI_29_), .ZN(n8944) );
  INV_X1 U5047 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5606) );
  INV_X1 U5048 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5597) );
  INV_X1 U5049 ( .A(n7309), .ZN(n7865) );
  OR2_X1 U5050 ( .A1(n7538), .A2(n7532), .ZN(n5624) );
  AOI21_X1 U5051 ( .B1(n7684), .B2(n4370), .A(n4428), .ZN(n7689) );
  INV_X1 U5052 ( .A(n7686), .ZN(n4428) );
  NAND2_X1 U5053 ( .A1(n4543), .A2(n7992), .ZN(n4542) );
  OR2_X1 U5054 ( .A1(n7993), .A2(n8120), .ZN(n4543) );
  OAI21_X1 U5055 ( .B1(n8015), .B2(n4568), .A(n8020), .ZN(n4567) );
  NAND2_X1 U5056 ( .A1(n8014), .A2(n8005), .ZN(n4568) );
  NAND2_X1 U5057 ( .A1(n4546), .A2(n9346), .ZN(n8051) );
  NAND2_X1 U5058 ( .A1(n4548), .A2(n4547), .ZN(n4546) );
  NAND2_X1 U5059 ( .A1(n8033), .A2(n8085), .ZN(n4547) );
  AOI21_X1 U5060 ( .B1(n8034), .B2(n8167), .A(n8041), .ZN(n4548) );
  AND2_X1 U5061 ( .A1(n8630), .A2(n7825), .ZN(n4426) );
  NAND2_X1 U5062 ( .A1(n4380), .A2(n9182), .ZN(n4562) );
  INV_X1 U5063 ( .A(n4855), .ZN(n4853) );
  INV_X1 U5064 ( .A(n5179), .ZN(n4627) );
  NOR2_X1 U5065 ( .A1(n4876), .A2(n4875), .ZN(n4874) );
  INV_X1 U5066 ( .A(n7498), .ZN(n4875) );
  NOR2_X1 U5067 ( .A1(n4877), .A2(n4879), .ZN(n4876) );
  OR2_X1 U5068 ( .A1(n4555), .A2(n7902), .ZN(n4554) );
  OAI21_X1 U5069 ( .B1(n5023), .B2(n4642), .A(n4640), .ZN(n7607) );
  AOI21_X1 U5070 ( .B1(n5487), .B2(n4641), .A(n4406), .ZN(n4640) );
  INV_X1 U5071 ( .A(n5487), .ZN(n4642) );
  INV_X1 U5072 ( .A(n4648), .ZN(n4647) );
  OAI21_X1 U5073 ( .B1(n5463), .B2(n4649), .A(n5474), .ZN(n4648) );
  NAND2_X1 U5074 ( .A1(n4665), .A2(n4660), .ZN(n4659) );
  INV_X1 U5075 ( .A(n4669), .ZN(n4660) );
  AND2_X1 U5076 ( .A1(n5290), .A2(n5293), .ZN(n4962) );
  NAND2_X1 U5077 ( .A1(n4959), .A2(n4958), .ZN(n5292) );
  AOI21_X1 U5078 ( .B1(n8264), .B2(n4820), .A(n4819), .ZN(n4818) );
  INV_X1 U5079 ( .A(n8258), .ZN(n4820) );
  INV_X1 U5080 ( .A(n8264), .ZN(n4821) );
  INV_X1 U5081 ( .A(n7234), .ZN(n4833) );
  AOI21_X1 U5082 ( .B1(n7739), .B2(n7653), .A(n4754), .ZN(n4753) );
  INV_X1 U5083 ( .A(n7743), .ZN(n4754) );
  INV_X1 U5084 ( .A(n7739), .ZN(n4755) );
  NAND2_X1 U5085 ( .A1(n4442), .A2(n4440), .ZN(n7742) );
  AND2_X1 U5086 ( .A1(n4441), .A2(n5272), .ZN(n4440) );
  NAND2_X1 U5087 ( .A1(n5149), .A2(n5148), .ZN(n5161) );
  NAND2_X1 U5088 ( .A1(n4840), .A2(n5571), .ZN(n6778) );
  OR2_X1 U5089 ( .A1(n6431), .A2(P2_D_REG_0__SCAN_IN), .ZN(n4840) );
  OR2_X1 U5090 ( .A1(n8883), .A2(n8441), .ZN(n7815) );
  OR2_X1 U5091 ( .A1(n8889), .A2(n8680), .ZN(n7813) );
  NOR2_X1 U5092 ( .A1(n5541), .A2(n4738), .ZN(n4737) );
  INV_X1 U5093 ( .A(n7800), .ZN(n4738) );
  INV_X1 U5094 ( .A(n7795), .ZN(n4735) );
  OR2_X1 U5095 ( .A1(n8804), .A2(n8382), .ZN(n7811) );
  AND2_X1 U5096 ( .A1(n8716), .A2(n5400), .ZN(n4603) );
  OR2_X1 U5097 ( .A1(n8927), .A2(n8250), .ZN(n7778) );
  INV_X1 U5098 ( .A(n4439), .ZN(n4437) );
  NOR2_X1 U5099 ( .A1(n4612), .A2(n5311), .ZN(n4606) );
  INV_X1 U5100 ( .A(n4613), .ZN(n4612) );
  AND4_X1 U5101 ( .A1(n5035), .A2(n5034), .A3(n5033), .A4(n5585), .ZN(n5559)
         );
  OAI21_X1 U5102 ( .B1(n8981), .B2(n4458), .A(n4457), .ZN(n6051) );
  INV_X1 U5103 ( .A(n8978), .ZN(n4458) );
  INV_X1 U5104 ( .A(n6047), .ZN(n4457) );
  NOR2_X1 U5105 ( .A1(n4885), .A2(n6889), .ZN(n4490) );
  AND2_X1 U5106 ( .A1(n9553), .A2(n9146), .ZN(n9147) );
  OR2_X1 U5107 ( .A1(n4584), .A2(n7596), .ZN(n4582) );
  NAND2_X1 U5108 ( .A1(n4586), .A2(n4585), .ZN(n4584) );
  INV_X1 U5109 ( .A(n8216), .ZN(n4586) );
  AND2_X1 U5110 ( .A1(n6270), .A2(n8066), .ZN(n4710) );
  INV_X1 U5111 ( .A(n9247), .ZN(n4709) );
  NOR2_X1 U5112 ( .A1(n6269), .A2(n4573), .ZN(n4572) );
  INV_X1 U5113 ( .A(n4574), .ZN(n4573) );
  INV_X1 U5114 ( .A(n7941), .ZN(n4726) );
  NOR2_X1 U5115 ( .A1(n4727), .A2(n4726), .ZN(n4725) );
  NOR2_X1 U5116 ( .A1(n7543), .A2(n7558), .ZN(n4588) );
  NAND2_X1 U5117 ( .A1(n4579), .A2(n7392), .ZN(n4578) );
  OR2_X1 U5118 ( .A1(n7024), .A2(n7454), .ZN(n8012) );
  OR2_X1 U5119 ( .A1(n7061), .A2(n7105), .ZN(n7996) );
  AND2_X1 U5120 ( .A1(n9182), .A2(n7939), .ZN(n8195) );
  NOR2_X1 U5121 ( .A1(n6240), .A2(n4807), .ZN(n4806) );
  INV_X1 U5122 ( .A(n6238), .ZN(n4807) );
  NAND2_X1 U5123 ( .A1(n9417), .A2(n9094), .ZN(n4513) );
  INV_X1 U5124 ( .A(n7954), .ZN(n4797) );
  INV_X1 U5125 ( .A(n9099), .ZN(n7466) );
  AND2_X1 U5126 ( .A1(n6459), .A2(n6247), .ZN(n6511) );
  NAND2_X1 U5127 ( .A1(n4810), .A2(n4809), .ZN(n5633) );
  NAND2_X1 U5128 ( .A1(n4987), .A2(n5401), .ZN(n4667) );
  OAI21_X1 U5129 ( .B1(n5370), .B2(n5369), .A(n4976), .ZN(n5358) );
  NAND2_X1 U5130 ( .A1(n4433), .A2(n4432), .ZN(n5243) );
  AOI21_X1 U5131 ( .B1(n4434), .B2(n4637), .A(n4634), .ZN(n4433) );
  NAND2_X1 U5132 ( .A1(n4434), .A2(n4934), .ZN(n4432) );
  INV_X1 U5133 ( .A(n4947), .ZN(n4634) );
  AND2_X1 U5134 ( .A1(n4947), .A2(n4946), .ZN(n5233) );
  NAND2_X1 U5135 ( .A1(n4919), .A2(n4418), .ZN(n4417) );
  INV_X1 U5136 ( .A(n5144), .ZN(n4418) );
  NAND2_X1 U5137 ( .A1(n4431), .A2(n4430), .ZN(n4910) );
  NAND2_X1 U5138 ( .A1(n4907), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4430) );
  XNOR2_X1 U5139 ( .A(n4910), .B(n4429), .ZN(n4909) );
  INV_X1 U5140 ( .A(SI_1_), .ZN(n4429) );
  NAND2_X1 U5141 ( .A1(n7228), .A2(n7227), .ZN(n4834) );
  OR2_X1 U5142 ( .A1(n5109), .A2(n6879), .ZN(n5099) );
  INV_X1 U5143 ( .A(n6927), .ZN(n4861) );
  INV_X1 U5144 ( .A(n7004), .ZN(n4859) );
  NAND2_X1 U5145 ( .A1(n4827), .A2(n4825), .ZN(n4824) );
  INV_X1 U5146 ( .A(n8242), .ZN(n4825) );
  AOI21_X1 U5147 ( .B1(n8401), .B2(n8242), .A(n4828), .ZN(n4827) );
  INV_X1 U5148 ( .A(n8283), .ZN(n4828) );
  NAND2_X1 U5149 ( .A1(n5565), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5045) );
  AND2_X1 U5150 ( .A1(n8610), .A2(n8607), .ZN(n7858) );
  AND3_X1 U5151 ( .A1(n5427), .A2(n5426), .A3(n5425), .ZN(n8417) );
  AND4_X1 U5152 ( .A1(n5356), .A2(n5355), .A3(n5354), .A4(n5353), .ZN(n8353)
         );
  NAND2_X1 U5153 ( .A1(n9696), .A2(n4699), .ZN(n4700) );
  NOR2_X1 U5154 ( .A1(n4354), .A2(n6660), .ZN(n4699) );
  OR2_X1 U5155 ( .A1(n9773), .A2(n5277), .ZN(n4690) );
  OR2_X1 U5156 ( .A1(n9839), .A2(n7525), .ZN(n4695) );
  NAND2_X1 U5157 ( .A1(n4696), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4693) );
  NAND2_X1 U5158 ( .A1(n8502), .A2(n4696), .ZN(n4692) );
  INV_X1 U5159 ( .A(n9859), .ZN(n4696) );
  NAND2_X1 U5160 ( .A1(n6291), .A2(n6767), .ZN(n6610) );
  OAI21_X1 U5161 ( .B1(n8643), .B2(n4388), .A(n4769), .ZN(n7605) );
  AND2_X1 U5162 ( .A1(n4398), .A2(n4770), .ZN(n4769) );
  OR2_X1 U5163 ( .A1(n5546), .A2(n7828), .ZN(n4772) );
  INV_X1 U5164 ( .A(n5466), .ZN(n5068) );
  NAND2_X1 U5165 ( .A1(n6438), .A2(n7635), .ZN(n4442) );
  OAI22_X1 U5166 ( .A1(n7174), .A2(n5242), .B1(n8466), .B2(n7239), .ZN(n7258)
         );
  NAND2_X1 U5167 ( .A1(n5534), .A2(n5533), .ZN(n7201) );
  NAND2_X1 U5168 ( .A1(n5051), .A2(n5050), .ZN(n5208) );
  INV_X1 U5169 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5050) );
  INV_X1 U5170 ( .A(n5195), .ZN(n5051) );
  NAND2_X1 U5171 ( .A1(n4760), .A2(n4759), .ZN(n6962) );
  AOI22_X1 U5172 ( .A1(n4761), .A2(n4763), .B1(n4764), .B2(n4758), .ZN(n4759)
         );
  INV_X1 U5173 ( .A(n4766), .ZN(n4763) );
  NAND2_X1 U5174 ( .A1(n4622), .A2(n4621), .ZN(n5119) );
  NAND2_X1 U5175 ( .A1(n5117), .A2(n4615), .ZN(n4621) );
  OAI21_X1 U5176 ( .B1(n5117), .B2(n4620), .A(n4617), .ZN(n4622) );
  NOR2_X1 U5177 ( .A1(n6297), .A2(n4616), .ZN(n4615) );
  INV_X1 U5178 ( .A(n8771), .ZN(n8838) );
  INV_X1 U5179 ( .A(n7827), .ZN(n4774) );
  NAND2_X1 U5180 ( .A1(n4776), .A2(n7824), .ZN(n8631) );
  NAND2_X1 U5181 ( .A1(n4768), .A2(n7823), .ZN(n4776) );
  INV_X1 U5182 ( .A(n8643), .ZN(n4768) );
  NAND2_X1 U5183 ( .A1(n6775), .A2(n7826), .ZN(n8840) );
  INV_X1 U5184 ( .A(n4597), .ZN(n4594) );
  AND2_X1 U5185 ( .A1(n7811), .A2(n8663), .ZN(n8676) );
  INV_X1 U5186 ( .A(n8730), .ZN(n4602) );
  NAND2_X1 U5187 ( .A1(n8730), .A2(n4603), .ZN(n8715) );
  NAND2_X1 U5188 ( .A1(n4742), .A2(n4740), .ZN(n8713) );
  AOI21_X1 U5189 ( .B1(n4743), .B2(n4746), .A(n4741), .ZN(n4740) );
  INV_X1 U5190 ( .A(n7790), .ZN(n4741) );
  NAND2_X1 U5191 ( .A1(n4589), .A2(n4381), .ZN(n8728) );
  NAND2_X1 U5192 ( .A1(n8742), .A2(n5383), .ZN(n4589) );
  NOR2_X1 U5193 ( .A1(n5539), .A2(n4748), .ZN(n4747) );
  INV_X1 U5194 ( .A(n7786), .ZN(n4748) );
  NAND2_X1 U5195 ( .A1(n5540), .A2(n7778), .ZN(n4749) );
  NOR2_X1 U5196 ( .A1(n7770), .A2(n4785), .ZN(n4784) );
  INV_X1 U5197 ( .A(n7768), .ZN(n4785) );
  AND2_X1 U5198 ( .A1(n4605), .A2(n4604), .ZN(n4607) );
  AND2_X1 U5199 ( .A1(n4611), .A2(n4394), .ZN(n4604) );
  OR2_X1 U5200 ( .A1(n8286), .A2(n8402), .ZN(n7768) );
  OR2_X1 U5201 ( .A1(n5289), .A2(n5311), .ZN(n4605) );
  NAND2_X1 U5202 ( .A1(n8408), .A2(n8465), .ZN(n4611) );
  NAND2_X1 U5203 ( .A1(n4606), .A2(n4614), .ZN(n4608) );
  INV_X1 U5204 ( .A(n7660), .ZN(n7762) );
  INV_X1 U5205 ( .A(n8840), .ZN(n8769) );
  AND2_X1 U5206 ( .A1(n5562), .A2(n4787), .ZN(n4786) );
  NOR2_X1 U5207 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4787) );
  NAND2_X1 U5208 ( .A1(n5551), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5553) );
  INV_X1 U5209 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U5210 ( .A1(n5553), .A2(n5552), .ZN(n5555) );
  INV_X1 U5211 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5201) );
  AND2_X1 U5212 ( .A1(n5038), .A2(n5039), .ZN(n4814) );
  INV_X1 U5213 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5039) );
  INV_X1 U5214 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U5215 ( .A1(n4864), .A2(n4863), .ZN(n8961) );
  INV_X1 U5216 ( .A(n4449), .ZN(n4863) );
  OAI21_X1 U5217 ( .B1(n4488), .B2(n4482), .A(n4480), .ZN(n5798) );
  AOI21_X1 U5218 ( .B1(n4410), .B2(n4487), .A(n4481), .ZN(n4480) );
  INV_X1 U5219 ( .A(n7099), .ZN(n4481) );
  OR2_X1 U5220 ( .A1(n6744), .A2(n4892), .ZN(n4886) );
  OR2_X1 U5221 ( .A1(n5952), .A2(n5951), .ZN(n5976) );
  OAI21_X1 U5222 ( .B1(n4469), .B2(n4468), .A(n4466), .ZN(n8181) );
  AOI21_X1 U5223 ( .B1(n4470), .B2(n4373), .A(n4467), .ZN(n4466) );
  INV_X1 U5224 ( .A(n8183), .ZN(n4467) );
  NOR2_X1 U5225 ( .A1(n4869), .A2(n4868), .ZN(n4867) );
  INV_X1 U5226 ( .A(n6052), .ZN(n4868) );
  INV_X1 U5227 ( .A(n6051), .ZN(n4869) );
  INV_X1 U5228 ( .A(n8976), .ZN(n4862) );
  INV_X1 U5229 ( .A(n5673), .ZN(n6049) );
  OR2_X1 U5230 ( .A1(n5819), .A2(n5818), .ZN(n4472) );
  NAND2_X1 U5231 ( .A1(n4475), .A2(n4474), .ZN(n4473) );
  INV_X1 U5232 ( .A(n7293), .ZN(n4474) );
  OR2_X1 U5233 ( .A1(n4353), .A2(n4490), .ZN(n4486) );
  NAND2_X1 U5234 ( .A1(n8987), .A2(n8988), .ZN(n4881) );
  OAI21_X1 U5235 ( .B1(n8096), .B2(n4551), .A(n4549), .ZN(n8165) );
  AND2_X1 U5236 ( .A1(n4556), .A2(n8101), .ZN(n4551) );
  INV_X1 U5237 ( .A(n4550), .ZN(n4549) );
  INV_X1 U5238 ( .A(n8099), .ZN(n8169) );
  INV_X1 U5239 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U5240 ( .A1(n5655), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5657) );
  OR2_X1 U5241 ( .A1(n6392), .A2(n6391), .ZN(n4532) );
  NOR2_X1 U5242 ( .A1(n9557), .A2(n4538), .ZN(n9127) );
  AND2_X1 U5243 ( .A1(n9562), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4538) );
  AND4_X1 U5244 ( .A1(n6115), .A2(n6114), .A3(n6113), .A4(n6112), .ZN(n9225)
         );
  INV_X1 U5245 ( .A(n4717), .ZN(n4718) );
  INV_X1 U5246 ( .A(n7923), .ZN(n4719) );
  INV_X1 U5247 ( .A(n6267), .ZN(n4721) );
  INV_X1 U5248 ( .A(n7971), .ZN(n4720) );
  NAND2_X1 U5249 ( .A1(n6267), .A2(n4722), .ZN(n9280) );
  AND2_X1 U5250 ( .A1(n5992), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U5251 ( .A1(n4508), .A2(n4507), .ZN(n4501) );
  INV_X1 U5252 ( .A(n9470), .ZN(n9317) );
  AND2_X1 U5253 ( .A1(n8043), .A2(n8052), .ZN(n9333) );
  NAND2_X1 U5254 ( .A1(n7574), .A2(n7575), .ZN(n7573) );
  INV_X1 U5255 ( .A(n8018), .ZN(n4423) );
  NAND2_X1 U5256 ( .A1(n7954), .A2(n4800), .ZN(n4796) );
  NAND2_X1 U5257 ( .A1(n4518), .A2(n4341), .ZN(n4795) );
  AND2_X1 U5258 ( .A1(n4795), .A2(n4793), .ZN(n7243) );
  NOR2_X1 U5259 ( .A1(n7245), .A2(n4794), .ZN(n4793) );
  INV_X1 U5260 ( .A(n4796), .ZN(n4794) );
  AND2_X1 U5261 ( .A1(n8018), .A2(n8133), .ZN(n7245) );
  NAND2_X1 U5262 ( .A1(n7019), .A2(n6223), .ZN(n7145) );
  OR2_X1 U5263 ( .A1(n7024), .A2(n9102), .ZN(n6223) );
  NAND2_X1 U5264 ( .A1(n6839), .A2(n6838), .ZN(n6837) );
  OR2_X1 U5265 ( .A1(n6306), .A2(n5703), .ZN(n5755) );
  INV_X1 U5266 ( .A(n9349), .ZN(n9337) );
  AND2_X1 U5267 ( .A1(n6562), .A2(n6501), .ZN(n6558) );
  NAND2_X1 U5268 ( .A1(n6324), .A2(n6403), .ZN(n9347) );
  NAND2_X1 U5269 ( .A1(n6324), .A2(n4324), .ZN(n9349) );
  INV_X1 U5270 ( .A(n9352), .ZN(n9299) );
  NOR2_X1 U5271 ( .A1(n6976), .A2(n6505), .ZN(n6501) );
  NAND2_X1 U5272 ( .A1(n6256), .A2(n8115), .ZN(n6502) );
  AOI22_X1 U5273 ( .A1(n8194), .A2(n8193), .B1(n8192), .B2(n9202), .ZN(n9176)
         );
  INV_X1 U5274 ( .A(n8195), .ZN(n9179) );
  NAND2_X1 U5275 ( .A1(n6310), .A2(n4791), .ZN(n4789) );
  AND4_X1 U5276 ( .A1(n6164), .A2(n6163), .A3(n6162), .A4(n6161), .ZN(n8196)
         );
  AND2_X1 U5277 ( .A1(n8093), .A2(n8094), .ZN(n8201) );
  AND2_X1 U5278 ( .A1(n8087), .A2(n9178), .ZN(n8191) );
  NAND2_X1 U5279 ( .A1(n7594), .A2(n7599), .ZN(n6286) );
  OR2_X1 U5280 ( .A1(n9246), .A2(n4348), .ZN(n6239) );
  NAND2_X1 U5281 ( .A1(n8070), .A2(n8071), .ZN(n9236) );
  AND2_X1 U5282 ( .A1(n8065), .A2(n8066), .ZN(n9247) );
  NAND2_X1 U5283 ( .A1(n4811), .A2(n4506), .ZN(n4505) );
  AND2_X1 U5284 ( .A1(n8044), .A2(n8150), .ZN(n9312) );
  OR2_X1 U5285 ( .A1(n4511), .A2(n4509), .ZN(n4507) );
  INV_X1 U5286 ( .A(n4513), .ZN(n4509) );
  AND2_X1 U5287 ( .A1(n6229), .A2(n4512), .ZN(n4511) );
  INV_X1 U5288 ( .A(n6227), .ZN(n4512) );
  NAND2_X1 U5289 ( .A1(n4513), .A2(n6228), .ZN(n4510) );
  AOI21_X1 U5290 ( .B1(n7568), .B2(n4727), .A(n6226), .ZN(n9344) );
  OR2_X1 U5291 ( .A1(n7428), .A2(n4522), .ZN(n4521) );
  AND2_X1 U5292 ( .A1(n7501), .A2(n8955), .ZN(n4522) );
  AOI21_X1 U5293 ( .B1(n7466), .B2(n7392), .A(n7243), .ZN(n7429) );
  NOR2_X1 U5294 ( .A1(n7429), .A2(n7955), .ZN(n7428) );
  OR2_X1 U5295 ( .A1(n6312), .A2(n5703), .ZN(n5723) );
  NOR2_X1 U5296 ( .A1(n4330), .A2(n6309), .ZN(n4730) );
  OAI22_X1 U5297 ( .A1(n5703), .A2(n5666), .B1(n6360), .B2(n5724), .ZN(n4731)
         );
  OR2_X1 U5298 ( .A1(n8103), .A2(n6273), .ZN(n9352) );
  NAND2_X1 U5299 ( .A1(n6135), .A2(n6134), .ZN(n6314) );
  XNOR2_X1 U5300 ( .A(n7620), .B(n7619), .ZN(n7894) );
  NAND2_X1 U5301 ( .A1(n7631), .A2(n7634), .ZN(n8220) );
  XNOR2_X1 U5302 ( .A(n5473), .B(n5474), .ZN(n7536) );
  NAND2_X1 U5303 ( .A1(n4646), .A2(n5012), .ZN(n5473) );
  NOR2_X1 U5304 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4889) );
  NAND2_X1 U5305 ( .A1(n4664), .A2(n4989), .ZN(n5431) );
  NAND2_X1 U5306 ( .A1(n4668), .A2(n4665), .ZN(n4664) );
  OAI21_X1 U5307 ( .B1(n5330), .B2(n4657), .A(n4656), .ZN(n5344) );
  AND2_X1 U5308 ( .A1(n5291), .A2(n5256), .ZN(n6475) );
  AND2_X1 U5309 ( .A1(n4940), .A2(n4939), .ZN(n5219) );
  NAND2_X1 U5310 ( .A1(n5204), .A2(n5203), .ZN(n4934) );
  NAND2_X1 U5311 ( .A1(n4445), .A2(n4926), .ZN(n5191) );
  OR2_X1 U5312 ( .A1(n5751), .A2(n9484), .ZN(n5705) );
  INV_X1 U5313 ( .A(n8655), .ZN(n8636) );
  AND3_X1 U5314 ( .A1(n5440), .A2(n5439), .A3(n5438), .ZN(n8700) );
  AND4_X1 U5315 ( .A1(n5414), .A2(n5413), .A3(n5412), .A4(n5411), .ZN(n8699)
         );
  NOR2_X1 U5316 ( .A1(n4342), .A2(n8410), .ZN(n4842) );
  NAND2_X1 U5317 ( .A1(n4845), .A2(n4850), .ZN(n4844) );
  NAND2_X1 U5318 ( .A1(n8327), .A2(n8325), .ZN(n4850) );
  AND4_X1 U5319 ( .A1(n5154), .A2(n5153), .A3(n5152), .A4(n5151), .ZN(n7007)
         );
  INV_X1 U5320 ( .A(n8469), .ZN(n7163) );
  AND4_X1 U5321 ( .A1(n5214), .A2(n5213), .A3(n5212), .A4(n5211), .ZN(n7237)
         );
  INV_X1 U5322 ( .A(n8470), .ZN(n7700) );
  NAND2_X1 U5323 ( .A1(n6771), .A2(n9869), .ZN(n9950) );
  OR2_X1 U5324 ( .A1(n6855), .A2(n7401), .ZN(n9948) );
  XNOR2_X1 U5325 ( .A(n5043), .B(n5072), .ZN(n7863) );
  NAND2_X1 U5326 ( .A1(n4335), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U5327 ( .A1(n5086), .A2(n5085), .ZN(n8461) );
  NAND2_X1 U5328 ( .A1(n5459), .A2(n5458), .ZN(n8462) );
  INV_X1 U5329 ( .A(n8426), .ZN(n8748) );
  INV_X1 U5330 ( .A(n8353), .ZN(n8757) );
  INV_X1 U5331 ( .A(n7007), .ZN(n8471) );
  INV_X1 U5332 ( .A(n8839), .ZN(n8472) );
  NAND2_X1 U5333 ( .A1(n8940), .A2(n5038), .ZN(n4674) );
  NAND2_X1 U5334 ( .A1(n5128), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n4675) );
  INV_X1 U5335 ( .A(n4686), .ZN(n4682) );
  OAI21_X1 U5336 ( .B1(n5527), .B2(n8679), .A(n5526), .ZN(n8615) );
  NOR2_X1 U5337 ( .A1(n5525), .A2(n5524), .ZN(n5526) );
  NOR2_X1 U5338 ( .A1(n7838), .A2(n8605), .ZN(n5524) );
  NAND2_X1 U5339 ( .A1(n5090), .A2(n5089), .ZN(n8791) );
  NAND2_X1 U5340 ( .A1(n5420), .A2(n5419), .ZN(n8810) );
  NAND2_X1 U5341 ( .A1(n5392), .A2(n5391), .ZN(n8738) );
  NAND2_X1 U5342 ( .A1(n5493), .A2(n5492), .ZN(n8619) );
  NAND2_X1 U5343 ( .A1(n5047), .A2(n5046), .ZN(n8867) );
  NAND2_X1 U5344 ( .A1(n5335), .A2(n5334), .ZN(n8243) );
  NAND2_X1 U5345 ( .A1(n5570), .A2(n5569), .ZN(n6753) );
  AND2_X1 U5346 ( .A1(n6757), .A2(n6856), .ZN(n6770) );
  INV_X1 U5347 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8940) );
  NAND2_X1 U5348 ( .A1(n5510), .A2(n4360), .ZN(n5505) );
  NOR2_X1 U5349 ( .A1(n4347), .A2(n4495), .ZN(n4494) );
  AOI21_X1 U5350 ( .B1(n6470), .B2(n6469), .A(n4463), .ZN(n6480) );
  AND2_X1 U5351 ( .A1(n5711), .A2(n5712), .ZN(n4463) );
  AND3_X1 U5352 ( .A1(n5980), .A2(n5979), .A3(n5978), .ZN(n9350) );
  AND2_X1 U5353 ( .A1(n6018), .A2(n6017), .ZN(n9313) );
  NAND2_X1 U5354 ( .A1(n5950), .A2(n5949), .ZN(n9360) );
  OR2_X1 U5355 ( .A1(n9257), .A2(n6058), .ZN(n6065) );
  AND2_X1 U5356 ( .A1(n6034), .A2(n6033), .ZN(n9301) );
  NAND2_X1 U5357 ( .A1(n6176), .A2(n9211), .ZN(n9035) );
  AND2_X1 U5358 ( .A1(n6001), .A2(n6000), .ZN(n9298) );
  AND4_X1 U5359 ( .A1(n6097), .A2(n6096), .A3(n6095), .A4(n6094), .ZN(n9240)
         );
  INV_X1 U5360 ( .A(n9238), .ZN(n9274) );
  INV_X1 U5361 ( .A(n6253), .ZN(n9336) );
  AND2_X1 U5362 ( .A1(n5698), .A2(n5697), .ZN(n5701) );
  NOR2_X1 U5363 ( .A1(n9544), .A2(n4539), .ZN(n9559) );
  AND2_X1 U5364 ( .A1(n9549), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4539) );
  INV_X1 U5365 ( .A(n7558), .ZN(n9081) );
  INV_X1 U5366 ( .A(n9368), .ZN(n9209) );
  OR2_X1 U5367 ( .A1(n9375), .A2(n9374), .ZN(n4899) );
  AND2_X1 U5368 ( .A1(n9373), .A2(n9430), .ZN(n9374) );
  INV_X1 U5369 ( .A(n9441), .ZN(n4421) );
  NAND2_X1 U5370 ( .A1(n6055), .A2(n6054), .ZN(n9458) );
  NAND2_X1 U5371 ( .A1(n5876), .A2(n5875), .ZN(n7446) );
  AND2_X1 U5372 ( .A1(n4397), .A2(n4809), .ZN(n4515) );
  INV_X1 U5373 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U5374 ( .A1(n4544), .A2(n4541), .ZN(n8000) );
  OR2_X1 U5375 ( .A1(n7994), .A2(n8167), .ZN(n4544) );
  NAND2_X1 U5376 ( .A1(n8021), .A2(n4566), .ZN(n8029) );
  NAND2_X1 U5377 ( .A1(n4567), .A2(n8085), .ZN(n4566) );
  NAND2_X1 U5378 ( .A1(n4545), .A2(n8149), .ZN(n8045) );
  NAND2_X1 U5379 ( .A1(n8051), .A2(n8042), .ZN(n4545) );
  MUX2_X1 U5380 ( .A(n7969), .B(n7968), .S(n8167), .Z(n8069) );
  INV_X1 U5381 ( .A(n5022), .ZN(n4641) );
  INV_X1 U5382 ( .A(n5342), .ZN(n4969) );
  NOR2_X1 U5383 ( .A1(n4454), .A2(n4953), .ZN(n4453) );
  INV_X1 U5384 ( .A(n4951), .ZN(n4454) );
  AND2_X1 U5385 ( .A1(n5267), .A2(SI_11_), .ZN(n4953) );
  OAI21_X1 U5386 ( .B1(n4365), .B2(n4427), .A(n4426), .ZN(n7831) );
  AOI21_X1 U5387 ( .B1(n7352), .B2(n5283), .A(n5285), .ZN(n5288) );
  NOR2_X1 U5388 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5026) );
  NAND2_X1 U5389 ( .A1(n4562), .A2(n8085), .ZN(n4557) );
  INV_X1 U5390 ( .A(n4562), .ZN(n4561) );
  AND2_X1 U5391 ( .A1(n4564), .A2(n9182), .ZN(n4563) );
  NOR2_X1 U5392 ( .A1(n8086), .A2(n4565), .ZN(n4564) );
  OAI22_X1 U5393 ( .A1(n8083), .A2(n8167), .B1(n8085), .B2(n8076), .ZN(n4565)
         );
  NAND2_X1 U5394 ( .A1(n8199), .A2(n8087), .ZN(n8086) );
  NOR2_X1 U5395 ( .A1(n6502), .A2(n6152), .ZN(n4788) );
  AND2_X1 U5396 ( .A1(n8066), .A2(n7922), .ZN(n7967) );
  AND2_X1 U5397 ( .A1(n6269), .A2(n9251), .ZN(n7919) );
  INV_X1 U5398 ( .A(n4507), .ZN(n4504) );
  INV_X1 U5399 ( .A(n5012), .ZN(n4649) );
  INV_X1 U5400 ( .A(n4989), .ZN(n4663) );
  INV_X1 U5401 ( .A(SI_19_), .ZN(n4981) );
  NAND2_X1 U5402 ( .A1(n4657), .A2(n4656), .ZN(n4652) );
  NOR2_X1 U5403 ( .A1(n4971), .A2(n4655), .ZN(n4654) );
  INV_X1 U5404 ( .A(n4656), .ZN(n4655) );
  INV_X1 U5405 ( .A(SI_17_), .ZN(n4972) );
  INV_X1 U5406 ( .A(SI_15_), .ZN(n4658) );
  INV_X1 U5407 ( .A(SI_12_), .ZN(n10052) );
  INV_X1 U5408 ( .A(n4636), .ZN(n4434) );
  OAI21_X1 U5409 ( .B1(n4638), .B2(n4637), .A(n5233), .ZN(n4636) );
  INV_X1 U5410 ( .A(n4940), .ZN(n4637) );
  INV_X1 U5411 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n4942) );
  INV_X1 U5412 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4902) );
  AND2_X1 U5413 ( .A1(n4852), .A2(n4854), .ZN(n4851) );
  NAND2_X1 U5414 ( .A1(n8324), .A2(n8646), .ZN(n4854) );
  NAND2_X1 U5415 ( .A1(n8325), .A2(n4853), .ZN(n4852) );
  NAND2_X1 U5416 ( .A1(n9747), .A2(n4414), .ZN(n8509) );
  OR2_X1 U5417 ( .A1(n9746), .A2(n8508), .ZN(n4414) );
  NAND2_X1 U5418 ( .A1(n9779), .A2(n4413), .ZN(n8511) );
  OR2_X1 U5419 ( .A1(n9778), .A2(n10029), .ZN(n4413) );
  NAND2_X1 U5420 ( .A1(n9813), .A2(n4415), .ZN(n8514) );
  OR2_X1 U5421 ( .A1(n9812), .A2(n8513), .ZN(n4415) );
  INV_X1 U5422 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5028) );
  OR2_X1 U5423 ( .A1(n5546), .A2(n4774), .ZN(n4773) );
  OR2_X1 U5424 ( .A1(n5546), .A2(n4771), .ZN(n4770) );
  NAND2_X1 U5425 ( .A1(n7644), .A2(n7645), .ZN(n4771) );
  INV_X1 U5426 ( .A(n5494), .ZN(n8608) );
  OR2_X1 U5427 ( .A1(n5274), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5276) );
  OR2_X1 U5428 ( .A1(n5248), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5274) );
  AOI21_X1 U5429 ( .B1(n4626), .B2(n5180), .A(n4336), .ZN(n4625) );
  NOR2_X1 U5430 ( .A1(n7700), .A2(n4758), .ZN(n4766) );
  AOI21_X1 U5431 ( .B1(n4766), .B2(n4762), .A(n7704), .ZN(n4761) );
  INV_X1 U5432 ( .A(n7710), .ZN(n4762) );
  INV_X1 U5433 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10017) );
  NAND2_X1 U5434 ( .A1(n5117), .A2(n4618), .ZN(n4617) );
  NAND2_X1 U5435 ( .A1(n4325), .A2(n4619), .ZN(n4618) );
  INV_X1 U5436 ( .A(n4623), .ZN(n4620) );
  INV_X1 U5437 ( .A(n5415), .ZN(n4600) );
  OAI21_X1 U5438 ( .B1(n4603), .B2(n4600), .A(n8709), .ZN(n4599) );
  AND2_X1 U5439 ( .A1(n7787), .A2(n4744), .ZN(n4743) );
  NAND2_X1 U5440 ( .A1(n4747), .A2(n4745), .ZN(n4744) );
  INV_X1 U5441 ( .A(n7778), .ZN(n4745) );
  INV_X1 U5442 ( .A(n4747), .ZN(n4746) );
  INV_X1 U5443 ( .A(n7769), .ZN(n4782) );
  INV_X1 U5444 ( .A(n4784), .ZN(n4779) );
  NOR2_X1 U5445 ( .A1(n5288), .A2(n7257), .ZN(n4613) );
  OR2_X1 U5446 ( .A1(n8408), .A2(n8238), .ZN(n7751) );
  OR2_X1 U5447 ( .A1(n6759), .A2(n6758), .ZN(n6773) );
  NOR2_X1 U5448 ( .A1(n6820), .A2(n6758), .ZN(n6768) );
  OAI21_X1 U5449 ( .B1(n4447), .B2(n4339), .A(n4446), .ZN(n4449) );
  INV_X1 U5450 ( .A(n6048), .ZN(n4447) );
  NAND2_X1 U5451 ( .A1(n4867), .A2(n6050), .ZN(n4446) );
  NAND2_X1 U5452 ( .A1(n4410), .A2(n4484), .ZN(n4483) );
  INV_X1 U5453 ( .A(n4490), .ZN(n4484) );
  AND2_X1 U5454 ( .A1(n5828), .A2(n5827), .ZN(n5861) );
  AND2_X1 U5455 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n5827) );
  NOR2_X1 U5456 ( .A1(n5809), .A2(n5808), .ZN(n5828) );
  NOR2_X1 U5457 ( .A1(n5938), .A2(n5937), .ZN(n5921) );
  OAI21_X1 U5458 ( .B1(n4556), .B2(n4384), .A(n4552), .ZN(n4550) );
  AOI21_X1 U5459 ( .B1(n4553), .B2(n4554), .A(n7937), .ZN(n4552) );
  INV_X1 U5460 ( .A(n8101), .ZN(n4553) );
  NOR2_X1 U5461 ( .A1(n9398), .A2(n9458), .ZN(n4574) );
  OR2_X1 U5462 ( .A1(n6027), .A2(n6026), .ZN(n6039) );
  INV_X1 U5463 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5975) );
  OR2_X1 U5464 ( .A1(n9429), .A2(n9348), .ZN(n8141) );
  NAND2_X1 U5465 ( .A1(n4588), .A2(n4587), .ZN(n7569) );
  NOR2_X1 U5466 ( .A1(n7484), .A2(n6277), .ZN(n4579) );
  NAND2_X1 U5467 ( .A1(n4392), .A2(n4704), .ZN(n8108) );
  NOR2_X1 U5468 ( .A1(n6262), .A2(n7986), .ZN(n4704) );
  NOR2_X1 U5469 ( .A1(n6841), .A2(n7107), .ZN(n6840) );
  NAND2_X1 U5470 ( .A1(n6551), .A2(n8118), .ZN(n6540) );
  INV_X1 U5471 ( .A(n7935), .ZN(n6324) );
  OR2_X1 U5472 ( .A1(n9458), .A2(n9238), .ZN(n8065) );
  INV_X1 U5473 ( .A(n4510), .ZN(n4506) );
  OR2_X1 U5474 ( .A1(n7022), .A2(n7024), .ZN(n7146) );
  NAND2_X1 U5475 ( .A1(n6562), .A2(n9108), .ZN(n8114) );
  OAI21_X1 U5476 ( .B1(n7610), .B2(n7609), .A(n7608), .ZN(n7633) );
  OR2_X1 U5477 ( .A1(n7607), .A2(n7606), .ZN(n7608) );
  INV_X1 U5478 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5592) );
  AND2_X1 U5479 ( .A1(n5022), .A2(n5021), .ZN(n5088) );
  AND2_X1 U5480 ( .A1(n5017), .A2(n5016), .ZN(n5474) );
  AND2_X1 U5481 ( .A1(n5006), .A2(n5005), .ZN(n5450) );
  NOR2_X1 U5482 ( .A1(n4990), .A2(n4666), .ZN(n4665) );
  INV_X1 U5483 ( .A(n4667), .ZN(n4666) );
  NAND2_X1 U5484 ( .A1(n4968), .A2(n4658), .ZN(n4656) );
  NOR2_X1 U5485 ( .A1(n4968), .A2(n4658), .ZN(n4657) );
  AND2_X1 U5486 ( .A1(n5594), .A2(n5593), .ZN(n5899) );
  INV_X1 U5487 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5595) );
  OR2_X1 U5488 ( .A1(n4963), .A2(n4962), .ZN(n4964) );
  OR2_X1 U5489 ( .A1(n5254), .A2(n4963), .ZN(n4965) );
  NAND2_X1 U5490 ( .A1(n4451), .A2(n4452), .ZN(n5255) );
  NOR2_X2 U5491 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5752) );
  OAI21_X1 U5492 ( .B1(n4986), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n4913), .ZN(
        n4914) );
  OR2_X1 U5493 ( .A1(n8277), .A2(n8636), .ZN(n4855) );
  INV_X1 U5494 ( .A(n4851), .ZN(n4849) );
  NAND2_X1 U5495 ( .A1(n4817), .A2(n4815), .ZN(n8334) );
  AOI21_X1 U5496 ( .B1(n4818), .B2(n4821), .A(n4816), .ZN(n4815) );
  INV_X1 U5497 ( .A(n8333), .ZN(n4816) );
  AOI21_X1 U5498 ( .B1(n4831), .B2(n4830), .A(n4367), .ZN(n4829) );
  INV_X1 U5499 ( .A(n7227), .ZN(n4830) );
  OR2_X1 U5500 ( .A1(n8400), .A2(n8401), .ZN(n8398) );
  XNOR2_X1 U5501 ( .A(n6784), .B(n8851), .ZN(n6781) );
  INV_X1 U5502 ( .A(n5522), .ZN(n6775) );
  NOR2_X1 U5503 ( .A1(n7605), .A2(n7604), .ZN(n7642) );
  AND2_X1 U5504 ( .A1(n4839), .A2(n7131), .ZN(n7856) );
  AND2_X1 U5505 ( .A1(n4839), .A2(n8592), .ZN(n7857) );
  AND4_X1 U5506 ( .A1(n5381), .A2(n5380), .A3(n5379), .A4(n5378), .ZN(n8250)
         );
  AND4_X1 U5507 ( .A1(n5140), .A2(n5139), .A3(n5138), .A4(n5137), .ZN(n8839)
         );
  XNOR2_X1 U5508 ( .A(n8483), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U5509 ( .A1(n8477), .A2(n8478), .ZN(n8476) );
  NAND2_X1 U5510 ( .A1(n6588), .A2(n9691), .ZN(n9696) );
  INV_X1 U5511 ( .A(n4698), .ZN(n4697) );
  OAI21_X1 U5512 ( .B1(n9691), .B2(n4354), .A(n6660), .ZN(n4698) );
  INV_X1 U5513 ( .A(n6908), .ZN(n4679) );
  AOI21_X1 U5514 ( .B1(n6908), .B2(n4678), .A(n4677), .ZN(n4676) );
  NAND2_X1 U5515 ( .A1(n6670), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6909) );
  NAND2_X1 U5516 ( .A1(n9748), .A2(n9749), .ZN(n9747) );
  NAND2_X1 U5517 ( .A1(n9780), .A2(n9781), .ZN(n9779) );
  OR2_X1 U5518 ( .A1(n5270), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5300) );
  OAI22_X1 U5519 ( .A1(n4691), .A2(n9789), .B1(n9773), .B2(n4689), .ZN(n9788)
         );
  NAND2_X1 U5520 ( .A1(n8496), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4689) );
  NOR2_X1 U5521 ( .A1(n5300), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U5522 ( .A1(n9814), .A2(n9815), .ZN(n9813) );
  INV_X1 U5523 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5331) );
  XNOR2_X1 U5524 ( .A(n8575), .B(n8566), .ZN(n8516) );
  NAND2_X1 U5525 ( .A1(n8516), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8577) );
  AND2_X1 U5526 ( .A1(n4409), .A2(n4688), .ZN(n4686) );
  INV_X1 U5527 ( .A(n8589), .ZN(n4688) );
  AOI21_X1 U5528 ( .B1(n8562), .B2(n4686), .A(n4685), .ZN(n4684) );
  NOR2_X1 U5529 ( .A1(n4688), .A2(n4409), .ZN(n4685) );
  NOR2_X1 U5530 ( .A1(n8461), .A2(n8867), .ZN(n4591) );
  NAND2_X1 U5531 ( .A1(n5070), .A2(n5069), .ZN(n5092) );
  INV_X1 U5532 ( .A(n8461), .ZN(n8635) );
  OR2_X1 U5533 ( .A1(n7827), .A2(n7828), .ZN(n8632) );
  NAND2_X1 U5534 ( .A1(n5066), .A2(n5065), .ZN(n5466) );
  NAND2_X1 U5535 ( .A1(n5064), .A2(n5063), .ZN(n5436) );
  INV_X1 U5536 ( .A(n5423), .ZN(n5064) );
  OR2_X1 U5537 ( .A1(n5436), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U5538 ( .A1(n5062), .A2(n5061), .ZN(n5407) );
  NAND2_X1 U5539 ( .A1(n5060), .A2(n5059), .ZN(n5377) );
  INV_X1 U5540 ( .A(n5375), .ZN(n5060) );
  INV_X1 U5541 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5057) );
  INV_X1 U5542 ( .A(n5336), .ZN(n5058) );
  OR2_X1 U5543 ( .A1(n5351), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5375) );
  OR2_X1 U5544 ( .A1(n5320), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U5545 ( .A1(n5054), .A2(n7417), .ZN(n5305) );
  INV_X1 U5546 ( .A(n5276), .ZN(n5054) );
  NAND2_X1 U5547 ( .A1(n5056), .A2(n5055), .ZN(n5320) );
  INV_X1 U5548 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5055) );
  INV_X1 U5549 ( .A(n5305), .ZN(n5056) );
  NAND2_X1 U5550 ( .A1(n4752), .A2(n4750), .ZN(n7348) );
  AOI21_X1 U5551 ( .B1(n4753), .B2(n4755), .A(n4751), .ZN(n4750) );
  INV_X1 U5552 ( .A(n7742), .ZN(n4751) );
  AND2_X1 U5553 ( .A1(n7758), .A2(n7755), .ZN(n7656) );
  NAND2_X1 U5554 ( .A1(n5053), .A2(n5052), .ZN(n5248) );
  INV_X1 U5555 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5052) );
  INV_X1 U5556 ( .A(n5227), .ZN(n5053) );
  OR2_X1 U5557 ( .A1(n5208), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5227) );
  OR2_X1 U5558 ( .A1(n5181), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5195) );
  AND2_X1 U5559 ( .A1(n4624), .A2(n4625), .ZN(n7034) );
  NAND2_X1 U5560 ( .A1(n4628), .A2(n5179), .ZN(n6964) );
  NAND2_X1 U5561 ( .A1(n4629), .A2(n4630), .ZN(n4628) );
  INV_X1 U5562 ( .A(n6810), .ZN(n4629) );
  INV_X1 U5563 ( .A(n5161), .ZN(n6849) );
  INV_X1 U5564 ( .A(n8837), .ZN(n8833) );
  NAND2_X1 U5565 ( .A1(n6822), .A2(n6821), .ZN(n6823) );
  AND2_X1 U5566 ( .A1(n6820), .A2(n6819), .ZN(n6821) );
  OR2_X1 U5567 ( .A1(n5528), .A2(n7682), .ZN(n6871) );
  NOR2_X1 U5568 ( .A1(n8846), .A2(n6872), .ZN(n6769) );
  INV_X1 U5569 ( .A(n8632), .ZN(n8630) );
  OAI21_X1 U5570 ( .B1(n8652), .B2(n5543), .A(n7816), .ZN(n8643) );
  OR2_X1 U5571 ( .A1(n7645), .A2(n7822), .ZN(n8644) );
  AND2_X1 U5572 ( .A1(n7815), .A2(n7816), .ZN(n8653) );
  AND2_X1 U5573 ( .A1(n7813), .A2(n7812), .ZN(n8666) );
  AOI21_X1 U5574 ( .B1(n4737), .B2(n4735), .A(n4734), .ZN(n4733) );
  INV_X1 U5575 ( .A(n7804), .ZN(n4734) );
  AND2_X1 U5576 ( .A1(n8724), .A2(n7786), .ZN(n8746) );
  INV_X1 U5577 ( .A(n8743), .ZN(n8755) );
  OAI21_X1 U5578 ( .B1(n5537), .B2(n4780), .A(n4777), .ZN(n8754) );
  INV_X1 U5579 ( .A(n4781), .ZN(n4780) );
  AOI21_X1 U5580 ( .B1(n4781), .B2(n4779), .A(n4778), .ZN(n4777) );
  NOR2_X1 U5581 ( .A1(n5538), .A2(n4782), .ZN(n4781) );
  OAI21_X1 U5582 ( .B1(n4607), .B2(n4439), .A(n4435), .ZN(n8768) );
  AOI21_X1 U5583 ( .B1(n4606), .B2(n4352), .A(n4436), .ZN(n4435) );
  NOR2_X1 U5584 ( .A1(n8459), .A2(n7507), .ZN(n4436) );
  AOI21_X1 U5585 ( .B1(n4614), .B2(n4613), .A(n4609), .ZN(n7274) );
  INV_X1 U5586 ( .A(n5289), .ZN(n4609) );
  AND2_X1 U5587 ( .A1(n7751), .A2(n7750), .ZN(n7760) );
  INV_X1 U5588 ( .A(n7420), .ZN(n7415) );
  NAND2_X1 U5589 ( .A1(n7309), .A2(n7857), .ZN(n8846) );
  NAND2_X1 U5590 ( .A1(n7826), .A2(n7856), .ZN(n7279) );
  INV_X1 U5591 ( .A(n8847), .ZN(n8852) );
  AND2_X1 U5592 ( .A1(n6767), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6856) );
  INV_X1 U5593 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5585) );
  XNOR2_X1 U5594 ( .A(n5078), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5081) );
  AND2_X1 U5595 ( .A1(n4360), .A2(n5506), .ZN(n4835) );
  INV_X1 U5596 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5506) );
  INV_X1 U5597 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5173) );
  INV_X1 U5598 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5040) );
  INV_X1 U5599 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10071) );
  AND2_X1 U5600 ( .A1(n5962), .A2(n5961), .ZN(n9011) );
  INV_X1 U5601 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U5602 ( .A1(n5921), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5952) );
  NAND2_X1 U5603 ( .A1(n5800), .A2(n5799), .ZN(n4476) );
  INV_X1 U5604 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U5605 ( .A1(n5688), .A2(n5686), .ZN(n6400) );
  NOR2_X1 U5606 ( .A1(n7389), .A2(n4880), .ZN(n4879) );
  INV_X1 U5607 ( .A(n5856), .ZN(n4880) );
  OAI22_X1 U5608 ( .A1(n7389), .A2(n4878), .B1(n5870), .B2(n5871), .ZN(n4877)
         );
  INV_X1 U5609 ( .A(n5855), .ZN(n4878) );
  NAND2_X1 U5610 ( .A1(n5861), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5878) );
  INV_X1 U5611 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U5612 ( .A1(n5709), .A2(n5708), .ZN(n5710) );
  OR2_X1 U5613 ( .A1(n6098), .A2(n6212), .ZN(n5708) );
  INV_X1 U5614 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5756) );
  INV_X1 U5615 ( .A(n9068), .ZN(n9076) );
  AND3_X1 U5616 ( .A1(n6282), .A2(n6512), .A3(n6247), .ZN(n6185) );
  INV_X1 U5617 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5937) );
  AOI21_X1 U5618 ( .B1(n8161), .B2(n8160), .A(n8169), .ZN(n8162) );
  AND4_X1 U5619 ( .A1(n6184), .A2(n6183), .A3(n6182), .A4(n6181), .ZN(n7929)
         );
  AND3_X1 U5620 ( .A1(n5956), .A2(n5955), .A3(n5954), .ZN(n6253) );
  AND2_X1 U5621 ( .A1(n5943), .A2(n5942), .ZN(n9001) );
  AND2_X1 U5622 ( .A1(n6447), .A2(n6446), .ZN(n6444) );
  OR2_X1 U5623 ( .A1(n6357), .A2(n6356), .ZN(n4530) );
  OR2_X1 U5624 ( .A1(n6377), .A2(n6376), .ZN(n4528) );
  NOR2_X1 U5625 ( .A1(n9512), .A2(n4536), .ZN(n9526) );
  AND2_X1 U5626 ( .A1(n9520), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4536) );
  NAND2_X1 U5627 ( .A1(n9526), .A2(n9527), .ZN(n9525) );
  XNOR2_X1 U5628 ( .A(n9127), .B(n9577), .ZN(n9573) );
  NOR2_X1 U5629 ( .A1(n9566), .A2(n9567), .ZN(n9568) );
  NAND2_X1 U5630 ( .A1(n9588), .A2(n9589), .ZN(n9587) );
  OR2_X1 U5631 ( .A1(n9583), .A2(n9582), .ZN(n4526) );
  AOI22_X1 U5632 ( .A1(n9598), .A2(n9597), .B1(n9149), .B2(n9425), .ZN(n9613)
         );
  NOR2_X1 U5633 ( .A1(n4582), .A2(n9169), .ZN(n4581) );
  INV_X1 U5634 ( .A(n4582), .ZN(n4580) );
  OR2_X1 U5635 ( .A1(n9373), .A2(n8196), .ZN(n9182) );
  INV_X1 U5636 ( .A(n7963), .ZN(n9207) );
  AOI21_X1 U5637 ( .B1(n9248), .B2(n4708), .A(n4707), .ZN(n4706) );
  NOR2_X1 U5638 ( .A1(n4710), .A2(n7918), .ZN(n4707) );
  NAND2_X1 U5639 ( .A1(n9221), .A2(n9222), .ZN(n9220) );
  NAND2_X1 U5640 ( .A1(n9265), .A2(n4338), .ZN(n9228) );
  NAND2_X1 U5641 ( .A1(n9265), .A2(n6278), .ZN(n9266) );
  INV_X1 U5642 ( .A(n9464), .ZN(n9288) );
  NAND2_X1 U5643 ( .A1(n6012), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6027) );
  OR2_X1 U5644 ( .A1(n4728), .A2(n4726), .ZN(n4723) );
  NOR2_X1 U5645 ( .A1(n8040), .A2(n4729), .ZN(n4728) );
  INV_X1 U5646 ( .A(n4588), .ZN(n7570) );
  INV_X1 U5647 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5650) );
  INV_X1 U5648 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5970) );
  NOR3_X1 U5649 ( .A1(n7146), .A2(n4578), .A3(n7446), .ZN(n7491) );
  NOR2_X1 U5650 ( .A1(n7146), .A2(n6277), .ZN(n7460) );
  NOR2_X1 U5651 ( .A1(n7146), .A2(n4577), .ZN(n7462) );
  INV_X1 U5652 ( .A(n4579), .ZN(n4577) );
  NAND2_X1 U5653 ( .A1(n8129), .A2(n8108), .ZN(n4703) );
  AND2_X1 U5654 ( .A1(n8005), .A2(n8010), .ZN(n7141) );
  INV_X1 U5655 ( .A(n7141), .ZN(n7951) );
  NAND2_X1 U5656 ( .A1(n6840), .A2(n7195), .ZN(n7022) );
  NAND2_X1 U5657 ( .A1(n4498), .A2(n4497), .ZN(n7021) );
  AOI21_X1 U5658 ( .B1(n6949), .B2(n4499), .A(n4343), .ZN(n4497) );
  INV_X1 U5659 ( .A(n6221), .ZN(n4499) );
  OR2_X1 U5660 ( .A1(n6222), .A2(n6263), .ZN(n7020) );
  INV_X1 U5661 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5787) );
  OR2_X1 U5662 ( .A1(n5788), .A2(n5787), .ZN(n5809) );
  NAND2_X1 U5663 ( .A1(n4570), .A2(n9632), .ZN(n6841) );
  INV_X1 U5664 ( .A(n7990), .ZN(n4714) );
  NAND2_X1 U5665 ( .A1(n6540), .A2(n7981), .ZN(n6539) );
  AND2_X1 U5666 ( .A1(n6136), .A2(n9482), .ZN(n6282) );
  OR2_X1 U5667 ( .A1(n6314), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U5668 ( .A1(n4808), .A2(n4383), .ZN(n4803) );
  NAND2_X1 U5669 ( .A1(n4524), .A2(n4523), .ZN(n9219) );
  AOI21_X1 U5670 ( .B1(n4806), .B2(n4348), .A(n4400), .ZN(n4523) );
  NAND2_X1 U5671 ( .A1(n5974), .A2(n5973), .ZN(n9417) );
  NAND2_X1 U5672 ( .A1(n7492), .A2(n9097), .ZN(n4520) );
  NOR2_X1 U5673 ( .A1(n7492), .A2(n9097), .ZN(n4519) );
  AND2_X1 U5674 ( .A1(n8137), .A2(n8134), .ZN(n7955) );
  INV_X1 U5675 ( .A(n9645), .ZN(n9430) );
  INV_X1 U5676 ( .A(n4798), .ZN(n7463) );
  OR2_X1 U5677 ( .A1(n7144), .A2(n4799), .ZN(n4798) );
  INV_X1 U5678 ( .A(n6259), .ZN(n7945) );
  NAND2_X1 U5679 ( .A1(n8114), .A2(n8118), .ZN(n7946) );
  NAND2_X1 U5680 ( .A1(n4569), .A2(n6215), .ZN(n6556) );
  INV_X1 U5681 ( .A(n6501), .ZN(n4569) );
  INV_X1 U5682 ( .A(n6282), .ZN(n6513) );
  AND2_X1 U5683 ( .A1(n6248), .A2(n6511), .ZN(n6283) );
  AND2_X1 U5684 ( .A1(n5631), .A2(n5606), .ZN(n5636) );
  XNOR2_X1 U5685 ( .A(n5488), .B(n5487), .ZN(n7565) );
  XNOR2_X1 U5686 ( .A(n5087), .B(n5088), .ZN(n7563) );
  INV_X1 U5687 ( .A(n5603), .ZN(n4516) );
  NAND2_X1 U5688 ( .A1(n4668), .A2(n4667), .ZN(n5416) );
  AND2_X1 U5689 ( .A1(n5299), .A2(n5298), .ZN(n6507) );
  OR2_X1 U5690 ( .A1(n5837), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5857) );
  OAI21_X1 U5691 ( .B1(n5243), .B2(n4952), .A(n4951), .ZN(n5269) );
  NAND2_X1 U5692 ( .A1(n4635), .A2(n4940), .ZN(n5234) );
  NAND2_X1 U5693 ( .A1(n4934), .A2(n4638), .ZN(n4635) );
  NAND2_X1 U5694 ( .A1(n4444), .A2(n4930), .ZN(n5204) );
  NAND2_X1 U5695 ( .A1(n4416), .A2(n4922), .ZN(n5176) );
  INV_X1 U5696 ( .A(n4918), .ZN(n4460) );
  INV_X1 U5697 ( .A(n4909), .ZN(n5104) );
  NAND2_X1 U5698 ( .A1(n8398), .A2(n8242), .ZN(n8284) );
  NAND2_X1 U5699 ( .A1(n4822), .A2(n4827), .ZN(n8447) );
  NAND2_X1 U5700 ( .A1(n8400), .A2(n8242), .ZN(n4822) );
  NAND2_X1 U5701 ( .A1(n8422), .A2(n8258), .ZN(n8391) );
  NAND2_X1 U5702 ( .A1(n7005), .A2(n7004), .ZN(n7044) );
  INV_X1 U5703 ( .A(n8691), .ZN(n8382) );
  NAND2_X1 U5704 ( .A1(n4834), .A2(n7231), .ZN(n7235) );
  NAND2_X1 U5705 ( .A1(n4834), .A2(n4831), .ZN(n7405) );
  AND4_X1 U5706 ( .A1(n5200), .A2(n5199), .A3(n5198), .A4(n5197), .ZN(n7216)
         );
  NAND2_X1 U5707 ( .A1(n4857), .A2(n4375), .ZN(n4856) );
  AND2_X1 U5708 ( .A1(n5472), .A2(n5471), .ZN(n8441) );
  INV_X1 U5709 ( .A(n9945), .ZN(n8440) );
  INV_X1 U5710 ( .A(n4827), .ZN(n4826) );
  AND2_X1 U5711 ( .A1(n8245), .A2(n4824), .ZN(n4823) );
  NAND2_X1 U5712 ( .A1(n5484), .A2(n5483), .ZN(n8655) );
  INV_X1 U5713 ( .A(n8441), .ZN(n8668) );
  INV_X1 U5714 ( .A(n8250), .ZN(n8772) );
  OR2_X2 U5715 ( .A1(n6610), .A2(P2_U3151), .ZN(n8474) );
  INV_X1 U5716 ( .A(n4690), .ZN(n9772) );
  INV_X1 U5717 ( .A(n4695), .ZN(n9838) );
  NAND2_X1 U5718 ( .A1(n6612), .A2(n6611), .ZN(n9846) );
  INV_X1 U5719 ( .A(n8502), .ZN(n4694) );
  INV_X1 U5720 ( .A(n9664), .ZN(n9856) );
  NAND2_X1 U5721 ( .A1(n4687), .A2(n4684), .ZN(n4683) );
  OR2_X1 U5722 ( .A1(n8562), .A2(n4688), .ZN(n4687) );
  AOI21_X1 U5723 ( .B1(n7894), .B2(n7635), .A(n7621), .ZN(n8610) );
  XNOR2_X1 U5724 ( .A(n7605), .B(n7643), .ZN(n8614) );
  NAND2_X1 U5725 ( .A1(n4595), .A2(n5441), .ZN(n8677) );
  NAND2_X1 U5726 ( .A1(n8690), .A2(n8689), .ZN(n4595) );
  NAND2_X1 U5727 ( .A1(n5445), .A2(n5444), .ZN(n8804) );
  NAND2_X1 U5728 ( .A1(n8715), .A2(n5415), .ZN(n8698) );
  NAND2_X1 U5729 ( .A1(n4442), .A2(n5272), .ZN(n9949) );
  NAND2_X1 U5730 ( .A1(n7201), .A2(n7739), .ZN(n7255) );
  NAND2_X1 U5731 ( .A1(n5531), .A2(n7706), .ZN(n7031) );
  OR2_X1 U5732 ( .A1(n6823), .A2(n9866), .ZN(n8613) );
  INV_X1 U5733 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7081) );
  INV_X1 U5734 ( .A(n9869), .ZN(n8777) );
  AND3_X1 U5735 ( .A1(n5131), .A2(n5130), .A3(n5129), .ZN(n9867) );
  NAND2_X1 U5736 ( .A1(n8852), .A2(n7861), .ZN(n9866) );
  INV_X1 U5737 ( .A(n5119), .ZN(n8851) );
  NAND2_X1 U5738 ( .A1(n7638), .A2(n7637), .ZN(n8861) );
  XNOR2_X1 U5739 ( .A(n4592), .B(n4356), .ZN(n8625) );
  AND2_X1 U5740 ( .A1(n4775), .A2(n4774), .ZN(n8623) );
  NAND2_X1 U5741 ( .A1(n8631), .A2(n7644), .ZN(n4775) );
  NAND2_X1 U5742 ( .A1(n5476), .A2(n5475), .ZN(n8877) );
  NAND2_X1 U5743 ( .A1(n5465), .A2(n5464), .ZN(n8883) );
  NAND2_X1 U5744 ( .A1(n5452), .A2(n5451), .ZN(n8889) );
  NAND2_X1 U5745 ( .A1(n5435), .A2(n5434), .ZN(n8899) );
  NAND2_X1 U5746 ( .A1(n8708), .A2(n7795), .ZN(n4739) );
  NOR2_X1 U5747 ( .A1(n4602), .A2(n4601), .ZN(n8717) );
  INV_X1 U5748 ( .A(n5400), .ZN(n4601) );
  NAND2_X1 U5749 ( .A1(n5406), .A2(n5405), .ZN(n8909) );
  NAND2_X1 U5750 ( .A1(n4749), .A2(n4747), .ZN(n8725) );
  NAND2_X1 U5751 ( .A1(n5362), .A2(n5361), .ZN(n8921) );
  NAND2_X1 U5752 ( .A1(n5374), .A2(n5373), .ZN(n8927) );
  NAND2_X1 U5753 ( .A1(n5350), .A2(n5349), .ZN(n8934) );
  NAND2_X1 U5754 ( .A1(n4783), .A2(n7769), .ZN(n8766) );
  NAND2_X1 U5755 ( .A1(n5537), .A2(n4784), .ZN(n4783) );
  NAND2_X1 U5756 ( .A1(n4438), .A2(n5327), .ZN(n7509) );
  NAND2_X1 U5757 ( .A1(n5537), .A2(n7768), .ZN(n7508) );
  NAND2_X1 U5758 ( .A1(n4608), .A2(n4610), .ZN(n7374) );
  AND2_X1 U5759 ( .A1(n4605), .A2(n4611), .ZN(n4610) );
  INV_X2 U5760 ( .A(n9898), .ZN(n9901) );
  CLKBUF_X2 U5761 ( .A(n6716), .Z(n6740) );
  XNOR2_X1 U5762 ( .A(n5584), .B(n5585), .ZN(n6767) );
  NAND2_X1 U5763 ( .A1(n5566), .A2(n5565), .ZN(n7541) );
  INV_X1 U5764 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5556) );
  INV_X1 U5765 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7225) );
  NAND2_X1 U5766 ( .A1(n5510), .A2(n5503), .ZN(n5508) );
  INV_X1 U5767 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7130) );
  INV_X1 U5768 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7014) );
  INV_X1 U5769 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6998) );
  INV_X1 U5770 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10068) );
  INV_X1 U5771 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6340) );
  INV_X1 U5772 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9984) );
  INV_X1 U5773 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6305) );
  OR2_X1 U5774 ( .A1(n5189), .A2(n5188), .ZN(n9714) );
  XNOR2_X1 U5775 ( .A(n6150), .B(n6149), .ZN(n6323) );
  OAI21_X1 U5776 ( .B1(n4488), .B2(n4486), .A(n5769), .ZN(n4485) );
  AND4_X1 U5777 ( .A1(n5883), .A2(n5882), .A3(n5881), .A4(n5880), .ZN(n8955)
         );
  INV_X1 U5778 ( .A(n6213), .ZN(n7877) );
  AND2_X1 U5779 ( .A1(n5996), .A2(n5995), .ZN(n9318) );
  NAND2_X1 U5780 ( .A1(n9066), .A2(n4455), .ZN(n6203) );
  NOR2_X1 U5781 ( .A1(n4347), .A2(n4456), .ZN(n4455) );
  INV_X1 U5782 ( .A(n6121), .ZN(n4456) );
  AND4_X1 U5783 ( .A1(n5814), .A2(n5813), .A3(n5812), .A4(n5811), .ZN(n7454)
         );
  INV_X1 U5784 ( .A(n4477), .ZN(n7190) );
  XNOR2_X1 U5785 ( .A(n6045), .B(n4459), .ZN(n8981) );
  AND4_X1 U5786 ( .A1(n5833), .A2(n5832), .A3(n5831), .A4(n5830), .ZN(n7391)
         );
  AOI21_X1 U5787 ( .B1(n9039), .B2(n5856), .A(n5855), .ZN(n7388) );
  INV_X1 U5788 ( .A(n4886), .ZN(n4884) );
  NAND2_X1 U5789 ( .A1(n4465), .A2(n4464), .ZN(n8182) );
  INV_X1 U5790 ( .A(n4469), .ZN(n4465) );
  NAND2_X1 U5791 ( .A1(n4468), .A2(n8962), .ZN(n4464) );
  NOR2_X1 U5792 ( .A1(n6745), .A2(n6746), .ZN(n6744) );
  INV_X1 U5793 ( .A(n4475), .ZN(n7292) );
  NAND2_X1 U5794 ( .A1(n6011), .A2(n6010), .ZN(n9408) );
  INV_X1 U5795 ( .A(n4873), .ZN(n7499) );
  AOI21_X1 U5796 ( .B1(n9039), .B2(n4879), .A(n4877), .ZN(n4873) );
  OAI21_X1 U5797 ( .B1(n8976), .B2(n6050), .A(n4867), .ZN(n9028) );
  AND2_X1 U5798 ( .A1(n4866), .A2(n6048), .ZN(n9029) );
  NAND2_X1 U5799 ( .A1(n4862), .A2(n4401), .ZN(n4866) );
  AND4_X1 U5800 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(n9046)
         );
  NAND2_X1 U5801 ( .A1(n5693), .A2(n5692), .ZN(n5694) );
  INV_X1 U5802 ( .A(n4486), .ZN(n4489) );
  NAND2_X1 U5803 ( .A1(n4881), .A2(n6106), .ZN(n9065) );
  AND2_X1 U5804 ( .A1(n6159), .A2(n6111), .ZN(n9210) );
  NAND2_X1 U5805 ( .A1(n6185), .A2(n8176), .ZN(n9078) );
  OR2_X1 U5806 ( .A1(n6191), .A2(n7399), .ZN(n9084) );
  NOR4_X1 U5807 ( .A1(n8169), .A2(n8107), .A3(n8156), .A4(n7965), .ZN(n8104)
         );
  OR2_X1 U5808 ( .A1(n5657), .A2(n5656), .ZN(n5658) );
  INV_X1 U5809 ( .A(n7934), .ZN(n8098) );
  INV_X1 U5810 ( .A(n9313), .ZN(n9093) );
  INV_X1 U5811 ( .A(n9350), .ZN(n9094) );
  INV_X1 U5812 ( .A(n9348), .ZN(n9095) );
  INV_X1 U5813 ( .A(n6216), .ZN(n9108) );
  NAND2_X1 U5814 ( .A1(n4329), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5671) );
  NOR2_X1 U5815 ( .A1(n6440), .A2(n4382), .ZN(n6392) );
  INV_X1 U5816 ( .A(n4532), .ZN(n6390) );
  NOR2_X1 U5817 ( .A1(n6407), .A2(n6406), .ZN(n6405) );
  AND2_X1 U5818 ( .A1(n4532), .A2(n4531), .ZN(n6407) );
  NAND2_X1 U5819 ( .A1(n6387), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4531) );
  INV_X1 U5820 ( .A(n4530), .ZN(n6375) );
  AND2_X1 U5821 ( .A1(n4530), .A2(n4529), .ZN(n6377) );
  NAND2_X1 U5822 ( .A1(n6379), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4529) );
  INV_X1 U5823 ( .A(n4528), .ZN(n6416) );
  AND2_X1 U5824 ( .A1(n4528), .A2(n4527), .ZN(n6420) );
  NAND2_X1 U5825 ( .A1(n6422), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4527) );
  NOR2_X1 U5826 ( .A1(n6493), .A2(n6492), .ZN(n6625) );
  NOR2_X1 U5827 ( .A1(n6490), .A2(n4535), .ZN(n6493) );
  AND2_X1 U5828 ( .A1(n6491), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4535) );
  NOR2_X1 U5829 ( .A1(n6625), .A2(n4534), .ZN(n6627) );
  AND2_X1 U5830 ( .A1(n6626), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4534) );
  NAND2_X1 U5831 ( .A1(n6627), .A2(n6628), .ZN(n9124) );
  NOR2_X1 U5832 ( .A1(n9514), .A2(n9513), .ZN(n9512) );
  NOR2_X1 U5833 ( .A1(n9497), .A2(n4537), .ZN(n9514) );
  AND2_X1 U5834 ( .A1(n9502), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4537) );
  NOR2_X1 U5835 ( .A1(n9559), .A2(n9558), .ZN(n9557) );
  INV_X1 U5836 ( .A(n4526), .ZN(n9581) );
  NAND2_X1 U5837 ( .A1(n5615), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U5838 ( .A1(n9596), .A2(n9595), .ZN(n9594) );
  AND2_X1 U5839 ( .A1(n4526), .A2(n4525), .ZN(n9596) );
  NAND2_X1 U5840 ( .A1(n9590), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4525) );
  OR2_X1 U5841 ( .A1(n9609), .A2(n9608), .ZN(n9618) );
  NAND2_X1 U5842 ( .A1(n9594), .A2(n9132), .ZN(n9609) );
  OR2_X1 U5843 ( .A1(n9510), .A2(n6355), .ZN(n9607) );
  INV_X1 U5844 ( .A(n9607), .ZN(n9602) );
  INV_X1 U5845 ( .A(n6274), .ZN(n6275) );
  NAND2_X1 U5846 ( .A1(n6108), .A2(n6107), .ZN(n9215) );
  NAND2_X1 U5847 ( .A1(n9250), .A2(n8066), .ZN(n9237) );
  NAND2_X1 U5848 ( .A1(n9280), .A2(n7923), .ZN(n9272) );
  NOR2_X1 U5849 ( .A1(n4721), .A2(n4720), .ZN(n9281) );
  NAND2_X1 U5850 ( .A1(n4813), .A2(n7975), .ZN(n9295) );
  NAND2_X1 U5851 ( .A1(n4501), .A2(n4500), .ZN(n4813) );
  AOI21_X1 U5852 ( .B1(n4510), .B2(n4507), .A(n6230), .ZN(n4500) );
  NOR2_X1 U5853 ( .A1(n4402), .A2(n6227), .ZN(n9324) );
  NAND2_X1 U5854 ( .A1(n7573), .A2(n8140), .ZN(n9345) );
  NAND2_X1 U5855 ( .A1(n4795), .A2(n4796), .ZN(n7244) );
  NAND2_X1 U5856 ( .A1(n6950), .A2(n6949), .ZN(n6948) );
  NAND2_X1 U5857 ( .A1(n6837), .A2(n6221), .ZN(n6950) );
  NAND2_X1 U5858 ( .A1(n6244), .A2(n6320), .ZN(n9211) );
  NAND2_X1 U5859 ( .A1(n9365), .A2(n6515), .ZN(n9368) );
  NOR2_X1 U5860 ( .A1(n6151), .A2(n6152), .ZN(n7584) );
  AND2_X1 U5861 ( .A1(n9365), .A2(n6522), .ZN(n9359) );
  INV_X1 U5862 ( .A(n9363), .ZN(n9342) );
  NAND2_X2 U5863 ( .A1(n6519), .A2(n9211), .ZN(n9365) );
  OR2_X1 U5864 ( .A1(n6327), .A2(n5703), .ZN(n5785) );
  INV_X1 U5865 ( .A(n9414), .ZN(n9384) );
  NAND2_X1 U5866 ( .A1(n4792), .A2(n5706), .ZN(n6505) );
  OAI211_X1 U5867 ( .C1(n4790), .C2(n4325), .A(n4789), .B(n5724), .ZN(n4792)
         );
  AND2_X1 U5868 ( .A1(n9659), .A2(n9430), .ZN(n9414) );
  AND2_X2 U5869 ( .A1(n6283), .A2(n6282), .ZN(n9659) );
  AOI21_X1 U5870 ( .B1(n7894), .B2(n7899), .A(n4671), .ZN(n9165) );
  INV_X1 U5871 ( .A(n7896), .ZN(n4671) );
  NAND2_X1 U5872 ( .A1(n7898), .A2(n7897), .ZN(n8216) );
  XNOR2_X1 U5873 ( .A(n8198), .B(n8197), .ZN(n8219) );
  INV_X1 U5874 ( .A(n9215), .ZN(n9446) );
  NAND2_X1 U5875 ( .A1(n6239), .A2(n6238), .ZN(n9235) );
  NAND2_X1 U5876 ( .A1(n5991), .A2(n5990), .ZN(n9470) );
  OAI21_X1 U5877 ( .B1(n4508), .B2(n4510), .A(n4507), .ZN(n9309) );
  NAND2_X1 U5878 ( .A1(n5936), .A2(n5935), .ZN(n7558) );
  INV_X1 U5879 ( .A(n4521), .ZN(n7487) );
  AND2_X1 U5880 ( .A1(n5860), .A2(n5859), .ZN(n7392) );
  INV_X1 U5881 ( .A(n6505), .ZN(n6212) );
  INV_X1 U5882 ( .A(n9471), .ZN(n9445) );
  AND2_X1 U5883 ( .A1(n6314), .A2(n6320), .ZN(n9623) );
  NAND2_X1 U5884 ( .A1(n9483), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5635) );
  INV_X1 U5885 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8222) );
  AND2_X1 U5886 ( .A1(n4889), .A2(n4395), .ZN(n4888) );
  INV_X1 U5887 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7312) );
  INV_X1 U5888 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7224) );
  INV_X1 U5889 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8190) );
  INV_X1 U5890 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7001) );
  INV_X1 U5891 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6997) );
  INV_X1 U5892 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6752) );
  AND2_X1 U5893 ( .A1(n5902), .A2(n5933), .ZN(n9562) );
  XNOR2_X1 U5894 ( .A(n5874), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9549) );
  XNOR2_X1 U5895 ( .A(n5220), .B(n5219), .ZN(n6327) );
  NAND2_X1 U5896 ( .A1(n4934), .A2(n4933), .ZN(n5220) );
  XNOR2_X1 U5897 ( .A(n5720), .B(n5719), .ZN(n6363) );
  NAND2_X1 U5898 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4533) );
  NOR2_X1 U5899 ( .A1(n7338), .A2(n10127), .ZN(n9936) );
  OAI21_X1 U5900 ( .B1(n9933), .B2(n9936), .A(n9932), .ZN(n9930) );
  AND2_X1 U5901 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7340) );
  NOR2_X1 U5902 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7341) );
  NAND2_X1 U5903 ( .A1(n4844), .A2(n9958), .ZN(n4843) );
  NAND2_X1 U5904 ( .A1(n6928), .A2(n6927), .ZN(n6930) );
  NOR2_X1 U5905 ( .A1(n7677), .A2(n4839), .ZN(n7870) );
  NAND2_X1 U5906 ( .A1(n9805), .A2(n4683), .ZN(n4681) );
  AOI211_X1 U5907 ( .C1(P2_ADDR_REG_19__SCAN_IN), .C2(n9845), .A(n8603), .B(
        n8602), .ZN(n8604) );
  NOR2_X1 U5908 ( .A1(n4896), .A2(n5589), .ZN(n5590) );
  NAND2_X1 U5909 ( .A1(n4347), .A2(n9056), .ZN(n4496) );
  AOI211_X1 U5910 ( .C1(n9458), .C2(n9035), .A(n8967), .B(n8966), .ZN(n8968)
         );
  NOR2_X1 U5911 ( .A1(n9650), .A2(n9440), .ZN(n4420) );
  AND2_X1 U5912 ( .A1(n6074), .A2(n6073), .ZN(n6268) );
  OAI211_X1 U5913 ( .C1(n5724), .C2(n6363), .A(n5723), .B(n5722), .ZN(n6215)
         );
  INV_X1 U5914 ( .A(n4333), .ZN(n6061) );
  NAND3_X1 U5915 ( .A1(n5702), .A2(n5701), .A3(n5700), .ZN(n6213) );
  AND2_X1 U5916 ( .A1(n9265), .A2(n4572), .ZN(n4334) );
  NAND2_X1 U5917 ( .A1(n5042), .A2(n4366), .ZN(n4335) );
  AND2_X1 U5918 ( .A1(n8469), .A2(n7074), .ZN(n4336) );
  AND2_X1 U5919 ( .A1(n5679), .A2(n6514), .ZN(n5695) );
  INV_X2 U5920 ( .A(n5695), .ZN(n6098) );
  NAND2_X1 U5921 ( .A1(n5773), .A2(n5772), .ZN(n7107) );
  AND2_X1 U5922 ( .A1(n6260), .A2(n8167), .ZN(n4337) );
  NAND2_X1 U5923 ( .A1(n5755), .A2(n5754), .ZN(n7112) );
  NAND2_X1 U5924 ( .A1(n4881), .A2(n4377), .ZN(n9066) );
  AND2_X1 U5925 ( .A1(n4572), .A2(n4571), .ZN(n4338) );
  OR2_X1 U5926 ( .A1(n4448), .A2(n4401), .ZN(n4339) );
  AND2_X1 U5927 ( .A1(n4705), .A2(n7948), .ZN(n4340) );
  AND2_X1 U5928 ( .A1(n4800), .A2(n4801), .ZN(n4341) );
  AND2_X1 U5929 ( .A1(n4845), .A2(n4363), .ZN(n4342) );
  AND2_X1 U5930 ( .A1(n7195), .A2(n7105), .ZN(n4343) );
  AND2_X1 U5931 ( .A1(n6780), .A2(n4839), .ZN(n4344) );
  NAND2_X1 U5932 ( .A1(n5303), .A2(n5302), .ZN(n8408) );
  AND2_X1 U5933 ( .A1(n7720), .A2(n7706), .ZN(n4345) );
  INV_X1 U5934 ( .A(n4832), .ZN(n4831) );
  NAND2_X1 U5935 ( .A1(n4833), .A2(n7231), .ZN(n4832) );
  NOR2_X1 U5936 ( .A1(n6872), .A2(n4839), .ZN(n4346) );
  XOR2_X1 U5937 ( .A(n6172), .B(n6174), .Z(n4347) );
  NOR2_X1 U5938 ( .A1(n9458), .A2(n9274), .ZN(n4348) );
  INV_X1 U5939 ( .A(n7492), .ZN(n8960) );
  NAND2_X1 U5940 ( .A1(n5904), .A2(n5903), .ZN(n7492) );
  AND2_X1 U5941 ( .A1(n4690), .A2(n4691), .ZN(n4349) );
  AND2_X1 U5942 ( .A1(n4749), .A2(n7785), .ZN(n4350) );
  INV_X1 U5943 ( .A(n5180), .ZN(n4630) );
  INV_X1 U5944 ( .A(n4485), .ZN(n7098) );
  AND2_X1 U5945 ( .A1(n4884), .A2(n5749), .ZN(n4351) );
  AND2_X1 U5946 ( .A1(n4614), .A2(n4437), .ZN(n4352) );
  NAND2_X1 U5947 ( .A1(n8950), .A2(n5917), .ZN(n8994) );
  INV_X1 U5948 ( .A(n7918), .ZN(n8070) );
  AND2_X1 U5949 ( .A1(n6148), .A2(n5658), .ZN(n6151) );
  AND2_X1 U5950 ( .A1(n4883), .A2(n6746), .ZN(n4353) );
  AND2_X1 U5951 ( .A1(n9683), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4354) );
  OR2_X1 U5952 ( .A1(n7569), .A2(n9360), .ZN(n4355) );
  AND4_X1 U5953 ( .A1(n5649), .A2(n5648), .A3(n5647), .A4(n5646), .ZN(n6542)
         );
  XOR2_X1 U5954 ( .A(n8867), .B(n8461), .Z(n4356) );
  OR2_X1 U5955 ( .A1(n7596), .A2(n9202), .ZN(n8087) );
  NOR2_X2 U5956 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5106) );
  BUF_X1 U5957 ( .A(n5106), .Z(n6590) );
  INV_X1 U5958 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9484) );
  NAND2_X1 U5959 ( .A1(n8804), .A2(n8691), .ZN(n4357) );
  OR2_X1 U5960 ( .A1(n8243), .A2(n8770), .ZN(n4358) );
  INV_X1 U5961 ( .A(n6046), .ZN(n4459) );
  XNOR2_X1 U5962 ( .A(n4478), .B(n5930), .ZN(n5691) );
  NAND2_X1 U5963 ( .A1(n9197), .A2(n4580), .ZN(n4359) );
  AND2_X1 U5964 ( .A1(n5503), .A2(n4836), .ZN(n4360) );
  AND4_X1 U5965 ( .A1(n5717), .A2(n5716), .A3(n5715), .A4(n5714), .ZN(n6216)
         );
  OR2_X1 U5966 ( .A1(n8804), .A2(n8691), .ZN(n4361) );
  AND2_X1 U5967 ( .A1(n5571), .A2(n4346), .ZN(n4362) );
  OR2_X1 U5968 ( .A1(n4731), .A2(n4730), .ZN(n6210) );
  OR2_X1 U5969 ( .A1(n8327), .A2(n4849), .ZN(n4363) );
  AND2_X1 U5970 ( .A1(n4885), .A2(n6889), .ZN(n4364) );
  AND4_X1 U5971 ( .A1(n7818), .A2(n7817), .A3(n7816), .A4(n7815), .ZN(n4365)
         );
  NAND2_X1 U5972 ( .A1(n6216), .A2(n6215), .ZN(n8118) );
  INV_X1 U5973 ( .A(n8118), .ZN(n4715) );
  AND2_X1 U5974 ( .A1(n5562), .A2(n5044), .ZN(n4366) );
  NAND2_X1 U5975 ( .A1(n6037), .A2(n6036), .ZN(n9398) );
  OR2_X1 U5976 ( .A1(n8877), .A2(n8636), .ZN(n7824) );
  AND2_X1 U5977 ( .A1(n7404), .A2(n8466), .ZN(n4367) );
  OR2_X1 U5978 ( .A1(n9408), .A2(n9093), .ZN(n4368) );
  AND2_X1 U5979 ( .A1(n4452), .A2(n4450), .ZN(n4369) );
  AND2_X1 U5980 ( .A1(n7685), .A2(n7683), .ZN(n4370) );
  AND2_X1 U5981 ( .A1(n4625), .A2(n5207), .ZN(n4371) );
  OAI21_X1 U5982 ( .B1(n8689), .B2(n4597), .A(n4357), .ZN(n4596) );
  OR2_X1 U5983 ( .A1(n8867), .A2(n8635), .ZN(n4372) );
  AND2_X1 U5984 ( .A1(n4471), .A2(n8964), .ZN(n4373) );
  INV_X1 U5985 ( .A(n7484), .ZN(n9047) );
  NAND2_X1 U5986 ( .A1(n5824), .A2(n5823), .ZN(n7484) );
  INV_X1 U5987 ( .A(n7115), .ZN(n9104) );
  AND4_X1 U5988 ( .A1(n5780), .A2(n5779), .A3(n5778), .A4(n5777), .ZN(n7115)
         );
  INV_X1 U5989 ( .A(n6892), .ZN(n9105) );
  AND4_X1 U5990 ( .A1(n5762), .A2(n5761), .A3(n5760), .A4(n5759), .ZN(n6892)
         );
  INV_X1 U5991 ( .A(n6243), .ZN(n4808) );
  NAND2_X1 U5992 ( .A1(n9265), .A2(n4574), .ZN(n4575) );
  AND2_X1 U5993 ( .A1(n8141), .A2(n8140), .ZN(n7575) );
  INV_X1 U5994 ( .A(n7575), .ZN(n4727) );
  AND2_X1 U5995 ( .A1(n8961), .A2(n8962), .ZN(n4374) );
  INV_X1 U5996 ( .A(n9169), .ZN(n7902) );
  NAND2_X1 U5997 ( .A1(n7901), .A2(n7900), .ZN(n9169) );
  NAND2_X1 U5998 ( .A1(n7042), .A2(n7700), .ZN(n4375) );
  NAND2_X1 U5999 ( .A1(n7118), .A2(n7117), .ZN(n4376) );
  INV_X1 U6000 ( .A(n4583), .ZN(n9190) );
  NOR2_X1 U6001 ( .A1(n9191), .A2(n9373), .ZN(n4583) );
  AND2_X1 U6002 ( .A1(n6117), .A2(n6106), .ZN(n4377) );
  AND2_X1 U6003 ( .A1(n7820), .A2(n7819), .ZN(n4378) );
  AND2_X1 U6004 ( .A1(n4695), .A2(n4694), .ZN(n4379) );
  AND2_X1 U6005 ( .A1(n8088), .A2(n8085), .ZN(n4380) );
  AND2_X1 U6006 ( .A1(n5386), .A2(n5387), .ZN(n4381) );
  AND2_X1 U6007 ( .A1(n6448), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4382) );
  INV_X1 U6008 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5038) );
  OR2_X1 U6009 ( .A1(n8934), .A2(n8353), .ZN(n7779) );
  INV_X1 U6010 ( .A(n7779), .ZN(n4778) );
  INV_X1 U6011 ( .A(n4791), .ZN(n4790) );
  NAND2_X1 U6012 ( .A1(n4907), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4791) );
  OR2_X1 U6013 ( .A1(n6241), .A2(n4400), .ZN(n4383) );
  INV_X1 U6014 ( .A(n4801), .ZN(n4799) );
  NAND2_X1 U6015 ( .A1(n9646), .A2(n9046), .ZN(n4801) );
  INV_X1 U6016 ( .A(n7944), .ZN(n7981) );
  INV_X1 U6017 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5622) );
  AND2_X1 U6018 ( .A1(n4554), .A2(n8095), .ZN(n4384) );
  OR2_X1 U6019 ( .A1(n5615), .A2(n5604), .ZN(n4385) );
  INV_X1 U6020 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5044) );
  NOR2_X1 U6021 ( .A1(n9011), .A2(n5969), .ZN(n4386) );
  INV_X1 U6022 ( .A(n6262), .ZN(n7995) );
  AND2_X1 U6023 ( .A1(n5890), .A2(n5889), .ZN(n4387) );
  OR2_X1 U6024 ( .A1(n4772), .A2(n7822), .ZN(n4388) );
  NAND2_X1 U6025 ( .A1(n5486), .A2(n5544), .ZN(n4389) );
  NOR2_X1 U6026 ( .A1(n5267), .A2(SI_11_), .ZN(n4390) );
  AND2_X1 U6027 ( .A1(n7722), .A2(n7086), .ZN(n7720) );
  NAND2_X1 U6028 ( .A1(n4460), .A2(SI_3_), .ZN(n4919) );
  AND4_X1 U6029 ( .A1(n5281), .A2(n5280), .A3(n5279), .A4(n5278), .ZN(n7408)
         );
  INV_X1 U6030 ( .A(n7408), .ZN(n4441) );
  NOR2_X1 U6031 ( .A1(n9008), .A2(n9011), .ZN(n4391) );
  AND2_X1 U6032 ( .A1(n8012), .A2(n7996), .ZN(n4392) );
  INV_X1 U6033 ( .A(n7596), .ZN(n8192) );
  NAND2_X1 U6034 ( .A1(n6123), .A2(n6122), .ZN(n7596) );
  OR2_X1 U6035 ( .A1(n4865), .A2(n4867), .ZN(n4393) );
  AND2_X1 U6036 ( .A1(n8877), .A2(n8636), .ZN(n7822) );
  NAND2_X1 U6037 ( .A1(n8286), .A2(n8464), .ZN(n4394) );
  AND2_X1 U6038 ( .A1(n5656), .A2(n6149), .ZN(n4395) );
  NAND3_X1 U6039 ( .A1(n7837), .A2(n7846), .A3(n7836), .ZN(n4396) );
  NOR2_X1 U6040 ( .A1(n4627), .A2(n5194), .ZN(n4626) );
  AND2_X1 U6041 ( .A1(n5636), .A2(n5632), .ZN(n4397) );
  INV_X1 U6042 ( .A(n4765), .ZN(n4764) );
  OAI21_X1 U6043 ( .B1(n7710), .B2(n4758), .A(n7700), .ZN(n4765) );
  AND2_X1 U6044 ( .A1(n7783), .A2(n7790), .ZN(n8727) );
  AND2_X1 U6045 ( .A1(n4773), .A2(n4372), .ZN(n4398) );
  INV_X1 U6046 ( .A(n4810), .ZN(n5615) );
  AND4_X2 U6047 ( .A1(n5599), .A2(n5899), .A3(n5898), .A4(n5598), .ZN(n4810)
         );
  INV_X1 U6048 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U6049 ( .A1(n6590), .A2(n5038), .ZN(n5141) );
  INV_X1 U6050 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5617) );
  INV_X1 U6051 ( .A(n4907), .ZN(n4616) );
  INV_X1 U6052 ( .A(n5687), .ZN(n6167) );
  NAND2_X1 U6053 ( .A1(n5651), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4492) );
  NAND2_X1 U6054 ( .A1(n6089), .A2(n6088), .ZN(n9449) );
  INV_X1 U6055 ( .A(n9449), .ZN(n4571) );
  AND2_X1 U6056 ( .A1(n8391), .A2(n8264), .ZN(n4399) );
  NAND2_X1 U6057 ( .A1(n6156), .A2(n6155), .ZN(n9373) );
  INV_X1 U6058 ( .A(n9373), .ZN(n4585) );
  INV_X1 U6059 ( .A(n8140), .ZN(n4729) );
  NAND2_X1 U6060 ( .A1(n4739), .A2(n7800), .ZN(n8687) );
  INV_X1 U6061 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4836) );
  INV_X1 U6062 ( .A(n8332), .ZN(n4819) );
  INV_X1 U6063 ( .A(n8465), .ZN(n8238) );
  AND2_X1 U6064 ( .A1(n6268), .A2(n9251), .ZN(n4400) );
  NAND2_X1 U6065 ( .A1(n5614), .A2(n5613), .ZN(n6520) );
  NOR2_X1 U6066 ( .A1(n6050), .A2(n6052), .ZN(n4401) );
  AND2_X1 U6067 ( .A1(n9344), .A2(n6228), .ZN(n4402) );
  AND4_X1 U6068 ( .A1(n5793), .A2(n5792), .A3(n5791), .A4(n5790), .ZN(n7105)
         );
  INV_X1 U6069 ( .A(n8962), .ZN(n4471) );
  AND2_X1 U6070 ( .A1(n4798), .A2(n4797), .ZN(n4403) );
  INV_X1 U6071 ( .A(n6230), .ZN(n4811) );
  AND2_X1 U6072 ( .A1(n4659), .A2(n4662), .ZN(n4404) );
  INV_X1 U6073 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4716) );
  XNOR2_X1 U6074 ( .A(n5512), .B(P2_IR_REG_20__SCAN_IN), .ZN(n6779) );
  INV_X1 U6075 ( .A(n6779), .ZN(n4839) );
  INV_X1 U6076 ( .A(n6784), .ZN(n7232) );
  NAND2_X1 U6077 ( .A1(n5550), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U6078 ( .A1(n4624), .A2(n4371), .ZN(n7033) );
  INV_X1 U6079 ( .A(n8566), .ZN(n8576) );
  NAND2_X1 U6080 ( .A1(n5920), .A2(n5919), .ZN(n9429) );
  INV_X1 U6081 ( .A(n9429), .ZN(n4587) );
  AND4_X1 U6082 ( .A1(n5910), .A2(n5909), .A3(n5908), .A4(n5907), .ZN(n9079)
         );
  INV_X1 U6083 ( .A(n4518), .ZN(n7144) );
  NAND2_X1 U6084 ( .A1(n7145), .A2(n7951), .ZN(n4518) );
  INV_X1 U6085 ( .A(n4570), .ZN(n6685) );
  NOR2_X1 U6086 ( .A1(n6537), .A2(n6520), .ZN(n4570) );
  NAND2_X1 U6087 ( .A1(n8495), .A2(n8527), .ZN(n4691) );
  NAND2_X1 U6088 ( .A1(n5359), .A2(n5562), .ZN(n4405) );
  AND2_X1 U6089 ( .A1(n5490), .A2(n5489), .ZN(n4406) );
  INV_X1 U6090 ( .A(n4576), .ZN(n7435) );
  NOR2_X1 U6091 ( .A1(n7146), .A2(n4578), .ZN(n4576) );
  AND2_X1 U6092 ( .A1(n4886), .A2(n4885), .ZN(n4407) );
  INV_X1 U6093 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n4678) );
  AND2_X1 U6094 ( .A1(n4701), .A2(n4703), .ZN(n4408) );
  INV_X1 U6095 ( .A(n8167), .ZN(n8085) );
  OR2_X1 U6096 ( .A1(n8586), .A2(n8557), .ZN(n4409) );
  OR2_X1 U6097 ( .A1(n5783), .A2(n5782), .ZN(n4410) );
  INV_X1 U6098 ( .A(n6907), .ZN(n4677) );
  INV_X1 U6099 ( .A(n5749), .ZN(n4885) );
  AND2_X1 U6100 ( .A1(n6185), .A2(n6154), .ZN(n9056) );
  NAND2_X1 U6101 ( .A1(n4684), .A2(n4682), .ZN(n4411) );
  INV_X1 U6102 ( .A(n5769), .ZN(n4487) );
  AND2_X1 U6103 ( .A1(n9805), .A2(n4411), .ZN(n4412) );
  NAND2_X1 U6104 ( .A1(n5108), .A2(n5107), .ZN(n6695) );
  INV_X1 U6105 ( .A(n6695), .ZN(n4623) );
  INV_X1 U6106 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4619) );
  OAI21_X1 U6107 ( .B1(n9524), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9529), .ZN(
        n9543) );
  NAND2_X1 U6108 ( .A1(n9555), .A2(n9554), .ZN(n9553) );
  AOI21_X1 U6109 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n9502), .A(n9494), .ZN(
        n9517) );
  AOI21_X1 U6110 ( .B1(n9520), .B2(P1_REG1_REG_11__SCAN_IN), .A(n9515), .ZN(
        n9530) );
  AOI21_X1 U6111 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6626), .A(n6618), .ZN(
        n6619) );
  AOI21_X1 U6112 ( .B1(n6387), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6393), .ZN(
        n6410) );
  AOI21_X1 U6113 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n6366), .A(n6408), .ZN(
        n6369) );
  AOI21_X1 U6114 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n6379), .A(n6378), .ZN(
        n6381) );
  AOI21_X1 U6115 ( .B1(n6422), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6421), .ZN(
        n6425) );
  NOR2_X1 U6116 ( .A1(n9568), .A2(n9148), .ZN(n9588) );
  NAND3_X1 U6117 ( .A1(n4632), .A2(n5156), .A3(n4417), .ZN(n4416) );
  NAND2_X1 U6118 ( .A1(n4422), .A2(n4419), .ZN(P1_U3518) );
  OR2_X1 U6119 ( .A1(n9439), .A2(n6284), .ZN(n4422) );
  NAND2_X1 U6120 ( .A1(n6264), .A2(n6261), .ZN(n8001) );
  NAND2_X1 U6121 ( .A1(n9310), .A2(n8150), .ZN(n9297) );
  OAI21_X2 U6122 ( .B1(n7489), .B2(n7488), .A(n8139), .ZN(n7545) );
  AOI21_X2 U6123 ( .B1(n7246), .B2(n7245), .A(n4423), .ZN(n7431) );
  NAND2_X1 U6124 ( .A1(n4724), .A2(n4723), .ZN(n9334) );
  NAND2_X1 U6125 ( .A1(n4905), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4431) );
  NAND3_X1 U6126 ( .A1(n4701), .A2(n4703), .A3(n7141), .ZN(n7464) );
  OAI21_X1 U6127 ( .B1(n7789), .B2(n7788), .A(n7787), .ZN(n7791) );
  NAND2_X1 U6128 ( .A1(n4424), .A2(n7697), .ZN(n7713) );
  MUX2_X2 U6129 ( .A(n7719), .B(n7718), .S(n7826), .Z(n7721) );
  OR2_X2 U6130 ( .A1(n7765), .A2(n7764), .ZN(n7767) );
  INV_X1 U6131 ( .A(n8475), .ZN(n6859) );
  MUX2_X2 U6132 ( .A(n7793), .B(n7792), .S(n7826), .Z(n7799) );
  OAI21_X2 U6133 ( .B1(n7799), .B2(n7798), .A(n7797), .ZN(n7803) );
  OAI21_X1 U6134 ( .B1(n4396), .B2(n4425), .A(n7843), .ZN(n7854) );
  OAI21_X2 U6135 ( .B1(n7776), .B2(n7775), .A(n8755), .ZN(n7780) );
  NAND2_X1 U6136 ( .A1(n4608), .A2(n4607), .ZN(n4438) );
  NAND2_X1 U6137 ( .A1(n7752), .A2(n7742), .ZN(n7261) );
  OAI21_X2 U6138 ( .B1(n8633), .B2(n4443), .A(n4389), .ZN(n4592) );
  NAND2_X1 U6139 ( .A1(n5191), .A2(n5190), .ZN(n4444) );
  NAND2_X1 U6140 ( .A1(n5176), .A2(n5175), .ZN(n4445) );
  AND2_X1 U6141 ( .A1(n6048), .A2(n9030), .ZN(n4865) );
  INV_X1 U6142 ( .A(n9030), .ZN(n4448) );
  AND2_X1 U6143 ( .A1(n9066), .A2(n6121), .ZN(n6204) );
  INV_X1 U6144 ( .A(n6203), .ZN(n6199) );
  MUX2_X1 U6145 ( .A(n6313), .B(n6300), .S(n4907), .Z(n4918) );
  NAND2_X1 U6146 ( .A1(n4462), .A2(n8970), .ZN(n6009) );
  XNOR2_X1 U6147 ( .A(n4462), .B(n4461), .ZN(n8975) );
  INV_X1 U6148 ( .A(n8970), .ZN(n4461) );
  NAND2_X1 U6149 ( .A1(n7873), .A2(n5694), .ZN(n6469) );
  NAND2_X1 U6150 ( .A1(n4470), .A2(n8964), .ZN(n4469) );
  NAND2_X2 U6151 ( .A1(n4473), .A2(n4472), .ZN(n9039) );
  NAND2_X2 U6152 ( .A1(n4477), .A2(n4476), .ZN(n4475) );
  NAND2_X2 U6153 ( .A1(n5673), .A2(n5687), .ZN(n5727) );
  NAND2_X1 U6154 ( .A1(n4489), .A2(n4882), .ZN(n7116) );
  XNOR2_X1 U6155 ( .A(n5986), .B(n5984), .ZN(n9053) );
  AOI21_X2 U6156 ( .B1(n8950), .B2(n4491), .A(n4386), .ZN(n5986) );
  NAND2_X1 U6157 ( .A1(n4492), .A2(n5652), .ZN(n5653) );
  NAND2_X1 U6158 ( .A1(n4492), .A2(n5970), .ZN(n5971) );
  XNOR2_X1 U6159 ( .A(n4492), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9600) );
  NAND2_X1 U6160 ( .A1(n6204), .A2(n4494), .ZN(n4493) );
  OAI211_X1 U6161 ( .C1(n6204), .C2(n4496), .A(n4493), .B(n4900), .ZN(P1_U3214) );
  NAND3_X1 U6162 ( .A1(n6839), .A2(n6838), .A3(n6949), .ZN(n4498) );
  INV_X1 U6163 ( .A(n9344), .ZN(n4508) );
  OAI21_X1 U6164 ( .B1(n4508), .B2(n4505), .A(n4502), .ZN(n6232) );
  NAND3_X1 U6165 ( .A1(n5601), .A2(n5600), .A3(n5602), .ZN(n4517) );
  NAND2_X1 U6166 ( .A1(n4515), .A2(n4810), .ZN(n9483) );
  NAND2_X1 U6167 ( .A1(n9246), .A2(n4806), .ZN(n4524) );
  INV_X2 U6168 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U6169 ( .A1(n4540), .A2(n6255), .ZN(n8117) );
  NOR2_X1 U6170 ( .A1(n9110), .A2(n7592), .ZN(n6977) );
  AOI21_X1 U6171 ( .B1(n4542), .B2(n4337), .A(n6262), .ZN(n4541) );
  INV_X1 U6172 ( .A(n8095), .ZN(n4555) );
  NAND2_X1 U6173 ( .A1(n8099), .A2(n8100), .ZN(n4556) );
  OR2_X1 U6174 ( .A1(n8084), .A2(n4557), .ZN(n4558) );
  OR2_X1 U6175 ( .A1(n8077), .A2(n4560), .ZN(n4559) );
  OAI211_X1 U6176 ( .C1(n4561), .C2(n4563), .A(n4559), .B(n4558), .ZN(n8091)
         );
  INV_X1 U6177 ( .A(n4575), .ZN(n9255) );
  NAND2_X1 U6178 ( .A1(n9197), .A2(n8192), .ZN(n9191) );
  NAND2_X1 U6179 ( .A1(n9197), .A2(n4581), .ZN(n9171) );
  NOR2_X2 U6180 ( .A1(n4355), .A2(n9417), .ZN(n9325) );
  XNOR2_X1 U6181 ( .A(n4590), .B(n7643), .ZN(n5527) );
  OAI22_X1 U6182 ( .A1(n4592), .A2(n4591), .B1(n5545), .B2(n8635), .ZN(n4590)
         );
  INV_X1 U6183 ( .A(n8690), .ZN(n4593) );
  AOI21_X1 U6184 ( .B1(n4593), .B2(n4594), .A(n4596), .ZN(n8667) );
  NAND2_X1 U6185 ( .A1(n6810), .A2(n4626), .ZN(n4624) );
  AND2_X2 U6186 ( .A1(n5560), .A2(n5037), .ZN(n5042) );
  NAND2_X1 U6187 ( .A1(n4631), .A2(n5450), .ZN(n5007) );
  XNOR2_X1 U6188 ( .A(n4631), .B(n5450), .ZN(n7911) );
  NAND2_X1 U6189 ( .A1(n5002), .A2(n5001), .ZN(n4631) );
  NAND3_X1 U6190 ( .A1(n4919), .A2(n4916), .A3(n4917), .ZN(n4632) );
  NAND2_X1 U6191 ( .A1(n4917), .A2(n4916), .ZN(n5145) );
  NAND2_X1 U6192 ( .A1(n4633), .A2(n4919), .ZN(n5157) );
  NAND2_X1 U6193 ( .A1(n5145), .A2(n5144), .ZN(n4633) );
  NAND2_X1 U6194 ( .A1(n5023), .A2(n5022), .ZN(n5488) );
  NAND2_X1 U6195 ( .A1(n5462), .A2(n4647), .ZN(n4643) );
  NAND2_X1 U6196 ( .A1(n4643), .A2(n4644), .ZN(n5087) );
  NAND2_X1 U6197 ( .A1(n5462), .A2(n5463), .ZN(n4646) );
  NAND2_X1 U6198 ( .A1(n5330), .A2(n4654), .ZN(n4653) );
  NAND2_X1 U6199 ( .A1(n7894), .A2(n4673), .ZN(n4670) );
  NAND2_X1 U6200 ( .A1(n4670), .A2(n4672), .ZN(n7937) );
  NAND2_X1 U6201 ( .A1(n8164), .A2(n8163), .ZN(n8173) );
  OAI22_X1 U6202 ( .A1(n8645), .A2(n5485), .B1(n8636), .B2(n8445), .ZN(n8633)
         );
  OAI22_X1 U6203 ( .A1(n8654), .A2(n8653), .B1(n8668), .B2(n8883), .ZN(n8645)
         );
  NAND2_X1 U6204 ( .A1(n8171), .A2(n8170), .ZN(n8172) );
  AND3_X2 U6205 ( .A1(n5141), .A2(n4675), .A3(n4674), .ZN(n8483) );
  OAI21_X2 U6206 ( .B1(n6670), .B2(n4679), .A(n4676), .ZN(n8492) );
  NAND2_X1 U6207 ( .A1(n8561), .A2(n4412), .ZN(n4680) );
  OAI211_X1 U6208 ( .C1(n8561), .C2(n4681), .A(n4680), .B(n8604), .ZN(P2_U3201) );
  NOR2_X1 U6209 ( .A1(n8561), .A2(n8562), .ZN(n8584) );
  OAI21_X1 U6210 ( .B1(n9839), .B2(n4693), .A(n4692), .ZN(n9858) );
  INV_X1 U6211 ( .A(n6833), .ZN(n4702) );
  NAND2_X1 U6212 ( .A1(n9248), .A2(n9247), .ZN(n9250) );
  INV_X1 U6213 ( .A(n4706), .ZN(n9221) );
  NOR2_X1 U6214 ( .A1(n4709), .A2(n7918), .ZN(n4708) );
  OAI21_X2 U6215 ( .B1(n8204), .B2(n9299), .A(n8203), .ZN(n4711) );
  NOR2_X1 U6216 ( .A1(n4711), .A2(n8208), .ZN(n8214) );
  OAI21_X1 U6217 ( .B1(n4711), .B2(n8211), .A(n9365), .ZN(n8212) );
  NAND2_X1 U6218 ( .A1(n4712), .A2(n6259), .ZN(n6517) );
  OAI21_X1 U6219 ( .B1(n6551), .B2(n7944), .A(n4713), .ZN(n4712) );
  AOI21_X1 U6220 ( .B1(n7981), .B2(n4715), .A(n4714), .ZN(n4713) );
  INV_X1 U6221 ( .A(n6254), .ZN(n7943) );
  OAI21_X1 U6222 ( .B1(n6254), .B2(n6975), .A(n6974), .ZN(n7884) );
  OAI21_X1 U6223 ( .B1(n4722), .B2(n4719), .A(n9271), .ZN(n4717) );
  OAI21_X2 U6224 ( .B1(n6267), .B2(n4719), .A(n4718), .ZN(n9270) );
  NAND2_X1 U6225 ( .A1(n7574), .A2(n4725), .ZN(n4724) );
  NAND2_X2 U6226 ( .A1(n4327), .A2(n4907), .ZN(n5721) );
  NAND2_X2 U6227 ( .A1(n4326), .A2(n4325), .ZN(n5703) );
  NAND2_X2 U6228 ( .A1(n6354), .A2(n4323), .ZN(n5724) );
  OR2_X1 U6229 ( .A1(n8708), .A2(n4736), .ZN(n4732) );
  NAND2_X1 U6230 ( .A1(n4732), .A2(n4733), .ZN(n8675) );
  NAND2_X1 U6231 ( .A1(n7030), .A2(n7724), .ZN(n5532) );
  NAND2_X1 U6232 ( .A1(n5531), .A2(n4345), .ZN(n7030) );
  NAND2_X1 U6233 ( .A1(n5540), .A2(n4743), .ZN(n4742) );
  NAND2_X1 U6234 ( .A1(n5534), .A2(n4753), .ZN(n4752) );
  NAND2_X1 U6235 ( .A1(n6848), .A2(n4756), .ZN(n4760) );
  NAND2_X1 U6236 ( .A1(n4757), .A2(n4765), .ZN(n4756) );
  INV_X1 U6237 ( .A(n4761), .ZN(n4757) );
  INV_X1 U6238 ( .A(n7702), .ZN(n4758) );
  NAND2_X1 U6239 ( .A1(n6848), .A2(n7710), .ZN(n4767) );
  NAND2_X1 U6240 ( .A1(n4767), .A2(n7702), .ZN(n6809) );
  NAND2_X1 U6241 ( .A1(n5042), .A2(n4786), .ZN(n5077) );
  INV_X1 U6242 ( .A(n5077), .ZN(n5074) );
  NAND3_X1 U6243 ( .A1(n7942), .A2(n7943), .A3(n4788), .ZN(n7947) );
  NAND2_X1 U6244 ( .A1(n6239), .A2(n4804), .ZN(n4802) );
  NAND2_X1 U6245 ( .A1(n4802), .A2(n4803), .ZN(n8194) );
  NAND3_X1 U6246 ( .A1(n4809), .A2(n4810), .A3(n5631), .ZN(n5605) );
  NAND2_X1 U6247 ( .A1(n8422), .A2(n4818), .ZN(n4817) );
  OAI21_X1 U6248 ( .B1(n8400), .B2(n4826), .A(n4823), .ZN(n8448) );
  OAI21_X1 U6249 ( .B1(n7228), .B2(n4832), .A(n4829), .ZN(n8306) );
  NAND2_X1 U6250 ( .A1(n5510), .A2(n4835), .ZN(n5550) );
  NAND2_X1 U6251 ( .A1(n6431), .A2(n4362), .ZN(n4838) );
  NAND2_X1 U6252 ( .A1(n8436), .A2(n4842), .ZN(n4841) );
  OAI211_X1 U6253 ( .C1(n8436), .C2(n4843), .A(n4841), .B(n8331), .ZN(P2_U3160) );
  NAND2_X1 U6254 ( .A1(n8436), .A2(n4855), .ZN(n8326) );
  NAND2_X1 U6255 ( .A1(n4859), .A2(n7043), .ZN(n4857) );
  AND2_X1 U6256 ( .A1(n4860), .A2(n7043), .ZN(n4858) );
  NOR2_X1 U6257 ( .A1(n6931), .A2(n4861), .ZN(n4860) );
  NAND2_X1 U6258 ( .A1(n8976), .A2(n4393), .ZN(n4864) );
  OAI21_X2 U6259 ( .B1(n4872), .B2(n4871), .A(n4870), .ZN(n5914) );
  NAND2_X1 U6260 ( .A1(n4883), .A2(n6745), .ZN(n4882) );
  NAND2_X1 U6261 ( .A1(n5626), .A2(n4889), .ZN(n5655) );
  NAND2_X1 U6262 ( .A1(n4887), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U6263 ( .A1(n5626), .A2(n4888), .ZN(n4887) );
  NAND2_X1 U6264 ( .A1(n5626), .A2(n5618), .ZN(n5630) );
  NOR2_X1 U6265 ( .A1(n8499), .A2(n9807), .ZN(n9824) );
  NAND4_X2 U6266 ( .A1(n5113), .A2(n5112), .A3(n5111), .A4(n5110), .ZN(n8475)
         );
  AOI21_X2 U6267 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8521), .A(n9822), .ZN(
        n8501) );
  NAND2_X1 U6268 ( .A1(n5433), .A2(n4995), .ZN(n5443) );
  NAND2_X1 U6269 ( .A1(n9439), .A2(n9659), .ZN(n9377) );
  INV_X1 U6270 ( .A(n8754), .ZN(n5540) );
  NAND2_X1 U6271 ( .A1(n6199), .A2(n4898), .ZN(n6200) );
  INV_X1 U6272 ( .A(n5109), .ZN(n5495) );
  NAND2_X1 U6273 ( .A1(n5584), .A2(n5585), .ZN(n5551) );
  NAND2_X1 U6274 ( .A1(n7414), .A2(n7413), .ZN(n8235) );
  XNOR2_X1 U6275 ( .A(n5620), .B(n5621), .ZN(n7538) );
  NAND2_X1 U6276 ( .A1(n5507), .A2(n5550), .ZN(n7309) );
  NOR2_X1 U6277 ( .A1(n7642), .A2(n7641), .ZN(n7670) );
  INV_X2 U6278 ( .A(n5721), .ZN(n5989) );
  XNOR2_X1 U6279 ( .A(n5745), .B(n5744), .ZN(n6746) );
  OR2_X1 U6280 ( .A1(n6431), .A2(n5583), .ZN(n6754) );
  NAND2_X1 U6281 ( .A1(n5914), .A2(n5916), .ZN(n5917) );
  NAND2_X2 U6282 ( .A1(n6009), .A2(n6008), .ZN(n8976) );
  OR3_X1 U6283 ( .A1(n7535), .A2(n7913), .A3(n7541), .ZN(n6757) );
  INV_X1 U6284 ( .A(n7161), .ZN(n7159) );
  NAND3_X2 U6285 ( .A1(n5679), .A2(n5664), .A3(n6249), .ZN(n5687) );
  OR2_X1 U6286 ( .A1(n6778), .A2(n6753), .ZN(n6820) );
  OAI22_X2 U6287 ( .A1(n6480), .A2(n6479), .B1(n5731), .B2(n5730), .ZN(n6745)
         );
  AND3_X2 U6288 ( .A1(n6817), .A2(n5587), .A3(n6759), .ZN(n8827) );
  INV_X2 U6289 ( .A(n9876), .ZN(n8693) );
  AND2_X1 U6290 ( .A1(n9446), .A2(n9225), .ZN(n4890) );
  AND2_X1 U6291 ( .A1(n5100), .A2(n5099), .ZN(n4891) );
  AND2_X1 U6292 ( .A1(n5747), .A2(n5746), .ZN(n4892) );
  OR2_X1 U6293 ( .A1(n9081), .A2(n9001), .ZN(n4893) );
  OR2_X1 U6294 ( .A1(n9446), .A2(n9225), .ZN(n4894) );
  NAND3_X1 U6295 ( .A1(n5617), .A2(n5970), .A3(n5650), .ZN(n4895) );
  NAND2_X1 U6296 ( .A1(n8693), .A2(n7068), .ZN(n8765) );
  AND2_X1 U6297 ( .A1(n8619), .A2(n8829), .ZN(n4896) );
  OR2_X1 U6298 ( .A1(n9659), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n4897) );
  AND2_X1 U6299 ( .A1(n6198), .A2(n9056), .ZN(n4898) );
  NAND2_X1 U6300 ( .A1(n7616), .A2(n7615), .ZN(n7631) );
  INV_X1 U6301 ( .A(n5699), .ZN(n5941) );
  INV_X1 U6302 ( .A(n9236), .ZN(n6270) );
  AND2_X1 U6303 ( .A1(n6283), .A2(n6513), .ZN(n9480) );
  OAI21_X1 U6304 ( .B1(n5255), .B2(n4965), .A(n4964), .ZN(n5312) );
  OAI21_X1 U6305 ( .B1(n5703), .B2(n6307), .A(n5742), .ZN(n6741) );
  AND2_X1 U6306 ( .A1(n6209), .A2(n6208), .ZN(n4900) );
  NAND2_X1 U6307 ( .A1(n8610), .A2(n8861), .ZN(n7639) );
  INV_X1 U6308 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5036) );
  INV_X1 U6309 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U6310 ( .A1(n7844), .A2(n7639), .ZN(n7640) );
  OR4_X1 U6311 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n5579) );
  MUX2_X1 U6312 ( .A(n8094), .B(n8093), .S(n8167), .Z(n8095) );
  OR2_X1 U6313 ( .A1(n7858), .A2(n7640), .ZN(n7641) );
  INV_X1 U6314 ( .A(n7720), .ZN(n5207) );
  INV_X1 U6315 ( .A(n5417), .ZN(n4988) );
  INV_X1 U6316 ( .A(SI_13_), .ZN(n4958) );
  INV_X1 U6317 ( .A(n8610), .ZN(n7672) );
  INV_X1 U6318 ( .A(n5394), .ZN(n5062) );
  INV_X1 U6319 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5059) );
  INV_X1 U6320 ( .A(n6754), .ZN(n6758) );
  NOR2_X1 U6321 ( .A1(n5976), .A2(n5975), .ZN(n5992) );
  AOI22_X1 U6322 ( .A1(n9089), .A2(n9337), .B1(n9335), .B2(n9090), .ZN(n6274)
         );
  INV_X1 U6323 ( .A(n9398), .ZN(n6278) );
  INV_X1 U6324 ( .A(SI_23_), .ZN(n4997) );
  INV_X1 U6325 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n4948) );
  INV_X1 U6326 ( .A(n7162), .ZN(n7158) );
  NAND2_X1 U6327 ( .A1(n7673), .A2(n7672), .ZN(n7674) );
  NOR2_X1 U6328 ( .A1(n8840), .A2(n8635), .ZN(n5525) );
  INV_X1 U6329 ( .A(n5453), .ZN(n5066) );
  NAND2_X1 U6330 ( .A1(n5058), .A2(n5057), .ZN(n5351) );
  INV_X1 U6331 ( .A(n8646), .ZN(n5544) );
  INV_X1 U6332 ( .A(n8758), .ZN(n8365) );
  OR2_X1 U6333 ( .A1(n6431), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U6334 ( .A1(n5560), .A2(n5562), .ZN(n5500) );
  AND2_X1 U6335 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5642) );
  INV_X1 U6336 ( .A(n5746), .ZN(n5744) );
  NAND2_X2 U6337 ( .A1(n5659), .A2(n5679), .ZN(n5673) );
  AND2_X1 U6338 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n6092), .ZN(n6109) );
  NOR2_X1 U6339 ( .A1(n6039), .A2(n6038), .ZN(n6056) );
  AND2_X1 U6340 ( .A1(n8210), .A2(n6160), .ZN(n9192) );
  AND2_X1 U6341 ( .A1(n6093), .A2(n6110), .ZN(n9229) );
  OR2_X1 U6342 ( .A1(n6314), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6137) );
  INV_X1 U6343 ( .A(n6215), .ZN(n6562) );
  INV_X1 U6344 ( .A(SI_20_), .ZN(n5401) );
  OAI21_X1 U6345 ( .B1(n5312), .B2(SI_14_), .A(n5313), .ZN(n4966) );
  OR2_X1 U6346 ( .A1(n5770), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U6347 ( .A1(n4986), .A2(n6311), .ZN(n4913) );
  NAND2_X1 U6348 ( .A1(n7159), .A2(n7158), .ZN(n7212) );
  NAND2_X1 U6349 ( .A1(n8412), .A2(n8270), .ZN(n8297) );
  INV_X1 U6350 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5048) );
  OR2_X1 U6351 ( .A1(n5407), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5423) );
  INV_X1 U6352 ( .A(n7626), .ZN(n5166) );
  INV_X1 U6353 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5072) );
  INV_X1 U6354 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7417) );
  OR2_X1 U6355 ( .A1(n5092), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U6356 ( .A1(n5068), .A2(n5067), .ZN(n5477) );
  INV_X1 U6357 ( .A(n7653), .ZN(n5533) );
  AND2_X1 U6358 ( .A1(n8614), .A2(n7371), .ZN(n5549) );
  OR2_X1 U6359 ( .A1(n8921), .A2(n8365), .ZN(n8724) );
  AND2_X1 U6360 ( .A1(n7826), .A2(n5522), .ZN(n8771) );
  INV_X1 U6361 ( .A(n9944), .ZN(n7409) );
  AND2_X1 U6362 ( .A1(n7706), .A2(n7714), .ZN(n7650) );
  NAND2_X1 U6363 ( .A1(n7309), .A2(n7681), .ZN(n8847) );
  NOR2_X1 U6364 ( .A1(n6773), .A2(n6772), .ZN(n7283) );
  NOR2_X1 U6365 ( .A1(n5238), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5258) );
  OR2_X1 U6366 ( .A1(n5905), .A2(n10071), .ZN(n5938) );
  INV_X1 U6367 ( .A(n9223), .ZN(n9251) );
  NOR2_X1 U6368 ( .A1(n6075), .A2(n6076), .ZN(n6092) );
  AOI22_X1 U6369 ( .A1(n5681), .A2(n5695), .B1(n5680), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5682) );
  OR2_X1 U6370 ( .A1(n5878), .A2(n5877), .ZN(n5905) );
  NAND2_X1 U6371 ( .A1(n6109), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6159) );
  INV_X1 U6372 ( .A(n9265), .ZN(n9287) );
  NOR2_X1 U6373 ( .A1(n9317), .A2(n9298), .ZN(n6230) );
  AND2_X1 U6374 ( .A1(n6137), .A2(n6315), .ZN(n6512) );
  INV_X1 U6375 ( .A(n9359), .ZN(n9330) );
  AND2_X1 U6376 ( .A1(n9429), .A2(n9095), .ZN(n6226) );
  INV_X1 U6377 ( .A(n7446), .ZN(n7501) );
  NAND2_X1 U6378 ( .A1(n5653), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5654) );
  INV_X1 U6379 ( .A(n8427), .ZN(n9952) );
  AND2_X1 U6380 ( .A1(n6774), .A2(n6775), .ZN(n9945) );
  INV_X1 U6381 ( .A(n8410), .ZN(n9958) );
  AND2_X1 U6382 ( .A1(n7630), .A2(n5499), .ZN(n8460) );
  NAND4_X1 U6383 ( .A1(n5125), .A2(n5124), .A3(n5123), .A4(n5122), .ZN(n5132)
         );
  INV_X1 U6384 ( .A(n9673), .ZN(n9855) );
  INV_X1 U6385 ( .A(n8679), .ZN(n8842) );
  NAND2_X1 U6386 ( .A1(n6770), .A2(n6769), .ZN(n9869) );
  INV_X1 U6387 ( .A(n8613), .ZN(n8778) );
  AND2_X1 U6388 ( .A1(n8827), .A2(n8852), .ZN(n8829) );
  NAND2_X1 U6389 ( .A1(n7178), .A2(n8846), .ZN(n7371) );
  INV_X1 U6390 ( .A(n6770), .ZN(n6772) );
  INV_X1 U6391 ( .A(n5514), .ZN(n6565) );
  XOR2_X1 U6392 ( .A(n5730), .B(n5729), .Z(n6479) );
  AND2_X1 U6393 ( .A1(n6065), .A2(n6064), .ZN(n9238) );
  OR2_X1 U6394 ( .A1(n9510), .A2(n6403), .ZN(n9616) );
  OR2_X1 U6395 ( .A1(n9510), .A2(n9507), .ZN(n9540) );
  INV_X1 U6396 ( .A(n9616), .ZN(n9599) );
  INV_X1 U6397 ( .A(n9540), .ZN(n9610) );
  AND2_X1 U6398 ( .A1(n7584), .A2(n8163), .ZN(n9354) );
  INV_X1 U6399 ( .A(n9347), .ZN(n9335) );
  INV_X1 U6400 ( .A(n9211), .ZN(n9356) );
  INV_X1 U6401 ( .A(n8201), .ZN(n8197) );
  INV_X1 U6402 ( .A(n7962), .ZN(n9222) );
  AND2_X1 U6403 ( .A1(n8057), .A2(n8046), .ZN(n9282) );
  AND2_X1 U6404 ( .A1(n9650), .A2(n9430), .ZN(n9471) );
  INV_X1 U6405 ( .A(n9480), .ZN(n6284) );
  NAND2_X1 U6406 ( .A1(n7467), .A2(n7480), .ZN(n9648) );
  AND2_X1 U6407 ( .A1(n5741), .A2(n5740), .ZN(n6366) );
  AND2_X1 U6408 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7337), .ZN(n7338) );
  OR2_X1 U6409 ( .A1(n6776), .A2(n6775), .ZN(n8427) );
  AND2_X1 U6410 ( .A1(n6793), .A2(n6792), .ZN(n8410) );
  INV_X1 U6411 ( .A(n9950), .ZN(n8458) );
  AND2_X1 U6412 ( .A1(n7630), .A2(n5521), .ZN(n7838) );
  INV_X1 U6413 ( .A(n8417), .ZN(n8718) );
  INV_X1 U6414 ( .A(n7216), .ZN(n8468) );
  INV_X1 U6415 ( .A(n9845), .ZN(n9745) );
  NAND2_X1 U6416 ( .A1(n6803), .A2(n6565), .ZN(n9860) );
  AND2_X1 U6417 ( .A1(n6823), .A2(n9869), .ZN(n9876) );
  INV_X1 U6418 ( .A(n8861), .ZN(n8786) );
  NAND2_X1 U6419 ( .A1(n8827), .A2(n7371), .ZN(n8832) );
  INV_X1 U6420 ( .A(n8827), .ZN(n8857) );
  NAND2_X1 U6421 ( .A1(n9901), .A2(n7371), .ZN(n8937) );
  AND2_X1 U6422 ( .A1(n7285), .A2(n7284), .ZN(n9898) );
  NOR2_X1 U6423 ( .A1(n6772), .A2(n6432), .ZN(n6716) );
  INV_X1 U6424 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7308) );
  INV_X1 U6425 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6342) );
  INV_X1 U6426 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6319) );
  INV_X1 U6427 ( .A(n9035), .ZN(n9080) );
  AND4_X1 U6428 ( .A1(n6127), .A2(n6126), .A3(n6125), .A4(n6124), .ZN(n9202)
         );
  INV_X1 U6429 ( .A(n9298), .ZN(n9338) );
  INV_X1 U6430 ( .A(n9586), .ZN(n9622) );
  OR2_X1 U6431 ( .A1(n6519), .A2(n4331), .ZN(n9363) );
  NAND2_X1 U6432 ( .A1(n9377), .A2(n4897), .ZN(n9378) );
  NAND2_X1 U6433 ( .A1(n9659), .A2(n9648), .ZN(n9427) );
  INV_X1 U6434 ( .A(n9659), .ZN(n9656) );
  NAND2_X1 U6435 ( .A1(n9650), .A2(n9648), .ZN(n9478) );
  INV_X1 U6436 ( .A(n6284), .ZN(n9650) );
  INV_X1 U6437 ( .A(n9623), .ZN(n9624) );
  INV_X1 U6438 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10062) );
  XNOR2_X1 U6439 ( .A(n5623), .B(n5622), .ZN(n7532) );
  INV_X1 U6440 ( .A(n5988), .ZN(n9203) );
  INV_X1 U6441 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6317) );
  NOR2_X1 U6442 ( .A1(n10129), .A2(n10128), .ZN(n10127) );
  INV_X1 U6443 ( .A(n8474), .ZN(P2_U3893) );
  AND2_X2 U6444 ( .A1(n6290), .A2(n6323), .ZN(P1_U3973) );
  NAND2_X1 U6445 ( .A1(n6281), .A2(n6280), .ZN(P1_U3549) );
  NAND2_X1 U6446 ( .A1(n6289), .A2(n6288), .ZN(P1_U3517) );
  NAND2_X1 U6447 ( .A1(n7341), .A2(n4901), .ZN(n4904) );
  INV_X1 U6448 ( .A(n4907), .ZN(n4905) );
  AND2_X1 U6449 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4906) );
  NAND2_X1 U6450 ( .A1(n4907), .A2(n4906), .ZN(n5116) );
  AND2_X1 U6451 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4908) );
  NAND2_X1 U6452 ( .A1(n4986), .A2(n4908), .ZN(n5677) );
  NAND2_X1 U6453 ( .A1(n5116), .A2(n5677), .ZN(n5103) );
  NAND2_X1 U6454 ( .A1(n4909), .A2(n5103), .ZN(n4912) );
  NAND2_X1 U6455 ( .A1(n4910), .A2(SI_1_), .ZN(n4911) );
  NAND2_X1 U6456 ( .A1(n4912), .A2(n4911), .ZN(n5127) );
  INV_X1 U6457 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6299) );
  INV_X1 U6458 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6311) );
  XNOR2_X1 U6459 ( .A(n4914), .B(SI_2_), .ZN(n5126) );
  NAND2_X1 U6460 ( .A1(n5127), .A2(n5126), .ZN(n4917) );
  INV_X1 U6461 ( .A(n4914), .ZN(n4915) );
  NAND2_X1 U6462 ( .A1(n4915), .A2(SI_2_), .ZN(n4916) );
  INV_X1 U6463 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6300) );
  INV_X1 U6464 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6313) );
  XNOR2_X1 U6465 ( .A(n4918), .B(SI_3_), .ZN(n5144) );
  INV_X1 U6466 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6298) );
  INV_X1 U6467 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6308) );
  MUX2_X1 U6468 ( .A(n6298), .B(n6308), .S(n4986), .Z(n4920) );
  XNOR2_X1 U6469 ( .A(n4920), .B(SI_4_), .ZN(n5156) );
  INV_X1 U6470 ( .A(n4920), .ZN(n4921) );
  NAND2_X1 U6471 ( .A1(n4921), .A2(SI_4_), .ZN(n4922) );
  INV_X1 U6472 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6301) );
  INV_X1 U6473 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4923) );
  MUX2_X1 U6474 ( .A(n6301), .B(n4923), .S(n4616), .Z(n4924) );
  XNOR2_X1 U6475 ( .A(n4924), .B(SI_5_), .ZN(n5175) );
  INV_X1 U6476 ( .A(n4924), .ZN(n4925) );
  NAND2_X1 U6477 ( .A1(n4925), .A2(SI_5_), .ZN(n4926) );
  INV_X1 U6478 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n4927) );
  MUX2_X1 U6479 ( .A(n6305), .B(n4927), .S(n4325), .Z(n4928) );
  XNOR2_X1 U6480 ( .A(n4928), .B(SI_6_), .ZN(n5190) );
  INV_X1 U6481 ( .A(n4928), .ZN(n4929) );
  NAND2_X1 U6482 ( .A1(n4929), .A2(SI_6_), .ZN(n4930) );
  MUX2_X1 U6483 ( .A(n6319), .B(n6317), .S(n4325), .Z(n4931) );
  XNOR2_X1 U6484 ( .A(n4931), .B(SI_7_), .ZN(n5203) );
  INV_X1 U6485 ( .A(n4931), .ZN(n4932) );
  NAND2_X1 U6486 ( .A1(n4932), .A2(SI_7_), .ZN(n4933) );
  INV_X1 U6487 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n4935) );
  MUX2_X1 U6488 ( .A(n9984), .B(n4935), .S(n4616), .Z(n4937) );
  INV_X1 U6489 ( .A(SI_8_), .ZN(n4936) );
  NAND2_X1 U6490 ( .A1(n4937), .A2(n4936), .ZN(n4940) );
  INV_X1 U6491 ( .A(n4937), .ZN(n4938) );
  NAND2_X1 U6492 ( .A1(n4938), .A2(SI_8_), .ZN(n4939) );
  INV_X1 U6493 ( .A(n5219), .ZN(n4941) );
  MUX2_X1 U6494 ( .A(n6340), .B(n4942), .S(n4325), .Z(n4944) );
  NAND2_X1 U6495 ( .A1(n4944), .A2(n4943), .ZN(n4947) );
  INV_X1 U6496 ( .A(n4944), .ZN(n4945) );
  NAND2_X1 U6497 ( .A1(n4945), .A2(SI_9_), .ZN(n4946) );
  MUX2_X1 U6498 ( .A(n6342), .B(n4948), .S(n4325), .Z(n4949) );
  XNOR2_X1 U6499 ( .A(n4949), .B(SI_10_), .ZN(n5244) );
  INV_X1 U6500 ( .A(n5244), .ZN(n4952) );
  INV_X1 U6501 ( .A(n4949), .ZN(n4950) );
  NAND2_X1 U6502 ( .A1(n4950), .A2(SI_10_), .ZN(n4951) );
  MUX2_X1 U6503 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n4325), .Z(n5267) );
  MUX2_X1 U6504 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n4325), .Z(n4954) );
  NAND2_X1 U6505 ( .A1(n4954), .A2(SI_12_), .ZN(n5290) );
  INV_X1 U6506 ( .A(n4954), .ZN(n4955) );
  NAND2_X1 U6507 ( .A1(n4955), .A2(n10052), .ZN(n4956) );
  NAND2_X1 U6508 ( .A1(n5290), .A2(n4956), .ZN(n5254) );
  MUX2_X1 U6509 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4325), .Z(n4957) );
  NAND2_X1 U6510 ( .A1(n4957), .A2(SI_13_), .ZN(n5293) );
  NAND2_X1 U6511 ( .A1(n5291), .A2(n4962), .ZN(n4961) );
  INV_X1 U6512 ( .A(n4957), .ZN(n4959) );
  NAND2_X1 U6513 ( .A1(n4961), .A2(n4960), .ZN(n4967) );
  INV_X1 U6514 ( .A(n5292), .ZN(n4963) );
  MUX2_X1 U6515 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4325), .Z(n5313) );
  NAND2_X1 U6516 ( .A1(n4967), .A2(n4966), .ZN(n5330) );
  MUX2_X1 U6517 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4325), .Z(n5328) );
  INV_X1 U6518 ( .A(n5328), .ZN(n4968) );
  MUX2_X1 U6519 ( .A(n10068), .B(n6752), .S(n4325), .Z(n5342) );
  NOR2_X1 U6520 ( .A1(n4969), .A2(SI_16_), .ZN(n4971) );
  NAND2_X1 U6521 ( .A1(n4969), .A2(SI_16_), .ZN(n4970) );
  MUX2_X1 U6522 ( .A(n6998), .B(n6997), .S(n4325), .Z(n4973) );
  NAND2_X1 U6523 ( .A1(n4973), .A2(n4972), .ZN(n4976) );
  INV_X1 U6524 ( .A(n4973), .ZN(n4974) );
  NAND2_X1 U6525 ( .A1(n4974), .A2(SI_17_), .ZN(n4975) );
  NAND2_X1 U6526 ( .A1(n4976), .A2(n4975), .ZN(n5369) );
  MUX2_X1 U6527 ( .A(n7014), .B(n7001), .S(n4325), .Z(n4977) );
  XNOR2_X1 U6528 ( .A(n4977), .B(SI_18_), .ZN(n5357) );
  INV_X1 U6529 ( .A(n5357), .ZN(n4980) );
  INV_X1 U6530 ( .A(n4977), .ZN(n4978) );
  NAND2_X1 U6531 ( .A1(n4978), .A2(SI_18_), .ZN(n4979) );
  MUX2_X1 U6532 ( .A(n7130), .B(n8190), .S(n4325), .Z(n4982) );
  NAND2_X1 U6533 ( .A1(n4982), .A2(n4981), .ZN(n4985) );
  INV_X1 U6534 ( .A(n4982), .ZN(n4983) );
  NAND2_X1 U6535 ( .A1(n4983), .A2(SI_19_), .ZN(n4984) );
  NAND2_X1 U6536 ( .A1(n4985), .A2(n4984), .ZN(n5388) );
  MUX2_X1 U6537 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n4616), .Z(n5402) );
  INV_X1 U6538 ( .A(n5402), .ZN(n4987) );
  MUX2_X1 U6539 ( .A(n7225), .B(n7224), .S(n4325), .Z(n5417) );
  NOR2_X1 U6540 ( .A1(n4988), .A2(SI_21_), .ZN(n4990) );
  NAND2_X1 U6541 ( .A1(n4988), .A2(SI_21_), .ZN(n4989) );
  MUX2_X1 U6542 ( .A(n7308), .B(n7312), .S(n4616), .Z(n4992) );
  INV_X1 U6543 ( .A(SI_22_), .ZN(n4991) );
  NAND2_X1 U6544 ( .A1(n4992), .A2(n4991), .ZN(n4995) );
  INV_X1 U6545 ( .A(n4992), .ZN(n4993) );
  NAND2_X1 U6546 ( .A1(n4993), .A2(SI_22_), .ZN(n4994) );
  NAND2_X1 U6547 ( .A1(n4995), .A2(n4994), .ZN(n5430) );
  INV_X1 U6548 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n4996) );
  INV_X1 U6549 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n6053) );
  MUX2_X1 U6550 ( .A(n4996), .B(n6053), .S(n4325), .Z(n4998) );
  NAND2_X1 U6551 ( .A1(n4998), .A2(n4997), .ZN(n5001) );
  INV_X1 U6552 ( .A(n4998), .ZN(n4999) );
  NAND2_X1 U6553 ( .A1(n4999), .A2(SI_23_), .ZN(n5000) );
  NAND2_X1 U6554 ( .A1(n5443), .A2(n5442), .ZN(n5002) );
  INV_X1 U6555 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7912) );
  MUX2_X1 U6556 ( .A(n7912), .B(n8222), .S(n4616), .Z(n5003) );
  INV_X1 U6557 ( .A(SI_24_), .ZN(n10018) );
  NAND2_X1 U6558 ( .A1(n5003), .A2(n10018), .ZN(n5006) );
  INV_X1 U6559 ( .A(n5003), .ZN(n5004) );
  NAND2_X1 U6560 ( .A1(n5004), .A2(SI_24_), .ZN(n5005) );
  NAND2_X1 U6561 ( .A1(n5007), .A2(n5006), .ZN(n5462) );
  INV_X1 U6562 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7533) );
  INV_X1 U6563 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7531) );
  MUX2_X1 U6564 ( .A(n7533), .B(n7531), .S(n4325), .Z(n5009) );
  INV_X1 U6565 ( .A(SI_25_), .ZN(n5008) );
  NAND2_X1 U6566 ( .A1(n5009), .A2(n5008), .ZN(n5012) );
  INV_X1 U6567 ( .A(n5009), .ZN(n5010) );
  NAND2_X1 U6568 ( .A1(n5010), .A2(SI_25_), .ZN(n5011) );
  INV_X1 U6569 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7539) );
  INV_X1 U6570 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7537) );
  MUX2_X1 U6571 ( .A(n7539), .B(n7537), .S(n4616), .Z(n5014) );
  INV_X1 U6572 ( .A(SI_26_), .ZN(n5013) );
  NAND2_X1 U6573 ( .A1(n5014), .A2(n5013), .ZN(n5017) );
  INV_X1 U6574 ( .A(n5014), .ZN(n5015) );
  NAND2_X1 U6575 ( .A1(n5015), .A2(SI_26_), .ZN(n5016) );
  INV_X1 U6576 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n10040) );
  INV_X1 U6577 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7582) );
  MUX2_X1 U6578 ( .A(n10040), .B(n7582), .S(n4325), .Z(n5019) );
  INV_X1 U6579 ( .A(SI_27_), .ZN(n5018) );
  NAND2_X1 U6580 ( .A1(n5019), .A2(n5018), .ZN(n5022) );
  INV_X1 U6581 ( .A(n5019), .ZN(n5020) );
  NAND2_X1 U6582 ( .A1(n5020), .A2(SI_27_), .ZN(n5021) );
  NAND2_X1 U6583 ( .A1(n5087), .A2(n5088), .ZN(n5023) );
  INV_X1 U6584 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5024) );
  INV_X1 U6585 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7580) );
  MUX2_X1 U6586 ( .A(n5024), .B(n7580), .S(n4616), .Z(n5490) );
  XNOR2_X1 U6587 ( .A(n5490), .B(SI_28_), .ZN(n5487) );
  NOR2_X1 U6588 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5027) );
  AND2_X1 U6589 ( .A1(n5027), .A2(n5026), .ZN(n5031) );
  NAND2_X1 U6590 ( .A1(n5331), .A2(n5028), .ZN(n5345) );
  INV_X1 U6591 ( .A(n5345), .ZN(n5030) );
  NOR3_X2 U6592 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .A3(
        P2_IR_REG_13__SCAN_IN), .ZN(n5029) );
  AND4_X2 U6593 ( .A1(n5235), .A2(n5031), .A3(n5030), .A4(n5029), .ZN(n5359)
         );
  AND2_X2 U6594 ( .A1(n5359), .A2(n5032), .ZN(n5560) );
  NOR2_X1 U6595 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5035) );
  NOR2_X1 U6596 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5034) );
  NOR2_X1 U6597 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5033) );
  NOR2_X4 U6598 ( .A1(n5171), .A2(n5041), .ZN(n5562) );
  XNOR2_X2 U6599 ( .A(n5045), .B(n5044), .ZN(n5514) );
  NAND2_X1 U6600 ( .A1(n7565), .A2(n7635), .ZN(n5047) );
  NAND2_X1 U6601 ( .A1(n5491), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5046) );
  INV_X1 U6602 ( .A(n8867), .ZN(n5545) );
  NAND2_X1 U6603 ( .A1(n7081), .A2(n10017), .ZN(n5164) );
  INV_X1 U6604 ( .A(n5164), .ZN(n5049) );
  NAND2_X1 U6605 ( .A1(n5049), .A2(n5048), .ZN(n5181) );
  INV_X1 U6606 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5061) );
  INV_X1 U6607 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5063) );
  INV_X1 U6608 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5065) );
  INV_X1 U6609 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5067) );
  INV_X1 U6610 ( .A(n5479), .ZN(n5070) );
  INV_X1 U6611 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5069) );
  NAND2_X1 U6612 ( .A1(n5092), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5071) );
  NAND2_X1 U6613 ( .A1(n5494), .A2(n5071), .ZN(n8627) );
  INV_X1 U6614 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5073) );
  NAND2_X1 U6615 ( .A1(n5074), .A2(n5073), .ZN(n8939) );
  XNOR2_X2 U6616 ( .A(n5076), .B(n5075), .ZN(n5080) );
  NAND2_X1 U6617 ( .A1(n5077), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U6618 ( .A1(n8627), .A2(n5495), .ZN(n5086) );
  INV_X1 U6619 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8626) );
  NAND2_X4 U6620 ( .A1(n5079), .A2(n8948), .ZN(n7626) );
  NAND2_X2 U6621 ( .A1(n5080), .A2(n8948), .ZN(n5135) );
  NAND2_X1 U6622 ( .A1(n5516), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5083) );
  AND2_X4 U6623 ( .A1(n5080), .A2(n5081), .ZN(n7622) );
  NAND2_X1 U6624 ( .A1(n7622), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5082) );
  OAI211_X1 U6625 ( .C1(n8626), .C2(n7626), .A(n5083), .B(n5082), .ZN(n5084)
         );
  INV_X1 U6626 ( .A(n5084), .ZN(n5085) );
  NAND2_X1 U6627 ( .A1(n7563), .A2(n7635), .ZN(n5090) );
  OR2_X1 U6628 ( .A1(n7636), .A2(n10040), .ZN(n5089) );
  INV_X1 U6629 ( .A(n8791), .ZN(n5486) );
  NAND2_X1 U6630 ( .A1(n5479), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5091) );
  NAND2_X1 U6631 ( .A1(n5092), .A2(n5091), .ZN(n8637) );
  NAND2_X1 U6632 ( .A1(n8637), .A2(n5495), .ZN(n5097) );
  INV_X1 U6633 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8639) );
  NAND2_X1 U6634 ( .A1(n7622), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U6635 ( .A1(n5516), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5093) );
  OAI211_X1 U6636 ( .C1(n8639), .C2(n7626), .A(n5094), .B(n5093), .ZN(n5095)
         );
  INV_X1 U6637 ( .A(n5095), .ZN(n5096) );
  NAND2_X2 U6638 ( .A1(n5097), .A2(n5096), .ZN(n8646) );
  NAND2_X1 U6639 ( .A1(n7622), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5102) );
  INV_X1 U6640 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6878) );
  OR2_X1 U6641 ( .A1(n7626), .A2(n6878), .ZN(n5101) );
  INV_X1 U6642 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5098) );
  OR2_X1 U6643 ( .A1(n5135), .A2(n5098), .ZN(n5100) );
  INV_X1 U6644 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6879) );
  AND3_X2 U6645 ( .A1(n5102), .A2(n5101), .A3(n4891), .ZN(n5118) );
  INV_X1 U6646 ( .A(n5118), .ZN(n8473) );
  XNOR2_X1 U6647 ( .A(n5104), .B(n5103), .ZN(n6297) );
  NAND2_X1 U6648 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5105) );
  MUX2_X1 U6649 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5105), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5108) );
  INV_X1 U6650 ( .A(n6590), .ZN(n5107) );
  NAND2_X1 U6651 ( .A1(n8473), .A2(n5119), .ZN(n7683) );
  NAND2_X1 U6652 ( .A1(n5118), .A2(n8851), .ZN(n7686) );
  NAND2_X1 U6653 ( .A1(n7683), .A2(n7686), .ZN(n5528) );
  INV_X1 U6654 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6824) );
  OR2_X1 U6655 ( .A1(n5364), .A2(n6824), .ZN(n5113) );
  NAND2_X1 U6656 ( .A1(n7622), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5112) );
  NAND2_X1 U6657 ( .A1(n5166), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5111) );
  NAND2_X1 U6658 ( .A1(n5516), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5110) );
  INV_X1 U6659 ( .A(SI_0_), .ZN(n5114) );
  INV_X1 U6660 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n10055) );
  OAI21_X1 U6661 ( .B1(n4325), .B2(n5114), .A(n10055), .ZN(n5115) );
  AND2_X1 U6662 ( .A1(n5116), .A2(n5115), .ZN(n8949) );
  MUX2_X1 U6663 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8949), .S(n5117), .Z(n8228) );
  NAND2_X1 U6664 ( .A1(n8475), .A2(n8228), .ZN(n6873) );
  NAND2_X1 U6665 ( .A1(n5528), .A2(n6873), .ZN(n5121) );
  NAND2_X1 U6666 ( .A1(n5118), .A2(n5119), .ZN(n5120) );
  NAND2_X1 U6667 ( .A1(n5121), .A2(n5120), .ZN(n8836) );
  NAND2_X1 U6668 ( .A1(n7622), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U6669 ( .A1(n4322), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5124) );
  NAND2_X1 U6670 ( .A1(n5516), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5123) );
  NAND2_X1 U6671 ( .A1(n5495), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5122) );
  XNOR2_X1 U6672 ( .A(n5127), .B(n5126), .ZN(n6310) );
  OR2_X1 U6673 ( .A1(n5221), .A2(n6310), .ZN(n5131) );
  OR2_X1 U6674 ( .A1(n7636), .A2(n6299), .ZN(n5130) );
  NOR2_X1 U6675 ( .A1(n6590), .A2(n8940), .ZN(n5128) );
  NAND2_X1 U6676 ( .A1(n6293), .A2(n8483), .ZN(n5129) );
  OR2_X1 U6677 ( .A1(n5132), .A2(n9867), .ZN(n7690) );
  NAND2_X1 U6678 ( .A1(n5132), .A2(n9867), .ZN(n7691) );
  NAND2_X1 U6679 ( .A1(n7690), .A2(n7691), .ZN(n8837) );
  NAND2_X1 U6680 ( .A1(n8836), .A2(n8837), .ZN(n5134) );
  INV_X1 U6681 ( .A(n9867), .ZN(n6865) );
  OR2_X1 U6682 ( .A1(n5132), .A2(n6865), .ZN(n5133) );
  NAND2_X1 U6683 ( .A1(n5134), .A2(n5133), .ZN(n6711) );
  NAND2_X1 U6684 ( .A1(n7622), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5140) );
  OR2_X1 U6685 ( .A1(n5364), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5139) );
  INV_X1 U6686 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7080) );
  OR2_X1 U6687 ( .A1(n7626), .A2(n7080), .ZN(n5138) );
  INV_X1 U6688 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5136) );
  OR2_X1 U6689 ( .A1(n5135), .A2(n5136), .ZN(n5137) );
  NAND2_X1 U6690 ( .A1(n5141), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5142) );
  MUX2_X1 U6691 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5142), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5143) );
  NAND2_X1 U6692 ( .A1(n5143), .A2(n5171), .ZN(n6599) );
  XNOR2_X1 U6693 ( .A(n5145), .B(n5144), .ZN(n6312) );
  OR2_X1 U6694 ( .A1(n5221), .A2(n6312), .ZN(n5147) );
  OR2_X1 U6695 ( .A1(n7636), .A2(n6300), .ZN(n5146) );
  OAI211_X1 U6696 ( .C1(n5117), .C2(n6599), .A(n5147), .B(n5146), .ZN(n7082)
         );
  NAND2_X1 U6697 ( .A1(n8839), .A2(n7082), .ZN(n7709) );
  INV_X1 U6698 ( .A(n7082), .ZN(n6789) );
  NAND2_X1 U6699 ( .A1(n8472), .A2(n6789), .ZN(n7698) );
  NAND2_X1 U6700 ( .A1(n7709), .A2(n7698), .ZN(n7647) );
  NAND2_X1 U6701 ( .A1(n6711), .A2(n7647), .ZN(n5149) );
  NAND2_X1 U6702 ( .A1(n8839), .A2(n6789), .ZN(n5148) );
  NAND2_X1 U6703 ( .A1(n5516), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5154) );
  INV_X1 U6704 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6603) );
  OR2_X1 U6705 ( .A1(n5409), .A2(n6603), .ZN(n5153) );
  NAND2_X1 U6706 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5150) );
  AND2_X1 U6707 ( .A1(n5164), .A2(n5150), .ZN(n6932) );
  OR2_X1 U6708 ( .A1(n5364), .A2(n6932), .ZN(n5152) );
  INV_X1 U6709 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7135) );
  OR2_X1 U6710 ( .A1(n7626), .A2(n7135), .ZN(n5151) );
  NAND2_X1 U6711 ( .A1(n5161), .A2(n7007), .ZN(n5160) );
  NAND2_X1 U6712 ( .A1(n5171), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5155) );
  XNOR2_X1 U6713 ( .A(n5155), .B(n5040), .ZN(n9683) );
  XNOR2_X1 U6714 ( .A(n5157), .B(n5156), .ZN(n6307) );
  OR2_X1 U6715 ( .A1(n5221), .A2(n6307), .ZN(n5159) );
  OR2_X1 U6716 ( .A1(n7636), .A2(n6298), .ZN(n5158) );
  OAI211_X1 U6717 ( .C1(n5117), .C2(n9683), .A(n5159), .B(n5158), .ZN(n7137)
         );
  NAND2_X1 U6718 ( .A1(n5160), .A2(n7137), .ZN(n5163) );
  NAND2_X1 U6719 ( .A1(n6849), .A2(n8471), .ZN(n5162) );
  NAND2_X1 U6720 ( .A1(n5163), .A2(n5162), .ZN(n6810) );
  NAND2_X1 U6721 ( .A1(n7622), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6722 ( .A1(n5164), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5165) );
  AND2_X1 U6723 ( .A1(n5181), .A2(n5165), .ZN(n7012) );
  OR2_X1 U6724 ( .A1(n5364), .A2(n7012), .ZN(n5169) );
  NAND2_X1 U6725 ( .A1(n5516), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U6726 ( .A1(n5166), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5167) );
  NAND4_X1 U6727 ( .A1(n5170), .A2(n5169), .A3(n5168), .A4(n5167), .ZN(n8470)
         );
  NOR2_X1 U6728 ( .A1(n5171), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5172) );
  OR2_X1 U6729 ( .A1(n5172), .A2(n8940), .ZN(n5174) );
  XNOR2_X1 U6730 ( .A(n5174), .B(n5173), .ZN(n6660) );
  XNOR2_X1 U6731 ( .A(n5176), .B(n5175), .ZN(n6303) );
  OR2_X1 U6732 ( .A1(n5221), .A2(n6303), .ZN(n5178) );
  OR2_X1 U6733 ( .A1(n7636), .A2(n6301), .ZN(n5177) );
  OAI211_X1 U6734 ( .C1(n5117), .C2(n6660), .A(n5178), .B(n5177), .ZN(n7699)
         );
  AND2_X1 U6735 ( .A1(n8470), .A2(n7699), .ZN(n5180) );
  INV_X1 U6736 ( .A(n7699), .ZN(n7704) );
  NAND2_X1 U6737 ( .A1(n7700), .A2(n7704), .ZN(n5179) );
  NAND2_X1 U6738 ( .A1(n5516), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6739 ( .A1(n5181), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5182) );
  AND2_X1 U6740 ( .A1(n5195), .A2(n5182), .ZN(n7072) );
  OR2_X1 U6741 ( .A1(n5364), .A2(n7072), .ZN(n5185) );
  NAND2_X1 U6742 ( .A1(n7622), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6743 ( .A1(n4322), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5183) );
  NAND4_X1 U6744 ( .A1(n5186), .A2(n5185), .A3(n5184), .A4(n5183), .ZN(n8469)
         );
  NOR2_X1 U6745 ( .A1(n5562), .A2(n8940), .ZN(n5187) );
  MUX2_X1 U6746 ( .A(n8940), .B(n5187), .S(P2_IR_REG_6__SCAN_IN), .Z(n5189) );
  AND2_X1 U6747 ( .A1(n5562), .A2(n5201), .ZN(n5188) );
  XNOR2_X1 U6748 ( .A(n5191), .B(n5190), .ZN(n6306) );
  OR2_X1 U6749 ( .A1(n5221), .A2(n6306), .ZN(n5193) );
  OR2_X1 U6750 ( .A1(n7636), .A2(n6305), .ZN(n5192) );
  OAI211_X1 U6751 ( .C1(n5117), .C2(n9714), .A(n5193), .B(n5192), .ZN(n7074)
         );
  NOR2_X1 U6752 ( .A1(n8469), .A2(n7074), .ZN(n5194) );
  NAND2_X1 U6753 ( .A1(n5516), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5200) );
  OR2_X1 U6754 ( .A1(n5409), .A2(n7039), .ZN(n5199) );
  NAND2_X1 U6755 ( .A1(n5195), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5196) );
  AND2_X1 U6756 ( .A1(n5208), .A2(n5196), .ZN(n7167) );
  OR2_X1 U6757 ( .A1(n5364), .A2(n7167), .ZN(n5198) );
  OR2_X1 U6758 ( .A1(n7626), .A2(n4678), .ZN(n5197) );
  NAND2_X1 U6759 ( .A1(n5562), .A2(n5201), .ZN(n5215) );
  NAND2_X1 U6760 ( .A1(n5215), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5202) );
  INV_X1 U6761 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n9971) );
  XNOR2_X1 U6762 ( .A(n5202), .B(n9971), .ZN(n6901) );
  OR2_X1 U6763 ( .A1(n7636), .A2(n6319), .ZN(n5206) );
  XNOR2_X1 U6764 ( .A(n5204), .B(n5203), .ZN(n6318) );
  OR2_X1 U6765 ( .A1(n5221), .A2(n6318), .ZN(n5205) );
  OAI211_X1 U6766 ( .C1(n5117), .C2(n6901), .A(n5206), .B(n5205), .ZN(n7166)
         );
  NAND2_X1 U6767 ( .A1(n7216), .A2(n7166), .ZN(n7722) );
  INV_X1 U6768 ( .A(n7166), .ZN(n7154) );
  NAND2_X1 U6769 ( .A1(n8468), .A2(n7154), .ZN(n7086) );
  NAND2_X1 U6770 ( .A1(n5516), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5214) );
  INV_X1 U6771 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6899) );
  OR2_X1 U6772 ( .A1(n5409), .A2(n6899), .ZN(n5213) );
  NAND2_X1 U6773 ( .A1(n5208), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5209) );
  AND2_X1 U6774 ( .A1(n5227), .A2(n5209), .ZN(n7222) );
  OR2_X1 U6775 ( .A1(n5364), .A2(n7222), .ZN(n5212) );
  INV_X1 U6776 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5210) );
  OR2_X1 U6777 ( .A1(n7626), .A2(n5210), .ZN(n5211) );
  OR2_X1 U6778 ( .A1(n5215), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6779 ( .A1(n5216), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5218) );
  INV_X1 U6780 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5217) );
  XNOR2_X1 U6781 ( .A(n5218), .B(n5217), .ZN(n8533) );
  OR2_X1 U6782 ( .A1(n5221), .A2(n6327), .ZN(n5223) );
  OR2_X1 U6783 ( .A1(n7636), .A2(n9984), .ZN(n5222) );
  OAI211_X1 U6784 ( .C1(n5117), .C2(n8533), .A(n5223), .B(n5222), .ZN(n7219)
         );
  NAND2_X1 U6785 ( .A1(n7237), .A2(n7219), .ZN(n7727) );
  INV_X1 U6786 ( .A(n7237), .ZN(n8467) );
  INV_X1 U6787 ( .A(n7219), .ZN(n7213) );
  NAND2_X1 U6788 ( .A1(n8467), .A2(n7213), .ZN(n7728) );
  NAND2_X1 U6789 ( .A1(n7727), .A2(n7728), .ZN(n7652) );
  NAND2_X1 U6790 ( .A1(n7216), .A2(n7154), .ZN(n7089) );
  AND2_X1 U6791 ( .A1(n7652), .A2(n7089), .ZN(n5224) );
  NAND2_X1 U6792 ( .A1(n7033), .A2(n5224), .ZN(n7088) );
  NAND2_X1 U6793 ( .A1(n8467), .A2(n7219), .ZN(n5225) );
  NAND2_X1 U6794 ( .A1(n7088), .A2(n5225), .ZN(n7174) );
  INV_X1 U6795 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5226) );
  OR2_X1 U6796 ( .A1(n5409), .A2(n5226), .ZN(n5232) );
  NAND2_X1 U6797 ( .A1(n5227), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5228) );
  AND2_X1 U6798 ( .A1(n5248), .A2(n5228), .ZN(n7242) );
  OR2_X1 U6799 ( .A1(n5364), .A2(n7242), .ZN(n5231) );
  NAND2_X1 U6800 ( .A1(n5516), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U6801 ( .A1(n4322), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5229) );
  NAND4_X1 U6802 ( .A1(n5232), .A2(n5231), .A3(n5230), .A4(n5229), .ZN(n8466)
         );
  NAND2_X1 U6803 ( .A1(n6336), .A2(n7635), .ZN(n5241) );
  NAND2_X1 U6804 ( .A1(n5562), .A2(n5235), .ZN(n5238) );
  NAND2_X1 U6805 ( .A1(n5238), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5236) );
  MUX2_X1 U6806 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5236), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n5237) );
  INV_X1 U6807 ( .A(n5237), .ZN(n5239) );
  NOR2_X1 U6808 ( .A1(n5239), .A2(n5258), .ZN(n9734) );
  AOI22_X1 U6809 ( .A1(n5491), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6293), .B2(
        n9734), .ZN(n5240) );
  NAND2_X1 U6810 ( .A1(n5241), .A2(n5240), .ZN(n7239) );
  AND2_X1 U6811 ( .A1(n8466), .A2(n7239), .ZN(n5242) );
  XNOR2_X1 U6812 ( .A(n5243), .B(n5244), .ZN(n6338) );
  NAND2_X1 U6813 ( .A1(n6338), .A2(n7635), .ZN(n5247) );
  OR2_X1 U6814 ( .A1(n5258), .A2(n8940), .ZN(n5245) );
  XNOR2_X1 U6815 ( .A(n5245), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9746) );
  AOI22_X1 U6816 ( .A1(n5491), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6293), .B2(
        n9746), .ZN(n5246) );
  NAND2_X1 U6817 ( .A1(n5247), .A2(n5246), .ZN(n8309) );
  NAND2_X1 U6818 ( .A1(n5516), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U6819 ( .A1(n5248), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5249) );
  AND2_X1 U6820 ( .A1(n5274), .A2(n5249), .ZN(n8310) );
  OR2_X1 U6821 ( .A1(n5364), .A2(n8310), .ZN(n5252) );
  NAND2_X1 U6822 ( .A1(n7622), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5251) );
  NAND2_X1 U6823 ( .A1(n5166), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5250) );
  NAND4_X1 U6824 ( .A1(n5253), .A2(n5252), .A3(n5251), .A4(n5250), .ZN(n9944)
         );
  NOR2_X1 U6825 ( .A1(n8309), .A2(n9944), .ZN(n7257) );
  NAND2_X1 U6826 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  NAND2_X1 U6827 ( .A1(n6475), .A2(n7635), .ZN(n5261) );
  INV_X1 U6828 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U6829 ( .A1(n5258), .A2(n5257), .ZN(n5270) );
  NAND2_X1 U6830 ( .A1(n5300), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5259) );
  XNOR2_X1 U6831 ( .A(n5259), .B(P2_IR_REG_12__SCAN_IN), .ZN(n9778) );
  AOI22_X1 U6832 ( .A1(n5491), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6293), .B2(
        n9778), .ZN(n5260) );
  NAND2_X1 U6833 ( .A1(n5261), .A2(n5260), .ZN(n7420) );
  NAND2_X1 U6834 ( .A1(n5276), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5262) );
  AND2_X1 U6835 ( .A1(n5305), .A2(n5262), .ZN(n7418) );
  OR2_X1 U6836 ( .A1(n5364), .A2(n7418), .ZN(n5266) );
  INV_X1 U6837 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7355) );
  OR2_X1 U6838 ( .A1(n7626), .A2(n7355), .ZN(n5265) );
  NAND2_X1 U6839 ( .A1(n5516), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5264) );
  NAND2_X1 U6840 ( .A1(n7622), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5263) );
  NAND4_X1 U6841 ( .A1(n5266), .A2(n5265), .A3(n5264), .A4(n5263), .ZN(n9951)
         );
  AND2_X1 U6842 ( .A1(n7420), .A2(n9951), .ZN(n5285) );
  INV_X1 U6843 ( .A(n9951), .ZN(n7263) );
  NAND2_X1 U6844 ( .A1(n7415), .A2(n7263), .ZN(n5283) );
  XNOR2_X1 U6845 ( .A(n5267), .B(SI_11_), .ZN(n5268) );
  XNOR2_X1 U6846 ( .A(n5269), .B(n5268), .ZN(n6438) );
  NAND2_X1 U6847 ( .A1(n5270), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5271) );
  XNOR2_X1 U6848 ( .A(n5271), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9764) );
  AOI22_X1 U6849 ( .A1(n5491), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6293), .B2(
        n9764), .ZN(n5272) );
  NAND2_X1 U6850 ( .A1(n5516), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5281) );
  INV_X1 U6851 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5273) );
  OR2_X1 U6852 ( .A1(n5409), .A2(n5273), .ZN(n5280) );
  NAND2_X1 U6853 ( .A1(n5274), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5275) );
  AND2_X1 U6854 ( .A1(n5276), .A2(n5275), .ZN(n9946) );
  OR2_X1 U6855 ( .A1(n5364), .A2(n9946), .ZN(n5279) );
  INV_X1 U6856 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5277) );
  OR2_X1 U6857 ( .A1(n7626), .A2(n5277), .ZN(n5278) );
  NAND2_X1 U6858 ( .A1(n9949), .A2(n4441), .ZN(n5284) );
  INV_X1 U6859 ( .A(n5284), .ZN(n5282) );
  NAND2_X1 U6860 ( .A1(n9949), .A2(n7408), .ZN(n7752) );
  OR2_X1 U6861 ( .A1(n5282), .A2(n7261), .ZN(n7352) );
  NAND2_X1 U6862 ( .A1(n8309), .A2(n9944), .ZN(n7259) );
  AND2_X1 U6863 ( .A1(n7259), .A2(n5284), .ZN(n7349) );
  INV_X1 U6864 ( .A(n5285), .ZN(n5286) );
  AND2_X1 U6865 ( .A1(n7349), .A2(n5286), .ZN(n5287) );
  OR2_X1 U6866 ( .A1(n5288), .A2(n5287), .ZN(n5289) );
  AND2_X1 U6867 ( .A1(n5291), .A2(n5290), .ZN(n5294) );
  NAND2_X1 U6868 ( .A1(n5293), .A2(n5292), .ZN(n5295) );
  NAND2_X1 U6869 ( .A1(n5294), .A2(n5295), .ZN(n5299) );
  INV_X1 U6870 ( .A(n5294), .ZN(n5297) );
  INV_X1 U6871 ( .A(n5295), .ZN(n5296) );
  NAND2_X1 U6872 ( .A1(n5297), .A2(n5296), .ZN(n5298) );
  NAND2_X1 U6873 ( .A1(n6507), .A2(n7635), .ZN(n5303) );
  OR2_X1 U6874 ( .A1(n5316), .A2(n8940), .ZN(n5301) );
  XNOR2_X1 U6875 ( .A(n5301), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9795) );
  AOI22_X1 U6876 ( .A1(n5491), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6293), .B2(
        n9795), .ZN(n5302) );
  INV_X1 U6877 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5304) );
  OR2_X1 U6878 ( .A1(n5409), .A2(n5304), .ZN(n5310) );
  NAND2_X1 U6879 ( .A1(n5305), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5306) );
  AND2_X1 U6880 ( .A1(n5320), .A2(n5306), .ZN(n8406) );
  OR2_X1 U6881 ( .A1(n5364), .A2(n8406), .ZN(n5309) );
  INV_X1 U6882 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8498) );
  OR2_X1 U6883 ( .A1(n7626), .A2(n8498), .ZN(n5308) );
  NAND2_X1 U6884 ( .A1(n5516), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5307) );
  NAND4_X1 U6885 ( .A1(n5310), .A2(n5309), .A3(n5308), .A4(n5307), .ZN(n8465)
         );
  NOR2_X1 U6886 ( .A1(n8408), .A2(n8465), .ZN(n5311) );
  INV_X1 U6887 ( .A(n8408), .ZN(n7289) );
  XNOR2_X1 U6888 ( .A(n5313), .B(SI_14_), .ZN(n5314) );
  XNOR2_X1 U6889 ( .A(n5312), .B(n5314), .ZN(n6533) );
  NAND2_X1 U6890 ( .A1(n6533), .A2(n7635), .ZN(n5319) );
  INV_X1 U6891 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6892 ( .A1(n5316), .A2(n5315), .ZN(n5317) );
  NAND2_X1 U6893 ( .A1(n5317), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5347) );
  XNOR2_X1 U6894 ( .A(n5347), .B(P2_IR_REG_14__SCAN_IN), .ZN(n9812) );
  AOI22_X1 U6895 ( .A1(n5491), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6293), .B2(
        n9812), .ZN(n5318) );
  INV_X1 U6896 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8513) );
  OR2_X1 U6897 ( .A1(n5409), .A2(n8513), .ZN(n5326) );
  NAND2_X1 U6898 ( .A1(n5320), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5321) );
  AND2_X1 U6899 ( .A1(n5336), .A2(n5321), .ZN(n8287) );
  OR2_X1 U6900 ( .A1(n5364), .A2(n8287), .ZN(n5325) );
  INV_X1 U6901 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5322) );
  OR2_X1 U6902 ( .A1(n7626), .A2(n5322), .ZN(n5324) );
  NAND2_X1 U6903 ( .A1(n5516), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5323) );
  NAND4_X1 U6904 ( .A1(n5326), .A2(n5325), .A3(n5324), .A4(n5323), .ZN(n8464)
         );
  OR2_X1 U6905 ( .A1(n8286), .A2(n8464), .ZN(n5327) );
  XNOR2_X1 U6906 ( .A(n5328), .B(SI_15_), .ZN(n5329) );
  XNOR2_X1 U6907 ( .A(n5330), .B(n5329), .ZN(n6691) );
  NAND2_X1 U6908 ( .A1(n6691), .A2(n7635), .ZN(n5335) );
  NAND2_X1 U6909 ( .A1(n5347), .A2(n5331), .ZN(n5332) );
  NAND2_X1 U6910 ( .A1(n5332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5333) );
  XNOR2_X1 U6911 ( .A(n5333), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9830) );
  AOI22_X1 U6912 ( .A1(n5491), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n9830), .B2(
        n6293), .ZN(n5334) );
  INV_X1 U6913 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9969) );
  OR2_X1 U6914 ( .A1(n5409), .A2(n9969), .ZN(n5341) );
  NAND2_X1 U6915 ( .A1(n5336), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5337) );
  AND2_X1 U6916 ( .A1(n5351), .A2(n5337), .ZN(n7526) );
  OR2_X1 U6917 ( .A1(n5364), .A2(n7526), .ZN(n5340) );
  NAND2_X1 U6918 ( .A1(n5516), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6919 ( .A1(n5166), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5338) );
  NAND4_X1 U6920 ( .A1(n5341), .A2(n5340), .A3(n5339), .A4(n5338), .ZN(n8770)
         );
  INV_X1 U6921 ( .A(n8770), .ZN(n7507) );
  INV_X1 U6922 ( .A(n8243), .ZN(n8459) );
  XNOR2_X1 U6923 ( .A(n5342), .B(SI_16_), .ZN(n5343) );
  XNOR2_X1 U6924 ( .A(n5344), .B(n5343), .ZN(n6751) );
  NAND2_X1 U6925 ( .A1(n6751), .A2(n7635), .ZN(n5350) );
  NAND2_X1 U6926 ( .A1(n5345), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6927 ( .A1(n5347), .A2(n5346), .ZN(n5371) );
  INV_X1 U6928 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5348) );
  XNOR2_X1 U6929 ( .A(n5371), .B(n5348), .ZN(n9847) );
  AOI22_X1 U6930 ( .A1(n5491), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6293), .B2(
        n9847), .ZN(n5349) );
  NAND2_X1 U6931 ( .A1(n5516), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5356) );
  INV_X1 U6932 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8828) );
  OR2_X1 U6933 ( .A1(n5409), .A2(n8828), .ZN(n5355) );
  NAND2_X1 U6934 ( .A1(n5351), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5352) );
  AND2_X1 U6935 ( .A1(n5375), .A2(n5352), .ZN(n8775) );
  OR2_X1 U6936 ( .A1(n5364), .A2(n8775), .ZN(n5354) );
  INV_X1 U6937 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8774) );
  OR2_X1 U6938 ( .A1(n7626), .A2(n8774), .ZN(n5353) );
  NAND2_X1 U6939 ( .A1(n8934), .A2(n8353), .ZN(n7777) );
  NAND2_X1 U6940 ( .A1(n7779), .A2(n7777), .ZN(n8767) );
  NAND2_X1 U6941 ( .A1(n8768), .A2(n8767), .ZN(n8742) );
  NAND2_X1 U6942 ( .A1(n8934), .A2(n8757), .ZN(n8741) );
  XNOR2_X1 U6943 ( .A(n5358), .B(n5357), .ZN(n7000) );
  NAND2_X1 U6944 ( .A1(n7000), .A2(n7635), .ZN(n5362) );
  NAND2_X1 U6945 ( .A1(n4405), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5360) );
  XNOR2_X1 U6946 ( .A(n5360), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8586) );
  AOI22_X1 U6947 ( .A1(n5491), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6293), .B2(
        n8586), .ZN(n5361) );
  NAND2_X1 U6948 ( .A1(n5516), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U6949 ( .A1(n5377), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5363) );
  AND2_X1 U6950 ( .A1(n5394), .A2(n5363), .ZN(n8750) );
  OR2_X1 U6951 ( .A1(n5364), .A2(n8750), .ZN(n5367) );
  NAND2_X1 U6952 ( .A1(n7622), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U6953 ( .A1(n4322), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5365) );
  NAND4_X1 U6954 ( .A1(n5368), .A2(n5367), .A3(n5366), .A4(n5365), .ZN(n8758)
         );
  NAND2_X1 U6955 ( .A1(n8921), .A2(n8758), .ZN(n5382) );
  XNOR2_X1 U6956 ( .A(n5370), .B(n5369), .ZN(n6996) );
  NAND2_X1 U6957 ( .A1(n6996), .A2(n7635), .ZN(n5374) );
  OAI21_X1 U6958 ( .B1(n5371), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5372) );
  XNOR2_X1 U6959 ( .A(n5372), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8566) );
  AOI22_X1 U6960 ( .A1(n8566), .A2(n6293), .B1(n5491), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6961 ( .A1(n5516), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5381) );
  INV_X1 U6962 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8824) );
  OR2_X1 U6963 ( .A1(n5409), .A2(n8824), .ZN(n5380) );
  NAND2_X1 U6964 ( .A1(n5375), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5376) );
  AND2_X1 U6965 ( .A1(n5377), .A2(n5376), .ZN(n8761) );
  OR2_X1 U6966 ( .A1(n5364), .A2(n8761), .ZN(n5379) );
  INV_X1 U6967 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8760) );
  OR2_X1 U6968 ( .A1(n7626), .A2(n8760), .ZN(n5378) );
  NAND2_X1 U6969 ( .A1(n8927), .A2(n8772), .ZN(n8744) );
  AND2_X1 U6970 ( .A1(n5382), .A2(n8744), .ZN(n5384) );
  AND2_X1 U6971 ( .A1(n8741), .A2(n5384), .ZN(n5383) );
  INV_X1 U6972 ( .A(n5384), .ZN(n5385) );
  NAND2_X1 U6973 ( .A1(n8927), .A2(n8250), .ZN(n7785) );
  NAND2_X1 U6974 ( .A1(n7778), .A2(n7785), .ZN(n8743) );
  OR2_X1 U6975 ( .A1(n5385), .A2(n8743), .ZN(n5386) );
  OR2_X1 U6976 ( .A1(n8921), .A2(n8758), .ZN(n5387) );
  XNOR2_X1 U6977 ( .A(n5389), .B(n5388), .ZN(n7129) );
  NAND2_X1 U6978 ( .A1(n7129), .A2(n7635), .ZN(n5392) );
  NAND2_X1 U6979 ( .A1(n5500), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5390) );
  AOI22_X1 U6980 ( .A1(n5491), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8592), .B2(
        n6293), .ZN(n5391) );
  NAND2_X1 U6981 ( .A1(n5516), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5399) );
  INV_X1 U6982 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5393) );
  OR2_X1 U6983 ( .A1(n5409), .A2(n5393), .ZN(n5398) );
  NAND2_X1 U6984 ( .A1(n5394), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5395) );
  AND2_X1 U6985 ( .A1(n5407), .A2(n5395), .ZN(n8736) );
  OR2_X1 U6986 ( .A1(n5364), .A2(n8736), .ZN(n5397) );
  INV_X1 U6987 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8734) );
  OR2_X1 U6988 ( .A1(n7626), .A2(n8734), .ZN(n5396) );
  OR2_X1 U6989 ( .A1(n8738), .A2(n8426), .ZN(n7783) );
  NAND2_X1 U6990 ( .A1(n8738), .A2(n8426), .ZN(n7790) );
  NAND2_X1 U6991 ( .A1(n8738), .A2(n8748), .ZN(n5400) );
  XNOR2_X1 U6992 ( .A(n5402), .B(n5401), .ZN(n5403) );
  XNOR2_X1 U6993 ( .A(n5404), .B(n5403), .ZN(n7183) );
  NAND2_X1 U6994 ( .A1(n7183), .A2(n7635), .ZN(n5406) );
  INV_X1 U6995 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10004) );
  OR2_X1 U6996 ( .A1(n7636), .A2(n10004), .ZN(n5405) );
  NAND2_X1 U6997 ( .A1(n5407), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U6998 ( .A1(n5423), .A2(n5408), .ZN(n8714) );
  NAND2_X1 U6999 ( .A1(n5495), .A2(n8714), .ZN(n5414) );
  INV_X1 U7000 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8908) );
  OR2_X1 U7001 ( .A1(n5135), .A2(n8908), .ZN(n5413) );
  INV_X1 U7002 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8815) );
  OR2_X1 U7003 ( .A1(n5409), .A2(n8815), .ZN(n5412) );
  INV_X1 U7004 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5410) );
  OR2_X1 U7005 ( .A1(n7626), .A2(n5410), .ZN(n5411) );
  NAND2_X1 U7006 ( .A1(n8909), .A2(n8699), .ZN(n8707) );
  NAND2_X1 U7007 ( .A1(n7794), .A2(n8707), .ZN(n8716) );
  INV_X1 U7008 ( .A(n8699), .ZN(n8731) );
  OR2_X1 U7009 ( .A1(n8731), .A2(n8909), .ZN(n5415) );
  XNOR2_X1 U7010 ( .A(n5417), .B(SI_21_), .ZN(n5418) );
  XNOR2_X1 U7011 ( .A(n5416), .B(n5418), .ZN(n7223) );
  NAND2_X1 U7012 ( .A1(n7223), .A2(n7635), .ZN(n5420) );
  NAND2_X1 U7013 ( .A1(n5491), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U7014 ( .A1(n5516), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U7015 ( .A1(n7622), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5421) );
  AND2_X1 U7016 ( .A1(n5422), .A2(n5421), .ZN(n5427) );
  NAND2_X1 U7017 ( .A1(n5423), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U7018 ( .A1(n5436), .A2(n5424), .ZN(n8703) );
  NAND2_X1 U7019 ( .A1(n8703), .A2(n5495), .ZN(n5426) );
  NAND2_X1 U7020 ( .A1(n5166), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U7021 ( .A1(n8810), .A2(n8417), .ZN(n7801) );
  NAND2_X1 U7022 ( .A1(n7800), .A2(n7801), .ZN(n8709) );
  OR2_X1 U7023 ( .A1(n8810), .A2(n8718), .ZN(n5428) );
  NAND2_X1 U7024 ( .A1(n5429), .A2(n5428), .ZN(n8690) );
  NAND2_X1 U7025 ( .A1(n5431), .A2(n5430), .ZN(n5432) );
  NAND2_X1 U7026 ( .A1(n5433), .A2(n5432), .ZN(n7307) );
  NAND2_X1 U7027 ( .A1(n7307), .A2(n7635), .ZN(n5435) );
  NAND2_X1 U7028 ( .A1(n5491), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U7029 ( .A1(n5436), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U7030 ( .A1(n5446), .A2(n5437), .ZN(n8695) );
  NAND2_X1 U7031 ( .A1(n8695), .A2(n5495), .ZN(n5440) );
  AOI22_X1 U7032 ( .A1(n5516), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n7622), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U7033 ( .A1(n4322), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5438) );
  NAND2_X1 U7034 ( .A1(n8899), .A2(n8700), .ZN(n7804) );
  NAND2_X1 U7035 ( .A1(n7805), .A2(n7804), .ZN(n8689) );
  INV_X1 U7036 ( .A(n8700), .ZN(n8463) );
  OR2_X1 U7037 ( .A1(n8899), .A2(n8463), .ZN(n5441) );
  XNOR2_X1 U7038 ( .A(n5443), .B(n5442), .ZN(n7398) );
  NAND2_X1 U7039 ( .A1(n7398), .A2(n7635), .ZN(n5445) );
  NAND2_X1 U7040 ( .A1(n5491), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5444) );
  INV_X1 U7041 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8894) );
  NAND2_X1 U7042 ( .A1(n5446), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U7043 ( .A1(n5453), .A2(n5447), .ZN(n8681) );
  NAND2_X1 U7044 ( .A1(n8681), .A2(n5495), .ZN(n5449) );
  AOI22_X1 U7045 ( .A1(n5166), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n7622), .B2(
        P2_REG1_REG_23__SCAN_IN), .ZN(n5448) );
  OAI211_X1 U7046 ( .C1(n5135), .C2(n8894), .A(n5449), .B(n5448), .ZN(n8691)
         );
  NAND2_X1 U7047 ( .A1(n7911), .A2(n7635), .ZN(n5452) );
  NAND2_X1 U7048 ( .A1(n5491), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U7049 ( .A1(n5453), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U7050 ( .A1(n5466), .A2(n5454), .ZN(n8671) );
  NAND2_X1 U7051 ( .A1(n8671), .A2(n5495), .ZN(n5459) );
  INV_X1 U7052 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8670) );
  NAND2_X1 U7053 ( .A1(n7622), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U7054 ( .A1(n5516), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5455) );
  OAI211_X1 U7055 ( .C1(n7626), .C2(n8670), .A(n5456), .B(n5455), .ZN(n5457)
         );
  INV_X1 U7056 ( .A(n5457), .ZN(n5458) );
  NAND2_X1 U7057 ( .A1(n8889), .A2(n8462), .ZN(n5461) );
  NOR2_X1 U7058 ( .A1(n8889), .A2(n8462), .ZN(n5460) );
  XNOR2_X1 U7059 ( .A(n5462), .B(n5463), .ZN(n7530) );
  NAND2_X1 U7060 ( .A1(n7530), .A2(n7635), .ZN(n5465) );
  NAND2_X1 U7061 ( .A1(n5491), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U7062 ( .A1(n5466), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U7063 ( .A1(n5477), .A2(n5467), .ZN(n8660) );
  NAND2_X1 U7064 ( .A1(n8660), .A2(n5495), .ZN(n5472) );
  INV_X1 U7065 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8659) );
  NAND2_X1 U7066 ( .A1(n5516), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U7067 ( .A1(n7622), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5468) );
  OAI211_X1 U7068 ( .C1(n8659), .C2(n7626), .A(n5469), .B(n5468), .ZN(n5470)
         );
  INV_X1 U7069 ( .A(n5470), .ZN(n5471) );
  NAND2_X1 U7070 ( .A1(n8883), .A2(n8441), .ZN(n7816) );
  NAND2_X1 U7071 ( .A1(n7536), .A2(n7635), .ZN(n5476) );
  NAND2_X1 U7072 ( .A1(n5491), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U7073 ( .A1(n5477), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U7074 ( .A1(n5479), .A2(n5478), .ZN(n8649) );
  NAND2_X1 U7075 ( .A1(n8649), .A2(n5495), .ZN(n5484) );
  INV_X1 U7076 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U7077 ( .A1(n5516), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U7078 ( .A1(n7622), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5480) );
  OAI211_X1 U7079 ( .C1(n8648), .C2(n7626), .A(n5481), .B(n5480), .ZN(n5482)
         );
  INV_X1 U7080 ( .A(n5482), .ZN(n5483) );
  NOR2_X1 U7081 ( .A1(n8877), .A2(n8655), .ZN(n5485) );
  INV_X1 U7082 ( .A(n8877), .ZN(n8445) );
  INV_X1 U7083 ( .A(SI_28_), .ZN(n5489) );
  INV_X1 U7084 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8946) );
  MUX2_X1 U7085 ( .A(n8946), .B(n10062), .S(n4325), .Z(n7606) );
  NAND2_X1 U7086 ( .A1(n8944), .A2(n7635), .ZN(n5493) );
  NAND2_X1 U7087 ( .A1(n5491), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U7088 ( .A1(n8608), .A2(n5495), .ZN(n7630) );
  INV_X1 U7089 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8617) );
  NAND2_X1 U7090 ( .A1(n5516), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U7091 ( .A1(n7622), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5496) );
  OAI211_X1 U7092 ( .C1(n8617), .C2(n7626), .A(n5497), .B(n5496), .ZN(n5498)
         );
  INV_X1 U7093 ( .A(n5498), .ZN(n5499) );
  NAND2_X1 U7094 ( .A1(n8619), .A2(n8460), .ZN(n7835) );
  NAND2_X1 U7095 ( .A1(n7846), .A2(n7835), .ZN(n7643) );
  INV_X1 U7096 ( .A(n5500), .ZN(n5502) );
  NAND2_X1 U7097 ( .A1(n5505), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5504) );
  MUX2_X1 U7098 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5504), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n5507) );
  NAND2_X1 U7099 ( .A1(n5508), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5509) );
  INV_X1 U7100 ( .A(n5510), .ZN(n5511) );
  NAND2_X1 U7101 ( .A1(n5511), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5512) );
  AND2_X1 U7102 ( .A1(n6872), .A2(n6779), .ZN(n5513) );
  INV_X1 U7103 ( .A(n7863), .ZN(n6581) );
  NAND2_X1 U7104 ( .A1(n6581), .A2(n6565), .ZN(n5515) );
  NAND2_X1 U7105 ( .A1(n5117), .A2(n5515), .ZN(n5522) );
  NOR2_X4 U7106 ( .A1(n7309), .A2(n7681), .ZN(n7826) );
  INV_X1 U7107 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7108 ( .A1(n5516), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U7109 ( .A1(n7622), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5517) );
  OAI211_X1 U7110 ( .C1(n5519), .C2(n7626), .A(n5518), .B(n5517), .ZN(n5520)
         );
  INV_X1 U7111 ( .A(n5520), .ZN(n5521) );
  NAND2_X1 U7112 ( .A1(n5117), .A2(P2_B_REG_SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7113 ( .A1(n8771), .A2(n5523), .ZN(n8605) );
  NAND2_X1 U7114 ( .A1(n6871), .A2(n7686), .ZN(n8834) );
  NAND2_X1 U7115 ( .A1(n8834), .A2(n8833), .ZN(n5529) );
  NAND2_X1 U7116 ( .A1(n5529), .A2(n7690), .ZN(n6710) );
  INV_X1 U7117 ( .A(n7647), .ZN(n6709) );
  NAND2_X1 U7118 ( .A1(n6710), .A2(n6709), .ZN(n5530) );
  NAND2_X1 U7119 ( .A1(n5530), .A2(n7709), .ZN(n6848) );
  INV_X1 U7120 ( .A(n7137), .ZN(n6934) );
  NAND2_X1 U7121 ( .A1(n8471), .A2(n6934), .ZN(n7710) );
  NAND2_X1 U7122 ( .A1(n7007), .A2(n7137), .ZN(n7702) );
  NAND2_X1 U7123 ( .A1(n7163), .A2(n7074), .ZN(n7706) );
  INV_X1 U7124 ( .A(n7074), .ZN(n7045) );
  NAND2_X1 U7125 ( .A1(n8469), .A2(n7045), .ZN(n7714) );
  NAND2_X1 U7126 ( .A1(n6962), .A2(n7650), .ZN(n5531) );
  AND2_X1 U7127 ( .A1(n7728), .A2(n7086), .ZN(n7724) );
  NAND2_X1 U7128 ( .A1(n5532), .A2(n7727), .ZN(n7172) );
  INV_X1 U7129 ( .A(n7172), .ZN(n5534) );
  INV_X1 U7130 ( .A(n8466), .ZN(n7215) );
  NAND2_X1 U7131 ( .A1(n7215), .A2(n7239), .ZN(n7736) );
  INV_X1 U7132 ( .A(n7239), .ZN(n7233) );
  NAND2_X1 U7133 ( .A1(n8466), .A2(n7233), .ZN(n7731) );
  NAND2_X1 U7134 ( .A1(n7736), .A2(n7731), .ZN(n7653) );
  INV_X1 U7135 ( .A(n8309), .ZN(n7268) );
  NAND2_X1 U7136 ( .A1(n7268), .A2(n9944), .ZN(n7740) );
  AND2_X1 U7137 ( .A1(n7740), .A2(n7731), .ZN(n7739) );
  NAND2_X1 U7138 ( .A1(n7409), .A2(n8309), .ZN(n7737) );
  AND2_X1 U7139 ( .A1(n7752), .A2(n7737), .ZN(n7743) );
  NAND2_X1 U7140 ( .A1(n7415), .A2(n9951), .ZN(n7758) );
  NAND2_X1 U7141 ( .A1(n7420), .A2(n7263), .ZN(n7755) );
  NAND2_X1 U7142 ( .A1(n7348), .A2(n7656), .ZN(n5535) );
  NAND2_X1 U7143 ( .A1(n5535), .A2(n7758), .ZN(n7286) );
  NAND2_X1 U7144 ( .A1(n8408), .A2(n8238), .ZN(n7750) );
  NAND2_X1 U7145 ( .A1(n7286), .A2(n7750), .ZN(n5536) );
  NAND2_X1 U7146 ( .A1(n5536), .A2(n7751), .ZN(n7373) );
  INV_X1 U7147 ( .A(n8464), .ZN(n8402) );
  NAND2_X1 U7148 ( .A1(n8286), .A2(n8402), .ZN(n7772) );
  NAND2_X1 U7149 ( .A1(n7373), .A2(n7772), .ZN(n5537) );
  NOR2_X1 U7150 ( .A1(n8243), .A2(n7507), .ZN(n7770) );
  NAND2_X1 U7151 ( .A1(n8243), .A2(n7507), .ZN(n7769) );
  INV_X1 U7152 ( .A(n7777), .ZN(n5538) );
  INV_X1 U7153 ( .A(n7785), .ZN(n5539) );
  NAND2_X1 U7154 ( .A1(n8921), .A2(n8365), .ZN(n7786) );
  AND2_X1 U7155 ( .A1(n7783), .A2(n8724), .ZN(n7787) );
  NAND2_X1 U7156 ( .A1(n8713), .A2(n7794), .ZN(n8708) );
  AND2_X1 U7157 ( .A1(n7801), .A2(n8707), .ZN(n7795) );
  INV_X1 U7158 ( .A(n7805), .ZN(n5541) );
  NAND2_X1 U7159 ( .A1(n8675), .A2(n7811), .ZN(n8664) );
  NAND2_X1 U7160 ( .A1(n8889), .A2(n8680), .ZN(n7812) );
  NAND2_X1 U7161 ( .A1(n8804), .A2(n8382), .ZN(n8663) );
  NAND3_X1 U7162 ( .A1(n8664), .A2(n7812), .A3(n8663), .ZN(n5542) );
  NAND2_X1 U7163 ( .A1(n5542), .A2(n7813), .ZN(n8652) );
  INV_X1 U7164 ( .A(n7815), .ZN(n5543) );
  NAND2_X1 U7165 ( .A1(n8791), .A2(n5544), .ZN(n7644) );
  NOR2_X1 U7166 ( .A1(n8791), .A2(n5544), .ZN(n7827) );
  NOR2_X1 U7167 ( .A1(n5545), .A2(n8461), .ZN(n5546) );
  INV_X1 U7168 ( .A(n8592), .ZN(n7131) );
  AOI21_X1 U7169 ( .B1(n7309), .B2(n6779), .A(n8592), .ZN(n5547) );
  AND2_X1 U7170 ( .A1(n8847), .A2(n5547), .ZN(n5548) );
  NAND2_X1 U7171 ( .A1(n7279), .A2(n5548), .ZN(n7178) );
  NOR2_X1 U7172 ( .A1(n8615), .A2(n5549), .ZN(n8224) );
  XNOR2_X1 U7173 ( .A(n7913), .B(P2_B_REG_SCAN_IN), .ZN(n5558) );
  AND2_X1 U7174 ( .A1(n5560), .A2(n5559), .ZN(n5561) );
  NAND2_X1 U7175 ( .A1(n5562), .A2(n5561), .ZN(n5563) );
  NAND2_X1 U7176 ( .A1(n5563), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5564) );
  MUX2_X1 U7177 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5564), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5566) );
  NAND2_X1 U7178 ( .A1(n7535), .A2(n7541), .ZN(n5569) );
  NAND2_X1 U7179 ( .A1(n7913), .A2(n7541), .ZN(n5571) );
  NAND3_X1 U7180 ( .A1(n7865), .A2(n6779), .A3(n7131), .ZN(n5572) );
  NAND2_X1 U7181 ( .A1(n5572), .A2(n7847), .ZN(n5573) );
  MUX2_X1 U7182 ( .A(n6753), .B(n6778), .S(n5573), .Z(n6817) );
  NOR4_X1 U7183 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n5582) );
  NOR4_X1 U7184 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5577) );
  NOR4_X1 U7185 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n5576) );
  NOR4_X1 U7186 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n5575) );
  NOR4_X1 U7187 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5574) );
  NAND4_X1 U7188 ( .A1(n5577), .A2(n5576), .A3(n5575), .A4(n5574), .ZN(n5578)
         );
  NOR4_X1 U7189 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        n5579), .A4(n5578), .ZN(n5581) );
  NOR4_X1 U7190 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5580) );
  AND3_X1 U7191 ( .A1(n5582), .A2(n5581), .A3(n5580), .ZN(n5583) );
  INV_X1 U7192 ( .A(n7856), .ZN(n5586) );
  NAND2_X1 U7193 ( .A1(n7826), .A2(n5586), .ZN(n6756) );
  NAND3_X1 U7194 ( .A1(n6754), .A2(n6770), .A3(n6756), .ZN(n6818) );
  NOR2_X1 U7195 ( .A1(n6818), .A2(n6769), .ZN(n5587) );
  NAND2_X1 U7196 ( .A1(n6778), .A2(n6753), .ZN(n6759) );
  OR2_X1 U7197 ( .A1(n8224), .A2(n8857), .ZN(n5591) );
  INV_X1 U7198 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5588) );
  NOR2_X1 U7199 ( .A1(n8827), .A2(n5588), .ZN(n5589) );
  NAND2_X1 U7200 ( .A1(n5591), .A2(n5590), .ZN(P2_U3488) );
  NOR2_X1 U7201 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5594) );
  NOR2_X1 U7202 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5593) );
  NOR2_X1 U7203 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5602) );
  NOR2_X1 U7204 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5601) );
  NOR2_X1 U7205 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5600) );
  NAND2_X1 U7206 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n5608) );
  NAND2_X1 U7207 ( .A1(n5620), .A2(n5608), .ZN(n5609) );
  XNOR2_X2 U7208 ( .A(n5609), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6354) );
  OR2_X1 U7209 ( .A1(n6303), .A2(n5703), .ZN(n5614) );
  NOR2_X1 U7210 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5751) );
  INV_X1 U7211 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5719) );
  OAI21_X1 U7212 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(P1_IR_REG_2__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5610) );
  AND2_X1 U7213 ( .A1(n5705), .A2(n5610), .ZN(n5738) );
  INV_X1 U7214 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7215 ( .A1(n5738), .A2(n5611), .ZN(n5741) );
  NAND2_X1 U7216 ( .A1(n5741), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5612) );
  XNOR2_X1 U7217 ( .A(n5612), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6379) );
  AOI22_X1 U7218 ( .A1(n5989), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6322), .B2(
        n6379), .ZN(n5613) );
  INV_X1 U7219 ( .A(n6520), .ZN(n6990) );
  NAND2_X1 U7220 ( .A1(n4810), .A2(n5616), .ZN(n5651) );
  NOR2_X2 U7221 ( .A1(n5651), .A2(n4895), .ZN(n5626) );
  XNOR2_X1 U7222 ( .A(n5619), .B(n4716), .ZN(n6132) );
  INV_X1 U7223 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U7224 ( .A1(n4385), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U7225 ( .A1(n5630), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5625) );
  INV_X1 U7226 ( .A(n5626), .ZN(n5627) );
  NAND2_X1 U7227 ( .A1(n5627), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5628) );
  MUX2_X1 U7228 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5628), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5629) );
  INV_X1 U7229 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5634) );
  XNOR2_X1 U7230 ( .A(n5635), .B(n5634), .ZN(n5640) );
  INV_X1 U7231 ( .A(n5640), .ZN(n5641) );
  NAND2_X1 U7232 ( .A1(n5637), .A2(n5636), .ZN(n5638) );
  NAND2_X1 U7233 ( .A1(n5696), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U7234 ( .A1(n5699), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U7235 ( .A1(n5642), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5757) );
  INV_X1 U7236 ( .A(n5642), .ZN(n5732) );
  INV_X1 U7237 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5643) );
  NAND2_X1 U7238 ( .A1(n5732), .A2(n5643), .ZN(n5644) );
  AND2_X1 U7239 ( .A1(n5757), .A2(n5644), .ZN(n6895) );
  NAND2_X1 U7240 ( .A1(n6180), .A2(n6895), .ZN(n5647) );
  NAND2_X1 U7241 ( .A1(n4333), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5646) );
  AND2_X1 U7242 ( .A1(n5970), .A2(n5650), .ZN(n5652) );
  NAND2_X1 U7243 ( .A1(n5657), .A2(n5656), .ZN(n6148) );
  OAI22_X1 U7244 ( .A1(n6990), .A2(n6098), .B1(n6542), .B2(n5673), .ZN(n6889)
         );
  NAND2_X1 U7245 ( .A1(n5696), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U7246 ( .A1(n4328), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7247 ( .A1(n5713), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7248 ( .A1(n5699), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5660) );
  NAND4_X2 U7249 ( .A1(n5663), .A2(n5662), .A3(n5661), .A4(n5660), .ZN(n9109)
         );
  NAND2_X1 U7250 ( .A1(n9109), .A2(n5695), .ZN(n5667) );
  INV_X1 U7251 ( .A(n6514), .ZN(n5664) );
  INV_X1 U7252 ( .A(n6297), .ZN(n5666) );
  INV_X1 U7253 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6309) );
  INV_X1 U7254 ( .A(n9109), .ZN(n6503) );
  OAI22_X1 U7255 ( .A1(n6503), .A2(n5673), .B1(n8110), .B2(n6098), .ZN(n5668)
         );
  INV_X1 U7256 ( .A(n5668), .ZN(n5692) );
  XNOR2_X1 U7257 ( .A(n5691), .B(n5692), .ZN(n7872) );
  NAND2_X1 U7258 ( .A1(n5699), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U7259 ( .A1(n4333), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U7260 ( .A1(n5696), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5669) );
  NAND4_X2 U7261 ( .A1(n5672), .A2(n5671), .A3(n5670), .A4(n5669), .ZN(n9110)
         );
  NAND2_X1 U7262 ( .A1(n9110), .A2(n6049), .ZN(n5683) );
  NAND2_X1 U7263 ( .A1(n4325), .A2(SI_0_), .ZN(n5676) );
  INV_X1 U7264 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5675) );
  NAND2_X1 U7265 ( .A1(n5676), .A2(n5675), .ZN(n5678) );
  NAND2_X1 U7266 ( .A1(n5678), .A2(n5677), .ZN(n6295) );
  MUX2_X1 U7267 ( .A(n5674), .B(n6295), .S(n5724), .Z(n7592) );
  INV_X1 U7268 ( .A(n7592), .ZN(n5681) );
  INV_X1 U7269 ( .A(n5679), .ZN(n5680) );
  NAND2_X1 U7270 ( .A1(n5683), .A2(n5682), .ZN(n6399) );
  NAND2_X1 U7271 ( .A1(n9110), .A2(n5695), .ZN(n5685) );
  NAND2_X1 U7272 ( .A1(n5727), .A2(n5681), .ZN(n5684) );
  AND2_X1 U7273 ( .A1(n5685), .A2(n5684), .ZN(n5688) );
  NAND2_X1 U7274 ( .A1(n5680), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U7275 ( .A1(n6399), .A2(n6400), .ZN(n5690) );
  NAND2_X1 U7276 ( .A1(n5688), .A2(n6167), .ZN(n5689) );
  AND2_X1 U7277 ( .A1(n5690), .A2(n5689), .ZN(n7874) );
  NAND2_X1 U7278 ( .A1(n7872), .A2(n7874), .ZN(n7873) );
  INV_X1 U7279 ( .A(n5691), .ZN(n5693) );
  NAND2_X1 U7280 ( .A1(n4333), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U7281 ( .A1(n4328), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5698) );
  NAND2_X1 U7282 ( .A1(n5696), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U7283 ( .A1(n5699), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7284 ( .A1(n5705), .A2(n5704), .ZN(n5718) );
  OR2_X1 U7285 ( .A1(n5724), .A2(n6358), .ZN(n5706) );
  AOI22_X1 U7286 ( .A1(n5695), .A2(n6213), .B1(n6505), .B2(n5727), .ZN(n5707)
         );
  XNOR2_X1 U7287 ( .A(n5707), .B(n5930), .ZN(n5712) );
  NAND2_X1 U7288 ( .A1(n6213), .A2(n6049), .ZN(n5709) );
  XNOR2_X1 U7289 ( .A(n5712), .B(n5710), .ZN(n6470) );
  INV_X1 U7290 ( .A(n5710), .ZN(n5711) );
  NAND2_X1 U7291 ( .A1(n5699), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5717) );
  INV_X1 U7292 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6649) );
  NAND2_X1 U7293 ( .A1(n4328), .A2(n6649), .ZN(n5716) );
  NAND2_X1 U7294 ( .A1(n4333), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U7295 ( .A1(n5696), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5714) );
  OR2_X1 U7296 ( .A1(n6216), .A2(n5673), .ZN(n5726) );
  NAND2_X1 U7297 ( .A1(n5718), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5720) );
  OR2_X1 U7298 ( .A1(n5721), .A2(n6313), .ZN(n5722) );
  NAND2_X1 U7299 ( .A1(n5695), .A2(n6215), .ZN(n5725) );
  NAND2_X1 U7300 ( .A1(n5726), .A2(n5725), .ZN(n5730) );
  XNOR2_X1 U7301 ( .A(n5728), .B(n5930), .ZN(n5729) );
  INV_X1 U7302 ( .A(n5729), .ZN(n5731) );
  NAND2_X1 U7303 ( .A1(n5696), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5737) );
  NAND2_X1 U7304 ( .A1(n5699), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5736) );
  OAI21_X1 U7305 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5732), .ZN(n5733) );
  INV_X1 U7306 ( .A(n5733), .ZN(n6749) );
  NAND2_X1 U7307 ( .A1(n6180), .A2(n6749), .ZN(n5735) );
  NAND2_X1 U7308 ( .A1(n4332), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5734) );
  INV_X1 U7309 ( .A(n5738), .ZN(n5739) );
  NAND2_X1 U7310 ( .A1(n5739), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5740) );
  AOI22_X1 U7311 ( .A1(n5989), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6322), .B2(
        n6366), .ZN(n5742) );
  AOI22_X1 U7312 ( .A1(n9107), .A2(n6066), .B1(n6741), .B2(n5786), .ZN(n5743)
         );
  XNOR2_X1 U7313 ( .A(n5743), .B(n5930), .ZN(n5745) );
  INV_X2 U7314 ( .A(n6741), .ZN(n9626) );
  OAI22_X1 U7315 ( .A1(n6555), .A2(n5673), .B1(n9626), .B2(n6098), .ZN(n5746)
         );
  INV_X1 U7316 ( .A(n5745), .ZN(n5747) );
  OAI22_X1 U7317 ( .A1(n6990), .A2(n6081), .B1(n6542), .B2(n6098), .ZN(n5748)
         );
  XOR2_X1 U7318 ( .A(n5930), .B(n5748), .Z(n5749) );
  NOR2_X1 U7319 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5750) );
  NAND3_X1 U7320 ( .A1(n5752), .A2(n5751), .A3(n5750), .ZN(n5770) );
  NAND2_X1 U7321 ( .A1(n5770), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5753) );
  XNOR2_X1 U7322 ( .A(n5753), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6422) );
  AOI22_X1 U7323 ( .A1(n5989), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6322), .B2(
        n6422), .ZN(n5754) );
  NAND2_X1 U7324 ( .A1(n7112), .A2(n5786), .ZN(n5764) );
  NAND2_X1 U7325 ( .A1(n5699), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U7326 ( .A1(n5696), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5761) );
  NOR2_X1 U7327 ( .A1(n5757), .A2(n5756), .ZN(n5774) );
  INV_X1 U7328 ( .A(n5774), .ZN(n5775) );
  NAND2_X1 U7329 ( .A1(n5757), .A2(n5756), .ZN(n5758) );
  AND2_X1 U7330 ( .A1(n5775), .A2(n5758), .ZN(n7123) );
  NAND2_X1 U7331 ( .A1(n6180), .A2(n7123), .ZN(n5760) );
  NAND2_X1 U7332 ( .A1(n4332), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5759) );
  OR2_X1 U7333 ( .A1(n6892), .A2(n6098), .ZN(n5763) );
  NAND2_X1 U7334 ( .A1(n5764), .A2(n5763), .ZN(n5765) );
  XNOR2_X1 U7335 ( .A(n5765), .B(n6167), .ZN(n7118) );
  NOR2_X1 U7336 ( .A1(n6892), .A2(n5673), .ZN(n5766) );
  AOI21_X1 U7337 ( .B1(n7112), .B2(n5695), .A(n5766), .ZN(n7117) );
  INV_X1 U7338 ( .A(n7118), .ZN(n5768) );
  INV_X1 U7339 ( .A(n7117), .ZN(n5767) );
  NAND2_X1 U7340 ( .A1(n5768), .A2(n5767), .ZN(n5769) );
  OR2_X1 U7341 ( .A1(n6318), .A2(n5703), .ZN(n5773) );
  NAND2_X1 U7342 ( .A1(n5896), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5771) );
  XNOR2_X1 U7343 ( .A(n5771), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6491) );
  AOI22_X1 U7344 ( .A1(n5989), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6322), .B2(
        n6491), .ZN(n5772) );
  NAND2_X1 U7345 ( .A1(n5696), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U7346 ( .A1(n5699), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U7347 ( .A1(n5774), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5788) );
  INV_X1 U7348 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10026) );
  NAND2_X1 U7349 ( .A1(n5775), .A2(n10026), .ZN(n5776) );
  AND2_X1 U7350 ( .A1(n5788), .A2(n5776), .ZN(n7101) );
  NAND2_X1 U7351 ( .A1(n6180), .A2(n7101), .ZN(n5778) );
  NAND2_X1 U7352 ( .A1(n4333), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5777) );
  AOI22_X1 U7353 ( .A1(n7107), .A2(n5786), .B1(n5695), .B2(n9104), .ZN(n5781)
         );
  XOR2_X1 U7354 ( .A(n5930), .B(n5781), .Z(n5783) );
  INV_X1 U7355 ( .A(n7107), .ZN(n6958) );
  OAI22_X1 U7356 ( .A1(n6958), .A2(n6098), .B1(n7115), .B2(n5673), .ZN(n5782)
         );
  NAND2_X1 U7357 ( .A1(n5783), .A2(n5782), .ZN(n7099) );
  INV_X1 U7358 ( .A(n5798), .ZN(n5800) );
  NOR2_X1 U7359 ( .A1(n5896), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5821) );
  OR2_X1 U7360 ( .A1(n5821), .A2(n9484), .ZN(n5802) );
  XNOR2_X1 U7361 ( .A(n5802), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6626) );
  AOI22_X1 U7362 ( .A1(n5989), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6322), .B2(
        n6626), .ZN(n5784) );
  NAND2_X1 U7363 ( .A1(n5785), .A2(n5784), .ZN(n7061) );
  NAND2_X1 U7364 ( .A1(n7061), .A2(n5786), .ZN(n5795) );
  NAND2_X1 U7365 ( .A1(n5699), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7366 ( .A1(n4332), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U7367 ( .A1(n5788), .A2(n5787), .ZN(n5789) );
  AND2_X1 U7368 ( .A1(n5809), .A2(n5789), .ZN(n7198) );
  NAND2_X1 U7369 ( .A1(n6180), .A2(n7198), .ZN(n5791) );
  NAND2_X1 U7370 ( .A1(n5696), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5790) );
  OR2_X1 U7371 ( .A1(n7105), .A2(n6098), .ZN(n5794) );
  NAND2_X1 U7372 ( .A1(n5795), .A2(n5794), .ZN(n5796) );
  XNOR2_X1 U7373 ( .A(n5796), .B(n5930), .ZN(n5797) );
  INV_X1 U7374 ( .A(n5797), .ZN(n5799) );
  XNOR2_X1 U7375 ( .A(n5798), .B(n5797), .ZN(n7192) );
  INV_X1 U7376 ( .A(n7061), .ZN(n7195) );
  OAI22_X1 U7377 ( .A1(n7195), .A2(n6098), .B1(n7105), .B2(n5673), .ZN(n7191)
         );
  NAND2_X1 U7378 ( .A1(n6336), .A2(n7899), .ZN(n5806) );
  NAND2_X1 U7379 ( .A1(n5802), .A2(n5801), .ZN(n5803) );
  NAND2_X1 U7380 ( .A1(n5803), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5804) );
  XNOR2_X1 U7381 ( .A(n5804), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9141) );
  AOI22_X1 U7382 ( .A1(n5989), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6322), .B2(
        n9141), .ZN(n5805) );
  NAND2_X1 U7383 ( .A1(n5806), .A2(n5805), .ZN(n7024) );
  NAND2_X1 U7384 ( .A1(n7024), .A2(n5786), .ZN(n5816) );
  NAND2_X1 U7385 ( .A1(n5699), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7386 ( .A1(n4333), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5813) );
  INV_X1 U7388 ( .A(n5828), .ZN(n5841) );
  NAND2_X1 U7389 ( .A1(n5809), .A2(n5808), .ZN(n5810) );
  AND2_X1 U7390 ( .A1(n5841), .A2(n5810), .ZN(n7298) );
  NAND2_X1 U7391 ( .A1(n6180), .A2(n7298), .ZN(n5812) );
  NAND2_X1 U7392 ( .A1(n5696), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5811) );
  OR2_X1 U7393 ( .A1(n7454), .A2(n6098), .ZN(n5815) );
  NAND2_X1 U7394 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  XNOR2_X1 U7395 ( .A(n5817), .B(n5930), .ZN(n5819) );
  INV_X1 U7396 ( .A(n7024), .ZN(n9638) );
  OAI22_X1 U7397 ( .A1(n9638), .A2(n6098), .B1(n7454), .B2(n5673), .ZN(n5818)
         );
  XNOR2_X1 U7398 ( .A(n5819), .B(n5818), .ZN(n7293) );
  NAND2_X1 U7399 ( .A1(n6438), .A2(n7899), .ZN(n5824) );
  NOR2_X1 U7400 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5820) );
  NAND2_X1 U7401 ( .A1(n5821), .A2(n5820), .ZN(n5837) );
  NAND2_X1 U7402 ( .A1(n5857), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5822) );
  XNOR2_X1 U7403 ( .A(n5822), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9520) );
  AOI22_X1 U7404 ( .A1(n5989), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6322), .B2(
        n9520), .ZN(n5823) );
  NAND2_X1 U7405 ( .A1(n7484), .A2(n5786), .ZN(n5835) );
  NAND2_X1 U7406 ( .A1(n5696), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7407 ( .A1(n5699), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5832) );
  INV_X1 U7408 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5826) );
  INV_X1 U7409 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5825) );
  OAI21_X1 U7410 ( .B1(n5841), .B2(n5826), .A(n5825), .ZN(n5829) );
  INV_X1 U7411 ( .A(n5861), .ZN(n5862) );
  AND2_X1 U7412 ( .A1(n5829), .A2(n5862), .ZN(n9050) );
  NAND2_X1 U7413 ( .A1(n6180), .A2(n9050), .ZN(n5831) );
  NAND2_X1 U7414 ( .A1(n4332), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5830) );
  OR2_X1 U7415 ( .A1(n7391), .A2(n6098), .ZN(n5834) );
  NAND2_X1 U7416 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  XNOR2_X1 U7417 ( .A(n5836), .B(n5930), .ZN(n9042) );
  INV_X1 U7418 ( .A(n7391), .ZN(n9100) );
  AOI22_X1 U7419 ( .A1(n7484), .A2(n6066), .B1(n6049), .B2(n9100), .ZN(n9041)
         );
  INV_X1 U7420 ( .A(n9041), .ZN(n5850) );
  NAND2_X1 U7421 ( .A1(n6338), .A2(n7899), .ZN(n5840) );
  NAND2_X1 U7422 ( .A1(n5837), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5838) );
  XNOR2_X1 U7423 ( .A(n5838), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9502) );
  AOI22_X1 U7424 ( .A1(n5989), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6322), .B2(
        n9502), .ZN(n5839) );
  NAND2_X1 U7425 ( .A1(n5840), .A2(n5839), .ZN(n6277) );
  NAND2_X1 U7426 ( .A1(n5699), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U7427 ( .A1(n5696), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5844) );
  XNOR2_X1 U7428 ( .A(n5841), .B(P1_REG3_REG_10__SCAN_IN), .ZN(n7457) );
  NAND2_X1 U7429 ( .A1(n6180), .A2(n7457), .ZN(n5843) );
  NAND2_X1 U7430 ( .A1(n4333), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5842) );
  NOR2_X1 U7431 ( .A1(n9046), .A2(n5673), .ZN(n5846) );
  AOI21_X1 U7432 ( .B1(n6277), .B2(n6066), .A(n5846), .ZN(n5851) );
  INV_X1 U7433 ( .A(n5851), .ZN(n7451) );
  NAND2_X1 U7434 ( .A1(n6277), .A2(n5786), .ZN(n5848) );
  OR2_X1 U7435 ( .A1(n9046), .A2(n6098), .ZN(n5847) );
  NAND2_X1 U7436 ( .A1(n5848), .A2(n5847), .ZN(n5849) );
  XNOR2_X1 U7437 ( .A(n5849), .B(n6167), .ZN(n9040) );
  INV_X1 U7438 ( .A(n9040), .ZN(n5853) );
  AOI22_X1 U7439 ( .A1(n9042), .A2(n5850), .B1(n7451), .B2(n5853), .ZN(n5856)
         );
  AOI21_X1 U7440 ( .B1(n9040), .B2(n5851), .A(n9041), .ZN(n5854) );
  NAND2_X1 U7441 ( .A1(n9041), .A2(n5851), .ZN(n5852) );
  OAI22_X1 U7442 ( .A1(n5854), .A2(n9042), .B1(n5853), .B2(n5852), .ZN(n5855)
         );
  NAND2_X1 U7443 ( .A1(n6475), .A2(n7899), .ZN(n5860) );
  INV_X1 U7444 ( .A(n5857), .ZN(n5858) );
  NAND2_X1 U7445 ( .A1(n5858), .A2(n5897), .ZN(n5894) );
  NAND2_X1 U7446 ( .A1(n5894), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5872) );
  XNOR2_X1 U7447 ( .A(n5872), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9524) );
  AOI22_X1 U7448 ( .A1(n5989), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6322), .B2(
        n9524), .ZN(n5859) );
  NAND2_X1 U7449 ( .A1(n5696), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U7450 ( .A1(n5699), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5866) );
  INV_X1 U7451 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10032) );
  NAND2_X1 U7452 ( .A1(n5862), .A2(n10032), .ZN(n5863) );
  AND2_X1 U7453 ( .A1(n5878), .A2(n5863), .ZN(n7395) );
  NAND2_X1 U7454 ( .A1(n4329), .A2(n7395), .ZN(n5865) );
  NAND2_X1 U7455 ( .A1(n4332), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5864) );
  NAND4_X1 U7456 ( .A1(n5867), .A2(n5866), .A3(n5865), .A4(n5864), .ZN(n9099)
         );
  OAI22_X1 U7457 ( .A1(n7392), .A2(n6098), .B1(n7466), .B2(n5673), .ZN(n5870)
         );
  INV_X1 U7458 ( .A(n7392), .ZN(n7249) );
  AOI22_X1 U7459 ( .A1(n7249), .A2(n5786), .B1(n5695), .B2(n9099), .ZN(n5868)
         );
  XNOR2_X1 U7460 ( .A(n5868), .B(n5930), .ZN(n5869) );
  XOR2_X1 U7461 ( .A(n5870), .B(n5869), .Z(n7389) );
  INV_X1 U7462 ( .A(n5869), .ZN(n5871) );
  NAND2_X1 U7463 ( .A1(n6507), .A2(n7899), .ZN(n5876) );
  NAND2_X1 U7464 ( .A1(n5872), .A2(n5892), .ZN(n5873) );
  NAND2_X1 U7465 ( .A1(n5873), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5874) );
  AOI22_X1 U7466 ( .A1(n6322), .A2(n9549), .B1(n5989), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7467 ( .A1(n7446), .A2(n5786), .ZN(n5885) );
  NAND2_X1 U7468 ( .A1(n5699), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U7469 ( .A1(n4332), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U7470 ( .A1(n5878), .A2(n5877), .ZN(n5879) );
  AND2_X1 U7471 ( .A1(n5905), .A2(n5879), .ZN(n7504) );
  NAND2_X1 U7472 ( .A1(n4328), .A2(n7504), .ZN(n5881) );
  NAND2_X1 U7473 ( .A1(n5696), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5880) );
  OR2_X1 U7474 ( .A1(n8955), .A2(n6098), .ZN(n5884) );
  NAND2_X1 U7475 ( .A1(n5885), .A2(n5884), .ZN(n5886) );
  XNOR2_X1 U7476 ( .A(n5886), .B(n5930), .ZN(n5887) );
  OAI22_X1 U7477 ( .A1(n7501), .A2(n6098), .B1(n8955), .B2(n5673), .ZN(n5888)
         );
  XOR2_X1 U7478 ( .A(n5887), .B(n5888), .Z(n7498) );
  INV_X1 U7479 ( .A(n5887), .ZN(n5890) );
  INV_X1 U7480 ( .A(n5888), .ZN(n5889) );
  NAND2_X1 U7481 ( .A1(n6533), .A2(n7899), .ZN(n5904) );
  INV_X1 U7482 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U7483 ( .A1(n5892), .A2(n5891), .ZN(n5893) );
  OAI21_X1 U7484 ( .B1(n5894), .B2(n5893), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5895) );
  MUX2_X1 U7485 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5895), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5902) );
  INV_X1 U7486 ( .A(n5896), .ZN(n5901) );
  AND3_X1 U7487 ( .A1(n5899), .A2(n5898), .A3(n5897), .ZN(n5900) );
  NAND2_X1 U7488 ( .A1(n5901), .A2(n5900), .ZN(n5933) );
  AOI22_X1 U7489 ( .A1(n5989), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n9562), .B2(
        n6322), .ZN(n5903) );
  NAND2_X1 U7490 ( .A1(n7492), .A2(n5727), .ZN(n5912) );
  NAND2_X1 U7491 ( .A1(n5696), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U7492 ( .A1(n5699), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7493 ( .A1(n5905), .A2(n10071), .ZN(n5906) );
  AND2_X1 U7494 ( .A1(n5938), .A2(n5906), .ZN(n8957) );
  NAND2_X1 U7495 ( .A1(n4328), .A2(n8957), .ZN(n5908) );
  NAND2_X1 U7496 ( .A1(n4333), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5907) );
  OR2_X1 U7497 ( .A1(n9079), .A2(n6098), .ZN(n5911) );
  NAND2_X1 U7498 ( .A1(n5912), .A2(n5911), .ZN(n5913) );
  XNOR2_X1 U7499 ( .A(n5913), .B(n5930), .ZN(n5915) );
  XNOR2_X1 U7500 ( .A(n5914), .B(n5915), .ZN(n8951) );
  INV_X1 U7501 ( .A(n9079), .ZN(n9097) );
  AOI22_X1 U7502 ( .A1(n7492), .A2(n6066), .B1(n6049), .B2(n9097), .ZN(n8952)
         );
  NAND2_X1 U7503 ( .A1(n8951), .A2(n8952), .ZN(n8950) );
  INV_X1 U7504 ( .A(n5915), .ZN(n5916) );
  NAND2_X1 U7505 ( .A1(n6751), .A2(n7899), .ZN(n5920) );
  XNOR2_X1 U7506 ( .A(n5918), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9590) );
  AOI22_X1 U7507 ( .A1(n5989), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6322), .B2(
        n9590), .ZN(n5919) );
  INV_X1 U7508 ( .A(n5921), .ZN(n5940) );
  INV_X1 U7509 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U7510 ( .A1(n5940), .A2(n5922), .ZN(n5923) );
  NAND2_X1 U7511 ( .A1(n5952), .A2(n5923), .ZN(n9004) );
  INV_X1 U7512 ( .A(n4329), .ZN(n6058) );
  OR2_X1 U7513 ( .A1(n9004), .A2(n6058), .ZN(n5928) );
  NAND2_X1 U7514 ( .A1(n5699), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U7515 ( .A1(n5696), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5924) );
  AND2_X1 U7516 ( .A1(n5925), .A2(n5924), .ZN(n5927) );
  NAND2_X1 U7517 ( .A1(n4333), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5926) );
  AOI22_X1 U7518 ( .A1(n9429), .A2(n5786), .B1(n6066), .B2(n9095), .ZN(n5929)
         );
  XOR2_X1 U7519 ( .A(n5930), .B(n5929), .Z(n8998) );
  NAND2_X1 U7520 ( .A1(n9429), .A2(n6066), .ZN(n5932) );
  NAND2_X1 U7521 ( .A1(n9095), .A2(n6049), .ZN(n5931) );
  NAND2_X1 U7522 ( .A1(n5932), .A2(n5931), .ZN(n5966) );
  NAND2_X1 U7523 ( .A1(n6691), .A2(n7899), .ZN(n5936) );
  NAND2_X1 U7524 ( .A1(n5933), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5934) );
  XNOR2_X1 U7525 ( .A(n5934), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9128) );
  AOI22_X1 U7526 ( .A1(n5989), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6322), .B2(
        n9128), .ZN(n5935) );
  NAND2_X1 U7527 ( .A1(n7558), .A2(n6066), .ZN(n5945) );
  NAND2_X1 U7528 ( .A1(n5938), .A2(n5937), .ZN(n5939) );
  AND2_X1 U7529 ( .A1(n5940), .A2(n5939), .ZN(n9085) );
  AOI22_X1 U7530 ( .A1(n9085), .A2(n4328), .B1(n5696), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n5943) );
  AOI22_X1 U7531 ( .A1(n4332), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n5699), .B2(
        P1_REG0_REG_15__SCAN_IN), .ZN(n5942) );
  OR2_X1 U7532 ( .A1(n9001), .A2(n5673), .ZN(n5944) );
  NAND2_X1 U7533 ( .A1(n5945), .A2(n5944), .ZN(n9074) );
  NAND2_X1 U7534 ( .A1(n7558), .A2(n5786), .ZN(n5947) );
  OR2_X1 U7535 ( .A1(n9001), .A2(n6098), .ZN(n5946) );
  NAND2_X1 U7536 ( .A1(n5947), .A2(n5946), .ZN(n5948) );
  XNOR2_X1 U7537 ( .A(n5948), .B(n5930), .ZN(n8995) );
  OAI22_X1 U7538 ( .A1(n8998), .A2(n5966), .B1(n9074), .B2(n8995), .ZN(n9008)
         );
  NAND2_X1 U7539 ( .A1(n6996), .A2(n7899), .ZN(n5950) );
  AOI22_X1 U7540 ( .A1(n5989), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6322), .B2(
        n9600), .ZN(n5949) );
  NAND2_X1 U7541 ( .A1(n9360), .A2(n5786), .ZN(n5958) );
  NAND2_X1 U7542 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  AND2_X1 U7543 ( .A1(n5976), .A2(n5953), .ZN(n9357) );
  NAND2_X1 U7544 ( .A1(n9357), .A2(n4329), .ZN(n5956) );
  AOI22_X1 U7545 ( .A1(n5696), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n5699), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7546 ( .A1(n4333), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5954) );
  OR2_X1 U7547 ( .A1(n6253), .A2(n6098), .ZN(n5957) );
  NAND2_X1 U7548 ( .A1(n5958), .A2(n5957), .ZN(n5959) );
  XNOR2_X1 U7549 ( .A(n5959), .B(n6167), .ZN(n5962) );
  NOR2_X1 U7550 ( .A1(n6253), .A2(n5673), .ZN(n5960) );
  AOI21_X1 U7551 ( .B1(n9360), .B2(n6066), .A(n5960), .ZN(n5961) );
  NOR2_X1 U7552 ( .A1(n5962), .A2(n5961), .ZN(n9012) );
  INV_X1 U7553 ( .A(n9012), .ZN(n5968) );
  NAND2_X1 U7554 ( .A1(n8995), .A2(n9074), .ZN(n5964) );
  INV_X1 U7555 ( .A(n5964), .ZN(n5967) );
  INV_X1 U7556 ( .A(n5966), .ZN(n8997) );
  INV_X1 U7557 ( .A(n8998), .ZN(n5963) );
  AOI21_X1 U7558 ( .B1(n8997), .B2(n5964), .A(n5963), .ZN(n5965) );
  AOI21_X1 U7559 ( .B1(n5967), .B2(n5966), .A(n5965), .ZN(n9009) );
  AND2_X1 U7560 ( .A1(n5968), .A2(n9009), .ZN(n5969) );
  NAND2_X1 U7561 ( .A1(n7000), .A2(n7899), .ZN(n5974) );
  NAND2_X1 U7562 ( .A1(n5971), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5972) );
  XNOR2_X1 U7563 ( .A(n5972), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9150) );
  AOI22_X1 U7564 ( .A1(n5989), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6322), .B2(
        n9150), .ZN(n5973) );
  NAND2_X1 U7565 ( .A1(n9417), .A2(n5727), .ZN(n5982) );
  INV_X1 U7566 ( .A(n5992), .ZN(n5994) );
  NAND2_X1 U7567 ( .A1(n5976), .A2(n5975), .ZN(n5977) );
  NAND2_X1 U7568 ( .A1(n5994), .A2(n5977), .ZN(n9327) );
  OR2_X1 U7569 ( .A1(n9327), .A2(n6058), .ZN(n5980) );
  AOI22_X1 U7570 ( .A1(n5696), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n5699), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7571 ( .A1(n4332), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U7572 ( .A1(n9094), .A2(n6066), .ZN(n5981) );
  NAND2_X1 U7573 ( .A1(n5982), .A2(n5981), .ZN(n5983) );
  XNOR2_X1 U7574 ( .A(n5983), .B(n5687), .ZN(n5984) );
  AOI22_X1 U7575 ( .A1(n9417), .A2(n6066), .B1(n6049), .B2(n9094), .ZN(n9055)
         );
  NAND2_X1 U7576 ( .A1(n9053), .A2(n9055), .ZN(n9054) );
  INV_X1 U7577 ( .A(n5984), .ZN(n5985) );
  NAND2_X1 U7578 ( .A1(n5986), .A2(n5985), .ZN(n5987) );
  NAND2_X1 U7579 ( .A1(n7129), .A2(n7899), .ZN(n5991) );
  AOI22_X1 U7580 ( .A1(n5989), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4331), .B2(
        n6322), .ZN(n5990) );
  NAND2_X1 U7581 ( .A1(n9470), .A2(n5727), .ZN(n6003) );
  INV_X1 U7582 ( .A(n6012), .ZN(n5996) );
  INV_X1 U7583 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7584 ( .A1(n5994), .A2(n5993), .ZN(n5995) );
  NAND2_X1 U7585 ( .A1(n9318), .A2(n4328), .ZN(n6001) );
  INV_X1 U7586 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9154) );
  NAND2_X1 U7587 ( .A1(n5696), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7588 ( .A1(n5699), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5997) );
  OAI211_X1 U7589 ( .C1(n9154), .C2(n6061), .A(n5998), .B(n5997), .ZN(n5999)
         );
  INV_X1 U7590 ( .A(n5999), .ZN(n6000) );
  NAND2_X1 U7591 ( .A1(n9338), .A2(n6066), .ZN(n6002) );
  NAND2_X1 U7592 ( .A1(n6003), .A2(n6002), .ZN(n6004) );
  XNOR2_X1 U7593 ( .A(n6004), .B(n5687), .ZN(n6005) );
  AOI22_X1 U7594 ( .A1(n9470), .A2(n6066), .B1(n6049), .B2(n9338), .ZN(n6006)
         );
  XNOR2_X1 U7595 ( .A(n6005), .B(n6006), .ZN(n8970) );
  INV_X1 U7596 ( .A(n6005), .ZN(n6007) );
  NAND2_X1 U7597 ( .A1(n6007), .A2(n6006), .ZN(n6008) );
  NAND2_X1 U7598 ( .A1(n7183), .A2(n7899), .ZN(n6011) );
  INV_X1 U7599 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7184) );
  OR2_X1 U7600 ( .A1(n5721), .A2(n7184), .ZN(n6010) );
  NAND2_X1 U7601 ( .A1(n9408), .A2(n5727), .ZN(n6020) );
  OR2_X1 U7602 ( .A1(n6012), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6013) );
  AND2_X1 U7603 ( .A1(n6027), .A2(n6013), .ZN(n9303) );
  NAND2_X1 U7604 ( .A1(n9303), .A2(n4328), .ZN(n6018) );
  INV_X1 U7605 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9986) );
  NAND2_X1 U7606 ( .A1(n4332), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7607 ( .A1(n5696), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6014) );
  OAI211_X1 U7608 ( .C1(n5941), .C2(n9986), .A(n6015), .B(n6014), .ZN(n6016)
         );
  INV_X1 U7609 ( .A(n6016), .ZN(n6017) );
  NAND2_X1 U7610 ( .A1(n9093), .A2(n6066), .ZN(n6019) );
  NAND2_X1 U7611 ( .A1(n6020), .A2(n6019), .ZN(n6021) );
  XNOR2_X1 U7612 ( .A(n6021), .B(n5687), .ZN(n9021) );
  NAND2_X1 U7613 ( .A1(n9408), .A2(n6066), .ZN(n6023) );
  NAND2_X1 U7614 ( .A1(n9093), .A2(n6049), .ZN(n6022) );
  NAND2_X1 U7615 ( .A1(n6023), .A2(n6022), .ZN(n9020) );
  NOR2_X1 U7616 ( .A1(n9021), .A2(n9020), .ZN(n8977) );
  NAND2_X1 U7617 ( .A1(n7223), .A2(n7899), .ZN(n6025) );
  OR2_X1 U7618 ( .A1(n5721), .A2(n7224), .ZN(n6024) );
  INV_X1 U7619 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U7620 ( .A1(n6027), .A2(n6026), .ZN(n6028) );
  AND2_X1 U7621 ( .A1(n6039), .A2(n6028), .ZN(n9289) );
  NAND2_X1 U7622 ( .A1(n9289), .A2(n4329), .ZN(n6034) );
  INV_X1 U7623 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7624 ( .A1(n5699), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7625 ( .A1(n5696), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6029) );
  OAI211_X1 U7626 ( .C1(n6031), .C2(n6061), .A(n6030), .B(n6029), .ZN(n6032)
         );
  INV_X1 U7627 ( .A(n6032), .ZN(n6033) );
  INV_X1 U7628 ( .A(n9301), .ZN(n9273) );
  AOI22_X1 U7629 ( .A1(n9464), .A2(n5727), .B1(n6066), .B2(n9273), .ZN(n6035)
         );
  XNOR2_X1 U7630 ( .A(n6035), .B(n5687), .ZN(n6045) );
  OAI22_X1 U7631 ( .A1(n9288), .A2(n6098), .B1(n9301), .B2(n5673), .ZN(n6046)
         );
  AND2_X1 U7632 ( .A1(n6045), .A2(n4459), .ZN(n6047) );
  OR2_X1 U7633 ( .A1(n8977), .A2(n6047), .ZN(n6050) );
  NAND2_X1 U7634 ( .A1(n7307), .A2(n7899), .ZN(n6037) );
  OR2_X1 U7635 ( .A1(n5721), .A2(n7312), .ZN(n6036) );
  INV_X1 U7636 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6038) );
  AND2_X1 U7637 ( .A1(n6039), .A2(n6038), .ZN(n6040) );
  NOR2_X1 U7638 ( .A1(n6040), .A2(n6056), .ZN(n9268) );
  INV_X1 U7639 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9966) );
  NAND2_X1 U7640 ( .A1(n5696), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U7641 ( .A1(n4332), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6041) );
  OAI211_X1 U7642 ( .C1(n5941), .C2(n9966), .A(n6042), .B(n6041), .ZN(n6043)
         );
  AOI21_X1 U7643 ( .B1(n9268), .B2(n4329), .A(n6043), .ZN(n9283) );
  INV_X1 U7644 ( .A(n9283), .ZN(n9092) );
  AOI22_X1 U7645 ( .A1(n9398), .A2(n5727), .B1(n5695), .B2(n9092), .ZN(n6044)
         );
  XNOR2_X1 U7646 ( .A(n6044), .B(n5687), .ZN(n6052) );
  NAND2_X1 U7647 ( .A1(n9021), .A2(n9020), .ZN(n8978) );
  OR2_X1 U7648 ( .A1(n6052), .A2(n6051), .ZN(n6048) );
  AOI22_X1 U7649 ( .A1(n9398), .A2(n6066), .B1(n6049), .B2(n9092), .ZN(n9030)
         );
  NAND2_X1 U7650 ( .A1(n7398), .A2(n7899), .ZN(n6055) );
  OR2_X1 U7651 ( .A1(n5721), .A2(n6053), .ZN(n6054) );
  NAND2_X1 U7652 ( .A1(n9458), .A2(n5727), .ZN(n6068) );
  OR2_X1 U7653 ( .A1(n6056), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7654 ( .A1(n6057), .A2(n6075), .ZN(n9257) );
  INV_X1 U7655 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7656 ( .A1(n5696), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7657 ( .A1(n5699), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6059) );
  OAI211_X1 U7658 ( .C1(n6062), .C2(n6061), .A(n6060), .B(n6059), .ZN(n6063)
         );
  INV_X1 U7659 ( .A(n6063), .ZN(n6064) );
  NAND2_X1 U7660 ( .A1(n9274), .A2(n6066), .ZN(n6067) );
  NAND2_X1 U7661 ( .A1(n6068), .A2(n6067), .ZN(n6069) );
  XNOR2_X1 U7662 ( .A(n6069), .B(n6167), .ZN(n6072) );
  NOR2_X1 U7663 ( .A1(n9238), .A2(n5673), .ZN(n6070) );
  AOI21_X1 U7664 ( .B1(n9458), .B2(n6066), .A(n6070), .ZN(n6071) );
  OR2_X1 U7665 ( .A1(n6072), .A2(n6071), .ZN(n8962) );
  NAND2_X1 U7666 ( .A1(n6072), .A2(n6071), .ZN(n8964) );
  NAND2_X1 U7667 ( .A1(n7911), .A2(n7899), .ZN(n6074) );
  OR2_X1 U7668 ( .A1(n5721), .A2(n8222), .ZN(n6073) );
  NAND2_X1 U7669 ( .A1(n5696), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7670 ( .A1(n5699), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6079) );
  INV_X1 U7671 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6076) );
  AOI21_X1 U7672 ( .B1(n6076), .B2(n6075), .A(n6092), .ZN(n9241) );
  NAND2_X1 U7673 ( .A1(n4329), .A2(n9241), .ZN(n6078) );
  NAND2_X1 U7674 ( .A1(n4333), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6077) );
  NAND4_X1 U7675 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n9223)
         );
  OAI22_X1 U7676 ( .A1(n6268), .A2(n6098), .B1(n9251), .B2(n5673), .ZN(n6084)
         );
  OAI22_X1 U7677 ( .A1(n6268), .A2(n6081), .B1(n9251), .B2(n6098), .ZN(n6082)
         );
  XNOR2_X1 U7678 ( .A(n6082), .B(n5687), .ZN(n6083) );
  XOR2_X1 U7679 ( .A(n6084), .B(n6083), .Z(n8183) );
  INV_X1 U7680 ( .A(n6083), .ZN(n6086) );
  INV_X1 U7681 ( .A(n6084), .ZN(n6085) );
  NAND2_X1 U7682 ( .A1(n6086), .A2(n6085), .ZN(n6087) );
  NAND2_X1 U7683 ( .A1(n8181), .A2(n6087), .ZN(n8987) );
  NAND2_X1 U7684 ( .A1(n7530), .A2(n7899), .ZN(n6089) );
  OR2_X1 U7685 ( .A1(n5721), .A2(n7531), .ZN(n6088) );
  NAND2_X1 U7686 ( .A1(n5696), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7687 ( .A1(n5699), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6096) );
  INV_X1 U7688 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6091) );
  INV_X1 U7689 ( .A(n6092), .ZN(n6090) );
  NAND2_X1 U7690 ( .A1(n6091), .A2(n6090), .ZN(n6093) );
  INV_X1 U7691 ( .A(n6109), .ZN(n6110) );
  NAND2_X1 U7692 ( .A1(n4328), .A2(n9229), .ZN(n6095) );
  NAND2_X1 U7693 ( .A1(n4332), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6094) );
  OAI22_X1 U7694 ( .A1(n4571), .A2(n6098), .B1(n9240), .B2(n5673), .ZN(n6103)
         );
  NAND2_X1 U7695 ( .A1(n9449), .A2(n5727), .ZN(n6100) );
  OR2_X1 U7696 ( .A1(n9240), .A2(n6098), .ZN(n6099) );
  NAND2_X1 U7697 ( .A1(n6100), .A2(n6099), .ZN(n6101) );
  XNOR2_X1 U7698 ( .A(n6101), .B(n5687), .ZN(n6102) );
  XOR2_X1 U7699 ( .A(n6103), .B(n6102), .Z(n8988) );
  INV_X1 U7700 ( .A(n6102), .ZN(n6105) );
  INV_X1 U7701 ( .A(n6103), .ZN(n6104) );
  NAND2_X1 U7702 ( .A1(n6105), .A2(n6104), .ZN(n6106) );
  NAND2_X1 U7703 ( .A1(n7536), .A2(n7899), .ZN(n6108) );
  OR2_X1 U7704 ( .A1(n5721), .A2(n7537), .ZN(n6107) );
  NAND2_X1 U7705 ( .A1(n5699), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7706 ( .A1(n4332), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6114) );
  INV_X1 U7707 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9981) );
  NAND2_X1 U7708 ( .A1(n6110), .A2(n9981), .ZN(n6111) );
  NAND2_X1 U7709 ( .A1(n4329), .A2(n9210), .ZN(n6113) );
  NAND2_X1 U7710 ( .A1(n5696), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6112) );
  OAI22_X1 U7711 ( .A1(n9446), .A2(n6098), .B1(n9225), .B2(n5673), .ZN(n6119)
         );
  INV_X1 U7712 ( .A(n9225), .ZN(n9090) );
  AOI22_X1 U7713 ( .A1(n9215), .A2(n5727), .B1(n6066), .B2(n9090), .ZN(n6116)
         );
  XNOR2_X1 U7714 ( .A(n6116), .B(n5687), .ZN(n6118) );
  XOR2_X1 U7715 ( .A(n6119), .B(n6118), .Z(n9064) );
  INV_X1 U7716 ( .A(n9064), .ZN(n6117) );
  INV_X1 U7717 ( .A(n6118), .ZN(n6120) );
  NAND2_X1 U7718 ( .A1(n6120), .A2(n6119), .ZN(n6121) );
  NAND2_X1 U7719 ( .A1(n7563), .A2(n7899), .ZN(n6123) );
  OR2_X1 U7720 ( .A1(n5721), .A2(n7582), .ZN(n6122) );
  NAND2_X1 U7721 ( .A1(n5696), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7722 ( .A1(n5699), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6126) );
  XNOR2_X1 U7723 ( .A(n6159), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n7595) );
  NAND2_X1 U7724 ( .A1(n6180), .A2(n7595), .ZN(n6125) );
  NAND2_X1 U7725 ( .A1(n4333), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6124) );
  NOR2_X1 U7726 ( .A1(n9202), .A2(n5673), .ZN(n6128) );
  AOI21_X1 U7727 ( .B1(n7596), .B2(n6066), .A(n6128), .ZN(n6172) );
  NAND2_X1 U7728 ( .A1(n7596), .A2(n5727), .ZN(n6130) );
  OR2_X1 U7729 ( .A1(n9202), .A2(n6098), .ZN(n6129) );
  NAND2_X1 U7730 ( .A1(n6130), .A2(n6129), .ZN(n6131) );
  XNOR2_X1 U7731 ( .A(n6131), .B(n5687), .ZN(n6174) );
  NAND2_X1 U7732 ( .A1(n7532), .A2(P1_B_REG_SCAN_IN), .ZN(n6133) );
  MUX2_X1 U7733 ( .A(P1_B_REG_SCAN_IN), .B(n6133), .S(n6132), .Z(n6135) );
  INV_X1 U7734 ( .A(n7538), .ZN(n6134) );
  NAND2_X1 U7735 ( .A1(n6132), .A2(n7538), .ZN(n9482) );
  NAND2_X1 U7736 ( .A1(n7538), .A2(n7532), .ZN(n6315) );
  NOR4_X1 U7737 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6146) );
  NOR4_X1 U7738 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6145) );
  OR4_X1 U7739 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6143) );
  NOR4_X1 U7740 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6141) );
  NOR4_X1 U7741 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6140) );
  NOR4_X1 U7742 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6139) );
  NOR4_X1 U7743 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6138) );
  NAND4_X1 U7744 ( .A1(n6141), .A2(n6140), .A3(n6139), .A4(n6138), .ZN(n6142)
         );
  NOR4_X1 U7745 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6143), .A4(n6142), .ZN(n6144) );
  AND3_X1 U7746 ( .A1(n6146), .A2(n6145), .A3(n6144), .ZN(n6147) );
  NAND2_X1 U7747 ( .A1(n6148), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7748 ( .A1(n6151), .A2(n6152), .ZN(n7935) );
  INV_X1 U7749 ( .A(n6250), .ZN(n6153) );
  NAND2_X1 U7750 ( .A1(n7584), .A2(n6153), .ZN(n9645) );
  AND3_X1 U7751 ( .A1(n6320), .A2(n7935), .A3(n9645), .ZN(n6154) );
  NAND2_X1 U7752 ( .A1(n7565), .A2(n7899), .ZN(n6156) );
  OR2_X1 U7753 ( .A1(n5721), .A2(n7580), .ZN(n6155) );
  NAND2_X1 U7754 ( .A1(n9373), .A2(n5727), .ZN(n6166) );
  NAND2_X1 U7755 ( .A1(n5696), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7756 ( .A1(n5699), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7757 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6157) );
  NOR2_X1 U7758 ( .A1(n6159), .A2(n6157), .ZN(n6179) );
  INV_X1 U7759 ( .A(n6179), .ZN(n8210) );
  INV_X1 U7760 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6205) );
  INV_X1 U7761 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6158) );
  OAI21_X1 U7762 ( .B1(n6159), .B2(n6205), .A(n6158), .ZN(n6160) );
  NAND2_X1 U7763 ( .A1(n4328), .A2(n9192), .ZN(n6162) );
  NAND2_X1 U7764 ( .A1(n4333), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6161) );
  OR2_X1 U7765 ( .A1(n8196), .A2(n6098), .ZN(n6165) );
  NAND2_X1 U7766 ( .A1(n6166), .A2(n6165), .ZN(n6168) );
  XNOR2_X1 U7767 ( .A(n6168), .B(n6167), .ZN(n6171) );
  NOR2_X1 U7768 ( .A1(n8196), .A2(n5673), .ZN(n6169) );
  AOI21_X1 U7769 ( .B1(n9373), .B2(n6066), .A(n6169), .ZN(n6170) );
  XNOR2_X1 U7770 ( .A(n6171), .B(n6170), .ZN(n6197) );
  INV_X1 U7771 ( .A(n6172), .ZN(n6173) );
  OR2_X1 U7772 ( .A1(n6174), .A2(n6173), .ZN(n6194) );
  NAND4_X1 U7773 ( .A1(n6203), .A2(n9056), .A3(n6197), .A4(n6194), .ZN(n6202)
         );
  INV_X1 U7774 ( .A(n8163), .ZN(n6272) );
  AND2_X1 U7775 ( .A1(n7584), .A2(n6272), .ZN(n6522) );
  AND2_X1 U7776 ( .A1(n6320), .A2(n6522), .ZN(n6175) );
  NAND2_X1 U7777 ( .A1(n6185), .A2(n6175), .ZN(n6176) );
  NAND2_X1 U7778 ( .A1(n6320), .A2(n6250), .ZN(n6246) );
  INV_X1 U7779 ( .A(n4324), .ZN(n6403) );
  NOR2_X1 U7780 ( .A1(n6246), .A2(n9347), .ZN(n8176) );
  NOR2_X1 U7781 ( .A1(n6246), .A2(n9349), .ZN(n6178) );
  NAND2_X1 U7782 ( .A1(n6185), .A2(n6178), .ZN(n9068) );
  NAND2_X1 U7783 ( .A1(n5699), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7784 ( .A1(n4332), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7785 ( .A1(n6180), .A2(n6179), .ZN(n6182) );
  NAND2_X1 U7786 ( .A1(n5696), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6181) );
  INV_X1 U7787 ( .A(n7929), .ZN(n9187) );
  AOI22_X1 U7788 ( .A1(n9076), .A2(n9187), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6193) );
  INV_X1 U7789 ( .A(n6185), .ZN(n6187) );
  INV_X1 U7790 ( .A(n6244), .ZN(n6186) );
  NAND2_X1 U7791 ( .A1(n6187), .A2(n6186), .ZN(n6460) );
  OAI21_X1 U7792 ( .B1(n7935), .B2(n6250), .A(n5679), .ZN(n6188) );
  INV_X1 U7793 ( .A(n6188), .ZN(n6189) );
  AOI21_X1 U7794 ( .B1(n6460), .B2(n6189), .A(P1_U3086), .ZN(n6191) );
  INV_X1 U7795 ( .A(n6323), .ZN(n6190) );
  NAND2_X1 U7796 ( .A1(n6190), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8179) );
  INV_X1 U7797 ( .A(n8179), .ZN(n7399) );
  NAND2_X1 U7798 ( .A1(n9084), .A2(n9192), .ZN(n6192) );
  OAI211_X1 U7799 ( .C1(n9202), .C2(n9078), .A(n6193), .B(n6192), .ZN(n6196)
         );
  NOR3_X1 U7800 ( .A1(n6197), .A2(n4495), .A3(n6194), .ZN(n6195) );
  AOI211_X1 U7801 ( .C1(n9373), .C2(n9035), .A(n6196), .B(n6195), .ZN(n6201)
         );
  INV_X1 U7802 ( .A(n6197), .ZN(n6198) );
  NAND3_X1 U7803 ( .A1(n6202), .A2(n6201), .A3(n6200), .ZN(P1_U3220) );
  NAND2_X1 U7804 ( .A1(n7596), .A2(n9035), .ZN(n6209) );
  NOR2_X1 U7805 ( .A1(n9068), .A2(n8196), .ZN(n6207) );
  OAI22_X1 U7806 ( .A1(n9078), .A2(n9225), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6205), .ZN(n6206) );
  AOI211_X1 U7807 ( .C1(n7595), .C2(n9084), .A(n6207), .B(n6206), .ZN(n6208)
         );
  INV_X1 U7808 ( .A(n6277), .ZN(n9646) );
  NAND2_X1 U7809 ( .A1(n9110), .A2(n5681), .ZN(n6975) );
  NAND2_X1 U7810 ( .A1(n6975), .A2(n6254), .ZN(n6974) );
  NAND2_X1 U7811 ( .A1(n6503), .A2(n8110), .ZN(n6211) );
  NAND2_X1 U7812 ( .A1(n6974), .A2(n6211), .ZN(n6500) );
  NAND2_X1 U7813 ( .A1(n6505), .A2(n7877), .ZN(n6256) );
  NAND2_X1 U7814 ( .A1(n6213), .A2(n6212), .ZN(n8115) );
  NAND2_X1 U7815 ( .A1(n6500), .A2(n6502), .ZN(n6499) );
  NAND2_X1 U7816 ( .A1(n7877), .A2(n6212), .ZN(n6214) );
  NAND2_X1 U7817 ( .A1(n6499), .A2(n6214), .ZN(n6559) );
  NAND2_X1 U7818 ( .A1(n6559), .A2(n7946), .ZN(n6561) );
  OR2_X1 U7819 ( .A1(n9108), .A2(n6215), .ZN(n6217) );
  NAND2_X1 U7820 ( .A1(n6561), .A2(n6217), .ZN(n6536) );
  NAND2_X1 U7821 ( .A1(n9626), .A2(n9107), .ZN(n8121) );
  NAND2_X1 U7822 ( .A1(n6555), .A2(n6741), .ZN(n7990) );
  NAND2_X1 U7823 ( .A1(n6536), .A2(n7944), .ZN(n6535) );
  NAND2_X1 U7824 ( .A1(n9626), .A2(n6555), .ZN(n6218) );
  NAND2_X1 U7825 ( .A1(n6535), .A2(n6218), .ZN(n6510) );
  NAND2_X1 U7826 ( .A1(n6520), .A2(n6542), .ZN(n7991) );
  OR2_X1 U7827 ( .A1(n6542), .A2(n6520), .ZN(n8123) );
  AND2_X1 U7828 ( .A1(n7991), .A2(n8123), .ZN(n6259) );
  NAND2_X1 U7829 ( .A1(n6510), .A2(n7945), .ZN(n6509) );
  INV_X1 U7830 ( .A(n6542), .ZN(n9106) );
  NAND2_X1 U7831 ( .A1(n6990), .A2(n6542), .ZN(n6219) );
  NAND2_X1 U7832 ( .A1(n6509), .A2(n6219), .ZN(n6684) );
  INV_X1 U7833 ( .A(n7112), .ZN(n9632) );
  AND2_X1 U7834 ( .A1(n9632), .A2(n9105), .ZN(n7986) );
  AND2_X1 U7835 ( .A1(n7112), .A2(n6892), .ZN(n7988) );
  OR2_X1 U7836 ( .A1(n7986), .A2(n7988), .ZN(n6683) );
  NAND2_X1 U7837 ( .A1(n6684), .A2(n6683), .ZN(n6682) );
  NAND2_X1 U7838 ( .A1(n9632), .A2(n6892), .ZN(n6220) );
  NAND2_X1 U7839 ( .A1(n6682), .A2(n6220), .ZN(n6839) );
  AND2_X1 U7840 ( .A1(n6958), .A2(n9104), .ZN(n6262) );
  NAND2_X1 U7841 ( .A1(n7107), .A2(n7115), .ZN(n6943) );
  NAND2_X1 U7842 ( .A1(n7995), .A2(n6943), .ZN(n6838) );
  NAND2_X1 U7843 ( .A1(n6958), .A2(n7115), .ZN(n6221) );
  NAND2_X1 U7844 ( .A1(n7061), .A2(n7105), .ZN(n7015) );
  NAND2_X1 U7845 ( .A1(n7996), .A2(n7015), .ZN(n6949) );
  INV_X1 U7846 ( .A(n7105), .ZN(n9103) );
  INV_X1 U7847 ( .A(n8012), .ZN(n6222) );
  AND2_X1 U7848 ( .A1(n7024), .A2(n7454), .ZN(n6263) );
  NAND2_X1 U7849 ( .A1(n7021), .A2(n7020), .ZN(n7019) );
  INV_X1 U7850 ( .A(n7454), .ZN(n9102) );
  OR2_X1 U7851 ( .A1(n6277), .A2(n9046), .ZN(n8005) );
  NAND2_X1 U7852 ( .A1(n6277), .A2(n9046), .ZN(n8010) );
  OR2_X1 U7853 ( .A1(n7484), .A2(n7391), .ZN(n8006) );
  NAND2_X1 U7854 ( .A1(n7484), .A2(n7391), .ZN(n8016) );
  AND2_X2 U7855 ( .A1(n8006), .A2(n8016), .ZN(n7954) );
  NAND2_X1 U7856 ( .A1(n7392), .A2(n9099), .ZN(n8018) );
  NAND2_X1 U7857 ( .A1(n7249), .A2(n7466), .ZN(n8133) );
  OR2_X1 U7858 ( .A1(n7446), .A2(n8955), .ZN(n8137) );
  NAND2_X1 U7859 ( .A1(n7446), .A2(n8955), .ZN(n8134) );
  INV_X1 U7860 ( .A(n9001), .ZN(n9096) );
  NAND2_X1 U7861 ( .A1(n7542), .A2(n6224), .ZN(n6225) );
  NAND2_X1 U7862 ( .A1(n9429), .A2(n9348), .ZN(n8140) );
  NAND2_X1 U7863 ( .A1(n9360), .A2(n9336), .ZN(n6228) );
  NOR2_X1 U7864 ( .A1(n9360), .A2(n9336), .ZN(n6227) );
  INV_X1 U7865 ( .A(n9417), .ZN(n9331) );
  NAND2_X1 U7866 ( .A1(n9331), .A2(n9350), .ZN(n6229) );
  OR2_X1 U7867 ( .A1(n9470), .A2(n9338), .ZN(n7975) );
  NAND2_X1 U7868 ( .A1(n9408), .A2(n9093), .ZN(n6231) );
  NAND2_X1 U7869 ( .A1(n6232), .A2(n6231), .ZN(n9279) );
  NOR2_X1 U7870 ( .A1(n9288), .A2(n9301), .ZN(n6234) );
  NAND2_X1 U7871 ( .A1(n9288), .A2(n9301), .ZN(n6233) );
  OAI21_X1 U7872 ( .B1(n9279), .B2(n6234), .A(n6233), .ZN(n9264) );
  NAND2_X1 U7873 ( .A1(n9398), .A2(n9092), .ZN(n6235) );
  NAND2_X1 U7874 ( .A1(n9264), .A2(n6235), .ZN(n6237) );
  NAND2_X1 U7875 ( .A1(n6278), .A2(n9283), .ZN(n6236) );
  NAND2_X1 U7876 ( .A1(n6237), .A2(n6236), .ZN(n9246) );
  NAND2_X1 U7877 ( .A1(n9458), .A2(n9274), .ZN(n6238) );
  NOR2_X1 U7878 ( .A1(n6268), .A2(n9251), .ZN(n6240) );
  INV_X1 U7879 ( .A(n9240), .ZN(n9091) );
  NOR2_X1 U7880 ( .A1(n9449), .A2(n9091), .ZN(n9204) );
  OR2_X1 U7881 ( .A1(n9204), .A2(n4890), .ZN(n6241) );
  NAND2_X1 U7882 ( .A1(n9449), .A2(n9091), .ZN(n9205) );
  AND2_X1 U7883 ( .A1(n4894), .A2(n9205), .ZN(n6242) );
  NOR2_X1 U7884 ( .A1(n4890), .A2(n6242), .ZN(n6243) );
  NAND2_X1 U7885 ( .A1(n7596), .A2(n9202), .ZN(n9178) );
  XNOR2_X1 U7886 ( .A(n8194), .B(n8191), .ZN(n7603) );
  NOR2_X1 U7887 ( .A1(n6512), .A2(n6244), .ZN(n6248) );
  NAND2_X1 U7888 ( .A1(n6320), .A2(n7935), .ZN(n6245) );
  NAND2_X1 U7889 ( .A1(n6246), .A2(n6245), .ZN(n6459) );
  INV_X1 U7890 ( .A(n6249), .ZN(n6251) );
  INV_X1 U7891 ( .A(n7584), .ZN(n7586) );
  NAND2_X1 U7892 ( .A1(n6324), .A2(n6250), .ZN(n7585) );
  OAI211_X1 U7893 ( .C1(n6251), .C2(n6250), .A(n7586), .B(n7585), .ZN(n7467)
         );
  INV_X1 U7894 ( .A(n6151), .ZN(n7310) );
  NAND2_X1 U7895 ( .A1(n8085), .A2(n8163), .ZN(n7480) );
  OAI22_X1 U7896 ( .A1(n7603), .A2(n9427), .B1(n8192), .B2(n9384), .ZN(n6252)
         );
  INV_X1 U7897 ( .A(n6252), .ZN(n6281) );
  OR2_X1 U7898 ( .A1(n9464), .A2(n9301), .ZN(n8057) );
  NAND2_X1 U7899 ( .A1(n9464), .A2(n9301), .ZN(n8046) );
  OR2_X1 U7900 ( .A1(n9360), .A2(n6253), .ZN(n7941) );
  NAND2_X1 U7901 ( .A1(n9360), .A2(n6253), .ZN(n7940) );
  NAND2_X1 U7902 ( .A1(n7941), .A2(n7940), .ZN(n8040) );
  NAND2_X1 U7903 ( .A1(n6503), .A2(n7888), .ZN(n6255) );
  NAND2_X1 U7904 ( .A1(n6257), .A2(n6256), .ZN(n7978) );
  INV_X1 U7905 ( .A(n7946), .ZN(n6258) );
  NAND2_X1 U7906 ( .A1(n7978), .A2(n6258), .ZN(n6551) );
  NAND2_X1 U7907 ( .A1(n6517), .A2(n7991), .ZN(n6833) );
  INV_X1 U7908 ( .A(n6263), .ZN(n6261) );
  INV_X1 U7909 ( .A(n7988), .ZN(n6260) );
  NAND2_X1 U7910 ( .A1(n7015), .A2(n6943), .ZN(n7997) );
  NAND2_X1 U7911 ( .A1(n7997), .A2(n7996), .ZN(n6264) );
  NAND2_X1 U7912 ( .A1(n8001), .A2(n8012), .ZN(n8129) );
  NAND3_X1 U7913 ( .A1(n7464), .A2(n7954), .A3(n8010), .ZN(n6265) );
  NAND2_X1 U7914 ( .A1(n6265), .A2(n8006), .ZN(n7246) );
  NAND2_X1 U7915 ( .A1(n7431), .A2(n7955), .ZN(n7430) );
  NAND2_X1 U7916 ( .A1(n7430), .A2(n8134), .ZN(n7489) );
  OR2_X1 U7917 ( .A1(n7492), .A2(n9079), .ZN(n8139) );
  NAND2_X1 U7918 ( .A1(n7492), .A2(n9079), .ZN(n8025) );
  NAND2_X1 U7919 ( .A1(n8139), .A2(n8025), .ZN(n7488) );
  OR2_X1 U7920 ( .A1(n7558), .A2(n9001), .ZN(n8142) );
  NAND2_X1 U7921 ( .A1(n7558), .A2(n9001), .ZN(n8035) );
  NAND2_X1 U7922 ( .A1(n8142), .A2(n8035), .ZN(n7957) );
  OR2_X2 U7923 ( .A1(n7545), .A2(n7957), .ZN(n7546) );
  NAND2_X1 U7924 ( .A1(n7546), .A2(n8035), .ZN(n7574) );
  OR2_X1 U7925 ( .A1(n9417), .A2(n9350), .ZN(n8043) );
  NAND2_X1 U7926 ( .A1(n9417), .A2(n9350), .ZN(n8052) );
  NAND2_X1 U7927 ( .A1(n9334), .A2(n9333), .ZN(n9332) );
  NAND2_X1 U7928 ( .A1(n9332), .A2(n8052), .ZN(n9311) );
  OR2_X1 U7929 ( .A1(n9470), .A2(n9298), .ZN(n8044) );
  NAND2_X1 U7930 ( .A1(n9470), .A2(n9298), .ZN(n8150) );
  NAND2_X1 U7931 ( .A1(n9311), .A2(n9312), .ZN(n9310) );
  NAND2_X1 U7932 ( .A1(n9408), .A2(n9313), .ZN(n7972) );
  INV_X1 U7933 ( .A(n7972), .ZN(n6266) );
  OR2_X2 U7934 ( .A1(n9297), .A2(n6266), .ZN(n6267) );
  OR2_X1 U7935 ( .A1(n9408), .A2(n9313), .ZN(n7971) );
  NAND2_X1 U7936 ( .A1(n8046), .A2(n7972), .ZN(n8056) );
  NAND2_X1 U7937 ( .A1(n8056), .A2(n8057), .ZN(n7923) );
  XNOR2_X1 U7938 ( .A(n9398), .B(n9092), .ZN(n9271) );
  NAND2_X1 U7939 ( .A1(n9398), .A2(n9283), .ZN(n7922) );
  NAND2_X1 U7940 ( .A1(n9270), .A2(n7922), .ZN(n9248) );
  AND2_X1 U7941 ( .A1(n6268), .A2(n9223), .ZN(n7918) );
  INV_X1 U7942 ( .A(n6268), .ZN(n6269) );
  INV_X1 U7943 ( .A(n7919), .ZN(n8071) );
  OR2_X1 U7944 ( .A1(n9449), .A2(n9240), .ZN(n8078) );
  NAND2_X1 U7945 ( .A1(n9449), .A2(n9240), .ZN(n8074) );
  NAND2_X1 U7946 ( .A1(n8078), .A2(n8074), .ZN(n7962) );
  NAND2_X1 U7947 ( .A1(n9220), .A2(n8074), .ZN(n9199) );
  NAND2_X1 U7948 ( .A1(n9215), .A2(n9225), .ZN(n8076) );
  NAND2_X1 U7949 ( .A1(n8083), .A2(n8076), .ZN(n7963) );
  NAND2_X1 U7950 ( .A1(n9199), .A2(n9207), .ZN(n9198) );
  NAND2_X1 U7951 ( .A1(n9198), .A2(n8076), .ZN(n6271) );
  OAI21_X1 U7952 ( .B1(n8191), .B2(n6271), .A(n9177), .ZN(n6276) );
  NOR2_X1 U7953 ( .A1(n7310), .A2(n9203), .ZN(n8103) );
  NAND2_X1 U7954 ( .A1(n6152), .A2(n6272), .ZN(n8168) );
  INV_X1 U7955 ( .A(n8168), .ZN(n6273) );
  INV_X1 U7956 ( .A(n8196), .ZN(n9089) );
  NAND2_X1 U7957 ( .A1(n8110), .A2(n7592), .ZN(n6976) );
  NAND2_X1 U7958 ( .A1(n6558), .A2(n9626), .ZN(n6537) );
  NAND2_X1 U7959 ( .A1(n8960), .A2(n7491), .ZN(n7543) );
  NAND2_X1 U7960 ( .A1(n9317), .A2(n9325), .ZN(n9316) );
  OR2_X1 U7961 ( .A1(n9408), .A2(n9316), .ZN(n9286) );
  NOR2_X2 U7962 ( .A1(n9286), .A2(n9464), .ZN(n9265) );
  NOR2_X2 U7963 ( .A1(n9215), .A2(n9228), .ZN(n9197) );
  OAI211_X1 U7964 ( .C1(n8192), .C2(n9197), .A(n9354), .B(n9191), .ZN(n7599)
         );
  MUX2_X1 U7965 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n6286), .S(n9659), .Z(n6279)
         );
  INV_X1 U7966 ( .A(n6279), .ZN(n6280) );
  OAI22_X1 U7967 ( .A1(n7603), .A2(n9478), .B1(n8192), .B2(n9445), .ZN(n6285)
         );
  INV_X1 U7968 ( .A(n6285), .ZN(n6289) );
  MUX2_X1 U7969 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n6286), .S(n9650), .Z(n6287)
         );
  INV_X1 U7970 ( .A(n6287), .ZN(n6288) );
  NOR2_X1 U7971 ( .A1(n5679), .A2(P1_U3086), .ZN(n6290) );
  INV_X1 U7972 ( .A(n6757), .ZN(n6291) );
  NAND2_X1 U7973 ( .A1(n7826), .A2(n6767), .ZN(n6292) );
  NAND2_X1 U7974 ( .A1(n6610), .A2(n6292), .ZN(n6609) );
  OR2_X1 U7975 ( .A1(n6609), .A2(n6293), .ZN(n6294) );
  NAND2_X1 U7976 ( .A1(n6294), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  XNOR2_X1 U7977 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  MUX2_X1 U7978 ( .A(n5674), .B(n6295), .S(P1_U3086), .Z(n6296) );
  INV_X1 U7979 ( .A(n6296), .ZN(P1_U3355) );
  AND2_X1 U7980 ( .A1(n4325), .A2(P2_U3151), .ZN(n8942) );
  INV_X2 U7981 ( .A(n8942), .ZN(n8945) );
  OAI222_X1 U7982 ( .A1(P2_U3151), .A2(n6695), .B1(n8947), .B2(n5666), .C1(
        n4619), .C2(n8945), .ZN(P2_U3294) );
  OAI222_X1 U7983 ( .A1(n8945), .A2(n6298), .B1(n8947), .B2(n6307), .C1(n9683), 
        .C2(P2_U3151), .ZN(P2_U3291) );
  INV_X1 U7984 ( .A(n8483), .ZN(n6570) );
  OAI222_X1 U7985 ( .A1(n6570), .A2(P2_U3151), .B1(n8947), .B2(n6310), .C1(
        n6299), .C2(n8945), .ZN(P2_U3293) );
  OAI222_X1 U7986 ( .A1(n6599), .A2(P2_U3151), .B1(n8947), .B2(n6312), .C1(
        n6300), .C2(n8945), .ZN(P2_U3292) );
  OAI222_X1 U7987 ( .A1(n6660), .A2(P2_U3151), .B1(n8947), .B2(n6303), .C1(
        n6301), .C2(n8945), .ZN(P2_U3290) );
  NAND2_X1 U7988 ( .A1(n4325), .A2(P1_U3086), .ZN(n9493) );
  CLKBUF_X1 U7989 ( .A(n9493), .Z(n9488) );
  OR2_X1 U7990 ( .A1(n4616), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9490) );
  INV_X1 U7991 ( .A(n9490), .ZN(n9486) );
  AOI22_X1 U7992 ( .A1(n6379), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9486), .ZN(n6302) );
  OAI21_X1 U7993 ( .B1(n6303), .B2(n9488), .A(n6302), .ZN(P1_U3350) );
  AOI22_X1 U7994 ( .A1(n6422), .A2(P1_STATE_REG_SCAN_IN), .B1(n9486), .B2(
        P2_DATAO_REG_6__SCAN_IN), .ZN(n6304) );
  OAI21_X1 U7995 ( .B1(n6306), .B2(n9488), .A(n6304), .ZN(P1_U3349) );
  OAI222_X1 U7996 ( .A1(n9714), .A2(P2_U3151), .B1(n8947), .B2(n6306), .C1(
        n6305), .C2(n8945), .ZN(P2_U3289) );
  INV_X1 U7997 ( .A(n6366), .ZN(n6412) );
  OAI222_X1 U7998 ( .A1(n9490), .A2(n6308), .B1(n9488), .B2(n6307), .C1(
        P1_U3086), .C2(n6412), .ZN(P1_U3351) );
  OAI222_X1 U7999 ( .A1(n9490), .A2(n6309), .B1(n9488), .B2(n5666), .C1(
        P1_U3086), .C2(n6360), .ZN(P1_U3354) );
  OAI222_X1 U8000 ( .A1(n9490), .A2(n6311), .B1(n9488), .B2(n6310), .C1(
        P1_U3086), .C2(n6358), .ZN(P1_U3353) );
  OAI222_X1 U8001 ( .A1(n9490), .A2(n6313), .B1(n9488), .B2(n6312), .C1(
        P1_U3086), .C2(n6363), .ZN(P1_U3352) );
  INV_X1 U8002 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10027) );
  NAND2_X1 U8003 ( .A1(n9623), .A2(n6315), .ZN(n6316) );
  OAI21_X1 U8004 ( .B1(n9623), .B2(n10027), .A(n6316), .ZN(P1_U3440) );
  INV_X1 U8005 ( .A(n6491), .ZN(n6427) );
  OAI222_X1 U8006 ( .A1(n9490), .A2(n6317), .B1(n9488), .B2(n6318), .C1(
        P1_U3086), .C2(n6427), .ZN(P1_U3348) );
  OAI222_X1 U8007 ( .A1(n8945), .A2(n6319), .B1(n8947), .B2(n6318), .C1(n6901), 
        .C2(P2_U3151), .ZN(P2_U3288) );
  INV_X1 U8008 ( .A(n6320), .ZN(n6321) );
  NAND2_X1 U8009 ( .A1(n6321), .A2(n8179), .ZN(n6353) );
  AOI21_X1 U8010 ( .B1(n6324), .B2(n6323), .A(n6322), .ZN(n6352) );
  INV_X1 U8011 ( .A(n6352), .ZN(n6325) );
  AND2_X1 U8012 ( .A1(n6353), .A2(n6325), .ZN(n9586) );
  NOR2_X1 U8013 ( .A1(n9586), .A2(P1_U3973), .ZN(P1_U3085) );
  AOI22_X1 U8014 ( .A1(n6626), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9486), .ZN(n6326) );
  OAI21_X1 U8015 ( .B1(n6327), .B2(n9488), .A(n6326), .ZN(P1_U3347) );
  OAI222_X1 U8016 ( .A1(n8533), .A2(P2_U3151), .B1(n8947), .B2(n6327), .C1(
        n9984), .C2(n8945), .ZN(P2_U3287) );
  INV_X1 U8017 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U8018 ( .A1(n4333), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U8019 ( .A1(n5696), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6329) );
  NAND2_X1 U8020 ( .A1(n5699), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6328) );
  AND3_X1 U8021 ( .A1(n6330), .A2(n6329), .A3(n6328), .ZN(n7934) );
  NAND2_X1 U8022 ( .A1(n8098), .A2(P1_U3973), .ZN(n6331) );
  OAI21_X1 U8023 ( .B1(P1_U3973), .B2(n6332), .A(n6331), .ZN(P1_U3585) );
  INV_X1 U8024 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6335) );
  INV_X1 U8025 ( .A(n6753), .ZN(n6333) );
  NAND2_X1 U8026 ( .A1(n6333), .A2(n6770), .ZN(n6334) );
  OAI21_X1 U8027 ( .B1(n6770), .B2(n6335), .A(n6334), .ZN(P2_U3377) );
  INV_X1 U8028 ( .A(n6336), .ZN(n6341) );
  AOI22_X1 U8029 ( .A1(n9141), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9486), .ZN(n6337) );
  OAI21_X1 U8030 ( .B1(n6341), .B2(n9488), .A(n6337), .ZN(P1_U3346) );
  INV_X1 U8031 ( .A(n6338), .ZN(n6343) );
  AOI22_X1 U8032 ( .A1(n9502), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9486), .ZN(n6339) );
  OAI21_X1 U8033 ( .B1(n6343), .B2(n9488), .A(n6339), .ZN(P1_U3345) );
  INV_X1 U8034 ( .A(n9734), .ZN(n8531) );
  OAI222_X1 U8035 ( .A1(P2_U3151), .A2(n8531), .B1(n8947), .B2(n6341), .C1(
        n6340), .C2(n8945), .ZN(P2_U3286) );
  INV_X1 U8036 ( .A(n9746), .ZN(n8529) );
  OAI222_X1 U8037 ( .A1(P2_U3151), .A2(n8529), .B1(n8947), .B2(n6343), .C1(
        n6342), .C2(n8945), .ZN(P2_U3285) );
  INV_X1 U8038 ( .A(n6363), .ZN(n6387) );
  INV_X1 U8039 ( .A(n6358), .ZN(n6448) );
  INV_X1 U8040 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6644) );
  MUX2_X1 U8041 ( .A(n6644), .B(P1_REG2_REG_2__SCAN_IN), .S(n6358), .Z(n6443)
         );
  INV_X1 U8042 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6344) );
  MUX2_X1 U8043 ( .A(n6344), .B(P1_REG2_REG_1__SCAN_IN), .S(n6360), .Z(n9113)
         );
  AND2_X1 U8044 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9112) );
  NAND2_X1 U8045 ( .A1(n9113), .A2(n9112), .ZN(n9111) );
  INV_X1 U8046 ( .A(n6360), .ZN(n9117) );
  NAND2_X1 U8047 ( .A1(n9117), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6345) );
  NAND2_X1 U8048 ( .A1(n9111), .A2(n6345), .ZN(n6442) );
  AND2_X1 U8049 ( .A1(n6443), .A2(n6442), .ZN(n6440) );
  INV_X1 U8050 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6346) );
  MUX2_X1 U8051 ( .A(n6346), .B(P1_REG2_REG_3__SCAN_IN), .S(n6363), .Z(n6347)
         );
  INV_X1 U8052 ( .A(n6347), .ZN(n6391) );
  INV_X1 U8053 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6348) );
  MUX2_X1 U8054 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6348), .S(n6366), .Z(n6349)
         );
  INV_X1 U8055 ( .A(n6349), .ZN(n6406) );
  AOI21_X1 U8056 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n6366), .A(n6405), .ZN(
        n6357) );
  INV_X1 U8057 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6350) );
  MUX2_X1 U8058 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6350), .S(n6379), .Z(n6351)
         );
  INV_X1 U8059 ( .A(n6351), .ZN(n6356) );
  NAND2_X1 U8060 ( .A1(n6353), .A2(n6352), .ZN(n9510) );
  OR2_X1 U8061 ( .A1(n4324), .A2(n6354), .ZN(n6355) );
  AOI211_X1 U8062 ( .C1(n6357), .C2(n6356), .A(n9607), .B(n6375), .ZN(n6374)
         );
  INV_X1 U8063 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6359) );
  MUX2_X1 U8064 ( .A(n6359), .B(P1_REG1_REG_2__SCAN_IN), .S(n6358), .Z(n6447)
         );
  INV_X1 U8065 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6361) );
  MUX2_X1 U8066 ( .A(n6361), .B(P1_REG1_REG_1__SCAN_IN), .S(n6360), .Z(n9116)
         );
  AND2_X1 U8067 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9115) );
  NAND2_X1 U8068 ( .A1(n9116), .A2(n9115), .ZN(n9114) );
  NAND2_X1 U8069 ( .A1(n9117), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6362) );
  NAND2_X1 U8070 ( .A1(n9114), .A2(n6362), .ZN(n6446) );
  AOI21_X1 U8071 ( .B1(n6448), .B2(P1_REG1_REG_2__SCAN_IN), .A(n6444), .ZN(
        n6395) );
  INV_X1 U8072 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6364) );
  MUX2_X1 U8073 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6364), .S(n6363), .Z(n6394)
         );
  NOR2_X1 U8074 ( .A1(n6395), .A2(n6394), .ZN(n6393) );
  INV_X1 U8075 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6365) );
  MUX2_X1 U8076 ( .A(n6365), .B(P1_REG1_REG_4__SCAN_IN), .S(n6366), .Z(n6409)
         );
  NOR2_X1 U8077 ( .A1(n6410), .A2(n6409), .ZN(n6408) );
  INV_X1 U8078 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6367) );
  MUX2_X1 U8079 ( .A(n6367), .B(P1_REG1_REG_5__SCAN_IN), .S(n6379), .Z(n6368)
         );
  INV_X1 U8080 ( .A(n6354), .ZN(n9507) );
  NOR2_X1 U8081 ( .A1(n6369), .A2(n6368), .ZN(n6378) );
  AOI211_X1 U8082 ( .C1(n6369), .C2(n6368), .A(n9540), .B(n6378), .ZN(n6373)
         );
  INV_X1 U8083 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6371) );
  NAND2_X1 U8084 ( .A1(n9599), .A2(n6379), .ZN(n6370) );
  NAND2_X1 U8085 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6891) );
  OAI211_X1 U8086 ( .C1(n6371), .C2(n9622), .A(n6370), .B(n6891), .ZN(n6372)
         );
  OR3_X1 U8087 ( .A1(n6374), .A2(n6373), .A3(n6372), .ZN(P1_U3248) );
  XNOR2_X1 U8088 ( .A(n6422), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n6376) );
  AOI211_X1 U8089 ( .C1(n6377), .C2(n6376), .A(n9607), .B(n6416), .ZN(n6386)
         );
  XNOR2_X1 U8090 ( .A(n6422), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n6380) );
  NOR2_X1 U8091 ( .A1(n6381), .A2(n6380), .ZN(n6421) );
  AOI211_X1 U8092 ( .C1(n6381), .C2(n6380), .A(n9540), .B(n6421), .ZN(n6385)
         );
  INV_X1 U8093 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6383) );
  NAND2_X1 U8094 ( .A1(n9599), .A2(n6422), .ZN(n6382) );
  NAND2_X1 U8095 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7110) );
  OAI211_X1 U8096 ( .C1(n6383), .C2(n9622), .A(n6382), .B(n7110), .ZN(n6384)
         );
  OR3_X1 U8097 ( .A1(n6386), .A2(n6385), .A3(n6384), .ZN(P1_U3249) );
  INV_X1 U8098 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U8099 ( .A1(n9599), .A2(n6387), .ZN(n6388) );
  NAND2_X1 U8100 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n6481) );
  OAI211_X1 U8101 ( .C1(n6389), .C2(n9622), .A(n6388), .B(n6481), .ZN(n6398)
         );
  AOI211_X1 U8102 ( .C1(n6392), .C2(n6391), .A(n6390), .B(n9607), .ZN(n6397)
         );
  AOI211_X1 U8103 ( .C1(n6395), .C2(n6394), .A(n6393), .B(n9540), .ZN(n6396)
         );
  OR3_X1 U8104 ( .A1(n6398), .A2(n6397), .A3(n6396), .ZN(P1_U3246) );
  XNOR2_X1 U8105 ( .A(n6400), .B(n6399), .ZN(n6463) );
  MUX2_X1 U8106 ( .A(n6463), .B(n9112), .S(n9507), .Z(n6404) );
  INV_X1 U8107 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6401) );
  AOI21_X1 U8108 ( .B1(n9507), .B2(n6401), .A(n4324), .ZN(n9506) );
  OAI21_X1 U8109 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n9506), .A(P1_U3973), .ZN(
        n6402) );
  AOI21_X1 U8110 ( .B1(n6404), .B2(n6403), .A(n6402), .ZN(n6454) );
  AOI211_X1 U8111 ( .C1(n6407), .C2(n6406), .A(n6405), .B(n9607), .ZN(n6415)
         );
  AOI211_X1 U8112 ( .C1(n6410), .C2(n6409), .A(n6408), .B(n9540), .ZN(n6414)
         );
  NAND2_X1 U8113 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n6742) );
  NAND2_X1 U8114 ( .A1(n9586), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n6411) );
  OAI211_X1 U8115 ( .C1(n9616), .C2(n6412), .A(n6742), .B(n6411), .ZN(n6413)
         );
  OR4_X1 U8116 ( .A1(n6454), .A2(n6415), .A3(n6414), .A4(n6413), .ZN(P1_U3247)
         );
  INV_X1 U8117 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6417) );
  MUX2_X1 U8118 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6417), .S(n6491), .Z(n6418)
         );
  INV_X1 U8119 ( .A(n6418), .ZN(n6419) );
  NOR2_X1 U8120 ( .A1(n6420), .A2(n6419), .ZN(n6490) );
  AOI211_X1 U8121 ( .C1(n6420), .C2(n6419), .A(n9607), .B(n6490), .ZN(n6430)
         );
  INV_X1 U8122 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6423) );
  MUX2_X1 U8123 ( .A(n6423), .B(P1_REG1_REG_7__SCAN_IN), .S(n6491), .Z(n6424)
         );
  NOR2_X1 U8124 ( .A1(n6425), .A2(n6424), .ZN(n6486) );
  AOI211_X1 U8125 ( .C1(n6425), .C2(n6424), .A(n9540), .B(n6486), .ZN(n6429)
         );
  NOR2_X1 U8126 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10026), .ZN(n7102) );
  AOI21_X1 U8127 ( .B1(n9586), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7102), .ZN(
        n6426) );
  OAI21_X1 U8128 ( .B1(n9616), .B2(n6427), .A(n6426), .ZN(n6428) );
  OR3_X1 U8129 ( .A1(n6430), .A2(n6429), .A3(n6428), .ZN(P1_U3250) );
  INV_X1 U8130 ( .A(n6431), .ZN(n6432) );
  INV_X1 U8131 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6433) );
  NOR2_X1 U8132 ( .A1(n6716), .A2(n6433), .ZN(P2_U3260) );
  INV_X1 U8133 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6434) );
  NOR2_X1 U8134 ( .A1(n6716), .A2(n6434), .ZN(P2_U3249) );
  INV_X1 U8135 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n6435) );
  NOR2_X1 U8136 ( .A1(n6716), .A2(n6435), .ZN(P2_U3261) );
  INV_X1 U8137 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6436) );
  NOR2_X1 U8138 ( .A1(n6716), .A2(n6436), .ZN(P2_U3259) );
  INV_X1 U8139 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6437) );
  NOR2_X1 U8140 ( .A1(n6716), .A2(n6437), .ZN(P2_U3258) );
  INV_X1 U8141 ( .A(n6438), .ZN(n6466) );
  AOI22_X1 U8142 ( .A1(n9520), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9486), .ZN(n6439) );
  OAI21_X1 U8143 ( .B1(n6466), .B2(n9488), .A(n6439), .ZN(P1_U3344) );
  INV_X1 U8144 ( .A(n6440), .ZN(n6441) );
  OAI211_X1 U8145 ( .C1(n6443), .C2(n6442), .A(n9602), .B(n6441), .ZN(n6452)
         );
  AOI22_X1 U8146 ( .A1(n9586), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6451) );
  INV_X1 U8147 ( .A(n6444), .ZN(n6445) );
  OAI211_X1 U8148 ( .C1(n6447), .C2(n6446), .A(n9610), .B(n6445), .ZN(n6450)
         );
  NAND2_X1 U8149 ( .A1(n9599), .A2(n6448), .ZN(n6449) );
  NAND4_X1 U8150 ( .A1(n6452), .A2(n6451), .A3(n6450), .A4(n6449), .ZN(n6453)
         );
  OR2_X1 U8151 ( .A1(n6454), .A2(n6453), .ZN(P1_U3245) );
  INV_X1 U8152 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6458) );
  AND2_X1 U8153 ( .A1(n9110), .A2(n7592), .ZN(n8109) );
  NOR2_X1 U8154 ( .A1(n8109), .A2(n6977), .ZN(n7942) );
  INV_X1 U8155 ( .A(n7942), .ZN(n6455) );
  OAI21_X1 U8156 ( .B1(n9352), .B2(n9648), .A(n6455), .ZN(n6456) );
  NAND2_X1 U8157 ( .A1(n9109), .A2(n9337), .ZN(n7587) );
  OAI211_X1 U8158 ( .C1(n7586), .C2(n7592), .A(n6456), .B(n7587), .ZN(n9435)
         );
  NAND2_X1 U8159 ( .A1(n9435), .A2(n9480), .ZN(n6457) );
  OAI21_X1 U8160 ( .B1(n9480), .B2(n6458), .A(n6457), .ZN(P1_U3453) );
  NAND2_X1 U8161 ( .A1(n6460), .A2(n6459), .ZN(n7871) );
  OAI22_X1 U8162 ( .A1(n9080), .A2(n7592), .B1(n6503), .B2(n9068), .ZN(n6461)
         );
  AOI21_X1 U8163 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n7871), .A(n6461), .ZN(
        n6462) );
  OAI21_X1 U8164 ( .B1(n4495), .B2(n6463), .A(n6462), .ZN(P1_U3232) );
  INV_X1 U8165 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U8166 ( .A1(P2_U3893), .A2(n8770), .ZN(n6464) );
  OAI21_X1 U8167 ( .B1(P2_U3893), .B2(n6692), .A(n6464), .ZN(P2_U3506) );
  INV_X1 U8168 ( .A(n9764), .ZN(n8527) );
  INV_X1 U8169 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6465) );
  OAI222_X1 U8170 ( .A1(n8527), .A2(P2_U3151), .B1(n8947), .B2(n6466), .C1(
        n6465), .C2(n8945), .ZN(P2_U3284) );
  NAND4_X1 U8171 ( .A1(n7913), .A2(P2_STATE_REG_SCAN_IN), .A3(n7541), .A4(
        n6767), .ZN(n6467) );
  OAI21_X1 U8172 ( .B1(n6716), .B2(P2_D_REG_0__SCAN_IN), .A(n6467), .ZN(n6468)
         );
  INV_X1 U8173 ( .A(n6468), .ZN(P2_U3376) );
  XOR2_X1 U8174 ( .A(n6469), .B(n6470), .Z(n6474) );
  INV_X1 U8175 ( .A(n9078), .ZN(n9061) );
  AOI22_X1 U8176 ( .A1(n9061), .A2(n9109), .B1(n9076), .B2(n9108), .ZN(n6471)
         );
  OAI21_X1 U8177 ( .B1(n6212), .B2(n9080), .A(n6471), .ZN(n6472) );
  AOI21_X1 U8178 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7871), .A(n6472), .ZN(
        n6473) );
  OAI21_X1 U8179 ( .B1(n6474), .B2(n4495), .A(n6473), .ZN(P1_U3237) );
  INV_X1 U8180 ( .A(n6475), .ZN(n6478) );
  AOI22_X1 U8181 ( .A1(n9524), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9486), .ZN(n6476) );
  OAI21_X1 U8182 ( .B1(n6478), .B2(n9488), .A(n6476), .ZN(P1_U3343) );
  INV_X1 U8183 ( .A(n9778), .ZN(n8525) );
  INV_X1 U8184 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6477) );
  OAI222_X1 U8185 ( .A1(P2_U3151), .A2(n8525), .B1(n8947), .B2(n6478), .C1(
        n6477), .C2(n8945), .ZN(P2_U3283) );
  XOR2_X1 U8186 ( .A(n6480), .B(n6479), .Z(n6485) );
  AOI22_X1 U8187 ( .A1(n9076), .A2(n9107), .B1(n9035), .B2(n6215), .ZN(n6482)
         );
  OAI211_X1 U8188 ( .C1(n7877), .C2(n9078), .A(n6482), .B(n6481), .ZN(n6483)
         );
  AOI21_X1 U8189 ( .B1(n6649), .B2(n9084), .A(n6483), .ZN(n6484) );
  OAI21_X1 U8190 ( .B1(n6485), .B2(n4495), .A(n6484), .ZN(P1_U3218) );
  AOI21_X1 U8191 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6491), .A(n6486), .ZN(
        n6489) );
  INV_X1 U8192 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6487) );
  MUX2_X1 U8193 ( .A(n6487), .B(P1_REG1_REG_8__SCAN_IN), .S(n6626), .Z(n6488)
         );
  NOR2_X1 U8194 ( .A1(n6489), .A2(n6488), .ZN(n6618) );
  AOI211_X1 U8195 ( .C1(n6489), .C2(n6488), .A(n9540), .B(n6618), .ZN(n6498)
         );
  XNOR2_X1 U8196 ( .A(n6626), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6492) );
  AOI211_X1 U8197 ( .C1(n6493), .C2(n6492), .A(n9607), .B(n6625), .ZN(n6497)
         );
  INV_X1 U8198 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6495) );
  NAND2_X1 U8199 ( .A1(n9599), .A2(n6626), .ZN(n6494) );
  NAND2_X1 U8200 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n7193) );
  OAI211_X1 U8201 ( .C1(n6495), .C2(n9622), .A(n6494), .B(n7193), .ZN(n6496)
         );
  OR3_X1 U8202 ( .A1(n6498), .A2(n6497), .A3(n6496), .ZN(P1_U3251) );
  OAI21_X1 U8203 ( .B1(n6500), .B2(n6502), .A(n6499), .ZN(n6646) );
  INV_X1 U8204 ( .A(n9354), .ZN(n9326) );
  AOI211_X1 U8205 ( .C1(n6505), .C2(n6976), .A(n9326), .B(n6501), .ZN(n6643)
         );
  XNOR2_X1 U8206 ( .A(n6502), .B(n8117), .ZN(n6504) );
  OAI222_X1 U8207 ( .A1(n9349), .A2(n6216), .B1(n6504), .B2(n9299), .C1(n9347), 
        .C2(n6503), .ZN(n6641) );
  AOI211_X1 U8208 ( .C1(n9648), .C2(n6646), .A(n6643), .B(n6641), .ZN(n6988)
         );
  AOI22_X1 U8209 ( .A1(n9414), .A2(n6505), .B1(n9656), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6506) );
  OAI21_X1 U8210 ( .B1(n6988), .B2(n9656), .A(n6506), .ZN(P1_U3524) );
  INV_X1 U8211 ( .A(n6507), .ZN(n6550) );
  AOI22_X1 U8212 ( .A1(n9549), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9486), .ZN(n6508) );
  OAI21_X1 U8213 ( .B1(n6550), .B2(n9488), .A(n6508), .ZN(P1_U3342) );
  OAI21_X1 U8214 ( .B1(n6510), .B2(n7945), .A(n6509), .ZN(n6993) );
  INV_X1 U8215 ( .A(n6993), .ZN(n6527) );
  NAND3_X1 U8216 ( .A1(n6513), .A2(n6512), .A3(n6511), .ZN(n6519) );
  NAND2_X1 U8217 ( .A1(n6514), .A2(n4331), .ZN(n7471) );
  NAND2_X1 U8218 ( .A1(n7467), .A2(n7471), .ZN(n6515) );
  NAND3_X1 U8219 ( .A1(n6539), .A2(n7990), .A3(n7945), .ZN(n6516) );
  NAND2_X1 U8220 ( .A1(n6517), .A2(n6516), .ZN(n6518) );
  AOI222_X1 U8221 ( .A1(n9352), .A2(n6518), .B1(n9105), .B2(n9337), .C1(n9107), 
        .C2(n9335), .ZN(n6632) );
  MUX2_X1 U8222 ( .A(n6350), .B(n6632), .S(n9365), .Z(n6526) );
  AOI21_X1 U8223 ( .B1(n6537), .B2(n6520), .A(n9326), .ZN(n6521) );
  AND2_X1 U8224 ( .A1(n6521), .A2(n6685), .ZN(n6633) );
  INV_X1 U8225 ( .A(n6895), .ZN(n6523) );
  OAI22_X1 U8226 ( .A1(n9330), .A2(n6990), .B1(n9211), .B2(n6523), .ZN(n6524)
         );
  AOI21_X1 U8227 ( .B1(n9342), .B2(n6633), .A(n6524), .ZN(n6525) );
  OAI211_X1 U8228 ( .C1(n6527), .C2(n9368), .A(n6526), .B(n6525), .ZN(P1_U3288) );
  NOR2_X1 U8229 ( .A1(n5118), .A2(n8838), .ZN(n6829) );
  AND2_X1 U8230 ( .A1(n8228), .A2(n8852), .ZN(n6528) );
  NOR2_X1 U8231 ( .A1(n6829), .A2(n6528), .ZN(n6531) );
  INV_X1 U8232 ( .A(n8228), .ZN(n6529) );
  NAND2_X1 U8233 ( .A1(n8475), .A2(n6529), .ZN(n7685) );
  NAND2_X1 U8234 ( .A1(n7682), .A2(n7685), .ZN(n8229) );
  OAI21_X1 U8235 ( .B1(n7371), .B2(n8842), .A(n8229), .ZN(n6530) );
  AND2_X1 U8236 ( .A1(n6531), .A2(n6530), .ZN(n9878) );
  NAND2_X1 U8237 ( .A1(n8857), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6532) );
  OAI21_X1 U8238 ( .B1(n8857), .B2(n9878), .A(n6532), .ZN(P2_U3459) );
  INV_X1 U8239 ( .A(n6533), .ZN(n6639) );
  AOI22_X1 U8240 ( .A1(n9562), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9486), .ZN(n6534) );
  OAI21_X1 U8241 ( .B1(n6639), .B2(n9488), .A(n6534), .ZN(P1_U3341) );
  OAI21_X1 U8242 ( .B1(n6536), .B2(n7944), .A(n6535), .ZN(n9629) );
  OAI211_X1 U8243 ( .C1(n6558), .C2(n9626), .A(n6537), .B(n9354), .ZN(n9625)
         );
  AOI22_X1 U8244 ( .A1(n9359), .A2(n6741), .B1(n9356), .B2(n6749), .ZN(n6538)
         );
  OAI21_X1 U8245 ( .B1(n9363), .B2(n9625), .A(n6538), .ZN(n6547) );
  OAI21_X1 U8246 ( .B1(n7981), .B2(n6540), .A(n6539), .ZN(n6541) );
  NAND2_X1 U8247 ( .A1(n6541), .A2(n9352), .ZN(n6545) );
  OAI22_X1 U8248 ( .A1(n6542), .A2(n9349), .B1(n6216), .B2(n9347), .ZN(n6543)
         );
  INV_X1 U8249 ( .A(n6543), .ZN(n6544) );
  NAND2_X1 U8250 ( .A1(n6545), .A2(n6544), .ZN(n9627) );
  MUX2_X1 U8251 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9627), .S(n9365), .Z(n6546)
         );
  AOI211_X1 U8252 ( .C1(n9209), .C2(n9629), .A(n6547), .B(n6546), .ZN(n6548)
         );
  INV_X1 U8253 ( .A(n6548), .ZN(P1_U3289) );
  INV_X1 U8254 ( .A(n9795), .ZN(n8523) );
  INV_X1 U8255 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6549) );
  OAI222_X1 U8256 ( .A1(P2_U3151), .A2(n8523), .B1(n8947), .B2(n6550), .C1(
        n6549), .C2(n8945), .ZN(P2_U3282) );
  INV_X1 U8257 ( .A(n7978), .ZN(n6553) );
  INV_X1 U8258 ( .A(n6551), .ZN(n6552) );
  AOI21_X1 U8259 ( .B1(n6553), .B2(n7946), .A(n6552), .ZN(n6554) );
  OAI222_X1 U8260 ( .A1(n9349), .A2(n6555), .B1(n9347), .B2(n7877), .C1(n9299), 
        .C2(n6554), .ZN(n6652) );
  NAND2_X1 U8261 ( .A1(n6556), .A2(n9354), .ZN(n6557) );
  NOR2_X1 U8262 ( .A1(n6558), .A2(n6557), .ZN(n6650) );
  NOR2_X1 U8263 ( .A1(n6652), .A2(n6650), .ZN(n6973) );
  INV_X1 U8264 ( .A(n9427), .ZN(n6636) );
  OR2_X1 U8265 ( .A1(n6559), .A2(n7946), .ZN(n6560) );
  NAND2_X1 U8266 ( .A1(n6561), .A2(n6560), .ZN(n6971) );
  OAI22_X1 U8267 ( .A1(n9384), .A2(n6562), .B1(n9659), .B2(n6364), .ZN(n6563)
         );
  AOI21_X1 U8268 ( .B1(n6636), .B2(n6971), .A(n6563), .ZN(n6564) );
  OAI21_X1 U8269 ( .B1(n6973), .B2(n9656), .A(n6564), .ZN(P1_U3525) );
  MUX2_X1 U8270 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8588), .Z(n6657) );
  XNOR2_X1 U8271 ( .A(n6657), .B(n6660), .ZN(n6579) );
  INV_X1 U8272 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6702) );
  MUX2_X1 U8273 ( .A(n6878), .B(n6702), .S(n5514), .Z(n6567) );
  XNOR2_X1 U8274 ( .A(n6567), .B(n6695), .ZN(n6697) );
  INV_X1 U8275 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6832) );
  INV_X1 U8276 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6566) );
  MUX2_X1 U8277 ( .A(n6832), .B(n6566), .S(n5514), .Z(n6801) );
  NAND2_X1 U8278 ( .A1(n6801), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6800) );
  NAND2_X1 U8279 ( .A1(n6697), .A2(n6800), .ZN(n6696) );
  INV_X1 U8280 ( .A(n6567), .ZN(n6568) );
  NAND2_X1 U8281 ( .A1(n6568), .A2(n6695), .ZN(n6569) );
  NAND2_X1 U8282 ( .A1(n6696), .A2(n6569), .ZN(n8485) );
  MUX2_X1 U8283 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n5514), .Z(n6571) );
  XNOR2_X1 U8284 ( .A(n6571), .B(n8483), .ZN(n8486) );
  NAND2_X1 U8285 ( .A1(n8485), .A2(n8486), .ZN(n8484) );
  NAND2_X1 U8286 ( .A1(n6571), .A2(n6570), .ZN(n6572) );
  NAND2_X1 U8287 ( .A1(n8484), .A2(n6572), .ZN(n9672) );
  MUX2_X1 U8288 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n5514), .Z(n6573) );
  XNOR2_X1 U8289 ( .A(n6573), .B(n6599), .ZN(n9671) );
  OR2_X1 U8290 ( .A1(n9672), .A2(n9671), .ZN(n9675) );
  INV_X1 U8291 ( .A(n6573), .ZN(n6574) );
  INV_X1 U8292 ( .A(n6599), .ZN(n9666) );
  NAND2_X1 U8293 ( .A1(n6574), .A2(n9666), .ZN(n6575) );
  AND2_X1 U8294 ( .A1(n9675), .A2(n6575), .ZN(n9689) );
  MUX2_X1 U8295 ( .A(n7135), .B(n6603), .S(n8588), .Z(n6576) );
  XNOR2_X1 U8296 ( .A(n6576), .B(n9683), .ZN(n9687) );
  INV_X1 U8297 ( .A(n6576), .ZN(n6577) );
  AOI22_X1 U8298 ( .A1(n9689), .A2(n9687), .B1(n6577), .B2(n9683), .ZN(n6578)
         );
  NAND2_X1 U8299 ( .A1(P2_U3893), .A2(n7863), .ZN(n9673) );
  NOR2_X1 U8300 ( .A1(n6578), .A2(n6579), .ZN(n6656) );
  AOI211_X1 U8301 ( .C1(n6579), .C2(n6578), .A(n9673), .B(n6656), .ZN(n6617)
         );
  INV_X1 U8302 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10125) );
  INV_X1 U8303 ( .A(n6610), .ZN(n6580) );
  NOR2_X2 U8304 ( .A1(P2_U3150), .A2(n6580), .ZN(n9845) );
  NAND2_X1 U8305 ( .A1(n6581), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7567) );
  NOR2_X1 U8306 ( .A1(n6609), .A2(n7567), .ZN(n6803) );
  INV_X1 U8307 ( .A(n9860), .ZN(n9805) );
  INV_X1 U8308 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10056) );
  AND2_X1 U8309 ( .A1(n10056), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6582) );
  NAND2_X1 U8310 ( .A1(n6590), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6583) );
  OAI21_X1 U8311 ( .B1(n6695), .B2(n6582), .A(n6583), .ZN(n6701) );
  OR2_X1 U8312 ( .A1(n6701), .A2(n6878), .ZN(n6699) );
  NAND2_X1 U8313 ( .A1(n6699), .A2(n6583), .ZN(n8477) );
  INV_X1 U8314 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6584) );
  OR2_X1 U8315 ( .A1(n8483), .A2(n6584), .ZN(n6585) );
  NAND2_X1 U8316 ( .A1(n8476), .A2(n6585), .ZN(n6586) );
  NAND2_X1 U8317 ( .A1(n6586), .A2(n6599), .ZN(n9692) );
  OR2_X1 U8318 ( .A1(n6586), .A2(n6599), .ZN(n6587) );
  AND2_X1 U8319 ( .A1(n9692), .A2(n6587), .ZN(n9660) );
  NAND2_X1 U8320 ( .A1(n9694), .A2(n9692), .ZN(n6588) );
  MUX2_X1 U8321 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7135), .S(n9683), .Z(n9691)
         );
  NAND2_X1 U8322 ( .A1(n6589), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9707) );
  OAI21_X1 U8323 ( .B1(n6589), .B2(P2_REG2_REG_5__SCAN_IN), .A(n9707), .ZN(
        n6606) );
  NAND2_X1 U8324 ( .A1(n6803), .A2(n8588), .ZN(n9664) );
  XNOR2_X1 U8325 ( .A(n8483), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n8480) );
  NAND2_X1 U8326 ( .A1(n6590), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6594) );
  NAND2_X1 U8327 ( .A1(n6695), .A2(n6594), .ZN(n6593) );
  NAND2_X1 U8328 ( .A1(n10056), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6591) );
  OR2_X1 U8329 ( .A1(n6591), .A2(n6590), .ZN(n6592) );
  NAND2_X1 U8330 ( .A1(n6593), .A2(n6592), .ZN(n6703) );
  NAND2_X1 U8331 ( .A1(n6703), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U8332 ( .A1(n6595), .A2(n6594), .ZN(n8479) );
  NAND2_X1 U8333 ( .A1(n8480), .A2(n8479), .ZN(n6598) );
  INV_X1 U8334 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6596) );
  OR2_X1 U8335 ( .A1(n8483), .A2(n6596), .ZN(n6597) );
  NAND2_X1 U8336 ( .A1(n6598), .A2(n6597), .ZN(n6600) );
  XNOR2_X1 U8337 ( .A(n6600), .B(n9666), .ZN(n9662) );
  NAND2_X1 U8338 ( .A1(n9662), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6602) );
  NAND2_X1 U8339 ( .A1(n6600), .A2(n6599), .ZN(n6601) );
  NAND2_X1 U8340 ( .A1(n6602), .A2(n6601), .ZN(n9680) );
  MUX2_X1 U8341 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6603), .S(n9683), .Z(n9681)
         );
  NAND2_X1 U8342 ( .A1(n9680), .A2(n9681), .ZN(n9679) );
  NAND2_X1 U8343 ( .A1(n9683), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U8344 ( .A1(n9679), .A2(n6604), .ZN(n6661) );
  INV_X1 U8345 ( .A(n6660), .ZN(n6613) );
  XNOR2_X1 U8346 ( .A(n6661), .B(n6613), .ZN(n6659) );
  XNOR2_X1 U8347 ( .A(n6659), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n6605) );
  AOI22_X1 U8348 ( .A1(n9805), .A2(n6606), .B1(n9856), .B2(n6605), .ZN(n6615)
         );
  NOR2_X1 U8349 ( .A1(n8588), .A2(P2_U3151), .ZN(n6607) );
  NAND2_X1 U8350 ( .A1(n6607), .A2(n7863), .ZN(n6608) );
  OR2_X1 U8351 ( .A1(n6609), .A2(n6608), .ZN(n6612) );
  OR2_X1 U8352 ( .A1(n6610), .A2(n7567), .ZN(n6611) );
  AND2_X1 U8353 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7009) );
  AOI21_X1 U8354 ( .B1(n9846), .B2(n6613), .A(n7009), .ZN(n6614) );
  OAI211_X1 U8355 ( .C1(n10125), .C2(n9745), .A(n6615), .B(n6614), .ZN(n6616)
         );
  OR2_X1 U8356 ( .A1(n6617), .A2(n6616), .ZN(P2_U3187) );
  XOR2_X1 U8357 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9141), .Z(n6620) );
  NAND2_X1 U8358 ( .A1(n6619), .A2(n6620), .ZN(n9140) );
  OAI21_X1 U8359 ( .B1(n6620), .B2(n6619), .A(n9140), .ZN(n6624) );
  INV_X1 U8360 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6622) );
  NAND2_X1 U8361 ( .A1(n9599), .A2(n9141), .ZN(n6621) );
  NAND2_X1 U8362 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n7294) );
  OAI211_X1 U8363 ( .C1(n6622), .C2(n9622), .A(n6621), .B(n7294), .ZN(n6623)
         );
  AOI21_X1 U8364 ( .B1(n6624), .B2(n9610), .A(n6623), .ZN(n6631) );
  XOR2_X1 U8365 ( .A(n9141), .B(P1_REG2_REG_9__SCAN_IN), .Z(n6628) );
  OAI21_X1 U8366 ( .B1(n6628), .B2(n6627), .A(n9124), .ZN(n6629) );
  NAND2_X1 U8367 ( .A1(n6629), .A2(n9602), .ZN(n6630) );
  NAND2_X1 U8368 ( .A1(n6631), .A2(n6630), .ZN(P1_U3252) );
  INV_X1 U8369 ( .A(n6632), .ZN(n6634) );
  NOR2_X1 U8370 ( .A1(n6634), .A2(n6633), .ZN(n6995) );
  OAI22_X1 U8371 ( .A1(n9384), .A2(n6990), .B1(n9659), .B2(n6367), .ZN(n6635)
         );
  AOI21_X1 U8372 ( .B1(n6993), .B2(n6636), .A(n6635), .ZN(n6637) );
  OAI21_X1 U8373 ( .B1(n6995), .B2(n9656), .A(n6637), .ZN(P1_U3527) );
  INV_X1 U8374 ( .A(n9812), .ZN(n8521) );
  INV_X1 U8375 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6638) );
  OAI222_X1 U8376 ( .A1(n8521), .A2(P2_U3151), .B1(n8947), .B2(n6639), .C1(
        n6638), .C2(n8945), .ZN(P2_U3281) );
  INV_X1 U8377 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6640) );
  NOR2_X1 U8378 ( .A1(n9211), .A2(n6640), .ZN(n6642) );
  AOI211_X1 U8379 ( .C1(n6643), .C2(n9203), .A(n6642), .B(n6641), .ZN(n6648)
         );
  OAI22_X1 U8380 ( .A1(n9330), .A2(n6212), .B1(n6644), .B2(n9365), .ZN(n6645)
         );
  AOI21_X1 U8381 ( .B1(n9209), .B2(n6646), .A(n6645), .ZN(n6647) );
  OAI21_X1 U8382 ( .B1(n6648), .B2(n9358), .A(n6647), .ZN(P1_U3291) );
  AOI22_X1 U8383 ( .A1(n9342), .A2(n6650), .B1(n9356), .B2(n6649), .ZN(n6651)
         );
  OAI21_X1 U8384 ( .B1(n9330), .B2(n6562), .A(n6651), .ZN(n6654) );
  MUX2_X1 U8385 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6652), .S(n9365), .Z(n6653)
         );
  AOI211_X1 U8386 ( .C1(n9209), .C2(n6971), .A(n6654), .B(n6653), .ZN(n6655)
         );
  INV_X1 U8387 ( .A(n6655), .ZN(P1_U3290) );
  MUX2_X1 U8388 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8588), .Z(n6916) );
  XOR2_X1 U8389 ( .A(n6901), .B(n6916), .Z(n6919) );
  MUX2_X1 U8390 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8588), .Z(n6658) );
  AOI21_X1 U8391 ( .B1(n6657), .B2(n6660), .A(n6656), .ZN(n9723) );
  XOR2_X1 U8392 ( .A(n9714), .B(n6658), .Z(n9722) );
  NAND2_X1 U8393 ( .A1(n9723), .A2(n9722), .ZN(n9721) );
  OAI21_X1 U8394 ( .B1(n6658), .B2(n9714), .A(n9721), .ZN(n6920) );
  XOR2_X1 U8395 ( .A(n6919), .B(n6920), .Z(n6678) );
  NAND2_X1 U8396 ( .A1(n6659), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U8397 ( .A1(n6661), .A2(n6660), .ZN(n6662) );
  NAND2_X1 U8398 ( .A1(n6663), .A2(n6662), .ZN(n9711) );
  INV_X1 U8399 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6664) );
  MUX2_X1 U8400 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6664), .S(n9714), .Z(n9712)
         );
  NAND2_X1 U8401 ( .A1(n9711), .A2(n9712), .ZN(n9710) );
  NAND2_X1 U8402 ( .A1(n9714), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6665) );
  NAND2_X1 U8403 ( .A1(n9710), .A2(n6665), .ZN(n6902) );
  INV_X1 U8404 ( .A(n6901), .ZN(n6918) );
  XNOR2_X1 U8405 ( .A(n6902), .B(n6918), .ZN(n6900) );
  XNOR2_X1 U8406 ( .A(n6900), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n6676) );
  NAND2_X1 U8407 ( .A1(n9707), .A2(n9705), .ZN(n6666) );
  INV_X1 U8408 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7071) );
  XNOR2_X1 U8409 ( .A(n9714), .B(n7071), .ZN(n9704) );
  NAND2_X1 U8410 ( .A1(n6666), .A2(n9704), .ZN(n9709) );
  NAND2_X1 U8411 ( .A1(n9714), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U8412 ( .A1(n9709), .A2(n6667), .ZN(n6668) );
  OR2_X1 U8413 ( .A1(n6668), .A2(n6901), .ZN(n6669) );
  NAND2_X1 U8414 ( .A1(n6668), .A2(n6901), .ZN(n6908) );
  OAI21_X1 U8415 ( .B1(n6670), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6909), .ZN(
        n6671) );
  INV_X1 U8416 ( .A(n6671), .ZN(n6674) );
  NAND2_X1 U8417 ( .A1(n9845), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6673) );
  AND2_X1 U8418 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7165) );
  AOI21_X1 U8419 ( .B1(n9846), .B2(n6918), .A(n7165), .ZN(n6672) );
  OAI211_X1 U8420 ( .C1(n6674), .C2(n9860), .A(n6673), .B(n6672), .ZN(n6675)
         );
  AOI21_X1 U8421 ( .B1(n9856), .B2(n6676), .A(n6675), .ZN(n6677) );
  OAI21_X1 U8422 ( .B1(n6678), .B2(n9673), .A(n6677), .ZN(P2_U3189) );
  INV_X1 U8423 ( .A(P1_U3973), .ZN(n6680) );
  NAND2_X1 U8424 ( .A1(n6680), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6679) );
  OAI21_X1 U8425 ( .B1(n9202), .B2(n6680), .A(n6679), .ZN(P1_U3581) );
  XNOR2_X1 U8426 ( .A(n6833), .B(n6683), .ZN(n6681) );
  OAI222_X1 U8427 ( .A1(n9349), .A2(n7115), .B1(n6681), .B2(n9299), .C1(n9347), 
        .C2(n6542), .ZN(n9633) );
  INV_X1 U8428 ( .A(n9633), .ZN(n6690) );
  OAI21_X1 U8429 ( .B1(n6684), .B2(n6683), .A(n6682), .ZN(n9635) );
  OAI211_X1 U8430 ( .C1(n4570), .C2(n9632), .A(n9354), .B(n6841), .ZN(n9631)
         );
  AOI22_X1 U8431 ( .A1(n9358), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7123), .B2(
        n9356), .ZN(n6687) );
  NAND2_X1 U8432 ( .A1(n9359), .A2(n7112), .ZN(n6686) );
  OAI211_X1 U8433 ( .C1(n9631), .C2(n9363), .A(n6687), .B(n6686), .ZN(n6688)
         );
  AOI21_X1 U8434 ( .B1(n9635), .B2(n9209), .A(n6688), .ZN(n6689) );
  OAI21_X1 U8435 ( .B1(n6690), .B2(n9358), .A(n6689), .ZN(P1_U3287) );
  INV_X1 U8436 ( .A(n9128), .ZN(n9577) );
  INV_X1 U8437 ( .A(n6691), .ZN(n6694) );
  OAI222_X1 U8438 ( .A1(n9577), .A2(P1_U3086), .B1(n9488), .B2(n6694), .C1(
        n9490), .C2(n6692), .ZN(P1_U3340) );
  INV_X1 U8439 ( .A(n9830), .ZN(n8519) );
  INV_X1 U8440 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6693) );
  OAI222_X1 U8441 ( .A1(n8519), .A2(P2_U3151), .B1(n8947), .B2(n6694), .C1(
        n6693), .C2(n8945), .ZN(P2_U3280) );
  INV_X1 U8442 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7319) );
  OAI21_X1 U8443 ( .B1(n6800), .B2(n6697), .A(n6696), .ZN(n6698) );
  OAI22_X1 U8444 ( .A1(n9673), .A2(n6698), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6879), .ZN(n6707) );
  INV_X1 U8445 ( .A(n6699), .ZN(n6700) );
  AOI21_X1 U8446 ( .B1(n6878), .B2(n6701), .A(n6700), .ZN(n6705) );
  XNOR2_X1 U8447 ( .A(n6703), .B(n6702), .ZN(n6704) );
  OAI22_X1 U8448 ( .A1(n6705), .A2(n9860), .B1(n9664), .B2(n6704), .ZN(n6706)
         );
  AOI211_X1 U8449 ( .C1(n4623), .C2(n9846), .A(n6707), .B(n6706), .ZN(n6708)
         );
  OAI21_X1 U8450 ( .B1(n7319), .B2(n9745), .A(n6708), .ZN(P2_U3183) );
  XNOR2_X1 U8451 ( .A(n6710), .B(n6709), .ZN(n7078) );
  XNOR2_X1 U8452 ( .A(n6711), .B(n7647), .ZN(n6712) );
  AOI222_X1 U8453 ( .A1(n8842), .A2(n6712), .B1(n8471), .B2(n8771), .C1(n5132), 
        .C2(n8769), .ZN(n7079) );
  OAI21_X1 U8454 ( .B1(n6789), .B2(n8847), .A(n7079), .ZN(n6713) );
  AOI21_X1 U8455 ( .B1(n7078), .B2(n7371), .A(n6713), .ZN(n9882) );
  INV_X1 U8456 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6714) );
  OR2_X1 U8457 ( .A1(n8827), .A2(n6714), .ZN(n6715) );
  OAI21_X1 U8458 ( .B1(n9882), .B2(n8857), .A(n6715), .ZN(P2_U3462) );
  INV_X1 U8459 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10063) );
  NOR2_X1 U8460 ( .A1(n6740), .A2(n10063), .ZN(P2_U3263) );
  INV_X1 U8461 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6717) );
  NOR2_X1 U8462 ( .A1(n6740), .A2(n6717), .ZN(P2_U3262) );
  INV_X1 U8463 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6718) );
  NOR2_X1 U8464 ( .A1(n6740), .A2(n6718), .ZN(P2_U3257) );
  INV_X1 U8465 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6719) );
  NOR2_X1 U8466 ( .A1(n6740), .A2(n6719), .ZN(P2_U3255) );
  INV_X1 U8467 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6720) );
  NOR2_X1 U8468 ( .A1(n6740), .A2(n6720), .ZN(P2_U3254) );
  INV_X1 U8469 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6721) );
  NOR2_X1 U8470 ( .A1(n6740), .A2(n6721), .ZN(P2_U3253) );
  INV_X1 U8471 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6722) );
  NOR2_X1 U8472 ( .A1(n6740), .A2(n6722), .ZN(P2_U3256) );
  INV_X1 U8473 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n6723) );
  NOR2_X1 U8474 ( .A1(n6740), .A2(n6723), .ZN(P2_U3252) );
  INV_X1 U8475 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6724) );
  NOR2_X1 U8476 ( .A1(n6740), .A2(n6724), .ZN(P2_U3251) );
  INV_X1 U8477 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6725) );
  NOR2_X1 U8478 ( .A1(n6740), .A2(n6725), .ZN(P2_U3244) );
  INV_X1 U8479 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n6726) );
  NOR2_X1 U8480 ( .A1(n6740), .A2(n6726), .ZN(P2_U3250) );
  INV_X1 U8481 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6727) );
  NOR2_X1 U8482 ( .A1(n6740), .A2(n6727), .ZN(P2_U3248) );
  INV_X1 U8483 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6728) );
  NOR2_X1 U8484 ( .A1(n6740), .A2(n6728), .ZN(P2_U3247) );
  INV_X1 U8485 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n6729) );
  NOR2_X1 U8486 ( .A1(n6740), .A2(n6729), .ZN(P2_U3246) );
  INV_X1 U8487 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n6730) );
  NOR2_X1 U8488 ( .A1(n6740), .A2(n6730), .ZN(P2_U3245) );
  INV_X1 U8489 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6731) );
  NOR2_X1 U8490 ( .A1(n6740), .A2(n6731), .ZN(P2_U3240) );
  INV_X1 U8491 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n6732) );
  NOR2_X1 U8492 ( .A1(n6740), .A2(n6732), .ZN(P2_U3243) );
  INV_X1 U8493 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6733) );
  NOR2_X1 U8494 ( .A1(n6740), .A2(n6733), .ZN(P2_U3242) );
  INV_X1 U8495 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n6734) );
  NOR2_X1 U8496 ( .A1(n6740), .A2(n6734), .ZN(P2_U3241) );
  INV_X1 U8497 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6735) );
  NOR2_X1 U8498 ( .A1(n6740), .A2(n6735), .ZN(P2_U3234) );
  INV_X1 U8499 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9996) );
  NOR2_X1 U8500 ( .A1(n6740), .A2(n9996), .ZN(P2_U3239) );
  INV_X1 U8501 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6736) );
  NOR2_X1 U8502 ( .A1(n6740), .A2(n6736), .ZN(P2_U3238) );
  INV_X1 U8503 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6737) );
  NOR2_X1 U8504 ( .A1(n6740), .A2(n6737), .ZN(P2_U3237) );
  INV_X1 U8505 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6738) );
  NOR2_X1 U8506 ( .A1(n6740), .A2(n6738), .ZN(P2_U3235) );
  INV_X1 U8507 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6739) );
  NOR2_X1 U8508 ( .A1(n6740), .A2(n6739), .ZN(P2_U3236) );
  AOI22_X1 U8509 ( .A1(n9076), .A2(n9106), .B1(n9035), .B2(n6741), .ZN(n6743)
         );
  OAI211_X1 U8510 ( .C1(n6216), .C2(n9078), .A(n6743), .B(n6742), .ZN(n6748)
         );
  AOI211_X1 U8511 ( .C1(n6746), .C2(n6745), .A(n4495), .B(n6744), .ZN(n6747)
         );
  AOI211_X1 U8512 ( .C1(n6749), .C2(n9084), .A(n6748), .B(n6747), .ZN(n6750)
         );
  INV_X1 U8513 ( .A(n6750), .ZN(P1_U3230) );
  INV_X1 U8514 ( .A(n6751), .ZN(n6799) );
  INV_X1 U8515 ( .A(n9590), .ZN(n9137) );
  OAI222_X1 U8516 ( .A1(n9493), .A2(n6799), .B1(n9137), .B2(P1_U3086), .C1(
        n6752), .C2(n9490), .ZN(P1_U3339) );
  NAND2_X1 U8517 ( .A1(n7681), .A2(n8592), .ZN(n6780) );
  NOR2_X1 U8518 ( .A1(n6780), .A2(n4839), .ZN(n6755) );
  NAND2_X1 U8519 ( .A1(n7865), .A2(n6755), .ZN(n7278) );
  NAND3_X1 U8520 ( .A1(n7847), .A2(n7278), .A3(n8847), .ZN(n6790) );
  INV_X1 U8521 ( .A(n7857), .ZN(n7861) );
  NAND2_X1 U8522 ( .A1(n6790), .A2(n9866), .ZN(n7282) );
  INV_X1 U8523 ( .A(n7282), .ZN(n6762) );
  AND2_X1 U8524 ( .A1(n6757), .A2(n6756), .ZN(n6761) );
  INV_X1 U8525 ( .A(n7278), .ZN(n6791) );
  NAND2_X1 U8526 ( .A1(n6773), .A2(n6791), .ZN(n6760) );
  OAI211_X1 U8527 ( .C1(n6768), .C2(n6762), .A(n6761), .B(n6760), .ZN(n6763)
         );
  NAND2_X1 U8528 ( .A1(n6763), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6766) );
  INV_X1 U8529 ( .A(n7279), .ZN(n6826) );
  NAND2_X1 U8530 ( .A1(n6770), .A2(n6826), .ZN(n7864) );
  INV_X1 U8531 ( .A(n7864), .ZN(n6764) );
  NAND2_X1 U8532 ( .A1(n6773), .A2(n6764), .ZN(n6765) );
  NAND2_X1 U8533 ( .A1(n6766), .A2(n6765), .ZN(n6855) );
  OR2_X1 U8534 ( .A1(n6767), .A2(P2_U3151), .ZN(n7866) );
  INV_X1 U8535 ( .A(n7866), .ZN(n7401) );
  INV_X1 U8536 ( .A(n9948), .ZN(n8428) );
  NAND2_X1 U8537 ( .A1(n6768), .A2(n6770), .ZN(n7281) );
  OR2_X1 U8538 ( .A1(n7281), .A2(n9866), .ZN(n6771) );
  AND2_X1 U8539 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9665) );
  AND2_X1 U8540 ( .A1(n7283), .A2(n6826), .ZN(n6774) );
  INV_X1 U8541 ( .A(n5132), .ZN(n6785) );
  INV_X1 U8542 ( .A(n6774), .ZN(n6776) );
  OAI22_X1 U8543 ( .A1(n8440), .A2(n6785), .B1(n7007), .B2(n8427), .ZN(n6777)
         );
  AOI211_X1 U8544 ( .C1(n7082), .C2(n9950), .A(n9665), .B(n6777), .ZN(n6798)
         );
  XNOR2_X1 U8545 ( .A(n6781), .B(n8473), .ZN(n6854) );
  OAI21_X1 U8546 ( .B1(n6784), .B2(n8228), .A(n7682), .ZN(n6853) );
  NAND2_X1 U8547 ( .A1(n6854), .A2(n6853), .ZN(n6783) );
  NAND2_X1 U8548 ( .A1(n6781), .A2(n5118), .ZN(n6782) );
  NAND2_X1 U8549 ( .A1(n6783), .A2(n6782), .ZN(n6864) );
  XNOR2_X1 U8550 ( .A(n6784), .B(n6865), .ZN(n6786) );
  XNOR2_X1 U8551 ( .A(n6786), .B(n5132), .ZN(n6863) );
  NAND2_X1 U8552 ( .A1(n6864), .A2(n6863), .ZN(n6788) );
  NAND2_X1 U8553 ( .A1(n6786), .A2(n6785), .ZN(n6787) );
  NAND2_X1 U8554 ( .A1(n6788), .A2(n6787), .ZN(n6795) );
  XNOR2_X1 U8555 ( .A(n6784), .B(n6789), .ZN(n6926) );
  XNOR2_X1 U8556 ( .A(n6926), .B(n8472), .ZN(n6794) );
  OR2_X1 U8557 ( .A1(n7281), .A2(n6790), .ZN(n6793) );
  NAND2_X1 U8558 ( .A1(n7283), .A2(n6791), .ZN(n6792) );
  AOI21_X1 U8559 ( .B1(n6795), .B2(n6794), .A(n8410), .ZN(n6796) );
  NAND2_X1 U8560 ( .A1(n6796), .A2(n6928), .ZN(n6797) );
  OAI211_X1 U8561 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8428), .A(n6798), .B(
        n6797), .ZN(P2_U3158) );
  INV_X1 U8562 ( .A(n9847), .ZN(n8517) );
  OAI222_X1 U8563 ( .A1(n8945), .A2(n10068), .B1(P2_U3151), .B2(n8517), .C1(
        n6799), .C2(n8947), .ZN(P2_U3279) );
  INV_X1 U8564 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6807) );
  OAI21_X1 U8565 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6801), .A(n6800), .ZN(n6802) );
  OAI21_X1 U8566 ( .B1(n9855), .B2(n6803), .A(n6802), .ZN(n6804) );
  OAI21_X1 U8567 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6824), .A(n6804), .ZN(n6805) );
  AOI21_X1 U8568 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9846), .A(n6805), .ZN(n6806) );
  OAI21_X1 U8569 ( .B1(n9745), .B2(n6807), .A(n6806), .ZN(P2_U3182) );
  XNOR2_X1 U8570 ( .A(n8470), .B(n7699), .ZN(n7649) );
  INV_X1 U8571 ( .A(n7649), .ZN(n6808) );
  XNOR2_X1 U8572 ( .A(n6809), .B(n6808), .ZN(n6888) );
  XNOR2_X1 U8573 ( .A(n6810), .B(n7649), .ZN(n6812) );
  OAI22_X1 U8574 ( .A1(n7163), .A2(n8838), .B1(n7007), .B2(n8840), .ZN(n6811)
         );
  AOI21_X1 U8575 ( .B1(n6812), .B2(n8842), .A(n6811), .ZN(n6813) );
  OAI21_X1 U8576 ( .B1(n6888), .B2(n7178), .A(n6813), .ZN(n6884) );
  OAI22_X1 U8577 ( .A1(n6888), .A2(n8846), .B1(n7704), .B2(n8847), .ZN(n6814)
         );
  NOR2_X1 U8578 ( .A1(n6884), .A2(n6814), .ZN(n9886) );
  INV_X1 U8579 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6815) );
  OR2_X1 U8580 ( .A1(n8827), .A2(n6815), .ZN(n6816) );
  OAI21_X1 U8581 ( .B1(n9886), .B2(n8857), .A(n6816), .ZN(P2_U3464) );
  INV_X1 U8582 ( .A(n6817), .ZN(n6822) );
  INV_X1 U8583 ( .A(n6818), .ZN(n6819) );
  NOR2_X1 U8584 ( .A1(n9869), .A2(n6824), .ZN(n6825) );
  AOI21_X1 U8585 ( .B1(n8778), .B2(n8228), .A(n6825), .ZN(n6831) );
  INV_X1 U8586 ( .A(n8229), .ZN(n6827) );
  NOR3_X1 U8587 ( .A1(n6827), .A2(n8852), .A3(n6826), .ZN(n6828) );
  OAI21_X1 U8588 ( .B1(n6829), .B2(n6828), .A(n8693), .ZN(n6830) );
  OAI211_X1 U8589 ( .C1(n6832), .C2(n8693), .A(n6831), .B(n6830), .ZN(P2_U3233) );
  INV_X1 U8590 ( .A(n6838), .ZN(n6835) );
  AOI21_X1 U8591 ( .B1(n4702), .B2(n6260), .A(n7986), .ZN(n6834) );
  NAND2_X1 U8592 ( .A1(n6834), .A2(n6835), .ZN(n6944) );
  OAI21_X1 U8593 ( .B1(n6835), .B2(n6834), .A(n6944), .ZN(n6836) );
  AOI222_X1 U8594 ( .A1(n9352), .A2(n6836), .B1(n9103), .B2(n9337), .C1(n9105), 
        .C2(n9335), .ZN(n6939) );
  OAI21_X1 U8595 ( .B1(n6839), .B2(n6838), .A(n6837), .ZN(n6941) );
  INV_X1 U8596 ( .A(n6840), .ZN(n6952) );
  AOI21_X1 U8597 ( .B1(n6841), .B2(n7107), .A(n9326), .ZN(n6842) );
  NAND2_X1 U8598 ( .A1(n6952), .A2(n6842), .ZN(n6938) );
  INV_X1 U8599 ( .A(n7101), .ZN(n6843) );
  OAI22_X1 U8600 ( .A1(n9365), .A2(n6417), .B1(n6843), .B2(n9211), .ZN(n6844)
         );
  AOI21_X1 U8601 ( .B1(n9359), .B2(n7107), .A(n6844), .ZN(n6845) );
  OAI21_X1 U8602 ( .B1(n6938), .B2(n9363), .A(n6845), .ZN(n6846) );
  AOI21_X1 U8603 ( .B1(n6941), .B2(n9209), .A(n6846), .ZN(n6847) );
  OAI21_X1 U8604 ( .B1(n6939), .B2(n9358), .A(n6847), .ZN(P1_U3286) );
  AND2_X1 U8605 ( .A1(n7702), .A2(n7710), .ZN(n7697) );
  XNOR2_X1 U8606 ( .A(n6848), .B(n7697), .ZN(n7133) );
  XNOR2_X1 U8607 ( .A(n6849), .B(n7697), .ZN(n6850) );
  AOI222_X1 U8608 ( .A1(n8842), .A2(n6850), .B1(n8470), .B2(n8771), .C1(n8472), 
        .C2(n8769), .ZN(n7134) );
  OAI21_X1 U8609 ( .B1(n6934), .B2(n8847), .A(n7134), .ZN(n6851) );
  AOI21_X1 U8610 ( .B1(n7133), .B2(n7371), .A(n6851), .ZN(n9884) );
  NAND2_X1 U8611 ( .A1(n8857), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6852) );
  OAI21_X1 U8612 ( .B1(n9884), .B2(n8857), .A(n6852), .ZN(P2_U3463) );
  XOR2_X1 U8613 ( .A(n6854), .B(n6853), .Z(n6862) );
  INV_X1 U8614 ( .A(n6855), .ZN(n6857) );
  NAND2_X1 U8615 ( .A1(n6857), .A2(n6856), .ZN(n8230) );
  AOI22_X1 U8616 ( .A1(n9952), .A2(n5132), .B1(n8851), .B2(n9950), .ZN(n6858)
         );
  OAI21_X1 U8617 ( .B1(n6859), .B2(n8440), .A(n6858), .ZN(n6860) );
  AOI21_X1 U8618 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n8230), .A(n6860), .ZN(
        n6861) );
  OAI21_X1 U8619 ( .B1(n8410), .B2(n6862), .A(n6861), .ZN(P2_U3162) );
  XOR2_X1 U8620 ( .A(n6864), .B(n6863), .Z(n6869) );
  AOI22_X1 U8621 ( .A1(n9952), .A2(n8472), .B1(n6865), .B2(n9950), .ZN(n6866)
         );
  OAI21_X1 U8622 ( .B1(n5118), .B2(n8440), .A(n6866), .ZN(n6867) );
  AOI21_X1 U8623 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n8230), .A(n6867), .ZN(
        n6868) );
  OAI21_X1 U8624 ( .B1(n6869), .B2(n8410), .A(n6868), .ZN(P2_U3177) );
  NAND2_X1 U8625 ( .A1(n5528), .A2(n7682), .ZN(n6870) );
  NAND2_X1 U8626 ( .A1(n6871), .A2(n6870), .ZN(n8854) );
  INV_X1 U8627 ( .A(n8854), .ZN(n6883) );
  NAND2_X1 U8628 ( .A1(n6872), .A2(n7857), .ZN(n7067) );
  INV_X1 U8629 ( .A(n7067), .ZN(n9874) );
  NAND2_X1 U8630 ( .A1(n8693), .A2(n9874), .ZN(n7182) );
  INV_X1 U8631 ( .A(n7178), .ZN(n8835) );
  NAND2_X1 U8632 ( .A1(n8854), .A2(n8835), .ZN(n6877) );
  AOI22_X1 U8633 ( .A1(n8769), .A2(n8475), .B1(n5132), .B2(n8771), .ZN(n6876)
         );
  XNOR2_X1 U8634 ( .A(n5528), .B(n6873), .ZN(n6874) );
  NAND2_X1 U8635 ( .A1(n6874), .A2(n8842), .ZN(n6875) );
  AND3_X1 U8636 ( .A1(n6877), .A2(n6876), .A3(n6875), .ZN(n8856) );
  MUX2_X1 U8637 ( .A(n8856), .B(n6878), .S(n9876), .Z(n6882) );
  NOR2_X1 U8638 ( .A1(n9869), .A2(n6879), .ZN(n6880) );
  AOI21_X1 U8639 ( .B1(n8778), .B2(n8851), .A(n6880), .ZN(n6881) );
  OAI211_X1 U8640 ( .C1(n6883), .C2(n7182), .A(n6882), .B(n6881), .ZN(P2_U3232) );
  NAND2_X1 U8641 ( .A1(n6884), .A2(n8693), .ZN(n6887) );
  OAI22_X1 U8642 ( .A1(n8613), .A2(n7704), .B1(n7012), .B2(n9869), .ZN(n6885)
         );
  AOI21_X1 U8643 ( .B1(n9876), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6885), .ZN(
        n6886) );
  OAI211_X1 U8644 ( .C1(n6888), .C2(n7182), .A(n6887), .B(n6886), .ZN(P2_U3228) );
  NOR2_X1 U8645 ( .A1(n4407), .A2(n4351), .ZN(n6890) );
  XNOR2_X1 U8646 ( .A(n6890), .B(n6889), .ZN(n6898) );
  INV_X1 U8647 ( .A(n6891), .ZN(n6894) );
  OAI22_X1 U8648 ( .A1(n9080), .A2(n6990), .B1(n6892), .B2(n9068), .ZN(n6893)
         );
  AOI211_X1 U8649 ( .C1(n9061), .C2(n9107), .A(n6894), .B(n6893), .ZN(n6897)
         );
  NAND2_X1 U8650 ( .A1(n9084), .A2(n6895), .ZN(n6896) );
  OAI211_X1 U8651 ( .C1(n6898), .C2(n4495), .A(n6897), .B(n6896), .ZN(P1_U3227) );
  MUX2_X1 U8652 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6899), .S(n8533), .Z(n6906)
         );
  NAND2_X1 U8653 ( .A1(n6900), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6904) );
  NAND2_X1 U8654 ( .A1(n6902), .A2(n6901), .ZN(n6903) );
  NAND2_X1 U8655 ( .A1(n6904), .A2(n6903), .ZN(n6905) );
  NAND2_X1 U8656 ( .A1(n6905), .A2(n6906), .ZN(n8505) );
  OAI21_X1 U8657 ( .B1(n6906), .B2(n6905), .A(n8505), .ZN(n6924) );
  MUX2_X1 U8658 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n5210), .S(n8533), .Z(n6907)
         );
  NAND3_X1 U8659 ( .A1(n6909), .A2(n4677), .A3(n6908), .ZN(n6910) );
  AND2_X1 U8660 ( .A1(n8492), .A2(n6910), .ZN(n6915) );
  NAND2_X1 U8661 ( .A1(n9845), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n6914) );
  INV_X1 U8662 ( .A(n8533), .ZN(n6912) );
  INV_X1 U8663 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6911) );
  NOR2_X1 U8664 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6911), .ZN(n7218) );
  AOI21_X1 U8665 ( .B1(n9846), .B2(n6912), .A(n7218), .ZN(n6913) );
  OAI211_X1 U8666 ( .C1(n6915), .C2(n9860), .A(n6914), .B(n6913), .ZN(n6923)
         );
  MUX2_X1 U8667 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8588), .Z(n8534) );
  XNOR2_X1 U8668 ( .A(n8534), .B(n8533), .ZN(n8535) );
  INV_X1 U8669 ( .A(n6916), .ZN(n6917) );
  AOI22_X1 U8670 ( .A1(n6920), .A2(n6919), .B1(n6918), .B2(n6917), .ZN(n8536)
         );
  XOR2_X1 U8671 ( .A(n8535), .B(n8536), .Z(n6921) );
  NOR2_X1 U8672 ( .A1(n6921), .A2(n9673), .ZN(n6922) );
  AOI211_X1 U8673 ( .C1(n9856), .C2(n6924), .A(n6923), .B(n6922), .ZN(n6925)
         );
  INV_X1 U8674 ( .A(n6925), .ZN(P2_U3190) );
  XNOR2_X1 U8675 ( .A(n6784), .B(n6934), .ZN(n7002) );
  XNOR2_X1 U8676 ( .A(n7002), .B(n8471), .ZN(n6931) );
  NAND2_X1 U8677 ( .A1(n6926), .A2(n8472), .ZN(n6927) );
  INV_X1 U8678 ( .A(n7005), .ZN(n6929) );
  AOI21_X1 U8679 ( .B1(n6931), .B2(n6930), .A(n6929), .ZN(n6937) );
  INV_X1 U8680 ( .A(n6932), .ZN(n7136) );
  AOI22_X1 U8681 ( .A1(n9952), .A2(n8470), .B1(n9945), .B2(n8472), .ZN(n6933)
         );
  NAND2_X1 U8682 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n9684) );
  OAI211_X1 U8683 ( .C1(n6934), .C2(n8458), .A(n6933), .B(n9684), .ZN(n6935)
         );
  AOI21_X1 U8684 ( .B1(n7136), .B2(n9948), .A(n6935), .ZN(n6936) );
  OAI21_X1 U8685 ( .B1(n6937), .B2(n8410), .A(n6936), .ZN(P2_U3170) );
  NAND2_X1 U8686 ( .A1(n6939), .A2(n6938), .ZN(n6940) );
  AOI21_X1 U8687 ( .B1(n9648), .B2(n6941), .A(n6940), .ZN(n6961) );
  AOI22_X1 U8688 ( .A1(n9414), .A2(n7107), .B1(n9656), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n6942) );
  OAI21_X1 U8689 ( .B1(n6961), .B2(n9656), .A(n6942), .ZN(P1_U3529) );
  INV_X1 U8690 ( .A(n6949), .ZN(n6946) );
  NAND2_X1 U8691 ( .A1(n6944), .A2(n6943), .ZN(n6945) );
  NAND2_X1 U8692 ( .A1(n6945), .A2(n6946), .ZN(n7016) );
  OAI21_X1 U8693 ( .B1(n6946), .B2(n6945), .A(n7016), .ZN(n6947) );
  AOI222_X1 U8694 ( .A1(n9352), .A2(n6947), .B1(n9102), .B2(n9337), .C1(n9104), 
        .C2(n9335), .ZN(n7057) );
  OAI21_X1 U8695 ( .B1(n6950), .B2(n6949), .A(n6948), .ZN(n7060) );
  INV_X1 U8696 ( .A(n7022), .ZN(n6951) );
  AOI211_X1 U8697 ( .C1(n7061), .C2(n6952), .A(n9326), .B(n6951), .ZN(n7059)
         );
  NAND2_X1 U8698 ( .A1(n7059), .A2(n9342), .ZN(n6954) );
  AOI22_X1 U8699 ( .A1(n9358), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7198), .B2(
        n9356), .ZN(n6953) );
  OAI211_X1 U8700 ( .C1(n7195), .C2(n9330), .A(n6954), .B(n6953), .ZN(n6955)
         );
  AOI21_X1 U8701 ( .B1(n7060), .B2(n9209), .A(n6955), .ZN(n6956) );
  OAI21_X1 U8702 ( .B1(n7057), .B2(n9358), .A(n6956), .ZN(P1_U3285) );
  INV_X1 U8703 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6957) );
  OAI22_X1 U8704 ( .A1(n9445), .A2(n6958), .B1(n9480), .B2(n6957), .ZN(n6959)
         );
  INV_X1 U8705 ( .A(n6959), .ZN(n6960) );
  OAI21_X1 U8706 ( .B1(n6961), .B2(n6284), .A(n6960), .ZN(P1_U3474) );
  XNOR2_X1 U8707 ( .A(n6962), .B(n7650), .ZN(n7069) );
  INV_X1 U8708 ( .A(n7650), .ZN(n6963) );
  XNOR2_X1 U8709 ( .A(n6964), .B(n6963), .ZN(n6967) );
  NAND2_X1 U8710 ( .A1(n8470), .A2(n8769), .ZN(n6965) );
  OAI21_X1 U8711 ( .B1(n7216), .B2(n8838), .A(n6965), .ZN(n6966) );
  AOI21_X1 U8712 ( .B1(n6967), .B2(n8842), .A(n6966), .ZN(n7070) );
  OAI21_X1 U8713 ( .B1(n7045), .B2(n8847), .A(n7070), .ZN(n6968) );
  AOI21_X1 U8714 ( .B1(n7069), .B2(n7371), .A(n6968), .ZN(n9888) );
  OR2_X1 U8715 ( .A1(n8827), .A2(n6664), .ZN(n6969) );
  OAI21_X1 U8716 ( .B1(n9888), .B2(n8857), .A(n6969), .ZN(P2_U3465) );
  INV_X1 U8717 ( .A(n9478), .ZN(n6992) );
  INV_X1 U8718 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10042) );
  OAI22_X1 U8719 ( .A1(n9445), .A2(n6562), .B1(n9480), .B2(n10042), .ZN(n6970)
         );
  AOI21_X1 U8720 ( .B1(n6992), .B2(n6971), .A(n6970), .ZN(n6972) );
  OAI21_X1 U8721 ( .B1(n6973), .B2(n6284), .A(n6972), .ZN(P1_U3462) );
  OAI211_X1 U8722 ( .C1(n8110), .C2(n7592), .A(n9354), .B(n6976), .ZN(n7886)
         );
  INV_X1 U8723 ( .A(n7886), .ZN(n6981) );
  XNOR2_X1 U8724 ( .A(n7943), .B(n6977), .ZN(n6978) );
  NAND2_X1 U8725 ( .A1(n6978), .A2(n9352), .ZN(n6980) );
  AOI22_X1 U8726 ( .A1(n9335), .A2(n9110), .B1(n6213), .B2(n9337), .ZN(n6979)
         );
  NAND2_X1 U8727 ( .A1(n6980), .A2(n6979), .ZN(n7889) );
  AOI211_X1 U8728 ( .C1(n9648), .C2(n7884), .A(n6981), .B(n7889), .ZN(n7883)
         );
  INV_X1 U8729 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6982) );
  OAI22_X1 U8730 ( .A1(n9445), .A2(n8110), .B1(n9480), .B2(n6982), .ZN(n6983)
         );
  INV_X1 U8731 ( .A(n6983), .ZN(n6984) );
  OAI21_X1 U8732 ( .B1(n7883), .B2(n6284), .A(n6984), .ZN(P1_U3456) );
  INV_X1 U8733 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6985) );
  OAI22_X1 U8734 ( .A1(n9445), .A2(n6212), .B1(n9480), .B2(n6985), .ZN(n6986)
         );
  INV_X1 U8735 ( .A(n6986), .ZN(n6987) );
  OAI21_X1 U8736 ( .B1(n6988), .B2(n6284), .A(n6987), .ZN(P1_U3459) );
  INV_X1 U8737 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6989) );
  OAI22_X1 U8738 ( .A1(n9445), .A2(n6990), .B1(n9650), .B2(n6989), .ZN(n6991)
         );
  AOI21_X1 U8739 ( .B1(n6993), .B2(n6992), .A(n6991), .ZN(n6994) );
  OAI21_X1 U8740 ( .B1(n6995), .B2(n6284), .A(n6994), .ZN(P1_U3468) );
  INV_X1 U8741 ( .A(n6996), .ZN(n6999) );
  INV_X1 U8742 ( .A(n9600), .ZN(n9149) );
  OAI222_X1 U8743 ( .A1(n9490), .A2(n6997), .B1(n9488), .B2(n6999), .C1(
        P1_U3086), .C2(n9149), .ZN(P1_U3338) );
  OAI222_X1 U8744 ( .A1(n8576), .A2(P2_U3151), .B1(n8947), .B2(n6999), .C1(
        n6998), .C2(n8945), .ZN(P2_U3278) );
  INV_X1 U8745 ( .A(n7000), .ZN(n7013) );
  INV_X1 U8746 ( .A(n9150), .ZN(n9615) );
  OAI222_X1 U8747 ( .A1(n9493), .A2(n7013), .B1(n9615), .B2(P1_U3086), .C1(
        n7001), .C2(n9490), .ZN(P1_U3337) );
  INV_X1 U8748 ( .A(n7002), .ZN(n7003) );
  NAND2_X1 U8749 ( .A1(n7003), .A2(n7007), .ZN(n7004) );
  XNOR2_X1 U8750 ( .A(n6784), .B(n7704), .ZN(n7041) );
  XNOR2_X1 U8751 ( .A(n7041), .B(n7700), .ZN(n7043) );
  XNOR2_X1 U8752 ( .A(n7044), .B(n7043), .ZN(n7006) );
  NAND2_X1 U8753 ( .A1(n7006), .A2(n9958), .ZN(n7011) );
  OAI22_X1 U8754 ( .A1(n8440), .A2(n7007), .B1(n7163), .B2(n8427), .ZN(n7008)
         );
  AOI211_X1 U8755 ( .C1(n7699), .C2(n9950), .A(n7009), .B(n7008), .ZN(n7010)
         );
  OAI211_X1 U8756 ( .C1(n7012), .C2(n8428), .A(n7011), .B(n7010), .ZN(P2_U3167) );
  INV_X1 U8757 ( .A(n8586), .ZN(n8596) );
  OAI222_X1 U8758 ( .A1(n8945), .A2(n7014), .B1(n8947), .B2(n7013), .C1(
        P2_U3151), .C2(n8596), .ZN(P2_U3277) );
  NAND2_X1 U8759 ( .A1(n7016), .A2(n7015), .ZN(n7017) );
  XNOR2_X1 U8760 ( .A(n7017), .B(n7020), .ZN(n7018) );
  OAI22_X1 U8761 ( .A1(n7018), .A2(n9299), .B1(n7105), .B2(n9347), .ZN(n9639)
         );
  INV_X1 U8762 ( .A(n9639), .ZN(n7029) );
  OAI21_X1 U8763 ( .B1(n7021), .B2(n7020), .A(n7019), .ZN(n9641) );
  XNOR2_X1 U8764 ( .A(n7022), .B(n9638), .ZN(n7023) );
  INV_X1 U8765 ( .A(n9046), .ZN(n9101) );
  AOI22_X1 U8766 ( .A1(n7023), .A2(n9354), .B1(n9337), .B2(n9101), .ZN(n9637)
         );
  AOI22_X1 U8767 ( .A1(n9358), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7298), .B2(
        n9356), .ZN(n7026) );
  NAND2_X1 U8768 ( .A1(n7024), .A2(n9359), .ZN(n7025) );
  OAI211_X1 U8769 ( .C1(n9637), .C2(n9363), .A(n7026), .B(n7025), .ZN(n7027)
         );
  AOI21_X1 U8770 ( .B1(n9641), .B2(n9209), .A(n7027), .ZN(n7028) );
  OAI21_X1 U8771 ( .B1(n9358), .B2(n7029), .A(n7028), .ZN(P1_U3284) );
  NAND2_X1 U8772 ( .A1(n7031), .A2(n5207), .ZN(n7032) );
  NAND2_X1 U8773 ( .A1(n7030), .A2(n7032), .ZN(n7056) );
  OAI21_X1 U8774 ( .B1(n7034), .B2(n5207), .A(n7033), .ZN(n7036) );
  OAI22_X1 U8775 ( .A1(n7163), .A2(n8840), .B1(n7237), .B2(n8838), .ZN(n7035)
         );
  AOI21_X1 U8776 ( .B1(n7036), .B2(n8842), .A(n7035), .ZN(n7037) );
  OAI21_X1 U8777 ( .B1(n7178), .B2(n7056), .A(n7037), .ZN(n7052) );
  OAI22_X1 U8778 ( .A1(n7056), .A2(n8846), .B1(n7154), .B2(n8847), .ZN(n7038)
         );
  NOR2_X1 U8779 ( .A1(n7052), .A2(n7038), .ZN(n9890) );
  INV_X1 U8780 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7039) );
  OR2_X1 U8781 ( .A1(n8827), .A2(n7039), .ZN(n7040) );
  OAI21_X1 U8782 ( .B1(n9890), .B2(n8857), .A(n7040), .ZN(P2_U3466) );
  INV_X1 U8783 ( .A(n7041), .ZN(n7042) );
  XNOR2_X1 U8784 ( .A(n6784), .B(n7045), .ZN(n7155) );
  XNOR2_X1 U8785 ( .A(n7155), .B(n7163), .ZN(n7046) );
  NAND2_X1 U8786 ( .A1(n7047), .A2(n7046), .ZN(n7157) );
  OAI211_X1 U8787 ( .C1(n7047), .C2(n7046), .A(n7157), .B(n9958), .ZN(n7051)
         );
  INV_X1 U8788 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7048) );
  NOR2_X1 U8789 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7048), .ZN(n9715) );
  OAI22_X1 U8790 ( .A1(n8440), .A2(n7700), .B1(n7216), .B2(n8427), .ZN(n7049)
         );
  AOI211_X1 U8791 ( .C1(n7074), .C2(n9950), .A(n9715), .B(n7049), .ZN(n7050)
         );
  OAI211_X1 U8792 ( .C1(n7072), .C2(n8428), .A(n7051), .B(n7050), .ZN(P2_U3179) );
  NAND2_X1 U8793 ( .A1(n7052), .A2(n8693), .ZN(n7055) );
  OAI22_X1 U8794 ( .A1(n8613), .A2(n7154), .B1(n7167), .B2(n9869), .ZN(n7053)
         );
  AOI21_X1 U8795 ( .B1(n9876), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7053), .ZN(
        n7054) );
  OAI211_X1 U8796 ( .C1(n7056), .C2(n7182), .A(n7055), .B(n7054), .ZN(P2_U3226) );
  INV_X1 U8797 ( .A(n7057), .ZN(n7058) );
  AOI211_X1 U8798 ( .C1(n9648), .C2(n7060), .A(n7059), .B(n7058), .ZN(n7066)
         );
  AOI22_X1 U8799 ( .A1(n9414), .A2(n7061), .B1(n9656), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7062) );
  OAI21_X1 U8800 ( .B1(n7066), .B2(n9656), .A(n7062), .ZN(P1_U3530) );
  INV_X1 U8801 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7063) );
  OAI22_X1 U8802 ( .A1(n9445), .A2(n7195), .B1(n9480), .B2(n7063), .ZN(n7064)
         );
  INV_X1 U8803 ( .A(n7064), .ZN(n7065) );
  OAI21_X1 U8804 ( .B1(n7066), .B2(n6284), .A(n7065), .ZN(P1_U3477) );
  NAND2_X1 U8805 ( .A1(n7178), .A2(n7067), .ZN(n7068) );
  INV_X1 U8806 ( .A(n7069), .ZN(n7077) );
  MUX2_X1 U8807 ( .A(n7071), .B(n7070), .S(n8693), .Z(n7076) );
  INV_X1 U8808 ( .A(n7072), .ZN(n7073) );
  AOI22_X1 U8809 ( .A1(n8778), .A2(n7074), .B1(n8777), .B2(n7073), .ZN(n7075)
         );
  OAI211_X1 U8810 ( .C1(n8765), .C2(n7077), .A(n7076), .B(n7075), .ZN(P2_U3227) );
  INV_X1 U8811 ( .A(n7078), .ZN(n7085) );
  MUX2_X1 U8812 ( .A(n7080), .B(n7079), .S(n8693), .Z(n7084) );
  AOI22_X1 U8813 ( .A1(n8778), .A2(n7082), .B1(n8777), .B2(n7081), .ZN(n7083)
         );
  OAI211_X1 U8814 ( .C1(n8765), .C2(n7085), .A(n7084), .B(n7083), .ZN(P2_U3230) );
  NAND2_X1 U8815 ( .A1(n7030), .A2(n7086), .ZN(n7087) );
  XNOR2_X1 U8816 ( .A(n7087), .B(n7652), .ZN(n7127) );
  INV_X1 U8817 ( .A(n7127), .ZN(n7097) );
  NAND2_X1 U8818 ( .A1(n7088), .A2(n8842), .ZN(n7092) );
  AOI21_X1 U8819 ( .B1(n7033), .B2(n7089), .A(n7652), .ZN(n7091) );
  AOI22_X1 U8820 ( .A1(n8468), .A2(n8769), .B1(n8771), .B2(n8466), .ZN(n7090)
         );
  OAI21_X1 U8821 ( .B1(n7092), .B2(n7091), .A(n7090), .ZN(n7125) );
  NOR2_X1 U8822 ( .A1(n8693), .A2(n5210), .ZN(n7095) );
  NAND2_X1 U8823 ( .A1(n8778), .A2(n7219), .ZN(n7093) );
  OAI21_X1 U8824 ( .B1(n7222), .B2(n9869), .A(n7093), .ZN(n7094) );
  AOI211_X1 U8825 ( .C1(n7125), .C2(n8693), .A(n7095), .B(n7094), .ZN(n7096)
         );
  OAI21_X1 U8826 ( .B1(n7097), .B2(n8765), .A(n7096), .ZN(P2_U3225) );
  NAND2_X1 U8827 ( .A1(n4410), .A2(n7099), .ZN(n7100) );
  XNOR2_X1 U8828 ( .A(n7098), .B(n7100), .ZN(n7109) );
  NAND2_X1 U8829 ( .A1(n9084), .A2(n7101), .ZN(n7104) );
  AOI21_X1 U8830 ( .B1(n9061), .B2(n9105), .A(n7102), .ZN(n7103) );
  OAI211_X1 U8831 ( .C1(n7105), .C2(n9068), .A(n7104), .B(n7103), .ZN(n7106)
         );
  AOI21_X1 U8832 ( .B1(n7107), .B2(n9035), .A(n7106), .ZN(n7108) );
  OAI21_X1 U8833 ( .B1(n7109), .B2(n4495), .A(n7108), .ZN(P1_U3213) );
  INV_X1 U8834 ( .A(n7110), .ZN(n7111) );
  AOI21_X1 U8835 ( .B1(n9061), .B2(n9106), .A(n7111), .ZN(n7114) );
  NAND2_X1 U8836 ( .A1(n9035), .A2(n7112), .ZN(n7113) );
  OAI211_X1 U8837 ( .C1(n7115), .C2(n9068), .A(n7114), .B(n7113), .ZN(n7122)
         );
  XNOR2_X1 U8838 ( .A(n7118), .B(n7117), .ZN(n7119) );
  XNOR2_X1 U8839 ( .A(n7116), .B(n7119), .ZN(n7120) );
  NOR2_X1 U8840 ( .A1(n7120), .A2(n4495), .ZN(n7121) );
  AOI211_X1 U8841 ( .C1(n7123), .C2(n9084), .A(n7122), .B(n7121), .ZN(n7124)
         );
  INV_X1 U8842 ( .A(n7124), .ZN(P1_U3239) );
  NOR2_X1 U8843 ( .A1(n7213), .A2(n8847), .ZN(n7126) );
  AOI211_X1 U8844 ( .C1(n7371), .C2(n7127), .A(n7126), .B(n7125), .ZN(n9891)
         );
  NAND2_X1 U8845 ( .A1(n8857), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7128) );
  OAI21_X1 U8846 ( .B1(n9891), .B2(n8857), .A(n7128), .ZN(P2_U3467) );
  INV_X1 U8847 ( .A(n7129), .ZN(n8189) );
  OAI222_X1 U8848 ( .A1(n7131), .A2(P2_U3151), .B1(n8947), .B2(n8189), .C1(
        n7130), .C2(n8945), .ZN(P2_U3276) );
  NAND2_X1 U8849 ( .A1(n8474), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7132) );
  OAI21_X1 U8850 ( .B1(n7838), .B2(n8474), .A(n7132), .ZN(P2_U3521) );
  INV_X1 U8851 ( .A(n7133), .ZN(n7140) );
  MUX2_X1 U8852 ( .A(n7135), .B(n7134), .S(n8693), .Z(n7139) );
  AOI22_X1 U8853 ( .A1(n8778), .A2(n7137), .B1(n8777), .B2(n7136), .ZN(n7138)
         );
  OAI211_X1 U8854 ( .C1(n8765), .C2(n7140), .A(n7139), .B(n7138), .ZN(P2_U3229) );
  OAI21_X1 U8855 ( .B1(n4408), .B2(n7141), .A(n7464), .ZN(n7143) );
  OAI22_X1 U8856 ( .A1(n7454), .A2(n9347), .B1(n7391), .B2(n9349), .ZN(n7142)
         );
  AOI21_X1 U8857 ( .B1(n7143), .B2(n9352), .A(n7142), .ZN(n9644) );
  OAI21_X1 U8858 ( .B1(n7145), .B2(n7951), .A(n4518), .ZN(n9649) );
  NAND2_X1 U8859 ( .A1(n9649), .A2(n9209), .ZN(n7153) );
  INV_X1 U8860 ( .A(n7146), .ZN(n7148) );
  INV_X1 U8861 ( .A(n7460), .ZN(n7147) );
  OAI211_X1 U8862 ( .C1(n9646), .C2(n7148), .A(n7147), .B(n9354), .ZN(n9643)
         );
  INV_X1 U8863 ( .A(n9643), .ZN(n7151) );
  AOI22_X1 U8864 ( .A1(n9358), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7457), .B2(
        n9356), .ZN(n7149) );
  OAI21_X1 U8865 ( .B1(n9646), .B2(n9330), .A(n7149), .ZN(n7150) );
  AOI21_X1 U8866 ( .B1(n7151), .B2(n9342), .A(n7150), .ZN(n7152) );
  OAI211_X1 U8867 ( .C1(n9358), .C2(n9644), .A(n7153), .B(n7152), .ZN(P1_U3283) );
  XNOR2_X1 U8868 ( .A(n6784), .B(n7154), .ZN(n7209) );
  XNOR2_X1 U8869 ( .A(n7209), .B(n8468), .ZN(n7162) );
  NAND2_X1 U8870 ( .A1(n7155), .A2(n8469), .ZN(n7156) );
  NAND2_X1 U8871 ( .A1(n7157), .A2(n7156), .ZN(n7161) );
  INV_X1 U8872 ( .A(n7212), .ZN(n7160) );
  AOI21_X1 U8873 ( .B1(n7162), .B2(n7161), .A(n7160), .ZN(n7171) );
  OAI22_X1 U8874 ( .A1(n8440), .A2(n7163), .B1(n7237), .B2(n8427), .ZN(n7164)
         );
  AOI211_X1 U8875 ( .C1(n7166), .C2(n9950), .A(n7165), .B(n7164), .ZN(n7170)
         );
  INV_X1 U8876 ( .A(n7167), .ZN(n7168) );
  NAND2_X1 U8877 ( .A1(n9948), .A2(n7168), .ZN(n7169) );
  OAI211_X1 U8878 ( .C1(n7171), .C2(n8410), .A(n7170), .B(n7169), .ZN(P2_U3153) );
  NAND2_X1 U8879 ( .A1(n7172), .A2(n7653), .ZN(n7173) );
  NAND2_X1 U8880 ( .A1(n7201), .A2(n7173), .ZN(n7185) );
  XOR2_X1 U8881 ( .A(n7174), .B(n7653), .Z(n7175) );
  NAND2_X1 U8882 ( .A1(n7175), .A2(n8842), .ZN(n7177) );
  AOI22_X1 U8883 ( .A1(n8467), .A2(n8769), .B1(n8771), .B2(n9944), .ZN(n7176)
         );
  OAI211_X1 U8884 ( .C1(n7178), .C2(n7185), .A(n7177), .B(n7176), .ZN(n7187)
         );
  NAND2_X1 U8885 ( .A1(n7187), .A2(n8693), .ZN(n7181) );
  INV_X1 U8886 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9728) );
  OAI22_X1 U8887 ( .A1(n8693), .A2(n9728), .B1(n7242), .B2(n9869), .ZN(n7179)
         );
  AOI21_X1 U8888 ( .B1(n8778), .B2(n7239), .A(n7179), .ZN(n7180) );
  OAI211_X1 U8889 ( .C1(n7185), .C2(n7182), .A(n7181), .B(n7180), .ZN(P2_U3224) );
  INV_X1 U8890 ( .A(n7183), .ZN(n7189) );
  OAI222_X1 U8891 ( .A1(n9493), .A2(n7189), .B1(n8163), .B2(P1_U3086), .C1(
        n7184), .C2(n9490), .ZN(P1_U3335) );
  OAI22_X1 U8892 ( .A1(n7185), .A2(n8846), .B1(n7233), .B2(n8847), .ZN(n7186)
         );
  NOR2_X1 U8893 ( .A1(n7187), .A2(n7186), .ZN(n9893) );
  OR2_X1 U8894 ( .A1(n8827), .A2(n5226), .ZN(n7188) );
  OAI21_X1 U8895 ( .B1(n9893), .B2(n8857), .A(n7188), .ZN(P2_U3468) );
  OAI222_X1 U8896 ( .A1(P2_U3151), .A2(n4839), .B1(n8947), .B2(n7189), .C1(
        n10004), .C2(n8945), .ZN(P2_U3275) );
  AOI21_X1 U8897 ( .B1(n7192), .B2(n7191), .A(n7190), .ZN(n7200) );
  NAND2_X1 U8898 ( .A1(n9061), .A2(n9104), .ZN(n7194) );
  OAI211_X1 U8899 ( .C1(n7454), .C2(n9068), .A(n7194), .B(n7193), .ZN(n7197)
         );
  NOR2_X1 U8900 ( .A1(n7195), .A2(n9080), .ZN(n7196) );
  AOI211_X1 U8901 ( .C1(n7198), .C2(n9084), .A(n7197), .B(n7196), .ZN(n7199)
         );
  OAI21_X1 U8902 ( .B1(n7200), .B2(n4495), .A(n7199), .ZN(P1_U3221) );
  NAND2_X1 U8903 ( .A1(n7201), .A2(n7731), .ZN(n7202) );
  NAND2_X1 U8904 ( .A1(n7740), .A2(n7737), .ZN(n7654) );
  XNOR2_X1 U8905 ( .A(n7202), .B(n7654), .ZN(n7271) );
  INV_X1 U8906 ( .A(n7271), .ZN(n7208) );
  XOR2_X1 U8907 ( .A(n7258), .B(n7654), .Z(n7203) );
  OAI222_X1 U8908 ( .A1(n8840), .A2(n7215), .B1(n8838), .B2(n7408), .C1(n8679), 
        .C2(n7203), .ZN(n7269) );
  NAND2_X1 U8909 ( .A1(n7269), .A2(n8693), .ZN(n7207) );
  INV_X1 U8910 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7204) );
  OAI22_X1 U8911 ( .A1(n8693), .A2(n7204), .B1(n8310), .B2(n9869), .ZN(n7205)
         );
  AOI21_X1 U8912 ( .B1(n8778), .B2(n8309), .A(n7205), .ZN(n7206) );
  OAI211_X1 U8913 ( .C1(n7208), .C2(n8765), .A(n7207), .B(n7206), .ZN(P2_U3223) );
  INV_X1 U8914 ( .A(n7209), .ZN(n7210) );
  NAND2_X1 U8915 ( .A1(n7210), .A2(n7216), .ZN(n7211) );
  NAND2_X1 U8916 ( .A1(n7212), .A2(n7211), .ZN(n7228) );
  XNOR2_X1 U8917 ( .A(n6784), .B(n7213), .ZN(n7229) );
  XNOR2_X1 U8918 ( .A(n7229), .B(n7237), .ZN(n7227) );
  XNOR2_X1 U8919 ( .A(n7228), .B(n7227), .ZN(n7214) );
  NAND2_X1 U8920 ( .A1(n7214), .A2(n9958), .ZN(n7221) );
  OAI22_X1 U8921 ( .A1(n8440), .A2(n7216), .B1(n7215), .B2(n8427), .ZN(n7217)
         );
  AOI211_X1 U8922 ( .C1(n7219), .C2(n9950), .A(n7218), .B(n7217), .ZN(n7220)
         );
  OAI211_X1 U8923 ( .C1(n7222), .C2(n8428), .A(n7221), .B(n7220), .ZN(P2_U3161) );
  INV_X1 U8924 ( .A(n7223), .ZN(n7226) );
  INV_X1 U8925 ( .A(n6152), .ZN(n8102) );
  OAI222_X1 U8926 ( .A1(n9493), .A2(n7226), .B1(P1_U3086), .B2(n8102), .C1(
        n7224), .C2(n9490), .ZN(P1_U3334) );
  OAI222_X1 U8927 ( .A1(P2_U3151), .A2(n7681), .B1(n8947), .B2(n7226), .C1(
        n7225), .C2(n8945), .ZN(P2_U3274) );
  INV_X1 U8928 ( .A(n7229), .ZN(n7230) );
  NAND2_X1 U8929 ( .A1(n7230), .A2(n7237), .ZN(n7231) );
  XNOR2_X1 U8930 ( .A(n6784), .B(n7233), .ZN(n7404) );
  XNOR2_X1 U8931 ( .A(n7404), .B(n8466), .ZN(n7234) );
  AOI21_X1 U8932 ( .B1(n7235), .B2(n7234), .A(n8410), .ZN(n7236) );
  NAND2_X1 U8933 ( .A1(n7236), .A2(n7405), .ZN(n7241) );
  AND2_X1 U8934 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n9733) );
  OAI22_X1 U8935 ( .A1(n8440), .A2(n7237), .B1(n7409), .B2(n8427), .ZN(n7238)
         );
  AOI211_X1 U8936 ( .C1(n7239), .C2(n9950), .A(n9733), .B(n7238), .ZN(n7240)
         );
  OAI211_X1 U8937 ( .C1(n7242), .C2(n8428), .A(n7241), .B(n7240), .ZN(P2_U3171) );
  AOI21_X1 U8938 ( .B1(n7244), .B2(n7245), .A(n7243), .ZN(n7362) );
  INV_X1 U8939 ( .A(n7245), .ZN(n7952) );
  XNOR2_X1 U8940 ( .A(n7952), .B(n7246), .ZN(n7248) );
  OAI22_X1 U8941 ( .A1(n7391), .A2(n9347), .B1(n8955), .B2(n9349), .ZN(n7247)
         );
  AOI21_X1 U8942 ( .B1(n7248), .B2(n9352), .A(n7247), .ZN(n7361) );
  INV_X1 U8943 ( .A(n7361), .ZN(n7253) );
  OAI211_X1 U8944 ( .C1(n7462), .C2(n7392), .A(n9354), .B(n7435), .ZN(n7360)
         );
  AOI22_X1 U8945 ( .A1(n9358), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7395), .B2(
        n9356), .ZN(n7251) );
  NAND2_X1 U8946 ( .A1(n7249), .A2(n9359), .ZN(n7250) );
  OAI211_X1 U8947 ( .C1(n7360), .C2(n9363), .A(n7251), .B(n7250), .ZN(n7252)
         );
  AOI21_X1 U8948 ( .B1(n7253), .B2(n9365), .A(n7252), .ZN(n7254) );
  OAI21_X1 U8949 ( .B1(n7362), .B2(n9368), .A(n7254), .ZN(P1_U3281) );
  NAND2_X1 U8950 ( .A1(n7255), .A2(n7737), .ZN(n7256) );
  INV_X1 U8951 ( .A(n7261), .ZN(n7657) );
  XNOR2_X1 U8952 ( .A(n7256), .B(n7657), .ZN(n7346) );
  INV_X1 U8953 ( .A(n7346), .ZN(n7267) );
  OR2_X1 U8954 ( .A1(n7258), .A2(n7257), .ZN(n7350) );
  NAND2_X1 U8955 ( .A1(n7350), .A2(n7259), .ZN(n7260) );
  XNOR2_X1 U8956 ( .A(n7261), .B(n7260), .ZN(n7262) );
  OAI222_X1 U8957 ( .A1(n8838), .A2(n7263), .B1(n8840), .B2(n7409), .C1(n7262), 
        .C2(n8679), .ZN(n7344) );
  NAND2_X1 U8958 ( .A1(n7344), .A2(n8693), .ZN(n7266) );
  OAI22_X1 U8959 ( .A1(n8693), .A2(n5277), .B1(n9946), .B2(n9869), .ZN(n7264)
         );
  AOI21_X1 U8960 ( .B1(n8778), .B2(n9949), .A(n7264), .ZN(n7265) );
  OAI211_X1 U8961 ( .C1(n7267), .C2(n8765), .A(n7266), .B(n7265), .ZN(P2_U3222) );
  NOR2_X1 U8962 ( .A1(n7268), .A2(n8847), .ZN(n7270) );
  AOI211_X1 U8963 ( .C1(n7371), .C2(n7271), .A(n7270), .B(n7269), .ZN(n9895)
         );
  NAND2_X1 U8964 ( .A1(n8857), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7272) );
  OAI21_X1 U8965 ( .B1(n9895), .B2(n8857), .A(n7272), .ZN(P2_U3469) );
  INV_X1 U8966 ( .A(n7760), .ZN(n7273) );
  XNOR2_X1 U8967 ( .A(n7274), .B(n7273), .ZN(n7275) );
  NAND2_X1 U8968 ( .A1(n7275), .A2(n8842), .ZN(n7277) );
  AOI22_X1 U8969 ( .A1(n8769), .A2(n9951), .B1(n8464), .B2(n8771), .ZN(n7276)
         );
  NAND2_X1 U8970 ( .A1(n7277), .A2(n7276), .ZN(n7301) );
  AND2_X1 U8971 ( .A1(n7279), .A2(n7278), .ZN(n7280) );
  OR2_X1 U8972 ( .A1(n7281), .A2(n7280), .ZN(n7285) );
  NAND2_X1 U8973 ( .A1(n7283), .A2(n7282), .ZN(n7284) );
  MUX2_X1 U8974 ( .A(n7301), .B(P2_REG0_REG_13__SCAN_IN), .S(n9898), .Z(n7288)
         );
  XNOR2_X1 U8975 ( .A(n7286), .B(n7760), .ZN(n7306) );
  NOR2_X2 U8976 ( .A1(n9898), .A2(n8847), .ZN(n8933) );
  INV_X1 U8977 ( .A(n8933), .ZN(n8914) );
  OAI22_X1 U8978 ( .A1(n7306), .A2(n8937), .B1(n7289), .B2(n8914), .ZN(n7287)
         );
  OR2_X1 U8979 ( .A1(n7288), .A2(n7287), .ZN(P2_U3429) );
  MUX2_X1 U8980 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n7301), .S(n8827), .Z(n7291)
         );
  INV_X1 U8981 ( .A(n8829), .ZN(n8818) );
  OAI22_X1 U8982 ( .A1(n7306), .A2(n8832), .B1(n7289), .B2(n8818), .ZN(n7290)
         );
  OR2_X1 U8983 ( .A1(n7291), .A2(n7290), .ZN(P2_U3472) );
  XOR2_X1 U8984 ( .A(n7293), .B(n7292), .Z(n7300) );
  NAND2_X1 U8985 ( .A1(n9061), .A2(n9103), .ZN(n7295) );
  OAI211_X1 U8986 ( .C1(n9046), .C2(n9068), .A(n7295), .B(n7294), .ZN(n7297)
         );
  NOR2_X1 U8987 ( .A1(n9638), .A2(n9080), .ZN(n7296) );
  AOI211_X1 U8988 ( .C1(n7298), .C2(n9084), .A(n7297), .B(n7296), .ZN(n7299)
         );
  OAI21_X1 U8989 ( .B1(n7300), .B2(n4495), .A(n7299), .ZN(P1_U3231) );
  MUX2_X1 U8990 ( .A(n7301), .B(P2_REG2_REG_13__SCAN_IN), .S(n9876), .Z(n7302)
         );
  INV_X1 U8991 ( .A(n7302), .ZN(n7305) );
  NOR2_X1 U8992 ( .A1(n9876), .A2(n9866), .ZN(n8672) );
  INV_X1 U8993 ( .A(n8406), .ZN(n7303) );
  AOI22_X1 U8994 ( .A1(n8672), .A2(n8408), .B1(n8777), .B2(n7303), .ZN(n7304)
         );
  OAI211_X1 U8995 ( .C1(n7306), .C2(n8765), .A(n7305), .B(n7304), .ZN(P2_U3220) );
  INV_X1 U8996 ( .A(n7307), .ZN(n7311) );
  OAI222_X1 U8997 ( .A1(n7309), .A2(P2_U3151), .B1(n8947), .B2(n7311), .C1(
        n7308), .C2(n8945), .ZN(P2_U3273) );
  OAI222_X1 U8998 ( .A1(n9490), .A2(n7312), .B1(n9488), .B2(n7311), .C1(n7310), 
        .C2(P1_U3086), .ZN(P1_U3333) );
  INV_X1 U8999 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9908) );
  NOR2_X1 U9000 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7313) );
  AOI21_X1 U9001 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7313), .ZN(n9912) );
  NOR2_X1 U9002 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7314) );
  AOI21_X1 U9003 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7314), .ZN(n9915) );
  NOR2_X1 U9004 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n7315) );
  AOI21_X1 U9005 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n7315), .ZN(n9918) );
  NOR2_X1 U9006 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7316) );
  AOI21_X1 U9007 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7316), .ZN(n9921) );
  NOR2_X1 U9008 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7317) );
  AOI21_X1 U9009 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7317), .ZN(n9924) );
  NOR2_X1 U9010 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7318) );
  AOI21_X1 U9011 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7318), .ZN(n9927) );
  OR2_X1 U9012 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9929) );
  NOR2_X1 U9013 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9933) );
  NOR2_X1 U9014 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n7325) );
  XNOR2_X1 U9015 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n10137) );
  NAND2_X1 U9016 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7323) );
  XOR2_X1 U9017 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10135) );
  NAND2_X1 U9018 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7321) );
  XOR2_X1 U9019 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10133) );
  AOI21_X1 U9020 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9902) );
  NAND3_X1 U9021 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9904) );
  OAI21_X1 U9022 ( .B1(n9902), .B2(n7319), .A(n9904), .ZN(n10132) );
  NAND2_X1 U9023 ( .A1(n10133), .A2(n10132), .ZN(n7320) );
  NAND2_X1 U9024 ( .A1(n7321), .A2(n7320), .ZN(n10134) );
  NAND2_X1 U9025 ( .A1(n10135), .A2(n10134), .ZN(n7322) );
  NAND2_X1 U9026 ( .A1(n7323), .A2(n7322), .ZN(n10136) );
  NOR2_X1 U9027 ( .A1(n10137), .A2(n10136), .ZN(n7324) );
  NOR2_X1 U9028 ( .A1(n7325), .A2(n7324), .ZN(n7326) );
  NOR2_X1 U9029 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7326), .ZN(n10123) );
  AND2_X1 U9030 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7326), .ZN(n10124) );
  NOR2_X1 U9031 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10124), .ZN(n7327) );
  NOR2_X1 U9032 ( .A1(n10123), .A2(n7327), .ZN(n7328) );
  NAND2_X1 U9033 ( .A1(n7328), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7330) );
  XOR2_X1 U9034 ( .A(n7328), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10122) );
  NAND2_X1 U9035 ( .A1(n10122), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7329) );
  NAND2_X1 U9036 ( .A1(n7330), .A2(n7329), .ZN(n7331) );
  NAND2_X1 U9037 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7331), .ZN(n7333) );
  XOR2_X1 U9038 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7331), .Z(n10130) );
  NAND2_X1 U9039 ( .A1(n10130), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7332) );
  NAND2_X1 U9040 ( .A1(n7333), .A2(n7332), .ZN(n7334) );
  NAND2_X1 U9041 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7334), .ZN(n7336) );
  XOR2_X1 U9042 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7334), .Z(n10131) );
  NAND2_X1 U9043 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10131), .ZN(n7335) );
  NAND2_X1 U9044 ( .A1(n7336), .A2(n7335), .ZN(n7337) );
  INV_X1 U9045 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10129) );
  XNOR2_X1 U9046 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n7337), .ZN(n10128) );
  NAND2_X1 U9047 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9932) );
  AOI22_X1 U9048 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .B1(n9929), .B2(n9930), .ZN(n9926) );
  NAND2_X1 U9049 ( .A1(n9927), .A2(n9926), .ZN(n9925) );
  OAI21_X1 U9050 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9925), .ZN(n9923) );
  NAND2_X1 U9051 ( .A1(n9924), .A2(n9923), .ZN(n9922) );
  OAI21_X1 U9052 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9922), .ZN(n9920) );
  NAND2_X1 U9053 ( .A1(n9921), .A2(n9920), .ZN(n9919) );
  OAI21_X1 U9054 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9919), .ZN(n9917) );
  NAND2_X1 U9055 ( .A1(n9918), .A2(n9917), .ZN(n9916) );
  OAI21_X1 U9056 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9916), .ZN(n9914) );
  NAND2_X1 U9057 ( .A1(n9915), .A2(n9914), .ZN(n9913) );
  OAI21_X1 U9058 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9913), .ZN(n9911) );
  NAND2_X1 U9059 ( .A1(n9912), .A2(n9911), .ZN(n9910) );
  OAI21_X1 U9060 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9910), .ZN(n9907) );
  NAND2_X1 U9061 ( .A1(n9908), .A2(n9907), .ZN(n7339) );
  NOR2_X1 U9062 ( .A1(n9908), .A2(n9907), .ZN(n9906) );
  AOI21_X1 U9063 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7339), .A(n9906), .ZN(
        n7343) );
  NOR2_X1 U9064 ( .A1(n7341), .A2(n7340), .ZN(n7342) );
  XNOR2_X1 U9065 ( .A(n7343), .B(n7342), .ZN(ADD_1068_U4) );
  INV_X1 U9066 ( .A(n9949), .ZN(n7754) );
  NOR2_X1 U9067 ( .A1(n7754), .A2(n8847), .ZN(n7345) );
  AOI211_X1 U9068 ( .C1(n7346), .C2(n7371), .A(n7345), .B(n7344), .ZN(n9897)
         );
  NAND2_X1 U9069 ( .A1(n8857), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7347) );
  OAI21_X1 U9070 ( .B1(n9897), .B2(n8857), .A(n7347), .ZN(P2_U3470) );
  XOR2_X1 U9071 ( .A(n7348), .B(n7656), .Z(n7370) );
  INV_X1 U9072 ( .A(n7370), .ZN(n7359) );
  NAND2_X1 U9073 ( .A1(n7350), .A2(n7349), .ZN(n7351) );
  AND2_X1 U9074 ( .A1(n7352), .A2(n7351), .ZN(n7353) );
  XOR2_X1 U9075 ( .A(n7656), .B(n7353), .Z(n7354) );
  OAI222_X1 U9076 ( .A1(n8838), .A2(n8238), .B1(n8840), .B2(n7408), .C1(n7354), 
        .C2(n8679), .ZN(n7368) );
  NAND2_X1 U9077 ( .A1(n7368), .A2(n8693), .ZN(n7358) );
  OAI22_X1 U9078 ( .A1(n8693), .A2(n7355), .B1(n7418), .B2(n9869), .ZN(n7356)
         );
  AOI21_X1 U9079 ( .B1(n8778), .B2(n7420), .A(n7356), .ZN(n7357) );
  OAI211_X1 U9080 ( .C1(n7359), .C2(n8765), .A(n7358), .B(n7357), .ZN(P2_U3221) );
  INV_X1 U9081 ( .A(n9648), .ZN(n9433) );
  OAI211_X1 U9082 ( .C1(n7362), .C2(n9433), .A(n7361), .B(n7360), .ZN(n7366)
         );
  INV_X1 U9083 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9143) );
  OAI22_X1 U9084 ( .A1(n7392), .A2(n9384), .B1(n9659), .B2(n9143), .ZN(n7363)
         );
  AOI21_X1 U9085 ( .B1(n7366), .B2(n9659), .A(n7363), .ZN(n7364) );
  INV_X1 U9086 ( .A(n7364), .ZN(P1_U3534) );
  INV_X1 U9087 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10011) );
  OAI22_X1 U9088 ( .A1(n7392), .A2(n9445), .B1(n9480), .B2(n10011), .ZN(n7365)
         );
  AOI21_X1 U9089 ( .B1(n7366), .B2(n9480), .A(n7365), .ZN(n7367) );
  INV_X1 U9090 ( .A(n7367), .ZN(P1_U3489) );
  NOR2_X1 U9091 ( .A1(n7415), .A2(n8847), .ZN(n7369) );
  AOI211_X1 U9092 ( .C1(n7371), .C2(n7370), .A(n7369), .B(n7368), .ZN(n9900)
         );
  NAND2_X1 U9093 ( .A1(n8857), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7372) );
  OAI21_X1 U9094 ( .B1(n9900), .B2(n8857), .A(n7372), .ZN(P2_U3471) );
  NAND2_X1 U9095 ( .A1(n7768), .A2(n7772), .ZN(n7660) );
  XNOR2_X1 U9096 ( .A(n7373), .B(n7762), .ZN(n7387) );
  XNOR2_X1 U9097 ( .A(n7374), .B(n7762), .ZN(n7375) );
  AOI222_X1 U9098 ( .A1(n8842), .A2(n7375), .B1(n8465), .B2(n8769), .C1(n8770), 
        .C2(n8771), .ZN(n7381) );
  MUX2_X1 U9099 ( .A(n8513), .B(n7381), .S(n8827), .Z(n7377) );
  NAND2_X1 U9100 ( .A1(n8286), .A2(n8829), .ZN(n7376) );
  OAI211_X1 U9101 ( .C1(n7387), .C2(n8832), .A(n7377), .B(n7376), .ZN(P2_U3473) );
  INV_X1 U9102 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7378) );
  MUX2_X1 U9103 ( .A(n7378), .B(n7381), .S(n9901), .Z(n7380) );
  NAND2_X1 U9104 ( .A1(n8933), .A2(n8286), .ZN(n7379) );
  OAI211_X1 U9105 ( .C1(n7387), .C2(n8937), .A(n7380), .B(n7379), .ZN(P2_U3432) );
  INV_X1 U9106 ( .A(n7381), .ZN(n7384) );
  INV_X1 U9107 ( .A(n8286), .ZN(n7382) );
  OAI22_X1 U9108 ( .A1(n7382), .A2(n9866), .B1(n8287), .B2(n9869), .ZN(n7383)
         );
  OAI21_X1 U9109 ( .B1(n7384), .B2(n7383), .A(n8693), .ZN(n7386) );
  NAND2_X1 U9110 ( .A1(n9876), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7385) );
  OAI211_X1 U9111 ( .C1(n7387), .C2(n8765), .A(n7386), .B(n7385), .ZN(P2_U3219) );
  XOR2_X1 U9112 ( .A(n7389), .B(n7388), .Z(n7397) );
  INV_X1 U9113 ( .A(n8955), .ZN(n9098) );
  NAND2_X1 U9114 ( .A1(n9076), .A2(n9098), .ZN(n7390) );
  NAND2_X1 U9115 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9537) );
  OAI211_X1 U9116 ( .C1(n7391), .C2(n9078), .A(n7390), .B(n9537), .ZN(n7394)
         );
  NOR2_X1 U9117 ( .A1(n7392), .A2(n9080), .ZN(n7393) );
  AOI211_X1 U9118 ( .C1(n7395), .C2(n9084), .A(n7394), .B(n7393), .ZN(n7396)
         );
  OAI21_X1 U9119 ( .B1(n7397), .B2(n4495), .A(n7396), .ZN(P1_U3224) );
  INV_X1 U9120 ( .A(n7398), .ZN(n7403) );
  AOI21_X1 U9121 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9486), .A(n7399), .ZN(
        n7400) );
  OAI21_X1 U9122 ( .B1(n7403), .B2(n9488), .A(n7400), .ZN(P1_U3332) );
  AOI21_X1 U9123 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8942), .A(n7401), .ZN(
        n7402) );
  OAI21_X1 U9124 ( .B1(n7403), .B2(n8947), .A(n7402), .ZN(P2_U3272) );
  XNOR2_X1 U9125 ( .A(n6784), .B(n8309), .ZN(n7407) );
  XNOR2_X1 U9126 ( .A(n6784), .B(n9949), .ZN(n9939) );
  AOI22_X1 U9127 ( .A1(n7409), .A2(n7407), .B1(n9939), .B2(n7408), .ZN(n7406)
         );
  NAND2_X1 U9128 ( .A1(n8306), .A2(n7406), .ZN(n7414) );
  OAI21_X1 U9129 ( .B1(n7407), .B2(n7409), .A(n7408), .ZN(n7412) );
  INV_X1 U9130 ( .A(n9939), .ZN(n7411) );
  INV_X1 U9131 ( .A(n7407), .ZN(n9937) );
  NOR2_X1 U9132 ( .A1(n7409), .A2(n7408), .ZN(n7410) );
  AOI22_X1 U9133 ( .A1(n7412), .A2(n7411), .B1(n9937), .B2(n7410), .ZN(n7413)
         );
  XNOR2_X1 U9134 ( .A(n6784), .B(n7415), .ZN(n8234) );
  XNOR2_X1 U9135 ( .A(n8234), .B(n9951), .ZN(n7416) );
  XNOR2_X1 U9136 ( .A(n8235), .B(n7416), .ZN(n7426) );
  NOR2_X1 U9137 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7417), .ZN(n9787) );
  AOI21_X1 U9138 ( .B1(n9945), .B2(n4441), .A(n9787), .ZN(n7424) );
  INV_X1 U9139 ( .A(n7418), .ZN(n7419) );
  NAND2_X1 U9140 ( .A1(n9948), .A2(n7419), .ZN(n7423) );
  NAND2_X1 U9141 ( .A1(n9950), .A2(n7420), .ZN(n7422) );
  NAND2_X1 U9142 ( .A1(n9952), .A2(n8465), .ZN(n7421) );
  NAND4_X1 U9143 ( .A1(n7424), .A2(n7423), .A3(n7422), .A4(n7421), .ZN(n7425)
         );
  AOI21_X1 U9144 ( .B1(n7426), .B2(n9958), .A(n7425), .ZN(n7427) );
  INV_X1 U9145 ( .A(n7427), .ZN(P2_U3164) );
  AOI21_X1 U9146 ( .B1(n7429), .B2(n7955), .A(n7428), .ZN(n7450) );
  OAI21_X1 U9147 ( .B1(n7955), .B2(n7431), .A(n7430), .ZN(n7434) );
  NAND2_X1 U9148 ( .A1(n9099), .A2(n9335), .ZN(n7432) );
  OAI21_X1 U9149 ( .B1(n9079), .B2(n9349), .A(n7432), .ZN(n7433) );
  AOI21_X1 U9150 ( .B1(n7434), .B2(n9352), .A(n7433), .ZN(n7443) );
  INV_X1 U9151 ( .A(n7443), .ZN(n7440) );
  INV_X1 U9152 ( .A(n7491), .ZN(n7436) );
  OAI211_X1 U9153 ( .C1(n7501), .C2(n4576), .A(n7436), .B(n9354), .ZN(n7442)
         );
  AOI22_X1 U9154 ( .A1(n9358), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7504), .B2(
        n9356), .ZN(n7438) );
  NAND2_X1 U9155 ( .A1(n7446), .A2(n9359), .ZN(n7437) );
  OAI211_X1 U9156 ( .C1(n7442), .C2(n9363), .A(n7438), .B(n7437), .ZN(n7439)
         );
  AOI21_X1 U9157 ( .B1(n7440), .B2(n9365), .A(n7439), .ZN(n7441) );
  OAI21_X1 U9158 ( .B1(n7450), .B2(n9368), .A(n7441), .ZN(P1_U3280) );
  AOI22_X1 U9159 ( .A1(n7446), .A2(n9471), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n6284), .ZN(n7445) );
  NAND2_X1 U9160 ( .A1(n7443), .A2(n7442), .ZN(n7447) );
  NAND2_X1 U9161 ( .A1(n7447), .A2(n9480), .ZN(n7444) );
  OAI211_X1 U9162 ( .C1(n7450), .C2(n9478), .A(n7445), .B(n7444), .ZN(P1_U3492) );
  AOI22_X1 U9163 ( .A1(n7446), .A2(n9414), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n9656), .ZN(n7449) );
  NAND2_X1 U9164 ( .A1(n7447), .A2(n9659), .ZN(n7448) );
  OAI211_X1 U9165 ( .C1(n7450), .C2(n9427), .A(n7449), .B(n7448), .ZN(P1_U3535) );
  XNOR2_X1 U9166 ( .A(n9039), .B(n9040), .ZN(n7452) );
  NOR2_X1 U9167 ( .A1(n7452), .A2(n7451), .ZN(n9038) );
  AOI21_X1 U9168 ( .B1(n7452), .B2(n7451), .A(n9038), .ZN(n7459) );
  NAND2_X1 U9169 ( .A1(n9076), .A2(n9100), .ZN(n7453) );
  NAND2_X1 U9170 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9503) );
  OAI211_X1 U9171 ( .C1(n7454), .C2(n9078), .A(n7453), .B(n9503), .ZN(n7456)
         );
  NOR2_X1 U9172 ( .A1(n9646), .A2(n9080), .ZN(n7455) );
  AOI211_X1 U9173 ( .C1(n7457), .C2(n9084), .A(n7456), .B(n7455), .ZN(n7458)
         );
  OAI21_X1 U9174 ( .B1(n7459), .B2(n4495), .A(n7458), .ZN(P1_U3217) );
  OAI21_X1 U9175 ( .B1(n7460), .B2(n9047), .A(n9354), .ZN(n7461) );
  OR2_X1 U9176 ( .A1(n7462), .A2(n7461), .ZN(n7478) );
  AOI21_X1 U9177 ( .B1(n7463), .B2(n7954), .A(n4403), .ZN(n7481) );
  NAND2_X1 U9178 ( .A1(n7464), .A2(n8010), .ZN(n7465) );
  XNOR2_X1 U9179 ( .A(n7465), .B(n7954), .ZN(n7470) );
  OAI22_X1 U9180 ( .A1(n7466), .A2(n9349), .B1(n9046), .B2(n9347), .ZN(n7469)
         );
  NOR2_X1 U9181 ( .A1(n7481), .A2(n7467), .ZN(n7468) );
  AOI211_X1 U9182 ( .C1(n7470), .C2(n9352), .A(n7469), .B(n7468), .ZN(n7479)
         );
  OAI21_X1 U9183 ( .B1(n7481), .B2(n7471), .A(n7479), .ZN(n7472) );
  NAND2_X1 U9184 ( .A1(n7472), .A2(n9365), .ZN(n7477) );
  INV_X1 U9185 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7474) );
  INV_X1 U9186 ( .A(n9050), .ZN(n7473) );
  OAI22_X1 U9187 ( .A1(n9365), .A2(n7474), .B1(n7473), .B2(n9211), .ZN(n7475)
         );
  AOI21_X1 U9188 ( .B1(n7484), .B2(n9359), .A(n7475), .ZN(n7476) );
  OAI211_X1 U9189 ( .C1(n7478), .C2(n9363), .A(n7477), .B(n7476), .ZN(P1_U3282) );
  OAI211_X1 U9190 ( .C1(n7481), .C2(n7480), .A(n7479), .B(n7478), .ZN(n7482)
         );
  INV_X1 U9191 ( .A(n7482), .ZN(n7486) );
  AOI22_X1 U9192 ( .A1(n7484), .A2(n9414), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n9656), .ZN(n7483) );
  OAI21_X1 U9193 ( .B1(n7486), .B2(n9656), .A(n7483), .ZN(P1_U3533) );
  AOI22_X1 U9194 ( .A1(n7484), .A2(n9471), .B1(P1_REG0_REG_11__SCAN_IN), .B2(
        n6284), .ZN(n7485) );
  OAI21_X1 U9195 ( .B1(n7486), .B2(n6284), .A(n7485), .ZN(P1_U3486) );
  XNOR2_X1 U9196 ( .A(n7487), .B(n7488), .ZN(n7520) );
  INV_X1 U9197 ( .A(n7488), .ZN(n8027) );
  XNOR2_X1 U9198 ( .A(n7489), .B(n8027), .ZN(n7490) );
  AOI222_X1 U9199 ( .A1(n9098), .A2(n9335), .B1(n9096), .B2(n9337), .C1(n9352), 
        .C2(n7490), .ZN(n7514) );
  INV_X1 U9200 ( .A(n7514), .ZN(n7496) );
  OAI211_X1 U9201 ( .C1(n8960), .C2(n7491), .A(n9354), .B(n7543), .ZN(n7513)
         );
  AOI22_X1 U9202 ( .A1(n9358), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8957), .B2(
        n9356), .ZN(n7494) );
  NAND2_X1 U9203 ( .A1(n7492), .A2(n9359), .ZN(n7493) );
  OAI211_X1 U9204 ( .C1(n7513), .C2(n9363), .A(n7494), .B(n7493), .ZN(n7495)
         );
  AOI21_X1 U9205 ( .B1(n7496), .B2(n9365), .A(n7495), .ZN(n7497) );
  OAI21_X1 U9206 ( .B1(n7520), .B2(n9368), .A(n7497), .ZN(P1_U3279) );
  XOR2_X1 U9207 ( .A(n7499), .B(n7498), .Z(n7506) );
  NAND2_X1 U9208 ( .A1(n9061), .A2(n9099), .ZN(n7500) );
  NAND2_X1 U9209 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9550) );
  OAI211_X1 U9210 ( .C1(n9079), .C2(n9068), .A(n7500), .B(n9550), .ZN(n7503)
         );
  NOR2_X1 U9211 ( .A1(n7501), .A2(n9080), .ZN(n7502) );
  AOI211_X1 U9212 ( .C1(n7504), .C2(n9084), .A(n7503), .B(n7502), .ZN(n7505)
         );
  OAI21_X1 U9213 ( .B1(n7506), .B2(n4495), .A(n7505), .ZN(P1_U3234) );
  XNOR2_X1 U9214 ( .A(n8243), .B(n7507), .ZN(n7661) );
  INV_X1 U9215 ( .A(n7661), .ZN(n7766) );
  XNOR2_X1 U9216 ( .A(n7508), .B(n7766), .ZN(n7529) );
  XNOR2_X1 U9217 ( .A(n7509), .B(n7661), .ZN(n7510) );
  AOI222_X1 U9218 ( .A1(n8842), .A2(n7510), .B1(n8757), .B2(n8771), .C1(n8464), 
        .C2(n8769), .ZN(n7524) );
  MUX2_X1 U9219 ( .A(n9969), .B(n7524), .S(n8827), .Z(n7512) );
  NAND2_X1 U9220 ( .A1(n8243), .A2(n8829), .ZN(n7511) );
  OAI211_X1 U9221 ( .C1(n8832), .C2(n7529), .A(n7512), .B(n7511), .ZN(P2_U3474) );
  OAI211_X1 U9222 ( .C1(n8960), .C2(n9645), .A(n7514), .B(n7513), .ZN(n7517)
         );
  NAND2_X1 U9223 ( .A1(n7517), .A2(n9480), .ZN(n7516) );
  NAND2_X1 U9224 ( .A1(n6284), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7515) );
  OAI211_X1 U9225 ( .C1(n7520), .C2(n9478), .A(n7516), .B(n7515), .ZN(P1_U3495) );
  NAND2_X1 U9226 ( .A1(n7517), .A2(n9659), .ZN(n7519) );
  NAND2_X1 U9227 ( .A1(n9656), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7518) );
  OAI211_X1 U9228 ( .C1(n7520), .C2(n9427), .A(n7519), .B(n7518), .ZN(P1_U3536) );
  INV_X1 U9229 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7521) );
  MUX2_X1 U9230 ( .A(n7521), .B(n7524), .S(n9901), .Z(n7523) );
  NAND2_X1 U9231 ( .A1(n8243), .A2(n8933), .ZN(n7522) );
  OAI211_X1 U9232 ( .C1(n7529), .C2(n8937), .A(n7523), .B(n7522), .ZN(P2_U3435) );
  INV_X1 U9233 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7525) );
  MUX2_X1 U9234 ( .A(n7525), .B(n7524), .S(n8693), .Z(n7528) );
  INV_X1 U9235 ( .A(n7526), .ZN(n8452) );
  AOI22_X1 U9236 ( .A1(n8243), .A2(n8778), .B1(n8777), .B2(n8452), .ZN(n7527)
         );
  OAI211_X1 U9237 ( .C1(n7529), .C2(n8765), .A(n7528), .B(n7527), .ZN(P2_U3218) );
  INV_X1 U9238 ( .A(n7530), .ZN(n7534) );
  OAI222_X1 U9239 ( .A1(n9493), .A2(n7534), .B1(n7532), .B2(P1_U3086), .C1(
        n7531), .C2(n9490), .ZN(P1_U3330) );
  OAI222_X1 U9240 ( .A1(n7535), .A2(P2_U3151), .B1(n8947), .B2(n7534), .C1(
        n7533), .C2(n8945), .ZN(P2_U3270) );
  INV_X1 U9241 ( .A(n7536), .ZN(n7540) );
  OAI222_X1 U9242 ( .A1(n9493), .A2(n7540), .B1(n7538), .B2(P1_U3086), .C1(
        n7537), .C2(n9490), .ZN(P1_U3329) );
  OAI222_X1 U9243 ( .A1(n7541), .A2(P2_U3151), .B1(n8947), .B2(n7540), .C1(
        n7539), .C2(n8945), .ZN(P2_U3269) );
  XNOR2_X1 U9244 ( .A(n7542), .B(n7957), .ZN(n7562) );
  INV_X1 U9245 ( .A(n7543), .ZN(n7544) );
  OAI211_X1 U9246 ( .C1(n9081), .C2(n7544), .A(n9354), .B(n7570), .ZN(n7554)
         );
  INV_X1 U9247 ( .A(n7545), .ZN(n7548) );
  INV_X1 U9248 ( .A(n7957), .ZN(n7547) );
  OAI21_X1 U9249 ( .B1(n7548), .B2(n7547), .A(n7546), .ZN(n7549) );
  AOI222_X1 U9250 ( .A1(n9352), .A2(n7549), .B1(n9095), .B2(n9337), .C1(n9097), 
        .C2(n9335), .ZN(n7555) );
  OAI21_X1 U9251 ( .B1(n4331), .B2(n7554), .A(n7555), .ZN(n7552) );
  AOI22_X1 U9252 ( .A1(n9358), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9085), .B2(
        n9356), .ZN(n7550) );
  OAI21_X1 U9253 ( .B1(n9081), .B2(n9330), .A(n7550), .ZN(n7551) );
  AOI21_X1 U9254 ( .B1(n7552), .B2(n9365), .A(n7551), .ZN(n7553) );
  OAI21_X1 U9255 ( .B1(n7562), .B2(n9368), .A(n7553), .ZN(P1_U3278) );
  AOI22_X1 U9256 ( .A1(n7558), .A2(n9471), .B1(P1_REG0_REG_15__SCAN_IN), .B2(
        n6284), .ZN(n7557) );
  NAND2_X1 U9257 ( .A1(n7555), .A2(n7554), .ZN(n7559) );
  NAND2_X1 U9258 ( .A1(n7559), .A2(n9480), .ZN(n7556) );
  OAI211_X1 U9259 ( .C1(n7562), .C2(n9478), .A(n7557), .B(n7556), .ZN(P1_U3498) );
  AOI22_X1 U9260 ( .A1(n7558), .A2(n9414), .B1(P1_REG1_REG_15__SCAN_IN), .B2(
        n9656), .ZN(n7561) );
  NAND2_X1 U9261 ( .A1(n7559), .A2(n9659), .ZN(n7560) );
  OAI211_X1 U9262 ( .C1(n7562), .C2(n9427), .A(n7561), .B(n7560), .ZN(P1_U3537) );
  INV_X1 U9263 ( .A(n7563), .ZN(n7583) );
  OAI222_X1 U9264 ( .A1(P2_U3151), .A2(n8588), .B1(n8947), .B2(n7583), .C1(
        n10040), .C2(n8945), .ZN(P2_U3268) );
  INV_X1 U9265 ( .A(n7565), .ZN(n7581) );
  NAND2_X1 U9266 ( .A1(n8942), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7566) );
  OAI211_X1 U9267 ( .C1(n7581), .C2(n8947), .A(n7567), .B(n7566), .ZN(P2_U3267) );
  XNOR2_X1 U9268 ( .A(n7568), .B(n4727), .ZN(n9434) );
  INV_X1 U9269 ( .A(n7569), .ZN(n9355) );
  AOI211_X1 U9270 ( .C1(n9429), .C2(n7570), .A(n9326), .B(n9355), .ZN(n9428)
         );
  INV_X1 U9271 ( .A(n9004), .ZN(n7571) );
  AOI22_X1 U9272 ( .A1(n9358), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7571), .B2(
        n9356), .ZN(n7572) );
  OAI21_X1 U9273 ( .B1(n4587), .B2(n9330), .A(n7572), .ZN(n7578) );
  OAI21_X1 U9274 ( .B1(n7575), .B2(n7574), .A(n7573), .ZN(n7576) );
  AOI222_X1 U9275 ( .A1(n9352), .A2(n7576), .B1(n9336), .B2(n9337), .C1(n9096), 
        .C2(n9335), .ZN(n9432) );
  NOR2_X1 U9276 ( .A1(n9432), .A2(n9358), .ZN(n7577) );
  AOI211_X1 U9277 ( .C1(n9428), .C2(n9342), .A(n7578), .B(n7577), .ZN(n7579)
         );
  OAI21_X1 U9278 ( .B1(n9434), .B2(n9368), .A(n7579), .ZN(P1_U3277) );
  OAI222_X1 U9279 ( .A1(n9493), .A2(n7581), .B1(P1_U3086), .B2(n4324), .C1(
        n7580), .C2(n9490), .ZN(P1_U3327) );
  AOI21_X1 U9280 ( .B1(n7584), .B2(n9342), .A(n9359), .ZN(n7593) );
  NAND2_X1 U9281 ( .A1(n7586), .A2(n7585), .ZN(n7588) );
  OAI21_X1 U9282 ( .B1(n7942), .B2(n7588), .A(n7587), .ZN(n7589) );
  AOI22_X1 U9283 ( .A1(n7589), .A2(n9365), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9356), .ZN(n7591) );
  NAND2_X1 U9284 ( .A1(n9358), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7590) );
  OAI211_X1 U9285 ( .C1(n7593), .C2(n7592), .A(n7591), .B(n7590), .ZN(P1_U3293) );
  INV_X1 U9286 ( .A(n7594), .ZN(n7601) );
  AOI22_X1 U9287 ( .A1(n9358), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n7595), .B2(
        n9356), .ZN(n7598) );
  NAND2_X1 U9288 ( .A1(n7596), .A2(n9359), .ZN(n7597) );
  OAI211_X1 U9289 ( .C1(n7599), .C2(n9363), .A(n7598), .B(n7597), .ZN(n7600)
         );
  AOI21_X1 U9290 ( .B1(n7601), .B2(n9365), .A(n7600), .ZN(n7602) );
  OAI21_X1 U9291 ( .B1(n7603), .B2(n9368), .A(n7602), .ZN(P1_U3266) );
  INV_X1 U9292 ( .A(n7846), .ZN(n7604) );
  INV_X1 U9293 ( .A(SI_29_), .ZN(n7609) );
  INV_X1 U9294 ( .A(n7633), .ZN(n7616) );
  INV_X1 U9295 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9995) );
  INV_X1 U9296 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8221) );
  MUX2_X1 U9297 ( .A(n9995), .B(n8221), .S(n4616), .Z(n7612) );
  INV_X1 U9298 ( .A(SI_30_), .ZN(n7611) );
  NAND2_X1 U9299 ( .A1(n7612), .A2(n7611), .ZN(n7617) );
  INV_X1 U9300 ( .A(n7612), .ZN(n7613) );
  NAND2_X1 U9301 ( .A1(n7613), .A2(SI_30_), .ZN(n7614) );
  NAND2_X1 U9302 ( .A1(n7617), .A2(n7614), .ZN(n7632) );
  INV_X1 U9303 ( .A(n7632), .ZN(n7615) );
  NAND2_X1 U9304 ( .A1(n7631), .A2(n7617), .ZN(n7620) );
  INV_X1 U9305 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7895) );
  MUX2_X1 U9306 ( .A(n6332), .B(n7895), .S(n4325), .Z(n7618) );
  XNOR2_X1 U9307 ( .A(n7618), .B(SI_31_), .ZN(n7619) );
  NOR2_X1 U9308 ( .A1(n7636), .A2(n6332), .ZN(n7621) );
  INV_X1 U9309 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7627) );
  NAND2_X1 U9310 ( .A1(n7622), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7625) );
  INV_X1 U9311 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7623) );
  OR2_X1 U9312 ( .A1(n5135), .A2(n7623), .ZN(n7624) );
  OAI211_X1 U9313 ( .C1(n7627), .C2(n7626), .A(n7625), .B(n7624), .ZN(n7628)
         );
  INV_X1 U9314 ( .A(n7628), .ZN(n7629) );
  NAND2_X1 U9315 ( .A1(n7630), .A2(n7629), .ZN(n8607) );
  NAND2_X1 U9316 ( .A1(n7633), .A2(n7632), .ZN(n7634) );
  NAND2_X1 U9317 ( .A1(n8220), .A2(n7635), .ZN(n7638) );
  OR2_X1 U9318 ( .A1(n7636), .A2(n9995), .ZN(n7637) );
  NAND2_X1 U9319 ( .A1(n8861), .A2(n7838), .ZN(n7666) );
  AND2_X1 U9320 ( .A1(n7666), .A2(n7835), .ZN(n7844) );
  INV_X1 U9321 ( .A(n7643), .ZN(n7668) );
  INV_X1 U9322 ( .A(n7644), .ZN(n7828) );
  INV_X1 U9323 ( .A(n7824), .ZN(n7645) );
  INV_X1 U9324 ( .A(n5528), .ZN(n7646) );
  NAND4_X1 U9325 ( .A1(n7646), .A2(n8833), .A3(n7697), .A4(n7681), .ZN(n7648)
         );
  NOR3_X1 U9326 ( .A1(n7648), .A2(n7647), .A3(n8229), .ZN(n7651) );
  NAND4_X1 U9327 ( .A1(n7651), .A2(n7720), .A3(n7650), .A4(n7649), .ZN(n7655)
         );
  NOR4_X1 U9328 ( .A1(n7655), .A2(n7654), .A3(n7653), .A4(n7652), .ZN(n7658)
         );
  NAND4_X1 U9329 ( .A1(n7658), .A2(n7760), .A3(n7657), .A4(n7656), .ZN(n7659)
         );
  NOR4_X1 U9330 ( .A1(n8767), .A2(n7661), .A3(n7660), .A4(n7659), .ZN(n7662)
         );
  NAND4_X1 U9331 ( .A1(n8727), .A2(n8746), .A3(n8755), .A4(n7662), .ZN(n7663)
         );
  NOR4_X1 U9332 ( .A1(n8689), .A2(n8709), .A3(n8716), .A4(n7663), .ZN(n7664)
         );
  NAND4_X1 U9333 ( .A1(n8653), .A2(n8666), .A3(n8676), .A4(n7664), .ZN(n7665)
         );
  NOR4_X1 U9334 ( .A1(n4356), .A2(n8632), .A3(n8644), .A4(n7665), .ZN(n7667)
         );
  OR2_X1 U9335 ( .A1(n8861), .A2(n7838), .ZN(n7837) );
  NAND4_X1 U9336 ( .A1(n7668), .A2(n7667), .A3(n7666), .A4(n7837), .ZN(n7669)
         );
  OAI22_X1 U9337 ( .A1(n7670), .A2(n7681), .B1(n7858), .B2(n7669), .ZN(n7675)
         );
  INV_X1 U9338 ( .A(n8607), .ZN(n7671) );
  NAND2_X1 U9339 ( .A1(n7672), .A2(n7671), .ZN(n7842) );
  INV_X1 U9340 ( .A(n7837), .ZN(n7673) );
  NAND3_X1 U9341 ( .A1(n7675), .A2(n7842), .A3(n7674), .ZN(n7676) );
  XNOR2_X1 U9342 ( .A(n7676), .B(n8592), .ZN(n7677) );
  MUX2_X1 U9343 ( .A(n7835), .B(n7846), .S(n7847), .Z(n7834) );
  INV_X1 U9344 ( .A(n8644), .ZN(n7821) );
  NAND4_X1 U9345 ( .A1(n7815), .A2(n8680), .A3(n7847), .A4(n8889), .ZN(n7679)
         );
  OR3_X1 U9346 ( .A1(n8883), .A2(n8441), .A3(n7847), .ZN(n7678) );
  OAI211_X1 U9347 ( .C1(n7826), .C2(n7816), .A(n7679), .B(n7678), .ZN(n7680)
         );
  INV_X1 U9348 ( .A(n7680), .ZN(n7820) );
  INV_X1 U9349 ( .A(n8889), .ZN(n8386) );
  NAND4_X1 U9350 ( .A1(n8653), .A2(n7826), .A3(n8386), .A4(n8462), .ZN(n7819)
         );
  NAND2_X1 U9351 ( .A1(n7682), .A2(n7681), .ZN(n7684) );
  INV_X1 U9352 ( .A(n7685), .ZN(n7687) );
  OAI21_X1 U9353 ( .B1(n5528), .B2(n7687), .A(n7686), .ZN(n7688) );
  MUX2_X1 U9354 ( .A(n7689), .B(n7688), .S(n7826), .Z(n7696) );
  NAND2_X1 U9355 ( .A1(n7709), .A2(n7690), .ZN(n7693) );
  NAND2_X1 U9356 ( .A1(n7698), .A2(n7691), .ZN(n7692) );
  MUX2_X1 U9357 ( .A(n7693), .B(n7692), .S(n7826), .Z(n7694) );
  INV_X1 U9358 ( .A(n7694), .ZN(n7695) );
  INV_X1 U9359 ( .A(n7698), .ZN(n7703) );
  NAND2_X1 U9360 ( .A1(n7700), .A2(n7699), .ZN(n7701) );
  AND2_X1 U9361 ( .A1(n7706), .A2(n7701), .ZN(n7716) );
  OAI211_X1 U9362 ( .C1(n7713), .C2(n7703), .A(n7716), .B(n7702), .ZN(n7708)
         );
  NAND2_X1 U9363 ( .A1(n8470), .A2(n7704), .ZN(n7711) );
  INV_X1 U9364 ( .A(n7711), .ZN(n7705) );
  NAND2_X1 U9365 ( .A1(n7706), .A2(n7705), .ZN(n7707) );
  NAND3_X1 U9366 ( .A1(n7708), .A2(n7714), .A3(n7707), .ZN(n7719) );
  INV_X1 U9367 ( .A(n7709), .ZN(n7712) );
  OAI211_X1 U9368 ( .C1(n7713), .C2(n7712), .A(n7711), .B(n7710), .ZN(n7717)
         );
  INV_X1 U9369 ( .A(n7714), .ZN(n7715) );
  AOI21_X1 U9370 ( .B1(n7717), .B2(n7716), .A(n7715), .ZN(n7718) );
  NAND2_X1 U9371 ( .A1(n7721), .A2(n7720), .ZN(n7726) );
  AND2_X1 U9372 ( .A1(n7727), .A2(n7722), .ZN(n7723) );
  MUX2_X1 U9373 ( .A(n7724), .B(n7723), .S(n7826), .Z(n7725) );
  NAND2_X1 U9374 ( .A1(n7726), .A2(n7725), .ZN(n7735) );
  NAND2_X1 U9375 ( .A1(n7727), .A2(n7736), .ZN(n7730) );
  INV_X1 U9376 ( .A(n7728), .ZN(n7729) );
  MUX2_X1 U9377 ( .A(n7730), .B(n7729), .S(n7826), .Z(n7733) );
  INV_X1 U9378 ( .A(n7731), .ZN(n7732) );
  NOR2_X1 U9379 ( .A1(n7733), .A2(n7732), .ZN(n7734) );
  NAND2_X1 U9380 ( .A1(n7735), .A2(n7734), .ZN(n7749) );
  AND2_X1 U9381 ( .A1(n7737), .A2(n7736), .ZN(n7738) );
  MUX2_X1 U9382 ( .A(n7739), .B(n7738), .S(n7826), .Z(n7748) );
  OR2_X1 U9383 ( .A1(n7740), .A2(n7847), .ZN(n7741) );
  NAND4_X1 U9384 ( .A1(n7758), .A2(n7742), .A3(n7755), .A4(n7741), .ZN(n7745)
         );
  NOR2_X1 U9385 ( .A1(n7743), .A2(n7826), .ZN(n7744) );
  NOR2_X1 U9386 ( .A1(n7745), .A2(n7744), .ZN(n7746) );
  NAND2_X1 U9387 ( .A1(n7760), .A2(n7746), .ZN(n7747) );
  AOI21_X1 U9388 ( .B1(n7749), .B2(n7748), .A(n7747), .ZN(n7765) );
  MUX2_X1 U9389 ( .A(n7751), .B(n7750), .S(n7826), .Z(n7763) );
  AOI21_X1 U9390 ( .B1(n7755), .B2(n7752), .A(n7847), .ZN(n7753) );
  NAND2_X1 U9391 ( .A1(n7753), .A2(n7758), .ZN(n7757) );
  NAND4_X1 U9392 ( .A1(n7755), .A2(n7754), .A3(n7847), .A4(n4441), .ZN(n7756)
         );
  OAI211_X1 U9393 ( .C1(n7826), .C2(n7758), .A(n7757), .B(n7756), .ZN(n7759)
         );
  NAND2_X1 U9394 ( .A1(n7760), .A2(n7759), .ZN(n7761) );
  NAND3_X1 U9395 ( .A1(n7763), .A2(n7762), .A3(n7761), .ZN(n7764) );
  OAI211_X1 U9396 ( .C1(n7847), .C2(n7768), .A(n7767), .B(n7766), .ZN(n7774)
         );
  NAND3_X1 U9397 ( .A1(n7774), .A2(n7777), .A3(n7769), .ZN(n7771) );
  MUX2_X1 U9398 ( .A(n7771), .B(n7770), .S(n7847), .Z(n7776) );
  INV_X1 U9399 ( .A(n7772), .ZN(n7773) );
  OAI21_X1 U9400 ( .B1(n7774), .B2(n7773), .A(n7779), .ZN(n7775) );
  OAI211_X1 U9401 ( .C1(n7780), .C2(n5538), .A(n8724), .B(n7778), .ZN(n7782)
         );
  NOR2_X1 U9402 ( .A1(n7780), .A2(n4778), .ZN(n7781) );
  MUX2_X1 U9403 ( .A(n7782), .B(n7781), .S(n7826), .Z(n7789) );
  NAND3_X1 U9404 ( .A1(n7789), .A2(n7790), .A3(n7786), .ZN(n7784) );
  NAND3_X1 U9405 ( .A1(n7784), .A2(n7794), .A3(n7783), .ZN(n7793) );
  NAND2_X1 U9406 ( .A1(n7786), .A2(n7785), .ZN(n7788) );
  NAND2_X1 U9407 ( .A1(n7791), .A2(n7790), .ZN(n7792) );
  INV_X1 U9408 ( .A(n8707), .ZN(n7798) );
  AND2_X1 U9409 ( .A1(n7800), .A2(n7794), .ZN(n7796) );
  MUX2_X1 U9410 ( .A(n7796), .B(n7795), .S(n7847), .Z(n7797) );
  INV_X1 U9411 ( .A(n8689), .ZN(n8688) );
  MUX2_X1 U9412 ( .A(n7801), .B(n7800), .S(n7847), .Z(n7802) );
  NAND3_X1 U9413 ( .A1(n7803), .A2(n8688), .A3(n7802), .ZN(n7810) );
  NAND2_X1 U9414 ( .A1(n8663), .A2(n7804), .ZN(n7807) );
  NAND2_X1 U9415 ( .A1(n7811), .A2(n7805), .ZN(n7806) );
  MUX2_X1 U9416 ( .A(n7807), .B(n7806), .S(n7826), .Z(n7808) );
  INV_X1 U9417 ( .A(n7808), .ZN(n7809) );
  NAND2_X1 U9418 ( .A1(n7810), .A2(n7809), .ZN(n7818) );
  MUX2_X1 U9419 ( .A(n7811), .B(n8663), .S(n7826), .Z(n7814) );
  AND3_X1 U9420 ( .A1(n7814), .A2(n7813), .A3(n7812), .ZN(n7817) );
  INV_X1 U9421 ( .A(n7822), .ZN(n7823) );
  MUX2_X1 U9422 ( .A(n7824), .B(n7823), .S(n7826), .Z(n7825) );
  MUX2_X1 U9423 ( .A(n7828), .B(n7827), .S(n7826), .Z(n7829) );
  INV_X1 U9424 ( .A(n7829), .ZN(n7830) );
  NAND2_X1 U9425 ( .A1(n7831), .A2(n7830), .ZN(n7845) );
  MUX2_X1 U9426 ( .A(n8461), .B(n8867), .S(n7847), .Z(n7832) );
  OR2_X1 U9427 ( .A1(n7845), .A2(n7832), .ZN(n7833) );
  NAND2_X1 U9428 ( .A1(n7834), .A2(n7833), .ZN(n7852) );
  NAND3_X1 U9429 ( .A1(n7835), .A2(n8461), .A3(n7845), .ZN(n7836) );
  NAND2_X1 U9430 ( .A1(n7838), .A2(n7847), .ZN(n7840) );
  NOR2_X1 U9431 ( .A1(n7838), .A2(n7847), .ZN(n7839) );
  AOI21_X1 U9432 ( .B1(n8786), .B2(n7840), .A(n7839), .ZN(n7841) );
  NAND2_X1 U9433 ( .A1(n7842), .A2(n7841), .ZN(n7843) );
  INV_X1 U9434 ( .A(n7844), .ZN(n7850) );
  NAND3_X1 U9435 ( .A1(n7846), .A2(n8867), .A3(n7845), .ZN(n7848) );
  NAND2_X1 U9436 ( .A1(n7848), .A2(n7847), .ZN(n7849) );
  NOR2_X1 U9437 ( .A1(n7850), .A2(n7849), .ZN(n7851) );
  OAI21_X1 U9438 ( .B1(n7852), .B2(n8461), .A(n7851), .ZN(n7853) );
  NAND2_X1 U9439 ( .A1(n7854), .A2(n7853), .ZN(n7862) );
  INV_X1 U9440 ( .A(n7858), .ZN(n7855) );
  NAND3_X1 U9441 ( .A1(n7862), .A2(n7856), .A3(n7855), .ZN(n7860) );
  AOI21_X1 U9442 ( .B1(n7858), .B2(n7857), .A(n7866), .ZN(n7859) );
  OAI211_X1 U9443 ( .C1(n7862), .C2(n7861), .A(n7860), .B(n7859), .ZN(n7869)
         );
  NOR3_X1 U9444 ( .A1(n7864), .A2(n6565), .A3(n7863), .ZN(n7868) );
  OAI21_X1 U9445 ( .B1(n7866), .B2(n7865), .A(P2_B_REG_SCAN_IN), .ZN(n7867) );
  OAI22_X1 U9446 ( .A1(n7870), .A2(n7869), .B1(n7868), .B2(n7867), .ZN(
        P2_U3296) );
  INV_X1 U9447 ( .A(n7871), .ZN(n7881) );
  INV_X1 U9448 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7885) );
  OAI21_X1 U9449 ( .B1(n7872), .B2(n7874), .A(n7873), .ZN(n7875) );
  NAND2_X1 U9450 ( .A1(n7875), .A2(n9056), .ZN(n7880) );
  INV_X1 U9451 ( .A(n9110), .ZN(n7876) );
  OAI22_X1 U9452 ( .A1(n7877), .A2(n9068), .B1(n9078), .B2(n7876), .ZN(n7878)
         );
  AOI21_X1 U9453 ( .B1(n7888), .B2(n9035), .A(n7878), .ZN(n7879) );
  OAI211_X1 U9454 ( .C1(n7881), .C2(n7885), .A(n7880), .B(n7879), .ZN(P1_U3222) );
  AOI22_X1 U9455 ( .A1(n9414), .A2(n7888), .B1(n9656), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n7882) );
  OAI21_X1 U9456 ( .B1(n7883), .B2(n9656), .A(n7882), .ZN(P1_U3523) );
  INV_X1 U9457 ( .A(n7884), .ZN(n7893) );
  OAI22_X1 U9458 ( .A1(n9363), .A2(n7886), .B1(n7885), .B2(n9211), .ZN(n7887)
         );
  AOI21_X1 U9459 ( .B1(n9359), .B2(n7888), .A(n7887), .ZN(n7892) );
  MUX2_X1 U9460 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n7889), .S(n9365), .Z(n7890)
         );
  INV_X1 U9461 ( .A(n7890), .ZN(n7891) );
  OAI211_X1 U9462 ( .C1(n7893), .C2(n9368), .A(n7892), .B(n7891), .ZN(P1_U3292) );
  OR2_X1 U9463 ( .A1(n5721), .A2(n7895), .ZN(n7896) );
  INV_X1 U9464 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n7906) );
  NAND2_X1 U9465 ( .A1(n8944), .A2(n7899), .ZN(n7898) );
  OR2_X1 U9466 ( .A1(n5721), .A2(n10062), .ZN(n7897) );
  NAND2_X1 U9467 ( .A1(n8220), .A2(n7899), .ZN(n7901) );
  OR2_X1 U9468 ( .A1(n5721), .A2(n8221), .ZN(n7900) );
  XNOR2_X1 U9469 ( .A(n9165), .B(n9171), .ZN(n7903) );
  NAND2_X1 U9470 ( .A1(n7903), .A2(n9354), .ZN(n9168) );
  INV_X1 U9471 ( .A(P1_B_REG_SCAN_IN), .ZN(n7904) );
  NOR2_X1 U9472 ( .A1(n6354), .A2(n7904), .ZN(n7905) );
  NOR2_X1 U9473 ( .A1(n9349), .A2(n7905), .ZN(n8202) );
  NAND2_X1 U9474 ( .A1(n8098), .A2(n8202), .ZN(n9369) );
  AND2_X1 U9475 ( .A1(n9168), .A2(n9369), .ZN(n7908) );
  MUX2_X1 U9476 ( .A(n7906), .B(n7908), .S(n9650), .Z(n7907) );
  OAI21_X1 U9477 ( .B1(n9165), .B2(n9445), .A(n7907), .ZN(P1_U3521) );
  INV_X1 U9478 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n7909) );
  MUX2_X1 U9479 ( .A(n7909), .B(n7908), .S(n9659), .Z(n7910) );
  OAI21_X1 U9480 ( .B1(n9165), .B2(n9384), .A(n7910), .ZN(P1_U3553) );
  INV_X1 U9481 ( .A(n7911), .ZN(n8223) );
  OAI222_X1 U9482 ( .A1(n7913), .A2(P2_U3151), .B1(n8947), .B2(n8223), .C1(
        n7912), .C2(n8945), .ZN(P2_U3271) );
  INV_X1 U9483 ( .A(n9165), .ZN(n8097) );
  NAND2_X1 U9484 ( .A1(n4332), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U9485 ( .A1(n5696), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7915) );
  NAND2_X1 U9486 ( .A1(n5699), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7914) );
  AND3_X1 U9487 ( .A1(n7916), .A2(n7915), .A3(n7914), .ZN(n7928) );
  INV_X1 U9488 ( .A(n7928), .ZN(n9088) );
  NAND2_X1 U9489 ( .A1(n7902), .A2(n9088), .ZN(n7938) );
  NAND2_X1 U9490 ( .A1(n8087), .A2(n8083), .ZN(n7926) );
  OR2_X1 U9491 ( .A1(n9398), .A2(n9283), .ZN(n7917) );
  NAND2_X1 U9492 ( .A1(n8065), .A2(n7917), .ZN(n7969) );
  AOI21_X1 U9493 ( .B1(n8066), .B2(n7969), .A(n7918), .ZN(n7920) );
  OAI21_X1 U9494 ( .B1(n7920), .B2(n7919), .A(n8078), .ZN(n7921) );
  NAND2_X1 U9495 ( .A1(n8057), .A2(n7971), .ZN(n7970) );
  NOR3_X1 U9496 ( .A1(n7926), .A2(n7921), .A3(n7970), .ZN(n8155) );
  INV_X1 U9497 ( .A(n7921), .ZN(n7925) );
  NAND3_X1 U9498 ( .A1(n8071), .A2(n7967), .A3(n7923), .ZN(n7924) );
  NAND2_X1 U9499 ( .A1(n8076), .A2(n8074), .ZN(n8079) );
  AOI21_X1 U9500 ( .B1(n7925), .B2(n7924), .A(n8079), .ZN(n7927) );
  NAND2_X1 U9501 ( .A1(n9373), .A2(n8196), .ZN(n7939) );
  AND2_X1 U9502 ( .A1(n7939), .A2(n9178), .ZN(n8199) );
  OAI21_X1 U9503 ( .B1(n7927), .B2(n7926), .A(n8199), .ZN(n8153) );
  AOI21_X1 U9504 ( .B1(n8155), .B2(n9297), .A(n8153), .ZN(n7932) );
  NAND2_X1 U9505 ( .A1(n8093), .A2(n9182), .ZN(n8158) );
  NAND2_X1 U9506 ( .A1(n9169), .A2(n7928), .ZN(n7930) );
  NAND2_X1 U9507 ( .A1(n8216), .A2(n7929), .ZN(n8094) );
  NAND2_X1 U9508 ( .A1(n7930), .A2(n8094), .ZN(n8156) );
  AOI21_X1 U9509 ( .B1(n7934), .B2(n9169), .A(n8156), .ZN(n7931) );
  OAI21_X1 U9510 ( .B1(n7932), .B2(n8158), .A(n7931), .ZN(n7933) );
  OAI21_X1 U9511 ( .B1(n7934), .B2(n7938), .A(n7933), .ZN(n7936) );
  AOI211_X1 U9512 ( .C1(n8099), .C2(n7936), .A(n7935), .B(n7937), .ZN(n7966)
         );
  INV_X1 U9513 ( .A(n7937), .ZN(n8166) );
  NAND2_X1 U9514 ( .A1(n8166), .A2(n7938), .ZN(n8107) );
  NAND2_X1 U9515 ( .A1(n7971), .A2(n7972), .ZN(n9296) );
  NAND2_X1 U9516 ( .A1(n8052), .A2(n7940), .ZN(n8147) );
  INV_X1 U9517 ( .A(n9312), .ZN(n7959) );
  NAND2_X1 U9518 ( .A1(n8043), .A2(n7941), .ZN(n8143) );
  NOR4_X1 U9519 ( .A1(n7947), .A2(n7946), .A3(n7945), .A4(n7944), .ZN(n7949)
         );
  INV_X1 U9520 ( .A(n7997), .ZN(n7948) );
  NAND4_X1 U9521 ( .A1(n7949), .A2(n7948), .A3(n6261), .A4(n6260), .ZN(n7950)
         );
  NOR4_X1 U9522 ( .A1(n7952), .A2(n8108), .A3(n7951), .A4(n7950), .ZN(n7953)
         );
  NAND4_X1 U9523 ( .A1(n8027), .A2(n7955), .A3(n7954), .A4(n7953), .ZN(n7956)
         );
  OR4_X1 U9524 ( .A1(n8143), .A2(n7957), .A3(n4727), .A4(n7956), .ZN(n7958) );
  NOR4_X1 U9525 ( .A1(n9296), .A2(n8147), .A3(n7959), .A4(n7958), .ZN(n7960)
         );
  NAND4_X1 U9526 ( .A1(n9247), .A2(n9282), .A3(n7960), .A4(n9271), .ZN(n7961)
         );
  NOR4_X1 U9527 ( .A1(n7963), .A2(n7962), .A3(n9236), .A4(n7961), .ZN(n7964)
         );
  NAND4_X1 U9528 ( .A1(n8093), .A2(n8195), .A3(n8191), .A4(n7964), .ZN(n7965)
         );
  NOR2_X1 U9529 ( .A1(n7966), .A2(n8104), .ZN(n8106) );
  INV_X1 U9530 ( .A(n7967), .ZN(n7968) );
  INV_X1 U9531 ( .A(n7970), .ZN(n8049) );
  NAND2_X1 U9532 ( .A1(n7971), .A2(n8044), .ZN(n7974) );
  NAND2_X1 U9533 ( .A1(n7972), .A2(n9338), .ZN(n7973) );
  MUX2_X1 U9534 ( .A(n7974), .B(n7973), .S(n8167), .Z(n7977) );
  OR2_X1 U9535 ( .A1(n9296), .A2(n7975), .ZN(n7976) );
  NAND2_X1 U9536 ( .A1(n7977), .A2(n7976), .ZN(n8055) );
  AND2_X1 U9537 ( .A1(n7978), .A2(n8114), .ZN(n7980) );
  NOR2_X1 U9538 ( .A1(n7978), .A2(n4715), .ZN(n7979) );
  MUX2_X1 U9539 ( .A(n7980), .B(n7979), .S(n8167), .Z(n7985) );
  MUX2_X1 U9540 ( .A(n8114), .B(n8118), .S(n8085), .Z(n7982) );
  NAND2_X1 U9541 ( .A1(n7982), .A2(n7981), .ZN(n7984) );
  NAND3_X1 U9542 ( .A1(n9626), .A2(n8085), .A3(n9107), .ZN(n7983) );
  OAI21_X1 U9543 ( .B1(n7985), .B2(n7984), .A(n7983), .ZN(n7993) );
  NAND2_X1 U9544 ( .A1(n7993), .A2(n7991), .ZN(n7989) );
  INV_X1 U9545 ( .A(n7986), .ZN(n7987) );
  AND2_X1 U9546 ( .A1(n7987), .A2(n8123), .ZN(n7992) );
  AOI21_X1 U9547 ( .B1(n7989), .B2(n7992), .A(n7988), .ZN(n7994) );
  NAND2_X1 U9548 ( .A1(n7991), .A2(n7990), .ZN(n8120) );
  AOI21_X1 U9549 ( .B1(n7996), .B2(n7995), .A(n8167), .ZN(n7998) );
  NOR2_X1 U9550 ( .A1(n7998), .A2(n7997), .ZN(n7999) );
  NAND2_X1 U9551 ( .A1(n8000), .A2(n7999), .ZN(n8004) );
  INV_X1 U9552 ( .A(n8001), .ZN(n8002) );
  MUX2_X1 U9553 ( .A(n8002), .B(n4392), .S(n8167), .Z(n8003) );
  NAND2_X1 U9554 ( .A1(n8004), .A2(n8003), .ZN(n8013) );
  INV_X1 U9555 ( .A(n8005), .ZN(n8128) );
  AOI21_X1 U9556 ( .B1(n8013), .B2(n6261), .A(n8128), .ZN(n8008) );
  NAND2_X1 U9557 ( .A1(n8016), .A2(n8010), .ZN(n8131) );
  OR2_X1 U9558 ( .A1(n8131), .A2(n8085), .ZN(n8007) );
  AND2_X1 U9559 ( .A1(n8018), .A2(n8006), .ZN(n8014) );
  OAI22_X1 U9560 ( .A1(n8008), .A2(n8007), .B1(n8014), .B2(n8085), .ZN(n8009)
         );
  NAND2_X1 U9561 ( .A1(n8009), .A2(n8133), .ZN(n8021) );
  INV_X1 U9562 ( .A(n8010), .ZN(n8011) );
  AOI21_X1 U9563 ( .B1(n8013), .B2(n8012), .A(n8011), .ZN(n8015) );
  INV_X1 U9564 ( .A(n8014), .ZN(n8136) );
  INV_X1 U9565 ( .A(n8016), .ZN(n8019) );
  INV_X1 U9566 ( .A(n8133), .ZN(n8017) );
  AOI21_X1 U9567 ( .B1(n8019), .B2(n8018), .A(n8017), .ZN(n8020) );
  INV_X1 U9568 ( .A(n8137), .ZN(n8022) );
  OAI211_X1 U9569 ( .C1(n8029), .C2(n8022), .A(n8134), .B(n8025), .ZN(n8023)
         );
  AND4_X1 U9570 ( .A1(n8023), .A2(n8139), .A3(n8142), .A4(n8141), .ZN(n8034)
         );
  NAND2_X1 U9571 ( .A1(n8140), .A2(n9096), .ZN(n8024) );
  NAND2_X1 U9572 ( .A1(n8024), .A2(n8085), .ZN(n8039) );
  NAND2_X1 U9573 ( .A1(n8039), .A2(n9081), .ZN(n8032) );
  AND2_X1 U9574 ( .A1(n8035), .A2(n8025), .ZN(n8026) );
  AND2_X1 U9575 ( .A1(n8140), .A2(n8026), .ZN(n8146) );
  INV_X1 U9576 ( .A(n8134), .ZN(n8028) );
  OAI211_X1 U9577 ( .C1(n8029), .C2(n8028), .A(n8027), .B(n8137), .ZN(n8030)
         );
  NAND2_X1 U9578 ( .A1(n8146), .A2(n8030), .ZN(n8031) );
  NAND3_X1 U9579 ( .A1(n8032), .A2(n8031), .A3(n8141), .ZN(n8033) );
  INV_X1 U9580 ( .A(n8035), .ZN(n8036) );
  NAND2_X1 U9581 ( .A1(n8141), .A2(n8036), .ZN(n8037) );
  NAND2_X1 U9582 ( .A1(n8037), .A2(n8140), .ZN(n8038) );
  AND2_X1 U9583 ( .A1(n8039), .A2(n8038), .ZN(n8041) );
  INV_X1 U9584 ( .A(n8040), .ZN(n9346) );
  INV_X1 U9585 ( .A(n8147), .ZN(n8042) );
  AND2_X1 U9586 ( .A1(n8044), .A2(n8043), .ZN(n8149) );
  NAND2_X1 U9587 ( .A1(n8055), .A2(n8045), .ZN(n8048) );
  INV_X1 U9588 ( .A(n8046), .ZN(n8047) );
  AOI21_X1 U9589 ( .B1(n8049), .B2(n8048), .A(n8047), .ZN(n8062) );
  INV_X1 U9590 ( .A(n8143), .ZN(n8050) );
  NAND2_X1 U9591 ( .A1(n8051), .A2(n8050), .ZN(n8053) );
  NAND3_X1 U9592 ( .A1(n8053), .A2(n8150), .A3(n8052), .ZN(n8054) );
  NAND2_X1 U9593 ( .A1(n8055), .A2(n8054), .ZN(n8060) );
  INV_X1 U9594 ( .A(n8056), .ZN(n8059) );
  INV_X1 U9595 ( .A(n8057), .ZN(n8058) );
  AOI21_X1 U9596 ( .B1(n8060), .B2(n8059), .A(n8058), .ZN(n8061) );
  MUX2_X1 U9597 ( .A(n8062), .B(n8061), .S(n8085), .Z(n8064) );
  INV_X1 U9598 ( .A(n9271), .ZN(n8063) );
  NOR2_X1 U9599 ( .A1(n8064), .A2(n8063), .ZN(n8068) );
  MUX2_X1 U9600 ( .A(n8066), .B(n8065), .S(n8167), .Z(n8067) );
  MUX2_X1 U9601 ( .A(n8071), .B(n8070), .S(n8085), .Z(n8072) );
  NAND2_X1 U9602 ( .A1(n8073), .A2(n8072), .ZN(n8082) );
  INV_X1 U9603 ( .A(n8074), .ZN(n8075) );
  OAI211_X1 U9604 ( .C1(n8082), .C2(n8075), .A(n8083), .B(n8078), .ZN(n8077)
         );
  INV_X1 U9605 ( .A(n8078), .ZN(n8081) );
  INV_X1 U9606 ( .A(n8079), .ZN(n8080) );
  OAI21_X1 U9607 ( .B1(n8082), .B2(n8081), .A(n8080), .ZN(n8084) );
  INV_X1 U9608 ( .A(n8199), .ZN(n8088) );
  OAI21_X1 U9609 ( .B1(n8088), .B2(n8087), .A(n9182), .ZN(n8089) );
  NAND2_X1 U9610 ( .A1(n8089), .A2(n8167), .ZN(n8090) );
  NAND2_X1 U9611 ( .A1(n8091), .A2(n8090), .ZN(n8092) );
  NAND2_X1 U9612 ( .A1(n8092), .A2(n8201), .ZN(n8096) );
  OAI211_X1 U9613 ( .C1(n9169), .C2(n8167), .A(n8097), .B(n9088), .ZN(n8101)
         );
  AOI22_X1 U9614 ( .A1(n9169), .A2(n8167), .B1(n8098), .B2(n9088), .ZN(n8100)
         );
  AOI22_X1 U9615 ( .A1(n8165), .A2(n8103), .B1(n4331), .B2(n8102), .ZN(n8105)
         );
  OAI22_X1 U9616 ( .A1(n4331), .A2(n8106), .B1(n8105), .B2(n8104), .ZN(n8175)
         );
  INV_X1 U9617 ( .A(n8107), .ZN(n8161) );
  INV_X1 U9618 ( .A(n8108), .ZN(n8127) );
  INV_X1 U9619 ( .A(n8109), .ZN(n8112) );
  NAND2_X1 U9620 ( .A1(n9109), .A2(n8110), .ZN(n8111) );
  NAND3_X1 U9621 ( .A1(n8112), .A2(n6152), .A3(n8111), .ZN(n8113) );
  NAND2_X1 U9622 ( .A1(n6256), .A2(n8113), .ZN(n8116) );
  OAI211_X1 U9623 ( .C1(n8117), .C2(n8116), .A(n8115), .B(n8114), .ZN(n8119)
         );
  NAND2_X1 U9624 ( .A1(n8119), .A2(n8118), .ZN(n8122) );
  AOI21_X1 U9625 ( .B1(n8122), .B2(n8121), .A(n8120), .ZN(n8125) );
  INV_X1 U9626 ( .A(n8123), .ZN(n8124) );
  OAI21_X1 U9627 ( .B1(n8125), .B2(n8124), .A(n6260), .ZN(n8126) );
  NAND2_X1 U9628 ( .A1(n8127), .A2(n8126), .ZN(n8130) );
  AOI21_X1 U9629 ( .B1(n8130), .B2(n8129), .A(n8128), .ZN(n8132) );
  NOR2_X1 U9630 ( .A1(n8132), .A2(n8131), .ZN(n8135) );
  OAI211_X1 U9631 ( .C1(n8136), .C2(n8135), .A(n8134), .B(n8133), .ZN(n8138)
         );
  NAND3_X1 U9632 ( .A1(n8139), .A2(n8138), .A3(n8137), .ZN(n8145) );
  OAI21_X1 U9633 ( .B1(n4729), .B2(n8142), .A(n8141), .ZN(n8144) );
  AOI211_X1 U9634 ( .C1(n8146), .C2(n8145), .A(n8144), .B(n8143), .ZN(n8148)
         );
  NOR2_X1 U9635 ( .A1(n8148), .A2(n8147), .ZN(n8152) );
  INV_X1 U9636 ( .A(n8149), .ZN(n8151) );
  OAI21_X1 U9637 ( .B1(n8152), .B2(n8151), .A(n8150), .ZN(n8154) );
  AOI21_X1 U9638 ( .B1(n8155), .B2(n8154), .A(n8153), .ZN(n8159) );
  INV_X1 U9639 ( .A(n8156), .ZN(n8157) );
  OAI21_X1 U9640 ( .B1(n8159), .B2(n8158), .A(n8157), .ZN(n8160) );
  XNOR2_X1 U9641 ( .A(n8162), .B(n4331), .ZN(n8164) );
  OAI21_X1 U9642 ( .B1(n8167), .B2(n8166), .A(n8165), .ZN(n8171) );
  AOI211_X1 U9643 ( .C1(n8169), .C2(n4331), .A(n6151), .B(n8168), .ZN(n8170)
         );
  NAND2_X1 U9644 ( .A1(n8173), .A2(n8172), .ZN(n8174) );
  AOI21_X1 U9645 ( .B1(n6272), .B2(n8175), .A(n8174), .ZN(n8180) );
  NAND2_X1 U9646 ( .A1(n8176), .A2(n9507), .ZN(n8177) );
  OAI211_X1 U9647 ( .C1(n6151), .C2(n8179), .A(n8177), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8178) );
  OAI21_X1 U9648 ( .B1(n8180), .B2(n8179), .A(n8178), .ZN(P1_U3242) );
  OAI21_X1 U9649 ( .B1(n8183), .B2(n8182), .A(n8181), .ZN(n8184) );
  NAND2_X1 U9650 ( .A1(n8184), .A2(n9056), .ZN(n8188) );
  AOI22_X1 U9651 ( .A1(n9076), .A2(n9091), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8185) );
  OAI21_X1 U9652 ( .B1(n9238), .B2(n9078), .A(n8185), .ZN(n8186) );
  AOI21_X1 U9653 ( .B1(n9241), .B2(n9084), .A(n8186), .ZN(n8187) );
  OAI211_X1 U9654 ( .C1(n6268), .C2(n9080), .A(n8188), .B(n8187), .ZN(P1_U3229) );
  OAI222_X1 U9655 ( .A1(n9490), .A2(n8190), .B1(n9493), .B2(n8189), .C1(
        P1_U3086), .C2(n9203), .ZN(P1_U3336) );
  INV_X1 U9656 ( .A(n8191), .ZN(n8193) );
  NAND2_X1 U9657 ( .A1(n9176), .A2(n9179), .ZN(n9175) );
  OAI21_X1 U9658 ( .B1(n8196), .B2(n4585), .A(n9175), .ZN(n8198) );
  INV_X1 U9659 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U9660 ( .A1(n9177), .A2(n8199), .ZN(n9184) );
  NAND2_X1 U9661 ( .A1(n9184), .A2(n9182), .ZN(n8200) );
  XNOR2_X1 U9662 ( .A(n8201), .B(n8200), .ZN(n8204) );
  AOI22_X1 U9663 ( .A1(n9089), .A2(n9335), .B1(n9088), .B2(n8202), .ZN(n8203)
         );
  AOI21_X1 U9664 ( .B1(n8216), .B2(n9190), .A(n9326), .ZN(n8205) );
  AND2_X1 U9665 ( .A1(n8205), .A2(n4359), .ZN(n8208) );
  MUX2_X1 U9666 ( .A(n9987), .B(n8214), .S(n9659), .Z(n8207) );
  NAND2_X1 U9667 ( .A1(n8216), .A2(n9414), .ZN(n8206) );
  OAI211_X1 U9668 ( .C1(n8219), .C2(n9427), .A(n8207), .B(n8206), .ZN(P1_U3551) );
  AOI22_X1 U9669 ( .A1(n8216), .A2(n9359), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9358), .ZN(n8213) );
  NAND2_X1 U9670 ( .A1(n8208), .A2(n9203), .ZN(n8209) );
  OAI21_X1 U9671 ( .B1(n9211), .B2(n8210), .A(n8209), .ZN(n8211) );
  OAI211_X1 U9672 ( .C1(n8219), .C2(n9368), .A(n8213), .B(n8212), .ZN(P1_U3356) );
  INV_X1 U9673 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8215) );
  MUX2_X1 U9674 ( .A(n8215), .B(n8214), .S(n9650), .Z(n8218) );
  NAND2_X1 U9675 ( .A1(n8216), .A2(n9471), .ZN(n8217) );
  OAI211_X1 U9676 ( .C1(n8219), .C2(n9478), .A(n8218), .B(n8217), .ZN(P1_U3519) );
  INV_X1 U9677 ( .A(n8220), .ZN(n8233) );
  OAI222_X1 U9678 ( .A1(n9490), .A2(n8221), .B1(n9493), .B2(n8233), .C1(
        P1_U3086), .C2(n5640), .ZN(P1_U3325) );
  OAI222_X1 U9679 ( .A1(n9493), .A2(n8223), .B1(n6132), .B2(P1_U3086), .C1(
        n8222), .C2(n9490), .ZN(P1_U3331) );
  INV_X1 U9680 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8225) );
  NAND2_X1 U9681 ( .A1(n8619), .A2(n8933), .ZN(n8226) );
  NAND2_X1 U9682 ( .A1(n8227), .A2(n8226), .ZN(P2_U3456) );
  AOI22_X1 U9683 ( .A1(n9958), .A2(n8229), .B1(n8228), .B2(n9950), .ZN(n8232)
         );
  NAND2_X1 U9684 ( .A1(n8230), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8231) );
  OAI211_X1 U9685 ( .C1(n5118), .C2(n8427), .A(n8232), .B(n8231), .ZN(P2_U3172) );
  OAI222_X1 U9686 ( .A1(n5080), .A2(P2_U3151), .B1(n8947), .B2(n8233), .C1(
        n9995), .C2(n8945), .ZN(P2_U3265) );
  XNOR2_X1 U9687 ( .A(n8877), .B(n6784), .ZN(n8277) );
  XNOR2_X1 U9688 ( .A(n8804), .B(n6784), .ZN(n8296) );
  OAI21_X1 U9689 ( .B1(n8235), .B2(n9951), .A(n8234), .ZN(n8237) );
  NAND2_X1 U9690 ( .A1(n8235), .A2(n9951), .ZN(n8236) );
  NAND2_X1 U9691 ( .A1(n8237), .A2(n8236), .ZN(n8400) );
  XNOR2_X1 U9692 ( .A(n8408), .B(n6784), .ZN(n8239) );
  NAND2_X1 U9693 ( .A1(n8239), .A2(n8238), .ZN(n8242) );
  INV_X1 U9694 ( .A(n8239), .ZN(n8240) );
  NAND2_X1 U9695 ( .A1(n8240), .A2(n8465), .ZN(n8241) );
  NAND2_X1 U9696 ( .A1(n8242), .A2(n8241), .ZN(n8401) );
  XNOR2_X1 U9697 ( .A(n8286), .B(n6784), .ZN(n8244) );
  XNOR2_X1 U9698 ( .A(n8244), .B(n8464), .ZN(n8283) );
  XNOR2_X1 U9699 ( .A(n8243), .B(n6784), .ZN(n8246) );
  XNOR2_X1 U9700 ( .A(n8246), .B(n8770), .ZN(n8449) );
  NAND2_X1 U9701 ( .A1(n8244), .A2(n8402), .ZN(n8446) );
  AND2_X1 U9702 ( .A1(n8449), .A2(n8446), .ZN(n8245) );
  INV_X1 U9703 ( .A(n8246), .ZN(n8247) );
  NAND2_X1 U9704 ( .A1(n8247), .A2(n8770), .ZN(n8248) );
  NAND2_X1 U9705 ( .A1(n8448), .A2(n8248), .ZN(n8359) );
  XNOR2_X1 U9706 ( .A(n8934), .B(n6784), .ZN(n8354) );
  NAND2_X1 U9707 ( .A1(n8354), .A2(n8353), .ZN(n8249) );
  NAND2_X1 U9708 ( .A1(n8359), .A2(n8249), .ZN(n8355) );
  XNOR2_X1 U9709 ( .A(n8927), .B(n6784), .ZN(n8251) );
  NAND2_X1 U9710 ( .A1(n8251), .A2(n8250), .ZN(n8256) );
  INV_X1 U9711 ( .A(n8251), .ZN(n8252) );
  NAND2_X1 U9712 ( .A1(n8252), .A2(n8772), .ZN(n8253) );
  NAND2_X1 U9713 ( .A1(n8256), .A2(n8253), .ZN(n8368) );
  INV_X1 U9714 ( .A(n8354), .ZN(n8254) );
  AND2_X1 U9715 ( .A1(n8254), .A2(n8757), .ZN(n8369) );
  NOR2_X1 U9716 ( .A1(n8368), .A2(n8369), .ZN(n8255) );
  NAND2_X1 U9717 ( .A1(n8355), .A2(n8255), .ZN(n8371) );
  NAND2_X1 U9718 ( .A1(n8371), .A2(n8256), .ZN(n8424) );
  XNOR2_X1 U9719 ( .A(n8921), .B(n6784), .ZN(n8257) );
  XNOR2_X1 U9720 ( .A(n8257), .B(n8758), .ZN(n8423) );
  NAND2_X1 U9721 ( .A1(n8424), .A2(n8423), .ZN(n8422) );
  XNOR2_X1 U9722 ( .A(n8738), .B(n6784), .ZN(n8262) );
  XNOR2_X1 U9723 ( .A(n8262), .B(n8748), .ZN(n8317) );
  NAND2_X1 U9724 ( .A1(n8257), .A2(n8365), .ZN(n8316) );
  AND2_X1 U9725 ( .A1(n8317), .A2(n8316), .ZN(n8258) );
  XNOR2_X1 U9726 ( .A(n8909), .B(n6784), .ZN(n8259) );
  NAND2_X1 U9727 ( .A1(n8259), .A2(n8699), .ZN(n8332) );
  INV_X1 U9728 ( .A(n8259), .ZN(n8260) );
  NAND2_X1 U9729 ( .A1(n8260), .A2(n8731), .ZN(n8261) );
  NAND2_X1 U9730 ( .A1(n8332), .A2(n8261), .ZN(n8388) );
  INV_X1 U9731 ( .A(n8262), .ZN(n8263) );
  AND2_X1 U9732 ( .A1(n8263), .A2(n8748), .ZN(n8387) );
  NOR2_X1 U9733 ( .A1(n8388), .A2(n8387), .ZN(n8264) );
  XNOR2_X1 U9734 ( .A(n8810), .B(n6784), .ZN(n8265) );
  NAND2_X1 U9735 ( .A1(n8265), .A2(n8417), .ZN(n8268) );
  INV_X1 U9736 ( .A(n8265), .ZN(n8266) );
  NAND2_X1 U9737 ( .A1(n8266), .A2(n8718), .ZN(n8267) );
  AND2_X1 U9738 ( .A1(n8268), .A2(n8267), .ZN(n8333) );
  NAND2_X1 U9739 ( .A1(n8334), .A2(n8268), .ZN(n8414) );
  XNOR2_X1 U9740 ( .A(n8899), .B(n6784), .ZN(n8269) );
  XNOR2_X1 U9741 ( .A(n8269), .B(n8463), .ZN(n8413) );
  NAND2_X1 U9742 ( .A1(n8414), .A2(n8413), .ZN(n8412) );
  NAND2_X1 U9743 ( .A1(n8269), .A2(n8700), .ZN(n8270) );
  XNOR2_X1 U9744 ( .A(n8889), .B(n7232), .ZN(n8271) );
  NAND2_X1 U9745 ( .A1(n8271), .A2(n8462), .ZN(n8342) );
  OAI211_X1 U9746 ( .C1(n8382), .C2(n8296), .A(n8297), .B(n8342), .ZN(n8274)
         );
  INV_X1 U9747 ( .A(n8271), .ZN(n8272) );
  NAND2_X1 U9748 ( .A1(n8272), .A2(n8680), .ZN(n8343) );
  NAND3_X1 U9749 ( .A1(n8342), .A2(n8382), .A3(n8296), .ZN(n8273) );
  NAND3_X1 U9750 ( .A1(n8274), .A2(n8343), .A3(n8273), .ZN(n8275) );
  XNOR2_X1 U9751 ( .A(n8883), .B(n6784), .ZN(n8276) );
  XNOR2_X1 U9752 ( .A(n8276), .B(n8668), .ZN(n8344) );
  NAND2_X1 U9753 ( .A1(n8275), .A2(n8344), .ZN(n8435) );
  NAND2_X1 U9754 ( .A1(n8276), .A2(n8441), .ZN(n8434) );
  XNOR2_X1 U9755 ( .A(n8277), .B(n8655), .ZN(n8437) );
  NAND3_X1 U9756 ( .A1(n8435), .A2(n8434), .A3(n8437), .ZN(n8436) );
  XNOR2_X1 U9757 ( .A(n8791), .B(n6784), .ZN(n8323) );
  XNOR2_X1 U9758 ( .A(n8323), .B(n8646), .ZN(n8325) );
  XNOR2_X1 U9759 ( .A(n8326), .B(n8325), .ZN(n8282) );
  AOI22_X1 U9760 ( .A1(n8461), .A2(n9952), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8279) );
  NAND2_X1 U9761 ( .A1(n9948), .A2(n8637), .ZN(n8278) );
  OAI211_X1 U9762 ( .C1(n8636), .C2(n8440), .A(n8279), .B(n8278), .ZN(n8280)
         );
  AOI21_X1 U9763 ( .B1(n8791), .B2(n9950), .A(n8280), .ZN(n8281) );
  OAI21_X1 U9764 ( .B1(n8282), .B2(n8410), .A(n8281), .ZN(P2_U3154) );
  OAI21_X1 U9765 ( .B1(n8284), .B2(n8283), .A(n8447), .ZN(n8294) );
  INV_X1 U9766 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8285) );
  NOR2_X1 U9767 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8285), .ZN(n9821) );
  AOI21_X1 U9768 ( .B1(n9952), .B2(n8770), .A(n9821), .ZN(n8292) );
  NAND2_X1 U9769 ( .A1(n8286), .A2(n9950), .ZN(n8291) );
  INV_X1 U9770 ( .A(n8287), .ZN(n8288) );
  NAND2_X1 U9771 ( .A1(n9948), .A2(n8288), .ZN(n8290) );
  NAND2_X1 U9772 ( .A1(n9945), .A2(n8465), .ZN(n8289) );
  NAND4_X1 U9773 ( .A1(n8292), .A2(n8291), .A3(n8290), .A4(n8289), .ZN(n8293)
         );
  AOI21_X1 U9774 ( .B1(n8294), .B2(n9958), .A(n8293), .ZN(n8295) );
  INV_X1 U9775 ( .A(n8295), .ZN(P2_U3155) );
  OR2_X1 U9776 ( .A1(n8297), .A2(n8296), .ZN(n8298) );
  NAND2_X1 U9777 ( .A1(n8298), .A2(n8382), .ZN(n8378) );
  INV_X1 U9778 ( .A(n8378), .ZN(n8300) );
  NAND2_X1 U9779 ( .A1(n8297), .A2(n8296), .ZN(n8377) );
  AOI21_X1 U9780 ( .B1(n8298), .B2(n8377), .A(n8382), .ZN(n8299) );
  AOI21_X1 U9781 ( .B1(n8300), .B2(n8377), .A(n8299), .ZN(n8305) );
  NAND2_X1 U9782 ( .A1(n9948), .A2(n8681), .ZN(n8302) );
  AOI22_X1 U9783 ( .A1(n9952), .A2(n8462), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8301) );
  OAI211_X1 U9784 ( .C1(n8700), .C2(n8440), .A(n8302), .B(n8301), .ZN(n8303)
         );
  AOI21_X1 U9785 ( .B1(n8804), .B2(n9950), .A(n8303), .ZN(n8304) );
  OAI21_X1 U9786 ( .B1(n8305), .B2(n8410), .A(n8304), .ZN(P2_U3156) );
  XNOR2_X1 U9787 ( .A(n8306), .B(n9944), .ZN(n9938) );
  XNOR2_X1 U9788 ( .A(n9938), .B(n9937), .ZN(n8307) );
  NAND2_X1 U9789 ( .A1(n8307), .A2(n9958), .ZN(n8315) );
  INV_X1 U9790 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8308) );
  NOR2_X1 U9791 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8308), .ZN(n9755) );
  AOI21_X1 U9792 ( .B1(n9945), .B2(n8466), .A(n9755), .ZN(n8314) );
  AOI22_X1 U9793 ( .A1(n9952), .A2(n4441), .B1(n8309), .B2(n9950), .ZN(n8313)
         );
  INV_X1 U9794 ( .A(n8310), .ZN(n8311) );
  NAND2_X1 U9795 ( .A1(n9948), .A2(n8311), .ZN(n8312) );
  NAND4_X1 U9796 ( .A1(n8315), .A2(n8314), .A3(n8313), .A4(n8312), .ZN(
        P2_U3157) );
  INV_X1 U9797 ( .A(n8738), .ZN(n8915) );
  AND2_X1 U9798 ( .A1(n8422), .A2(n8316), .ZN(n8318) );
  OAI211_X1 U9799 ( .C1(n8318), .C2(n8317), .A(n9958), .B(n8391), .ZN(n8322)
         );
  NAND2_X1 U9800 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8594) );
  OAI21_X1 U9801 ( .B1(n8427), .B2(n8699), .A(n8594), .ZN(n8320) );
  NOR2_X1 U9802 ( .A1(n8428), .A2(n8736), .ZN(n8319) );
  AOI211_X1 U9803 ( .C1(n9945), .C2(n8758), .A(n8320), .B(n8319), .ZN(n8321)
         );
  OAI211_X1 U9804 ( .C1(n8915), .C2(n8458), .A(n8322), .B(n8321), .ZN(P2_U3159) );
  INV_X1 U9805 ( .A(n8323), .ZN(n8324) );
  XNOR2_X1 U9806 ( .A(n4356), .B(n6784), .ZN(n8327) );
  AOI22_X1 U9807 ( .A1(n9945), .A2(n8646), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8329) );
  NAND2_X1 U9808 ( .A1(n9948), .A2(n8627), .ZN(n8328) );
  OAI211_X1 U9809 ( .C1(n8460), .C2(n8427), .A(n8329), .B(n8328), .ZN(n8330)
         );
  AOI21_X1 U9810 ( .B1(n8867), .B2(n9950), .A(n8330), .ZN(n8331) );
  INV_X1 U9811 ( .A(n8810), .ZN(n8341) );
  NOR3_X1 U9812 ( .A1(n4399), .A2(n4819), .A3(n8333), .ZN(n8336) );
  INV_X1 U9813 ( .A(n8334), .ZN(n8335) );
  OAI21_X1 U9814 ( .B1(n8336), .B2(n8335), .A(n9958), .ZN(n8340) );
  AOI22_X1 U9815 ( .A1(n9952), .A2(n8463), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8337) );
  OAI21_X1 U9816 ( .B1(n8699), .B2(n8440), .A(n8337), .ZN(n8338) );
  AOI21_X1 U9817 ( .B1(n8703), .B2(n9948), .A(n8338), .ZN(n8339) );
  OAI211_X1 U9818 ( .C1(n8341), .C2(n8458), .A(n8340), .B(n8339), .ZN(P2_U3163) );
  INV_X1 U9819 ( .A(n8883), .ZN(n8352) );
  NAND2_X1 U9820 ( .A1(n8342), .A2(n8343), .ZN(n8376) );
  AOI21_X1 U9821 ( .B1(n8378), .B2(n8377), .A(n8376), .ZN(n8380) );
  INV_X1 U9822 ( .A(n8343), .ZN(n8345) );
  NOR3_X1 U9823 ( .A1(n8380), .A2(n8345), .A3(n8344), .ZN(n8347) );
  INV_X1 U9824 ( .A(n8435), .ZN(n8346) );
  OAI21_X1 U9825 ( .B1(n8347), .B2(n8346), .A(n9958), .ZN(n8351) );
  AOI22_X1 U9826 ( .A1(n9952), .A2(n8655), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8348) );
  OAI21_X1 U9827 ( .B1(n8680), .B2(n8440), .A(n8348), .ZN(n8349) );
  AOI21_X1 U9828 ( .B1(n8660), .B2(n9948), .A(n8349), .ZN(n8350) );
  OAI211_X1 U9829 ( .C1(n8352), .C2(n8458), .A(n8351), .B(n8350), .ZN(P2_U3165) );
  INV_X1 U9830 ( .A(n8359), .ZN(n8357) );
  XNOR2_X1 U9831 ( .A(n8354), .B(n8353), .ZN(n8356) );
  INV_X1 U9832 ( .A(n8355), .ZN(n8370) );
  AOI21_X1 U9833 ( .B1(n8357), .B2(n8356), .A(n8370), .ZN(n8358) );
  AOI21_X1 U9834 ( .B1(n8369), .B2(n8359), .A(n8358), .ZN(n8364) );
  AOI22_X1 U9835 ( .A1(n9952), .A2(n8772), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3151), .ZN(n8361) );
  NAND2_X1 U9836 ( .A1(n9945), .A2(n8770), .ZN(n8360) );
  OAI211_X1 U9837 ( .C1(n8428), .C2(n8775), .A(n8361), .B(n8360), .ZN(n8362)
         );
  AOI21_X1 U9838 ( .B1(n8934), .B2(n9950), .A(n8362), .ZN(n8363) );
  OAI21_X1 U9839 ( .B1(n8364), .B2(n8410), .A(n8363), .ZN(P2_U3166) );
  AND2_X1 U9840 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8549) );
  NOR2_X1 U9841 ( .A1(n8427), .A2(n8365), .ZN(n8366) );
  AOI211_X1 U9842 ( .C1(n9945), .C2(n8757), .A(n8549), .B(n8366), .ZN(n8367)
         );
  OAI21_X1 U9843 ( .B1(n8761), .B2(n8428), .A(n8367), .ZN(n8374) );
  OAI21_X1 U9844 ( .B1(n8370), .B2(n8369), .A(n8368), .ZN(n8372) );
  AOI21_X1 U9845 ( .B1(n8372), .B2(n8371), .A(n8410), .ZN(n8373) );
  AOI211_X1 U9846 ( .C1(n8927), .C2(n9950), .A(n8374), .B(n8373), .ZN(n8375)
         );
  INV_X1 U9847 ( .A(n8375), .ZN(P2_U3168) );
  AND3_X1 U9848 ( .A1(n8378), .A2(n8377), .A3(n8376), .ZN(n8379) );
  OAI21_X1 U9849 ( .B1(n8380), .B2(n8379), .A(n9958), .ZN(n8385) );
  AOI22_X1 U9850 ( .A1(n9952), .A2(n8668), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8381) );
  OAI21_X1 U9851 ( .B1(n8382), .B2(n8440), .A(n8381), .ZN(n8383) );
  AOI21_X1 U9852 ( .B1(n8671), .B2(n9948), .A(n8383), .ZN(n8384) );
  OAI211_X1 U9853 ( .C1(n8386), .C2(n8458), .A(n8385), .B(n8384), .ZN(P2_U3169) );
  INV_X1 U9854 ( .A(n8909), .ZN(n8397) );
  INV_X1 U9855 ( .A(n8387), .ZN(n8390) );
  INV_X1 U9856 ( .A(n8388), .ZN(n8389) );
  AOI21_X1 U9857 ( .B1(n8391), .B2(n8390), .A(n8389), .ZN(n8392) );
  OAI21_X1 U9858 ( .B1(n4399), .B2(n8392), .A(n9958), .ZN(n8396) );
  AOI22_X1 U9859 ( .A1(n9952), .A2(n8718), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8393) );
  OAI21_X1 U9860 ( .B1(n8426), .B2(n8440), .A(n8393), .ZN(n8394) );
  AOI21_X1 U9861 ( .B1(n8714), .B2(n9948), .A(n8394), .ZN(n8395) );
  OAI211_X1 U9862 ( .C1(n8397), .C2(n8458), .A(n8396), .B(n8395), .ZN(P2_U3173) );
  INV_X1 U9863 ( .A(n8398), .ZN(n8399) );
  AOI21_X1 U9864 ( .B1(n8401), .B2(n8400), .A(n8399), .ZN(n8411) );
  NAND2_X1 U9865 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9809) );
  INV_X1 U9866 ( .A(n9809), .ZN(n8404) );
  NOR2_X1 U9867 ( .A1(n8427), .A2(n8402), .ZN(n8403) );
  AOI211_X1 U9868 ( .C1(n9945), .C2(n9951), .A(n8404), .B(n8403), .ZN(n8405)
         );
  OAI21_X1 U9869 ( .B1(n8406), .B2(n8428), .A(n8405), .ZN(n8407) );
  AOI21_X1 U9870 ( .B1(n8408), .B2(n9950), .A(n8407), .ZN(n8409) );
  OAI21_X1 U9871 ( .B1(n8411), .B2(n8410), .A(n8409), .ZN(P2_U3174) );
  INV_X1 U9872 ( .A(n8899), .ZN(n8421) );
  OAI21_X1 U9873 ( .B1(n8414), .B2(n8413), .A(n8412), .ZN(n8415) );
  NAND2_X1 U9874 ( .A1(n8415), .A2(n9958), .ZN(n8420) );
  AOI22_X1 U9875 ( .A1(n9952), .A2(n8691), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8416) );
  OAI21_X1 U9876 ( .B1(n8417), .B2(n8440), .A(n8416), .ZN(n8418) );
  AOI21_X1 U9877 ( .B1(n8695), .B2(n9948), .A(n8418), .ZN(n8419) );
  OAI211_X1 U9878 ( .C1(n8421), .C2(n8458), .A(n8420), .B(n8419), .ZN(P2_U3175) );
  INV_X1 U9879 ( .A(n8921), .ZN(n8433) );
  OAI21_X1 U9880 ( .B1(n8424), .B2(n8423), .A(n8422), .ZN(n8425) );
  NAND2_X1 U9881 ( .A1(n8425), .A2(n9958), .ZN(n8432) );
  NAND2_X1 U9882 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8573) );
  OAI21_X1 U9883 ( .B1(n8427), .B2(n8426), .A(n8573), .ZN(n8430) );
  NOR2_X1 U9884 ( .A1(n8428), .A2(n8750), .ZN(n8429) );
  AOI211_X1 U9885 ( .C1(n9945), .C2(n8772), .A(n8430), .B(n8429), .ZN(n8431)
         );
  OAI211_X1 U9886 ( .C1(n8433), .C2(n8458), .A(n8432), .B(n8431), .ZN(P2_U3178) );
  AND2_X1 U9887 ( .A1(n8435), .A2(n8434), .ZN(n8438) );
  OAI211_X1 U9888 ( .C1(n8438), .C2(n8437), .A(n9958), .B(n8436), .ZN(n8444)
         );
  AOI22_X1 U9889 ( .A1(n9952), .A2(n8646), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8439) );
  OAI21_X1 U9890 ( .B1(n8441), .B2(n8440), .A(n8439), .ZN(n8442) );
  AOI21_X1 U9891 ( .B1(n8649), .B2(n9948), .A(n8442), .ZN(n8443) );
  OAI211_X1 U9892 ( .C1(n8445), .C2(n8458), .A(n8444), .B(n8443), .ZN(P2_U3180) );
  AND2_X1 U9893 ( .A1(n8447), .A2(n8446), .ZN(n8450) );
  OAI211_X1 U9894 ( .C1(n8450), .C2(n8449), .A(n9958), .B(n8448), .ZN(n8457)
         );
  NAND2_X1 U9895 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9842) );
  INV_X1 U9896 ( .A(n9842), .ZN(n8451) );
  AOI21_X1 U9897 ( .B1(n9952), .B2(n8757), .A(n8451), .ZN(n8455) );
  NAND2_X1 U9898 ( .A1(n9948), .A2(n8452), .ZN(n8454) );
  NAND2_X1 U9899 ( .A1(n9945), .A2(n8464), .ZN(n8453) );
  AND3_X1 U9900 ( .A1(n8455), .A2(n8454), .A3(n8453), .ZN(n8456) );
  OAI211_X1 U9901 ( .C1(n8459), .C2(n8458), .A(n8457), .B(n8456), .ZN(P2_U3181) );
  MUX2_X1 U9902 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8607), .S(P2_U3893), .Z(
        P2_U3522) );
  INV_X1 U9903 ( .A(n8460), .ZN(n8624) );
  MUX2_X1 U9904 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8624), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9905 ( .A(n8461), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8474), .Z(
        P2_U3519) );
  MUX2_X1 U9906 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8646), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9907 ( .A(n8655), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8474), .Z(
        P2_U3517) );
  MUX2_X1 U9908 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8668), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9909 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8462), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9910 ( .A(n8691), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8474), .Z(
        P2_U3514) );
  MUX2_X1 U9911 ( .A(n8463), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8474), .Z(
        P2_U3513) );
  MUX2_X1 U9912 ( .A(n8718), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8474), .Z(
        P2_U3512) );
  MUX2_X1 U9913 ( .A(n8731), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8474), .Z(
        P2_U3511) );
  MUX2_X1 U9914 ( .A(n8748), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8474), .Z(
        P2_U3510) );
  MUX2_X1 U9915 ( .A(n8758), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8474), .Z(
        P2_U3509) );
  MUX2_X1 U9916 ( .A(n8772), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8474), .Z(
        P2_U3508) );
  MUX2_X1 U9917 ( .A(n8757), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8474), .Z(
        P2_U3507) );
  MUX2_X1 U9918 ( .A(n8464), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8474), .Z(
        P2_U3505) );
  MUX2_X1 U9919 ( .A(n8465), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8474), .Z(
        P2_U3504) );
  MUX2_X1 U9920 ( .A(n9951), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8474), .Z(
        P2_U3503) );
  MUX2_X1 U9921 ( .A(n4441), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8474), .Z(
        P2_U3502) );
  MUX2_X1 U9922 ( .A(n9944), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8474), .Z(
        P2_U3501) );
  MUX2_X1 U9923 ( .A(n8466), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8474), .Z(
        P2_U3500) );
  MUX2_X1 U9924 ( .A(n8467), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8474), .Z(
        P2_U3499) );
  MUX2_X1 U9925 ( .A(n8468), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8474), .Z(
        P2_U3498) );
  MUX2_X1 U9926 ( .A(n8469), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8474), .Z(
        P2_U3497) );
  MUX2_X1 U9927 ( .A(n8470), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8474), .Z(
        P2_U3496) );
  MUX2_X1 U9928 ( .A(n8471), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8474), .Z(
        P2_U3495) );
  MUX2_X1 U9929 ( .A(n8472), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8474), .Z(
        P2_U3494) );
  MUX2_X1 U9930 ( .A(n5132), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8474), .Z(
        P2_U3493) );
  MUX2_X1 U9931 ( .A(n8473), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8474), .Z(
        P2_U3492) );
  MUX2_X1 U9932 ( .A(n8475), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8474), .Z(
        P2_U3491) );
  OAI21_X1 U9933 ( .B1(n8478), .B2(n8477), .A(n8476), .ZN(n8482) );
  XNOR2_X1 U9934 ( .A(n8480), .B(n8479), .ZN(n8481) );
  AOI22_X1 U9935 ( .A1(n9805), .A2(n8482), .B1(n9856), .B2(n8481), .ZN(n8490)
         );
  AOI22_X1 U9936 ( .A1(n9846), .A2(n8483), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n8489) );
  OAI211_X1 U9937 ( .C1(n8486), .C2(n8485), .A(n9855), .B(n8484), .ZN(n8488)
         );
  NAND2_X1 U9938 ( .A1(n9845), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n8487) );
  NAND4_X1 U9939 ( .A1(n8490), .A2(n8489), .A3(n8488), .A4(n8487), .ZN(
        P2_U3184) );
  NAND2_X1 U9940 ( .A1(n8533), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8491) );
  NAND2_X1 U9941 ( .A1(n8492), .A2(n8491), .ZN(n8493) );
  XNOR2_X1 U9942 ( .A(n8493), .B(n8531), .ZN(n9729) );
  NOR2_X1 U9943 ( .A1(n9728), .A2(n9729), .ZN(n9727) );
  AOI21_X1 U9944 ( .B1(n8493), .B2(n8531), .A(n9727), .ZN(n9758) );
  MUX2_X1 U9945 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7204), .S(n9746), .Z(n9757)
         );
  NOR2_X1 U9946 ( .A1(n9758), .A2(n9757), .ZN(n9756) );
  INV_X1 U9947 ( .A(n8494), .ZN(n8495) );
  MUX2_X1 U9948 ( .A(n7355), .B(P2_REG2_REG_12__SCAN_IN), .S(n9778), .Z(n8496)
         );
  INV_X1 U9949 ( .A(n8496), .ZN(n9789) );
  NOR2_X1 U9950 ( .A1(n9795), .A2(n8497), .ZN(n8499) );
  XNOR2_X1 U9951 ( .A(n9795), .B(n8497), .ZN(n9803) );
  NOR2_X1 U9952 ( .A1(n8498), .A2(n9803), .ZN(n9807) );
  MUX2_X1 U9953 ( .A(n5322), .B(P2_REG2_REG_14__SCAN_IN), .S(n9812), .Z(n8500)
         );
  INV_X1 U9954 ( .A(n8500), .ZN(n9823) );
  NOR2_X1 U9955 ( .A1(n9824), .A2(n9823), .ZN(n9822) );
  NOR2_X1 U9956 ( .A1(n9830), .A2(n8501), .ZN(n8502) );
  MUX2_X1 U9957 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n8774), .S(n9847), .Z(n9859)
         );
  AOI21_X1 U9958 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8517), .A(n9858), .ZN(
        n8558) );
  XOR2_X1 U9959 ( .A(n8558), .B(n8576), .Z(n8503) );
  NOR2_X1 U9960 ( .A1(n8760), .A2(n8503), .ZN(n8559) );
  AOI21_X1 U9961 ( .B1(n8760), .B2(n8503), .A(n8559), .ZN(n8555) );
  AOI22_X1 U9962 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8517), .B1(n9847), .B2(
        n8828), .ZN(n9850) );
  AOI22_X1 U9963 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8521), .B1(n9812), .B2(
        n8513), .ZN(n9815) );
  INV_X1 U9964 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10029) );
  AOI22_X1 U9965 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8525), .B1(n9778), .B2(
        n10029), .ZN(n9781) );
  INV_X1 U9966 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8508) );
  AOI22_X1 U9967 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n8529), .B1(n9746), .B2(
        n8508), .ZN(n9749) );
  NAND2_X1 U9968 ( .A1(n8533), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8504) );
  NAND2_X1 U9969 ( .A1(n8505), .A2(n8504), .ZN(n8506) );
  NAND2_X1 U9970 ( .A1(n8506), .A2(n8531), .ZN(n8507) );
  XNOR2_X1 U9971 ( .A(n8506), .B(n9734), .ZN(n9731) );
  NAND2_X1 U9972 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n9731), .ZN(n9730) );
  NAND2_X1 U9973 ( .A1(n8507), .A2(n9730), .ZN(n9748) );
  NAND2_X1 U9974 ( .A1(n8509), .A2(n8527), .ZN(n8510) );
  XNOR2_X1 U9975 ( .A(n8509), .B(n9764), .ZN(n9766) );
  NAND2_X1 U9976 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n9766), .ZN(n9765) );
  NAND2_X1 U9977 ( .A1(n8510), .A2(n9765), .ZN(n9780) );
  NAND2_X1 U9978 ( .A1(n8523), .A2(n8511), .ZN(n8512) );
  XNOR2_X1 U9979 ( .A(n8511), .B(n9795), .ZN(n9797) );
  NAND2_X1 U9980 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n9797), .ZN(n9796) );
  NAND2_X1 U9981 ( .A1(n8512), .A2(n9796), .ZN(n9814) );
  NAND2_X1 U9982 ( .A1(n8519), .A2(n8514), .ZN(n8515) );
  XNOR2_X1 U9983 ( .A(n8514), .B(n9830), .ZN(n9832) );
  NAND2_X1 U9984 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n9832), .ZN(n9831) );
  NAND2_X1 U9985 ( .A1(n8515), .A2(n9831), .ZN(n9849) );
  NAND2_X1 U9986 ( .A1(n9850), .A2(n9849), .ZN(n9848) );
  OAI21_X1 U9987 ( .B1(n9847), .B2(n8828), .A(n9848), .ZN(n8575) );
  OAI21_X1 U9988 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8516), .A(n8577), .ZN(
        n8553) );
  INV_X1 U9989 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9974) );
  MUX2_X1 U9990 ( .A(n8760), .B(n8824), .S(n8588), .Z(n8565) );
  XNOR2_X1 U9991 ( .A(n8576), .B(n8565), .ZN(n8546) );
  MUX2_X1 U9992 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8588), .Z(n8518) );
  OR2_X1 U9993 ( .A1(n8517), .A2(n8518), .ZN(n8544) );
  XNOR2_X1 U9994 ( .A(n8518), .B(n9847), .ZN(n9853) );
  MUX2_X1 U9995 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8588), .Z(n8520) );
  OR2_X1 U9996 ( .A1(n8520), .A2(n8519), .ZN(n8543) );
  XNOR2_X1 U9997 ( .A(n8520), .B(n9830), .ZN(n9835) );
  MUX2_X1 U9998 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8588), .Z(n8522) );
  OR2_X1 U9999 ( .A1(n8522), .A2(n8521), .ZN(n8542) );
  XNOR2_X1 U10000 ( .A(n8522), .B(n9812), .ZN(n9818) );
  MUX2_X1 U10001 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8588), .Z(n8524) );
  OR2_X1 U10002 ( .A1(n8524), .A2(n8523), .ZN(n8541) );
  XNOR2_X1 U10003 ( .A(n8524), .B(n9795), .ZN(n9800) );
  MUX2_X1 U10004 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8588), .Z(n8526) );
  OR2_X1 U10005 ( .A1(n8526), .A2(n8525), .ZN(n8540) );
  XNOR2_X1 U10006 ( .A(n8526), .B(n9778), .ZN(n9784) );
  MUX2_X1 U10007 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8588), .Z(n8528) );
  OR2_X1 U10008 ( .A1(n8528), .A2(n8527), .ZN(n8539) );
  XNOR2_X1 U10009 ( .A(n8528), .B(n9764), .ZN(n9769) );
  MUX2_X1 U10010 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8588), .Z(n8530) );
  OR2_X1 U10011 ( .A1(n8530), .A2(n8529), .ZN(n8538) );
  XNOR2_X1 U10012 ( .A(n8530), .B(n9746), .ZN(n9752) );
  MUX2_X1 U10013 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8588), .Z(n8532) );
  OR2_X1 U10014 ( .A1(n8532), .A2(n8531), .ZN(n8537) );
  XNOR2_X1 U10015 ( .A(n8532), .B(n9734), .ZN(n9740) );
  OAI22_X1 U10016 ( .A1(n8536), .A2(n8535), .B1(n8534), .B2(n8533), .ZN(n9741)
         );
  NAND2_X1 U10017 ( .A1(n9740), .A2(n9741), .ZN(n9739) );
  NAND2_X1 U10018 ( .A1(n8537), .A2(n9739), .ZN(n9751) );
  NAND2_X1 U10019 ( .A1(n9752), .A2(n9751), .ZN(n9750) );
  NAND2_X1 U10020 ( .A1(n8538), .A2(n9750), .ZN(n9768) );
  NAND2_X1 U10021 ( .A1(n9769), .A2(n9768), .ZN(n9767) );
  NAND2_X1 U10022 ( .A1(n8539), .A2(n9767), .ZN(n9783) );
  NAND2_X1 U10023 ( .A1(n9784), .A2(n9783), .ZN(n9782) );
  NAND2_X1 U10024 ( .A1(n8540), .A2(n9782), .ZN(n9799) );
  NAND2_X1 U10025 ( .A1(n9800), .A2(n9799), .ZN(n9798) );
  NAND2_X1 U10026 ( .A1(n8541), .A2(n9798), .ZN(n9817) );
  NAND2_X1 U10027 ( .A1(n9818), .A2(n9817), .ZN(n9816) );
  NAND2_X1 U10028 ( .A1(n8542), .A2(n9816), .ZN(n9834) );
  NAND2_X1 U10029 ( .A1(n9835), .A2(n9834), .ZN(n9833) );
  NAND2_X1 U10030 ( .A1(n8543), .A2(n9833), .ZN(n9852) );
  NAND2_X1 U10031 ( .A1(n9853), .A2(n9852), .ZN(n9851) );
  NAND2_X1 U10032 ( .A1(n8544), .A2(n9851), .ZN(n8545) );
  NAND2_X1 U10033 ( .A1(n8546), .A2(n8545), .ZN(n8563) );
  OAI21_X1 U10034 ( .B1(n8546), .B2(n8545), .A(n8563), .ZN(n8550) );
  INV_X1 U10035 ( .A(n9846), .ZN(n8547) );
  NOR2_X1 U10036 ( .A1(n8547), .A2(n8576), .ZN(n8548) );
  AOI211_X1 U10037 ( .C1(n9855), .C2(n8550), .A(n8549), .B(n8548), .ZN(n8551)
         );
  OAI21_X1 U10038 ( .B1(n9745), .B2(n9974), .A(n8551), .ZN(n8552) );
  AOI21_X1 U10039 ( .B1(n8553), .B2(n9856), .A(n8552), .ZN(n8554) );
  OAI21_X1 U10040 ( .B1(n8555), .B2(n9860), .A(n8554), .ZN(P2_U3199) );
  INV_X1 U10041 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8557) );
  NOR2_X1 U10042 ( .A1(n8596), .A2(n8557), .ZN(n8556) );
  AOI21_X1 U10043 ( .B1(n8557), .B2(n8596), .A(n8556), .ZN(n8562) );
  NOR2_X1 U10044 ( .A1(n8566), .A2(n8558), .ZN(n8560) );
  NOR2_X2 U10045 ( .A1(n8560), .A2(n8559), .ZN(n8561) );
  AOI21_X1 U10046 ( .B1(n8562), .B2(n8561), .A(n8584), .ZN(n8583) );
  INV_X1 U10047 ( .A(n8563), .ZN(n8564) );
  AOI21_X1 U10048 ( .B1(n8566), .B2(n8565), .A(n8564), .ZN(n8568) );
  MUX2_X1 U10049 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8588), .Z(n8567) );
  NOR2_X1 U10050 ( .A1(n8568), .A2(n8567), .ZN(n8587) );
  NAND2_X1 U10051 ( .A1(n8568), .A2(n8567), .ZN(n8585) );
  INV_X1 U10052 ( .A(n8585), .ZN(n8569) );
  NOR2_X1 U10053 ( .A1(n8587), .A2(n8569), .ZN(n8570) );
  AOI21_X1 U10054 ( .B1(P2_U3893), .B2(n8570), .A(n9846), .ZN(n8574) );
  INV_X1 U10055 ( .A(n8570), .ZN(n8571) );
  NAND3_X1 U10056 ( .A1(n9855), .A2(n8596), .A3(n8571), .ZN(n8572) );
  OAI211_X1 U10057 ( .C1(n8574), .C2(n8596), .A(n8573), .B(n8572), .ZN(n8581)
         );
  XNOR2_X1 U10058 ( .A(n8586), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U10059 ( .A1(n8576), .A2(n8575), .ZN(n8578) );
  NAND2_X1 U10060 ( .A1(n8578), .A2(n8577), .ZN(n8598) );
  XOR2_X1 U10061 ( .A(n8597), .B(n8598), .Z(n8579) );
  NOR2_X1 U10062 ( .A1(n8579), .A2(n9664), .ZN(n8580) );
  AOI211_X1 U10063 ( .C1(n9845), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8581), .B(
        n8580), .ZN(n8582) );
  OAI21_X1 U10064 ( .B1(n8583), .B2(n9860), .A(n8582), .ZN(P2_U3200) );
  MUX2_X1 U10065 ( .A(n8734), .B(P2_REG2_REG_19__SCAN_IN), .S(n8592), .Z(n8589) );
  OAI21_X1 U10066 ( .B1(n8587), .B2(n8586), .A(n8585), .ZN(n8591) );
  XNOR2_X1 U10067 ( .A(n8592), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8599) );
  MUX2_X1 U10068 ( .A(n8589), .B(n8599), .S(n8588), .Z(n8590) );
  XNOR2_X1 U10069 ( .A(n8591), .B(n8590), .ZN(n8595) );
  NAND2_X1 U10070 ( .A1(n9846), .A2(n8592), .ZN(n8593) );
  OAI211_X1 U10071 ( .C1(n9673), .C2(n8595), .A(n8594), .B(n8593), .ZN(n8603)
         );
  AOI22_X1 U10072 ( .A1(n8598), .A2(n8597), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8596), .ZN(n8600) );
  XNOR2_X1 U10073 ( .A(n8600), .B(n8599), .ZN(n8601) );
  NOR2_X1 U10074 ( .A1(n8601), .A2(n9664), .ZN(n8602) );
  INV_X1 U10075 ( .A(n8605), .ZN(n8606) );
  NAND2_X1 U10076 ( .A1(n8607), .A2(n8606), .ZN(n8859) );
  NAND2_X1 U10077 ( .A1(n8608), .A2(n8777), .ZN(n8616) );
  OAI21_X1 U10078 ( .B1(n9876), .B2(n8859), .A(n8616), .ZN(n8611) );
  AOI21_X1 U10079 ( .B1(n9876), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8611), .ZN(
        n8609) );
  OAI21_X1 U10080 ( .B1(n8610), .B2(n8613), .A(n8609), .ZN(P2_U3202) );
  AOI21_X1 U10081 ( .B1(n9876), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8611), .ZN(
        n8612) );
  OAI21_X1 U10082 ( .B1(n8786), .B2(n8613), .A(n8612), .ZN(P2_U3203) );
  INV_X1 U10083 ( .A(n8614), .ZN(n8622) );
  NAND2_X1 U10084 ( .A1(n8615), .A2(n8693), .ZN(n8621) );
  OAI21_X1 U10085 ( .B1(n8693), .B2(n8617), .A(n8616), .ZN(n8618) );
  AOI21_X1 U10086 ( .B1(n8619), .B2(n8778), .A(n8618), .ZN(n8620) );
  OAI211_X1 U10087 ( .C1(n8622), .C2(n8765), .A(n8621), .B(n8620), .ZN(
        P2_U3204) );
  XNOR2_X1 U10088 ( .A(n8623), .B(n4356), .ZN(n8870) );
  AOI222_X1 U10089 ( .A1(n8842), .A2(n8625), .B1(n8646), .B2(n8769), .C1(n8624), .C2(n8771), .ZN(n8865) );
  MUX2_X1 U10090 ( .A(n8626), .B(n8865), .S(n8693), .Z(n8629) );
  AOI22_X1 U10091 ( .A1(n8867), .A2(n8778), .B1(n8777), .B2(n8627), .ZN(n8628)
         );
  OAI211_X1 U10092 ( .C1(n8870), .C2(n8765), .A(n8629), .B(n8628), .ZN(
        P2_U3205) );
  XNOR2_X1 U10093 ( .A(n8631), .B(n8630), .ZN(n8874) );
  XNOR2_X1 U10094 ( .A(n8633), .B(n8632), .ZN(n8634) );
  OAI222_X1 U10095 ( .A1(n8840), .A2(n8636), .B1(n8838), .B2(n8635), .C1(n8634), .C2(n8679), .ZN(n8790) );
  NAND2_X1 U10096 ( .A1(n8790), .A2(n8693), .ZN(n8642) );
  NAND2_X1 U10097 ( .A1(n8637), .A2(n8777), .ZN(n8638) );
  OAI21_X1 U10098 ( .B1(n8693), .B2(n8639), .A(n8638), .ZN(n8640) );
  AOI21_X1 U10099 ( .B1(n8791), .B2(n8778), .A(n8640), .ZN(n8641) );
  OAI211_X1 U10100 ( .C1(n8874), .C2(n8765), .A(n8642), .B(n8641), .ZN(
        P2_U3206) );
  XNOR2_X1 U10101 ( .A(n8643), .B(n8644), .ZN(n8880) );
  XNOR2_X1 U10102 ( .A(n8645), .B(n8644), .ZN(n8647) );
  AOI222_X1 U10103 ( .A1(n8842), .A2(n8647), .B1(n8668), .B2(n8769), .C1(n8646), .C2(n8771), .ZN(n8875) );
  MUX2_X1 U10104 ( .A(n8648), .B(n8875), .S(n8693), .Z(n8651) );
  AOI22_X1 U10105 ( .A1(n8877), .A2(n8778), .B1(n8777), .B2(n8649), .ZN(n8650)
         );
  OAI211_X1 U10106 ( .C1(n8880), .C2(n8765), .A(n8651), .B(n8650), .ZN(
        P2_U3207) );
  XNOR2_X1 U10107 ( .A(n8652), .B(n8653), .ZN(n8886) );
  XNOR2_X1 U10108 ( .A(n8654), .B(n8653), .ZN(n8658) );
  NAND2_X1 U10109 ( .A1(n8655), .A2(n8771), .ZN(n8656) );
  OAI21_X1 U10110 ( .B1(n8680), .B2(n8840), .A(n8656), .ZN(n8657) );
  AOI21_X1 U10111 ( .B1(n8658), .B2(n8842), .A(n8657), .ZN(n8881) );
  MUX2_X1 U10112 ( .A(n8659), .B(n8881), .S(n8693), .Z(n8662) );
  AOI22_X1 U10113 ( .A1(n8883), .A2(n8672), .B1(n8777), .B2(n8660), .ZN(n8661)
         );
  OAI211_X1 U10114 ( .C1(n8886), .C2(n8765), .A(n8662), .B(n8661), .ZN(
        P2_U3208) );
  NAND2_X1 U10115 ( .A1(n8664), .A2(n8663), .ZN(n8665) );
  XOR2_X1 U10116 ( .A(n8666), .B(n8665), .Z(n8892) );
  XOR2_X1 U10117 ( .A(n8667), .B(n8666), .Z(n8669) );
  AOI222_X1 U10118 ( .A1(n8842), .A2(n8669), .B1(n8668), .B2(n8771), .C1(n8691), .C2(n8769), .ZN(n8887) );
  MUX2_X1 U10119 ( .A(n8670), .B(n8887), .S(n8693), .Z(n8674) );
  AOI22_X1 U10120 ( .A1(n8889), .A2(n8672), .B1(n8777), .B2(n8671), .ZN(n8673)
         );
  OAI211_X1 U10121 ( .C1(n8892), .C2(n8765), .A(n8674), .B(n8673), .ZN(
        P2_U3209) );
  XOR2_X1 U10122 ( .A(n8675), .B(n8676), .Z(n8896) );
  XNOR2_X1 U10123 ( .A(n8677), .B(n8676), .ZN(n8678) );
  OAI222_X1 U10124 ( .A1(n8840), .A2(n8700), .B1(n8838), .B2(n8680), .C1(n8679), .C2(n8678), .ZN(n8803) );
  NAND2_X1 U10125 ( .A1(n8803), .A2(n8693), .ZN(n8686) );
  INV_X1 U10126 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8683) );
  INV_X1 U10127 ( .A(n8681), .ZN(n8682) );
  OAI22_X1 U10128 ( .A1(n8693), .A2(n8683), .B1(n8682), .B2(n9869), .ZN(n8684)
         );
  AOI21_X1 U10129 ( .B1(n8804), .B2(n8778), .A(n8684), .ZN(n8685) );
  OAI211_X1 U10130 ( .C1(n8896), .C2(n8765), .A(n8686), .B(n8685), .ZN(
        P2_U3210) );
  XNOR2_X1 U10131 ( .A(n8687), .B(n8688), .ZN(n8902) );
  INV_X1 U10132 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8694) );
  XNOR2_X1 U10133 ( .A(n8690), .B(n8689), .ZN(n8692) );
  AOI222_X1 U10134 ( .A1(n8842), .A2(n8692), .B1(n8718), .B2(n8769), .C1(n8691), .C2(n8771), .ZN(n8897) );
  MUX2_X1 U10135 ( .A(n8694), .B(n8897), .S(n8693), .Z(n8697) );
  AOI22_X1 U10136 ( .A1(n8899), .A2(n8778), .B1(n8777), .B2(n8695), .ZN(n8696)
         );
  OAI211_X1 U10137 ( .C1(n8902), .C2(n8765), .A(n8697), .B(n8696), .ZN(
        P2_U3211) );
  XNOR2_X1 U10138 ( .A(n8698), .B(n8709), .ZN(n8702) );
  OAI22_X1 U10139 ( .A1(n8700), .A2(n8838), .B1(n8699), .B2(n8840), .ZN(n8701)
         );
  AOI21_X1 U10140 ( .B1(n8702), .B2(n8842), .A(n8701), .ZN(n8812) );
  INV_X1 U10141 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8705) );
  INV_X1 U10142 ( .A(n8703), .ZN(n8704) );
  OAI22_X1 U10143 ( .A1(n8693), .A2(n8705), .B1(n8704), .B2(n9869), .ZN(n8706)
         );
  AOI21_X1 U10144 ( .B1(n8810), .B2(n8778), .A(n8706), .ZN(n8712) );
  NAND2_X1 U10145 ( .A1(n8708), .A2(n8707), .ZN(n8710) );
  XNOR2_X1 U10146 ( .A(n8710), .B(n8709), .ZN(n8906) );
  OR2_X1 U10147 ( .A1(n8906), .A2(n8765), .ZN(n8711) );
  OAI211_X1 U10148 ( .C1(n8812), .C2(n9876), .A(n8712), .B(n8711), .ZN(
        P2_U3212) );
  XNOR2_X1 U10149 ( .A(n8713), .B(n8716), .ZN(n8912) );
  INV_X1 U10150 ( .A(n8714), .ZN(n8720) );
  OAI21_X1 U10151 ( .B1(n8717), .B2(n8716), .A(n8715), .ZN(n8719) );
  AOI222_X1 U10152 ( .A1(n8842), .A2(n8719), .B1(n8718), .B2(n8771), .C1(n8748), .C2(n8769), .ZN(n8907) );
  OAI21_X1 U10153 ( .B1(n8720), .B2(n9869), .A(n8907), .ZN(n8721) );
  NAND2_X1 U10154 ( .A1(n8721), .A2(n8693), .ZN(n8723) );
  AOI22_X1 U10155 ( .A1(n8909), .A2(n8778), .B1(P2_REG2_REG_20__SCAN_IN), .B2(
        n9876), .ZN(n8722) );
  OAI211_X1 U10156 ( .C1(n8912), .C2(n8765), .A(n8723), .B(n8722), .ZN(
        P2_U3213) );
  NAND2_X1 U10157 ( .A1(n8725), .A2(n8724), .ZN(n8726) );
  XNOR2_X1 U10158 ( .A(n8726), .B(n8727), .ZN(n8916) );
  NAND2_X1 U10159 ( .A1(n8728), .A2(n8727), .ZN(n8729) );
  NAND3_X1 U10160 ( .A1(n8730), .A2(n8842), .A3(n8729), .ZN(n8733) );
  AOI22_X1 U10161 ( .A1(n8731), .A2(n8771), .B1(n8769), .B2(n8758), .ZN(n8732)
         );
  NAND2_X1 U10162 ( .A1(n8733), .A2(n8732), .ZN(n8913) );
  INV_X1 U10163 ( .A(n8913), .ZN(n8735) );
  MUX2_X1 U10164 ( .A(n8735), .B(n8734), .S(n9876), .Z(n8740) );
  INV_X1 U10165 ( .A(n8736), .ZN(n8737) );
  AOI22_X1 U10166 ( .A1(n8738), .A2(n8778), .B1(n8777), .B2(n8737), .ZN(n8739)
         );
  OAI211_X1 U10167 ( .C1(n8916), .C2(n8765), .A(n8740), .B(n8739), .ZN(
        P2_U3214) );
  XNOR2_X1 U10168 ( .A(n4350), .B(n8746), .ZN(n8924) );
  NAND2_X1 U10169 ( .A1(n8742), .A2(n8741), .ZN(n8756) );
  NAND2_X1 U10170 ( .A1(n8756), .A2(n8743), .ZN(n8745) );
  NAND2_X1 U10171 ( .A1(n8745), .A2(n8744), .ZN(n8747) );
  XNOR2_X1 U10172 ( .A(n8747), .B(n8746), .ZN(n8749) );
  AOI222_X1 U10173 ( .A1(n8842), .A2(n8749), .B1(n8772), .B2(n8769), .C1(n8748), .C2(n8771), .ZN(n8919) );
  MUX2_X1 U10174 ( .A(n8557), .B(n8919), .S(n8693), .Z(n8753) );
  INV_X1 U10175 ( .A(n8750), .ZN(n8751) );
  AOI22_X1 U10176 ( .A1(n8921), .A2(n8778), .B1(n8777), .B2(n8751), .ZN(n8752)
         );
  OAI211_X1 U10177 ( .C1(n8924), .C2(n8765), .A(n8753), .B(n8752), .ZN(
        P2_U3215) );
  XNOR2_X1 U10178 ( .A(n8754), .B(n8755), .ZN(n8930) );
  XNOR2_X1 U10179 ( .A(n8756), .B(n8755), .ZN(n8759) );
  AOI222_X1 U10180 ( .A1(n8842), .A2(n8759), .B1(n8758), .B2(n8771), .C1(n8757), .C2(n8769), .ZN(n8925) );
  MUX2_X1 U10181 ( .A(n8760), .B(n8925), .S(n8693), .Z(n8764) );
  INV_X1 U10182 ( .A(n8761), .ZN(n8762) );
  AOI22_X1 U10183 ( .A1(n8927), .A2(n8778), .B1(n8777), .B2(n8762), .ZN(n8763)
         );
  OAI211_X1 U10184 ( .C1(n8930), .C2(n8765), .A(n8764), .B(n8763), .ZN(
        P2_U3216) );
  XNOR2_X1 U10185 ( .A(n8766), .B(n8767), .ZN(n8938) );
  XOR2_X1 U10186 ( .A(n8768), .B(n8767), .Z(n8773) );
  AOI222_X1 U10187 ( .A1(n8842), .A2(n8773), .B1(n8772), .B2(n8771), .C1(n8770), .C2(n8769), .ZN(n8931) );
  MUX2_X1 U10188 ( .A(n8774), .B(n8931), .S(n8693), .Z(n8780) );
  INV_X1 U10189 ( .A(n8775), .ZN(n8776) );
  AOI22_X1 U10190 ( .A1(n8934), .A2(n8778), .B1(n8777), .B2(n8776), .ZN(n8779)
         );
  OAI211_X1 U10191 ( .C1(n8938), .C2(n8765), .A(n8780), .B(n8779), .ZN(
        P2_U3217) );
  INV_X1 U10192 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8783) );
  NAND2_X1 U10193 ( .A1(n7672), .A2(n8829), .ZN(n8782) );
  INV_X1 U10194 ( .A(n8859), .ZN(n8781) );
  NAND2_X1 U10195 ( .A1(n8781), .A2(n8827), .ZN(n8784) );
  OAI211_X1 U10196 ( .C1(n8827), .C2(n8783), .A(n8782), .B(n8784), .ZN(
        P2_U3490) );
  NAND2_X1 U10197 ( .A1(n8857), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8785) );
  OAI211_X1 U10198 ( .C1(n8786), .C2(n8818), .A(n8785), .B(n8784), .ZN(
        P2_U3489) );
  INV_X1 U10199 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8787) );
  MUX2_X1 U10200 ( .A(n8787), .B(n8865), .S(n8827), .Z(n8789) );
  NAND2_X1 U10201 ( .A1(n8867), .A2(n8829), .ZN(n8788) );
  OAI211_X1 U10202 ( .C1(n8870), .C2(n8832), .A(n8789), .B(n8788), .ZN(
        P2_U3487) );
  INV_X1 U10203 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8792) );
  AOI21_X1 U10204 ( .B1(n8852), .B2(n8791), .A(n8790), .ZN(n8871) );
  MUX2_X1 U10205 ( .A(n8792), .B(n8871), .S(n8827), .Z(n8793) );
  OAI21_X1 U10206 ( .B1(n8874), .B2(n8832), .A(n8793), .ZN(P2_U3486) );
  INV_X1 U10207 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8794) );
  MUX2_X1 U10208 ( .A(n8794), .B(n8875), .S(n8827), .Z(n8796) );
  NAND2_X1 U10209 ( .A1(n8877), .A2(n8829), .ZN(n8795) );
  OAI211_X1 U10210 ( .C1(n8832), .C2(n8880), .A(n8796), .B(n8795), .ZN(
        P2_U3485) );
  INV_X1 U10211 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8797) );
  MUX2_X1 U10212 ( .A(n8797), .B(n8881), .S(n8827), .Z(n8799) );
  NAND2_X1 U10213 ( .A1(n8883), .A2(n8829), .ZN(n8798) );
  OAI211_X1 U10214 ( .C1(n8886), .C2(n8832), .A(n8799), .B(n8798), .ZN(
        P2_U3484) );
  INV_X1 U10215 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8800) );
  MUX2_X1 U10216 ( .A(n8800), .B(n8887), .S(n8827), .Z(n8802) );
  NAND2_X1 U10217 ( .A1(n8889), .A2(n8829), .ZN(n8801) );
  OAI211_X1 U10218 ( .C1(n8832), .C2(n8892), .A(n8802), .B(n8801), .ZN(
        P2_U3483) );
  INV_X1 U10219 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8805) );
  AOI21_X1 U10220 ( .B1(n8852), .B2(n8804), .A(n8803), .ZN(n8893) );
  MUX2_X1 U10221 ( .A(n8805), .B(n8893), .S(n8827), .Z(n8806) );
  OAI21_X1 U10222 ( .B1(n8832), .B2(n8896), .A(n8806), .ZN(P2_U3482) );
  INV_X1 U10223 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8807) );
  MUX2_X1 U10224 ( .A(n8807), .B(n8897), .S(n8827), .Z(n8809) );
  NAND2_X1 U10225 ( .A1(n8899), .A2(n8829), .ZN(n8808) );
  OAI211_X1 U10226 ( .C1(n8902), .C2(n8832), .A(n8809), .B(n8808), .ZN(
        P2_U3481) );
  INV_X1 U10227 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8813) );
  NAND2_X1 U10228 ( .A1(n8810), .A2(n8852), .ZN(n8811) );
  AND2_X1 U10229 ( .A1(n8812), .A2(n8811), .ZN(n8903) );
  MUX2_X1 U10230 ( .A(n8813), .B(n8903), .S(n8827), .Z(n8814) );
  OAI21_X1 U10231 ( .B1(n8832), .B2(n8906), .A(n8814), .ZN(P2_U3480) );
  MUX2_X1 U10232 ( .A(n8815), .B(n8907), .S(n8827), .Z(n8817) );
  NAND2_X1 U10233 ( .A1(n8909), .A2(n8829), .ZN(n8816) );
  OAI211_X1 U10234 ( .C1(n8832), .C2(n8912), .A(n8817), .B(n8816), .ZN(
        P2_U3479) );
  MUX2_X1 U10235 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8913), .S(n8827), .Z(n8820) );
  OAI22_X1 U10236 ( .A1(n8916), .A2(n8832), .B1(n8915), .B2(n8818), .ZN(n8819)
         );
  OR2_X1 U10237 ( .A1(n8820), .A2(n8819), .ZN(P2_U3478) );
  INV_X1 U10238 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8821) );
  MUX2_X1 U10239 ( .A(n8821), .B(n8919), .S(n8827), .Z(n8823) );
  NAND2_X1 U10240 ( .A1(n8921), .A2(n8829), .ZN(n8822) );
  OAI211_X1 U10241 ( .C1(n8832), .C2(n8924), .A(n8823), .B(n8822), .ZN(
        P2_U3477) );
  MUX2_X1 U10242 ( .A(n8824), .B(n8925), .S(n8827), .Z(n8826) );
  NAND2_X1 U10243 ( .A1(n8927), .A2(n8829), .ZN(n8825) );
  OAI211_X1 U10244 ( .C1(n8930), .C2(n8832), .A(n8826), .B(n8825), .ZN(
        P2_U3476) );
  MUX2_X1 U10245 ( .A(n8828), .B(n8931), .S(n8827), .Z(n8831) );
  NAND2_X1 U10246 ( .A1(n8934), .A2(n8829), .ZN(n8830) );
  OAI211_X1 U10247 ( .C1(n8832), .C2(n8938), .A(n8831), .B(n8830), .ZN(
        P2_U3475) );
  XNOR2_X1 U10248 ( .A(n8834), .B(n8833), .ZN(n9873) );
  NAND2_X1 U10249 ( .A1(n9873), .A2(n8835), .ZN(n8845) );
  XNOR2_X1 U10250 ( .A(n8837), .B(n8836), .ZN(n8843) );
  OAI22_X1 U10251 ( .A1(n5118), .A2(n8840), .B1(n8839), .B2(n8838), .ZN(n8841)
         );
  AOI21_X1 U10252 ( .B1(n8843), .B2(n8842), .A(n8841), .ZN(n8844) );
  AND2_X1 U10253 ( .A1(n8845), .A2(n8844), .ZN(n9870) );
  INV_X1 U10254 ( .A(n8846), .ZN(n8853) );
  NOR2_X1 U10255 ( .A1(n9867), .A2(n8847), .ZN(n8848) );
  AOI21_X1 U10256 ( .B1(n9873), .B2(n8853), .A(n8848), .ZN(n8849) );
  AND2_X1 U10257 ( .A1(n9870), .A2(n8849), .ZN(n9881) );
  INV_X1 U10258 ( .A(n9881), .ZN(n8850) );
  MUX2_X1 U10259 ( .A(n8850), .B(P2_REG1_REG_2__SCAN_IN), .S(n8857), .Z(
        P2_U3461) );
  AOI22_X1 U10260 ( .A1(n8854), .A2(n8853), .B1(n8852), .B2(n8851), .ZN(n8855)
         );
  AND2_X1 U10261 ( .A1(n8856), .A2(n8855), .ZN(n9879) );
  INV_X1 U10262 ( .A(n9879), .ZN(n8858) );
  MUX2_X1 U10263 ( .A(n8858), .B(P2_REG1_REG_1__SCAN_IN), .S(n8857), .Z(
        P2_U3460) );
  NAND2_X1 U10264 ( .A1(n7672), .A2(n8933), .ZN(n8860) );
  OR2_X1 U10265 ( .A1(n8859), .A2(n9898), .ZN(n8862) );
  OAI211_X1 U10266 ( .C1(n7623), .C2(n9901), .A(n8860), .B(n8862), .ZN(
        P2_U3458) );
  INV_X1 U10267 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8864) );
  NAND2_X1 U10268 ( .A1(n8861), .A2(n8933), .ZN(n8863) );
  OAI211_X1 U10269 ( .C1(n8864), .C2(n9901), .A(n8863), .B(n8862), .ZN(
        P2_U3457) );
  INV_X1 U10270 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8866) );
  MUX2_X1 U10271 ( .A(n8866), .B(n8865), .S(n9901), .Z(n8869) );
  NAND2_X1 U10272 ( .A1(n8867), .A2(n8933), .ZN(n8868) );
  OAI211_X1 U10273 ( .C1(n8870), .C2(n8937), .A(n8869), .B(n8868), .ZN(
        P2_U3455) );
  INV_X1 U10274 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8872) );
  MUX2_X1 U10275 ( .A(n8872), .B(n8871), .S(n9901), .Z(n8873) );
  OAI21_X1 U10276 ( .B1(n8874), .B2(n8937), .A(n8873), .ZN(P2_U3454) );
  INV_X1 U10277 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8876) );
  MUX2_X1 U10278 ( .A(n8876), .B(n8875), .S(n9901), .Z(n8879) );
  NAND2_X1 U10279 ( .A1(n8877), .A2(n8933), .ZN(n8878) );
  OAI211_X1 U10280 ( .C1(n8880), .C2(n8937), .A(n8879), .B(n8878), .ZN(
        P2_U3453) );
  INV_X1 U10281 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8882) );
  MUX2_X1 U10282 ( .A(n8882), .B(n8881), .S(n9901), .Z(n8885) );
  NAND2_X1 U10283 ( .A1(n8883), .A2(n8933), .ZN(n8884) );
  OAI211_X1 U10284 ( .C1(n8886), .C2(n8937), .A(n8885), .B(n8884), .ZN(
        P2_U3452) );
  INV_X1 U10285 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8888) );
  MUX2_X1 U10286 ( .A(n8888), .B(n8887), .S(n9901), .Z(n8891) );
  NAND2_X1 U10287 ( .A1(n8889), .A2(n8933), .ZN(n8890) );
  OAI211_X1 U10288 ( .C1(n8892), .C2(n8937), .A(n8891), .B(n8890), .ZN(
        P2_U3451) );
  MUX2_X1 U10289 ( .A(n8894), .B(n8893), .S(n9901), .Z(n8895) );
  OAI21_X1 U10290 ( .B1(n8896), .B2(n8937), .A(n8895), .ZN(P2_U3450) );
  INV_X1 U10291 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8898) );
  MUX2_X1 U10292 ( .A(n8898), .B(n8897), .S(n9901), .Z(n8901) );
  NAND2_X1 U10293 ( .A1(n8899), .A2(n8933), .ZN(n8900) );
  OAI211_X1 U10294 ( .C1(n8902), .C2(n8937), .A(n8901), .B(n8900), .ZN(
        P2_U3449) );
  INV_X1 U10295 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8904) );
  MUX2_X1 U10296 ( .A(n8904), .B(n8903), .S(n9901), .Z(n8905) );
  OAI21_X1 U10297 ( .B1(n8906), .B2(n8937), .A(n8905), .ZN(P2_U3448) );
  MUX2_X1 U10298 ( .A(n8908), .B(n8907), .S(n9901), .Z(n8911) );
  NAND2_X1 U10299 ( .A1(n8909), .A2(n8933), .ZN(n8910) );
  OAI211_X1 U10300 ( .C1(n8912), .C2(n8937), .A(n8911), .B(n8910), .ZN(
        P2_U3447) );
  MUX2_X1 U10301 ( .A(n8913), .B(P2_REG0_REG_19__SCAN_IN), .S(n9898), .Z(n8918) );
  OAI22_X1 U10302 ( .A1(n8916), .A2(n8937), .B1(n8915), .B2(n8914), .ZN(n8917)
         );
  OR2_X1 U10303 ( .A1(n8918), .A2(n8917), .ZN(P2_U3446) );
  INV_X1 U10304 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8920) );
  MUX2_X1 U10305 ( .A(n8920), .B(n8919), .S(n9901), .Z(n8923) );
  NAND2_X1 U10306 ( .A1(n8921), .A2(n8933), .ZN(n8922) );
  OAI211_X1 U10307 ( .C1(n8924), .C2(n8937), .A(n8923), .B(n8922), .ZN(
        P2_U3444) );
  INV_X1 U10308 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8926) );
  MUX2_X1 U10309 ( .A(n8926), .B(n8925), .S(n9901), .Z(n8929) );
  NAND2_X1 U10310 ( .A1(n8927), .A2(n8933), .ZN(n8928) );
  OAI211_X1 U10311 ( .C1(n8930), .C2(n8937), .A(n8929), .B(n8928), .ZN(
        P2_U3441) );
  INV_X1 U10312 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8932) );
  MUX2_X1 U10313 ( .A(n8932), .B(n8931), .S(n9901), .Z(n8936) );
  NAND2_X1 U10314 ( .A1(n8934), .A2(n8933), .ZN(n8935) );
  OAI211_X1 U10315 ( .C1(n8938), .C2(n8937), .A(n8936), .B(n8935), .ZN(
        P2_U3438) );
  INV_X1 U10316 ( .A(n7894), .ZN(n9489) );
  NOR4_X1 U10317 ( .A1(n8939), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n8940), .ZN(n8941) );
  AOI21_X1 U10318 ( .B1(n8942), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8941), .ZN(
        n8943) );
  OAI21_X1 U10319 ( .B1(n9489), .B2(n8947), .A(n8943), .ZN(P2_U3264) );
  INV_X1 U10320 ( .A(n8944), .ZN(n9492) );
  OAI222_X1 U10321 ( .A1(P2_U3151), .A2(n8948), .B1(n8947), .B2(n9492), .C1(
        n8946), .C2(n8945), .ZN(P2_U3266) );
  MUX2_X1 U10322 ( .A(n8949), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  OAI21_X1 U10323 ( .B1(n8952), .B2(n8951), .A(n8950), .ZN(n8953) );
  NAND2_X1 U10324 ( .A1(n8953), .A2(n9056), .ZN(n8959) );
  NAND2_X1 U10325 ( .A1(n9076), .A2(n9096), .ZN(n8954) );
  NAND2_X1 U10326 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9563) );
  OAI211_X1 U10327 ( .C1(n8955), .C2(n9078), .A(n8954), .B(n9563), .ZN(n8956)
         );
  AOI21_X1 U10328 ( .B1(n8957), .B2(n9084), .A(n8956), .ZN(n8958) );
  OAI211_X1 U10329 ( .C1(n8960), .C2(n9080), .A(n8959), .B(n8958), .ZN(
        P1_U3215) );
  AOI21_X1 U10330 ( .B1(n8962), .B2(n8964), .A(n8961), .ZN(n8963) );
  AOI21_X1 U10331 ( .B1(n4374), .B2(n8964), .A(n8963), .ZN(n8969) );
  INV_X1 U10332 ( .A(n9084), .ZN(n9058) );
  NOR2_X1 U10333 ( .A1(n9257), .A2(n9058), .ZN(n8967) );
  AOI22_X1 U10334 ( .A1(n9076), .A2(n9223), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n8965) );
  OAI21_X1 U10335 ( .B1(n9283), .B2(n9078), .A(n8965), .ZN(n8966) );
  OAI21_X1 U10336 ( .B1(n8969), .B2(n4495), .A(n8968), .ZN(P1_U3216) );
  NAND2_X1 U10337 ( .A1(n9093), .A2(n9076), .ZN(n8971) );
  NAND2_X1 U10338 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9162) );
  OAI211_X1 U10339 ( .C1(n9350), .C2(n9078), .A(n8971), .B(n9162), .ZN(n8973)
         );
  NOR2_X1 U10340 ( .A1(n9317), .A2(n9080), .ZN(n8972) );
  AOI211_X1 U10341 ( .C1(n9318), .C2(n9084), .A(n8973), .B(n8972), .ZN(n8974)
         );
  OAI21_X1 U10342 ( .B1(n8975), .B2(n4495), .A(n8974), .ZN(P1_U3219) );
  OR2_X1 U10343 ( .A1(n8976), .A2(n8977), .ZN(n8979) );
  NAND2_X1 U10344 ( .A1(n8979), .A2(n8978), .ZN(n8980) );
  XOR2_X1 U10345 ( .A(n8981), .B(n8980), .Z(n8986) );
  AOI22_X1 U10346 ( .A1(n9092), .A2(n9076), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n8983) );
  NAND2_X1 U10347 ( .A1(n9084), .A2(n9289), .ZN(n8982) );
  OAI211_X1 U10348 ( .C1(n9313), .C2(n9078), .A(n8983), .B(n8982), .ZN(n8984)
         );
  AOI21_X1 U10349 ( .B1(n9464), .B2(n9035), .A(n8984), .ZN(n8985) );
  OAI21_X1 U10350 ( .B1(n8986), .B2(n4495), .A(n8985), .ZN(P1_U3223) );
  XOR2_X1 U10351 ( .A(n8988), .B(n8987), .Z(n8993) );
  AOI22_X1 U10352 ( .A1(n9076), .A2(n9090), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n8990) );
  NAND2_X1 U10353 ( .A1(n9084), .A2(n9229), .ZN(n8989) );
  OAI211_X1 U10354 ( .C1(n9251), .C2(n9078), .A(n8990), .B(n8989), .ZN(n8991)
         );
  AOI21_X1 U10355 ( .B1(n9449), .B2(n9035), .A(n8991), .ZN(n8992) );
  OAI21_X1 U10356 ( .B1(n8993), .B2(n4495), .A(n8992), .ZN(P1_U3225) );
  INV_X1 U10357 ( .A(n8995), .ZN(n8996) );
  XOR2_X1 U10358 ( .A(n8994), .B(n8995), .Z(n9075) );
  NOR2_X1 U10359 ( .A1(n9075), .A2(n9074), .ZN(n9073) );
  AOI21_X1 U10360 ( .B1(n8996), .B2(n8994), .A(n9073), .ZN(n9000) );
  XNOR2_X1 U10361 ( .A(n8998), .B(n8997), .ZN(n8999) );
  XNOR2_X1 U10362 ( .A(n9000), .B(n8999), .ZN(n9007) );
  AND2_X1 U10363 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9585) );
  NOR2_X1 U10364 ( .A1(n9078), .A2(n9001), .ZN(n9002) );
  AOI211_X1 U10365 ( .C1(n9076), .C2(n9336), .A(n9585), .B(n9002), .ZN(n9003)
         );
  OAI21_X1 U10366 ( .B1(n9058), .B2(n9004), .A(n9003), .ZN(n9005) );
  AOI21_X1 U10367 ( .B1(n9429), .B2(n9035), .A(n9005), .ZN(n9006) );
  OAI21_X1 U10368 ( .B1(n9007), .B2(n4495), .A(n9006), .ZN(P1_U3226) );
  OR2_X1 U10369 ( .A1(n8994), .A2(n9008), .ZN(n9010) );
  NAND2_X1 U10370 ( .A1(n9010), .A2(n9009), .ZN(n9014) );
  NOR2_X1 U10371 ( .A1(n9012), .A2(n9011), .ZN(n9013) );
  XNOR2_X1 U10372 ( .A(n9014), .B(n9013), .ZN(n9019) );
  NAND2_X1 U10373 ( .A1(n9061), .A2(n9095), .ZN(n9015) );
  NAND2_X1 U10374 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9604) );
  OAI211_X1 U10375 ( .C1(n9350), .C2(n9068), .A(n9015), .B(n9604), .ZN(n9016)
         );
  AOI21_X1 U10376 ( .B1(n9357), .B2(n9084), .A(n9016), .ZN(n9018) );
  NAND2_X1 U10377 ( .A1(n9360), .A2(n9035), .ZN(n9017) );
  OAI211_X1 U10378 ( .C1(n9019), .C2(n4495), .A(n9018), .B(n9017), .ZN(
        P1_U3228) );
  XNOR2_X1 U10379 ( .A(n9021), .B(n9020), .ZN(n9022) );
  XNOR2_X1 U10380 ( .A(n8976), .B(n9022), .ZN(n9027) );
  AOI22_X1 U10381 ( .A1(n9273), .A2(n9076), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9024) );
  NAND2_X1 U10382 ( .A1(n9084), .A2(n9303), .ZN(n9023) );
  OAI211_X1 U10383 ( .C1(n9298), .C2(n9078), .A(n9024), .B(n9023), .ZN(n9025)
         );
  AOI21_X1 U10384 ( .B1(n9408), .B2(n9035), .A(n9025), .ZN(n9026) );
  OAI21_X1 U10385 ( .B1(n9027), .B2(n4495), .A(n9026), .ZN(P1_U3233) );
  NAND2_X1 U10386 ( .A1(n9029), .A2(n9028), .ZN(n9031) );
  XNOR2_X1 U10387 ( .A(n9031), .B(n9030), .ZN(n9037) );
  AOI22_X1 U10388 ( .A1(n9274), .A2(n9076), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9033) );
  NAND2_X1 U10389 ( .A1(n9268), .A2(n9084), .ZN(n9032) );
  OAI211_X1 U10390 ( .C1(n9301), .C2(n9078), .A(n9033), .B(n9032), .ZN(n9034)
         );
  AOI21_X1 U10391 ( .B1(n9398), .B2(n9035), .A(n9034), .ZN(n9036) );
  OAI21_X1 U10392 ( .B1(n9037), .B2(n4495), .A(n9036), .ZN(P1_U3235) );
  AOI21_X1 U10393 ( .B1(n9040), .B2(n9039), .A(n9038), .ZN(n9044) );
  XNOR2_X1 U10394 ( .A(n9042), .B(n9041), .ZN(n9043) );
  XNOR2_X1 U10395 ( .A(n9044), .B(n9043), .ZN(n9052) );
  NAND2_X1 U10396 ( .A1(n9076), .A2(n9099), .ZN(n9045) );
  NAND2_X1 U10397 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9521) );
  OAI211_X1 U10398 ( .C1(n9046), .C2(n9078), .A(n9045), .B(n9521), .ZN(n9049)
         );
  NOR2_X1 U10399 ( .A1(n9047), .A2(n9080), .ZN(n9048) );
  AOI211_X1 U10400 ( .C1(n9050), .C2(n9084), .A(n9049), .B(n9048), .ZN(n9051)
         );
  OAI21_X1 U10401 ( .B1(n9052), .B2(n4495), .A(n9051), .ZN(P1_U3236) );
  OAI21_X1 U10402 ( .B1(n9055), .B2(n9053), .A(n9054), .ZN(n9057) );
  NAND2_X1 U10403 ( .A1(n9057), .A2(n9056), .ZN(n9063) );
  NAND2_X1 U10404 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9620) );
  OAI21_X1 U10405 ( .B1(n9298), .B2(n9068), .A(n9620), .ZN(n9060) );
  NOR2_X1 U10406 ( .A1(n9058), .A2(n9327), .ZN(n9059) );
  AOI211_X1 U10407 ( .C1(n9061), .C2(n9336), .A(n9060), .B(n9059), .ZN(n9062)
         );
  OAI211_X1 U10408 ( .C1(n9331), .C2(n9080), .A(n9063), .B(n9062), .ZN(
        P1_U3238) );
  AOI21_X1 U10409 ( .B1(n9065), .B2(n9064), .A(n4495), .ZN(n9067) );
  NAND2_X1 U10410 ( .A1(n9067), .A2(n9066), .ZN(n9072) );
  NOR2_X1 U10411 ( .A1(n9068), .A2(n9202), .ZN(n9070) );
  OAI22_X1 U10412 ( .A1(n9078), .A2(n9240), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9981), .ZN(n9069) );
  AOI211_X1 U10413 ( .C1(n9210), .C2(n9084), .A(n9070), .B(n9069), .ZN(n9071)
         );
  OAI211_X1 U10414 ( .C1(n9446), .C2(n9080), .A(n9072), .B(n9071), .ZN(
        P1_U3240) );
  AOI21_X1 U10415 ( .B1(n9075), .B2(n9074), .A(n9073), .ZN(n9087) );
  NAND2_X1 U10416 ( .A1(n9076), .A2(n9095), .ZN(n9077) );
  NAND2_X1 U10417 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9579) );
  OAI211_X1 U10418 ( .C1(n9079), .C2(n9078), .A(n9077), .B(n9579), .ZN(n9083)
         );
  NOR2_X1 U10419 ( .A1(n9081), .A2(n9080), .ZN(n9082) );
  AOI211_X1 U10420 ( .C1(n9085), .C2(n9084), .A(n9083), .B(n9082), .ZN(n9086)
         );
  OAI21_X1 U10421 ( .B1(n9087), .B2(n4495), .A(n9086), .ZN(P1_U3241) );
  MUX2_X1 U10422 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9088), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10423 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9187), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10424 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9089), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10425 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9090), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10426 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9091), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10427 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9223), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10428 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9274), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10429 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9092), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10430 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9273), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10431 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9093), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10432 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9338), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10433 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9094), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10434 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9336), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10435 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9095), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10436 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9096), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10437 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9097), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10438 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9098), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10439 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9099), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10440 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9100), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10441 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9101), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10442 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9102), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10443 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9103), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10444 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9104), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10445 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9105), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10446 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9106), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10447 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9107), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10448 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9108), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10449 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n6213), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10450 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9109), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10451 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9110), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI211_X1 U10452 ( .C1(n9113), .C2(n9112), .A(n9602), .B(n9111), .ZN(n9121)
         );
  OAI211_X1 U10453 ( .C1(n9116), .C2(n9115), .A(n9610), .B(n9114), .ZN(n9120)
         );
  AOI22_X1 U10454 ( .A1(n9586), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9119) );
  NAND2_X1 U10455 ( .A1(n9599), .A2(n9117), .ZN(n9118) );
  NAND4_X1 U10456 ( .A1(n9121), .A2(n9120), .A3(n9119), .A4(n9118), .ZN(
        P1_U3244) );
  INV_X1 U10457 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9164) );
  XNOR2_X1 U10458 ( .A(n9562), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n9558) );
  NAND2_X1 U10459 ( .A1(n9549), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9122) );
  OAI21_X1 U10460 ( .B1(n9549), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9122), .ZN(
        n9545) );
  NOR2_X1 U10461 ( .A1(n9524), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9123) );
  AOI21_X1 U10462 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9524), .A(n9123), .ZN(
        n9527) );
  OAI21_X1 U10463 ( .B1(n9141), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9124), .ZN(
        n9499) );
  NAND2_X1 U10464 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n9502), .ZN(n9125) );
  OAI21_X1 U10465 ( .B1(n9502), .B2(P1_REG2_REG_10__SCAN_IN), .A(n9125), .ZN(
        n9498) );
  NOR2_X1 U10466 ( .A1(n9499), .A2(n9498), .ZN(n9497) );
  NAND2_X1 U10467 ( .A1(n9520), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9126) );
  OAI21_X1 U10468 ( .B1(n9520), .B2(P1_REG2_REG_11__SCAN_IN), .A(n9126), .ZN(
        n9513) );
  OAI21_X1 U10469 ( .B1(n9524), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9525), .ZN(
        n9546) );
  NOR2_X1 U10470 ( .A1(n9545), .A2(n9546), .ZN(n9544) );
  NOR2_X1 U10471 ( .A1(n9127), .A2(n9577), .ZN(n9129) );
  INV_X1 U10472 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9572) );
  NOR2_X1 U10473 ( .A1(n9572), .A2(n9573), .ZN(n9571) );
  NOR2_X1 U10474 ( .A1(n9129), .A2(n9571), .ZN(n9583) );
  NAND2_X1 U10475 ( .A1(n9590), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9130) );
  OAI21_X1 U10476 ( .B1(n9590), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9130), .ZN(
        n9582) );
  OR2_X1 U10477 ( .A1(n9600), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U10478 ( .A1(n9600), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9131) );
  AND2_X1 U10479 ( .A1(n9132), .A2(n9131), .ZN(n9595) );
  NAND2_X1 U10480 ( .A1(n9150), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9134) );
  OR2_X1 U10481 ( .A1(n9150), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9133) );
  NAND2_X1 U10482 ( .A1(n9134), .A2(n9133), .ZN(n9608) );
  NAND2_X1 U10483 ( .A1(n9618), .A2(n9134), .ZN(n9136) );
  INV_X1 U10484 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9135) );
  XNOR2_X1 U10485 ( .A(n9136), .B(n9135), .ZN(n9156) );
  INV_X1 U10486 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9138) );
  AOI22_X1 U10487 ( .A1(n9590), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9138), .B2(
        n9137), .ZN(n9589) );
  INV_X1 U10488 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9139) );
  XNOR2_X1 U10489 ( .A(n9562), .B(n9139), .ZN(n9555) );
  NAND2_X1 U10490 ( .A1(n9549), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9145) );
  XNOR2_X1 U10491 ( .A(n9549), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9542) );
  OAI21_X1 U10492 ( .B1(n9141), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9140), .ZN(
        n9496) );
  NAND2_X1 U10493 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n9502), .ZN(n9142) );
  OAI21_X1 U10494 ( .B1(n9502), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9142), .ZN(
        n9495) );
  NOR2_X1 U10495 ( .A1(n9496), .A2(n9495), .ZN(n9494) );
  XNOR2_X1 U10496 ( .A(n9520), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n9516) );
  NOR2_X1 U10497 ( .A1(n9517), .A2(n9516), .ZN(n9515) );
  XNOR2_X1 U10498 ( .A(n9524), .B(n9143), .ZN(n9531) );
  NAND2_X1 U10499 ( .A1(n9530), .A2(n9531), .ZN(n9529) );
  NOR2_X1 U10500 ( .A1(n9542), .A2(n9543), .ZN(n9541) );
  INV_X1 U10501 ( .A(n9541), .ZN(n9144) );
  NAND2_X1 U10502 ( .A1(n9145), .A2(n9144), .ZN(n9554) );
  NAND2_X1 U10503 ( .A1(n9562), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9146) );
  NOR2_X1 U10504 ( .A1(n9147), .A2(n9577), .ZN(n9148) );
  INV_X1 U10505 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9566) );
  XNOR2_X1 U10506 ( .A(n9147), .B(n9577), .ZN(n9567) );
  OAI21_X1 U10507 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n9590), .A(n9587), .ZN(
        n9598) );
  INV_X1 U10508 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9425) );
  XNOR2_X1 U10509 ( .A(n9600), .B(n9425), .ZN(n9597) );
  INV_X1 U10510 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9151) );
  AND2_X1 U10511 ( .A1(n9150), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9152) );
  AOI21_X1 U10512 ( .B1(n9151), .B2(n9615), .A(n9152), .ZN(n9612) );
  NAND2_X1 U10513 ( .A1(n9613), .A2(n9612), .ZN(n9611) );
  INV_X1 U10514 ( .A(n9152), .ZN(n9153) );
  NAND2_X1 U10515 ( .A1(n9611), .A2(n9153), .ZN(n9155) );
  XNOR2_X1 U10516 ( .A(n9155), .B(n9154), .ZN(n9157) );
  AOI22_X1 U10517 ( .A1(n9156), .A2(n9602), .B1(n9610), .B2(n9157), .ZN(n9161)
         );
  INV_X1 U10518 ( .A(n9156), .ZN(n9159) );
  OAI21_X1 U10519 ( .B1(n9157), .B2(n9540), .A(n9616), .ZN(n9158) );
  AOI21_X1 U10520 ( .B1(n9159), .B2(n9602), .A(n9158), .ZN(n9160) );
  MUX2_X1 U10521 ( .A(n9161), .B(n9160), .S(n4331), .Z(n9163) );
  OAI211_X1 U10522 ( .C1(n9164), .C2(n9622), .A(n9163), .B(n9162), .ZN(
        P1_U3262) );
  NOR2_X1 U10523 ( .A1(n9358), .A2(n9369), .ZN(n9173) );
  NOR2_X1 U10524 ( .A1(n9165), .A2(n9330), .ZN(n9166) );
  AOI211_X1 U10525 ( .C1(n9358), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9173), .B(
        n9166), .ZN(n9167) );
  OAI21_X1 U10526 ( .B1(n9168), .B2(n9363), .A(n9167), .ZN(P1_U3263) );
  NAND2_X1 U10527 ( .A1(n9169), .A2(n4359), .ZN(n9170) );
  NAND3_X1 U10528 ( .A1(n9171), .A2(n9354), .A3(n9170), .ZN(n9370) );
  NOR2_X1 U10529 ( .A1(n7902), .A2(n9330), .ZN(n9172) );
  AOI211_X1 U10530 ( .C1(n9358), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9173), .B(
        n9172), .ZN(n9174) );
  OAI21_X1 U10531 ( .B1(n9363), .B2(n9370), .A(n9174), .ZN(P1_U3264) );
  OAI21_X1 U10532 ( .B1(n9176), .B2(n9179), .A(n9175), .ZN(n9441) );
  INV_X1 U10533 ( .A(n9177), .ZN(n9181) );
  INV_X1 U10534 ( .A(n9178), .ZN(n9180) );
  OAI21_X1 U10535 ( .B1(n9181), .B2(n9180), .A(n9179), .ZN(n9186) );
  INV_X1 U10536 ( .A(n9182), .ZN(n9183) );
  OR2_X2 U10537 ( .A1(n9184), .A2(n9183), .ZN(n9185) );
  NAND3_X1 U10538 ( .A1(n9186), .A2(n9352), .A3(n9185), .ZN(n9189) );
  NAND2_X1 U10539 ( .A1(n9187), .A2(n9337), .ZN(n9188) );
  OAI211_X1 U10540 ( .C1(n9202), .C2(n9347), .A(n9189), .B(n9188), .ZN(n9376)
         );
  AOI211_X1 U10541 ( .C1(n9373), .C2(n9191), .A(n9326), .B(n4583), .ZN(n9375)
         );
  NAND2_X1 U10542 ( .A1(n9375), .A2(n9342), .ZN(n9194) );
  AOI22_X1 U10543 ( .A1(n9358), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9192), .B2(
        n9356), .ZN(n9193) );
  OAI211_X1 U10544 ( .C1(n4585), .C2(n9330), .A(n9194), .B(n9193), .ZN(n9195)
         );
  AOI21_X1 U10545 ( .B1(n9365), .B2(n9376), .A(n9195), .ZN(n9196) );
  OAI21_X1 U10546 ( .B1(n9441), .B2(n9368), .A(n9196), .ZN(P1_U3265) );
  AOI211_X1 U10547 ( .C1(n9215), .C2(n9228), .A(n9326), .B(n9197), .ZN(n9380)
         );
  OAI21_X1 U10548 ( .B1(n9207), .B2(n9199), .A(n9198), .ZN(n9200) );
  INV_X1 U10549 ( .A(n9200), .ZN(n9201) );
  OAI222_X1 U10550 ( .A1(n9349), .A2(n9202), .B1(n9347), .B2(n9240), .C1(n9299), .C2(n9201), .ZN(n9379) );
  AOI21_X1 U10551 ( .B1(n9380), .B2(n9203), .A(n9379), .ZN(n9218) );
  OR2_X1 U10552 ( .A1(n9219), .A2(n9204), .ZN(n9206) );
  NAND2_X1 U10553 ( .A1(n9206), .A2(n9205), .ZN(n9208) );
  XNOR2_X1 U10554 ( .A(n9208), .B(n9207), .ZN(n9381) );
  NAND2_X1 U10555 ( .A1(n9381), .A2(n9209), .ZN(n9217) );
  INV_X1 U10556 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9213) );
  INV_X1 U10557 ( .A(n9210), .ZN(n9212) );
  OAI22_X1 U10558 ( .A1(n9365), .A2(n9213), .B1(n9212), .B2(n9211), .ZN(n9214)
         );
  AOI21_X1 U10559 ( .B1(n9215), .B2(n9359), .A(n9214), .ZN(n9216) );
  OAI211_X1 U10560 ( .C1(n9358), .C2(n9218), .A(n9217), .B(n9216), .ZN(
        P1_U3267) );
  XNOR2_X1 U10561 ( .A(n9219), .B(n9222), .ZN(n9451) );
  OAI21_X1 U10562 ( .B1(n9222), .B2(n9221), .A(n9220), .ZN(n9227) );
  NAND2_X1 U10563 ( .A1(n9223), .A2(n9335), .ZN(n9224) );
  OAI21_X1 U10564 ( .B1(n9225), .B2(n9349), .A(n9224), .ZN(n9226) );
  AOI21_X1 U10565 ( .B1(n9227), .B2(n9352), .A(n9226), .ZN(n9386) );
  INV_X1 U10566 ( .A(n9386), .ZN(n9233) );
  OAI211_X1 U10567 ( .C1(n4571), .C2(n4334), .A(n9354), .B(n9228), .ZN(n9385)
         );
  AOI22_X1 U10568 ( .A1(n9358), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9229), .B2(
        n9356), .ZN(n9231) );
  NAND2_X1 U10569 ( .A1(n9449), .A2(n9359), .ZN(n9230) );
  OAI211_X1 U10570 ( .C1(n9385), .C2(n9363), .A(n9231), .B(n9230), .ZN(n9232)
         );
  AOI21_X1 U10571 ( .B1(n9233), .B2(n9365), .A(n9232), .ZN(n9234) );
  OAI21_X1 U10572 ( .B1(n9451), .B2(n9368), .A(n9234), .ZN(P1_U3268) );
  XNOR2_X1 U10573 ( .A(n9235), .B(n9236), .ZN(n9455) );
  XNOR2_X1 U10574 ( .A(n9237), .B(n9236), .ZN(n9239) );
  OAI222_X1 U10575 ( .A1(n9349), .A2(n9240), .B1(n9239), .B2(n9299), .C1(n9347), .C2(n9238), .ZN(n9389) );
  AOI211_X1 U10576 ( .C1(n6269), .C2(n4575), .A(n9326), .B(n4334), .ZN(n9390)
         );
  NAND2_X1 U10577 ( .A1(n9390), .A2(n9342), .ZN(n9243) );
  AOI22_X1 U10578 ( .A1(n9358), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9241), .B2(
        n9356), .ZN(n9242) );
  OAI211_X1 U10579 ( .C1(n6268), .C2(n9330), .A(n9243), .B(n9242), .ZN(n9244)
         );
  AOI21_X1 U10580 ( .B1(n9365), .B2(n9389), .A(n9244), .ZN(n9245) );
  OAI21_X1 U10581 ( .B1(n9455), .B2(n9368), .A(n9245), .ZN(P1_U3269) );
  XNOR2_X1 U10582 ( .A(n9246), .B(n9247), .ZN(n9460) );
  OR2_X1 U10583 ( .A1(n9248), .A2(n9247), .ZN(n9249) );
  NAND2_X1 U10584 ( .A1(n9250), .A2(n9249), .ZN(n9253) );
  OAI22_X1 U10585 ( .A1(n9283), .A2(n9347), .B1(n9251), .B2(n9349), .ZN(n9252)
         );
  AOI21_X1 U10586 ( .B1(n9253), .B2(n9352), .A(n9252), .ZN(n9394) );
  INV_X1 U10587 ( .A(n9394), .ZN(n9262) );
  NAND2_X1 U10588 ( .A1(n9458), .A2(n9266), .ZN(n9254) );
  NAND2_X1 U10589 ( .A1(n9254), .A2(n9354), .ZN(n9256) );
  OR2_X1 U10590 ( .A1(n9256), .A2(n9255), .ZN(n9393) );
  INV_X1 U10591 ( .A(n9257), .ZN(n9258) );
  AOI22_X1 U10592 ( .A1(n9258), .A2(n9356), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9358), .ZN(n9260) );
  NAND2_X1 U10593 ( .A1(n9458), .A2(n9359), .ZN(n9259) );
  OAI211_X1 U10594 ( .C1(n9393), .C2(n9363), .A(n9260), .B(n9259), .ZN(n9261)
         );
  AOI21_X1 U10595 ( .B1(n9262), .B2(n9365), .A(n9261), .ZN(n9263) );
  OAI21_X1 U10596 ( .B1(n9460), .B2(n9368), .A(n9263), .ZN(P1_U3270) );
  XNOR2_X1 U10597 ( .A(n9264), .B(n9271), .ZN(n9401) );
  INV_X1 U10598 ( .A(n9266), .ZN(n9267) );
  AOI211_X1 U10599 ( .C1(n9398), .C2(n9287), .A(n9326), .B(n9267), .ZN(n9397)
         );
  AOI22_X1 U10600 ( .A1(n9268), .A2(n9356), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9358), .ZN(n9269) );
  OAI21_X1 U10601 ( .B1(n6278), .B2(n9330), .A(n9269), .ZN(n9277) );
  OAI21_X1 U10602 ( .B1(n9272), .B2(n9271), .A(n9270), .ZN(n9275) );
  AOI222_X1 U10603 ( .A1(n9352), .A2(n9275), .B1(n9274), .B2(n9337), .C1(n9273), .C2(n9335), .ZN(n9400) );
  NOR2_X1 U10604 ( .A1(n9400), .A2(n9358), .ZN(n9276) );
  AOI211_X1 U10605 ( .C1(n9397), .C2(n9342), .A(n9277), .B(n9276), .ZN(n9278)
         );
  OAI21_X1 U10606 ( .B1(n9401), .B2(n9368), .A(n9278), .ZN(P1_U3271) );
  XOR2_X1 U10607 ( .A(n9282), .B(n9279), .Z(n9466) );
  OAI21_X1 U10608 ( .B1(n9282), .B2(n9281), .A(n9280), .ZN(n9285) );
  OAI22_X1 U10609 ( .A1(n9283), .A2(n9349), .B1(n9313), .B2(n9347), .ZN(n9284)
         );
  AOI21_X1 U10610 ( .B1(n9285), .B2(n9352), .A(n9284), .ZN(n9403) );
  INV_X1 U10611 ( .A(n9403), .ZN(n9293) );
  INV_X1 U10612 ( .A(n9286), .ZN(n9302) );
  OAI211_X1 U10613 ( .C1(n9288), .C2(n9302), .A(n9354), .B(n9287), .ZN(n9402)
         );
  AOI22_X1 U10614 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(n9358), .B1(n9289), .B2(
        n9356), .ZN(n9291) );
  NAND2_X1 U10615 ( .A1(n9464), .A2(n9359), .ZN(n9290) );
  OAI211_X1 U10616 ( .C1(n9402), .C2(n9363), .A(n9291), .B(n9290), .ZN(n9292)
         );
  AOI21_X1 U10617 ( .B1(n9293), .B2(n9365), .A(n9292), .ZN(n9294) );
  OAI21_X1 U10618 ( .B1(n9466), .B2(n9368), .A(n9294), .ZN(P1_U3272) );
  XOR2_X1 U10619 ( .A(n9295), .B(n9296), .Z(n9410) );
  XNOR2_X1 U10620 ( .A(n9297), .B(n9296), .ZN(n9300) );
  OAI222_X1 U10621 ( .A1(n9349), .A2(n9301), .B1(n9300), .B2(n9299), .C1(n9347), .C2(n9298), .ZN(n9406) );
  INV_X1 U10622 ( .A(n9408), .ZN(n9306) );
  AOI211_X1 U10623 ( .C1(n9408), .C2(n9316), .A(n9326), .B(n9302), .ZN(n9407)
         );
  NAND2_X1 U10624 ( .A1(n9407), .A2(n9342), .ZN(n9305) );
  AOI22_X1 U10625 ( .A1(n9358), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9303), .B2(
        n9356), .ZN(n9304) );
  OAI211_X1 U10626 ( .C1(n9306), .C2(n9330), .A(n9305), .B(n9304), .ZN(n9307)
         );
  AOI21_X1 U10627 ( .B1(n9365), .B2(n9406), .A(n9307), .ZN(n9308) );
  OAI21_X1 U10628 ( .B1(n9410), .B2(n9368), .A(n9308), .ZN(P1_U3273) );
  XNOR2_X1 U10629 ( .A(n9309), .B(n9312), .ZN(n9473) );
  OAI21_X1 U10630 ( .B1(n9312), .B2(n9311), .A(n9310), .ZN(n9315) );
  OAI22_X1 U10631 ( .A1(n9313), .A2(n9349), .B1(n9350), .B2(n9347), .ZN(n9314)
         );
  AOI21_X1 U10632 ( .B1(n9315), .B2(n9352), .A(n9314), .ZN(n9412) );
  INV_X1 U10633 ( .A(n9412), .ZN(n9322) );
  OAI211_X1 U10634 ( .C1(n9317), .C2(n9325), .A(n9354), .B(n9316), .ZN(n9411)
         );
  AOI22_X1 U10635 ( .A1(n9358), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9318), .B2(
        n9356), .ZN(n9320) );
  NAND2_X1 U10636 ( .A1(n9470), .A2(n9359), .ZN(n9319) );
  OAI211_X1 U10637 ( .C1(n9411), .C2(n9363), .A(n9320), .B(n9319), .ZN(n9321)
         );
  AOI21_X1 U10638 ( .B1(n9322), .B2(n9365), .A(n9321), .ZN(n9323) );
  OAI21_X1 U10639 ( .B1(n9473), .B2(n9368), .A(n9323), .ZN(P1_U3274) );
  XOR2_X1 U10640 ( .A(n9333), .B(n9324), .Z(n9420) );
  AOI211_X1 U10641 ( .C1(n9417), .C2(n4355), .A(n9326), .B(n9325), .ZN(n9416)
         );
  INV_X1 U10642 ( .A(n9327), .ZN(n9328) );
  AOI22_X1 U10643 ( .A1(n9358), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9328), .B2(
        n9356), .ZN(n9329) );
  OAI21_X1 U10644 ( .B1(n9331), .B2(n9330), .A(n9329), .ZN(n9341) );
  OAI21_X1 U10645 ( .B1(n9334), .B2(n9333), .A(n9332), .ZN(n9339) );
  AOI222_X1 U10646 ( .A1(n9352), .A2(n9339), .B1(n9338), .B2(n9337), .C1(n9336), .C2(n9335), .ZN(n9419) );
  NOR2_X1 U10647 ( .A1(n9419), .A2(n9358), .ZN(n9340) );
  AOI211_X1 U10648 ( .C1(n9416), .C2(n9342), .A(n9341), .B(n9340), .ZN(n9343)
         );
  OAI21_X1 U10649 ( .B1(n9420), .B2(n9368), .A(n9343), .ZN(P1_U3275) );
  XNOR2_X1 U10650 ( .A(n9344), .B(n9346), .ZN(n9479) );
  XNOR2_X1 U10651 ( .A(n9346), .B(n9345), .ZN(n9353) );
  OAI22_X1 U10652 ( .A1(n9350), .A2(n9349), .B1(n9348), .B2(n9347), .ZN(n9351)
         );
  AOI21_X1 U10653 ( .B1(n9353), .B2(n9352), .A(n9351), .ZN(n9422) );
  INV_X1 U10654 ( .A(n9422), .ZN(n9366) );
  INV_X1 U10655 ( .A(n9360), .ZN(n9423) );
  OAI211_X1 U10656 ( .C1(n9423), .C2(n9355), .A(n4355), .B(n9354), .ZN(n9421)
         );
  AOI22_X1 U10657 ( .A1(n9358), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9357), .B2(
        n9356), .ZN(n9362) );
  NAND2_X1 U10658 ( .A1(n9360), .A2(n9359), .ZN(n9361) );
  OAI211_X1 U10659 ( .C1(n9421), .C2(n9363), .A(n9362), .B(n9361), .ZN(n9364)
         );
  AOI21_X1 U10660 ( .B1(n9366), .B2(n9365), .A(n9364), .ZN(n9367) );
  OAI21_X1 U10661 ( .B1(n9479), .B2(n9368), .A(n9367), .ZN(P1_U3276) );
  AND2_X1 U10662 ( .A1(n9370), .A2(n9369), .ZN(n9436) );
  INV_X1 U10663 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9371) );
  MUX2_X1 U10664 ( .A(n9436), .B(n9371), .S(n9656), .Z(n9372) );
  OAI21_X1 U10665 ( .B1(n7902), .B2(n9384), .A(n9372), .ZN(P1_U3552) );
  NOR2_X2 U10666 ( .A1(n9376), .A2(n4899), .ZN(n9439) );
  OAI21_X1 U10667 ( .B1(n9441), .B2(n9427), .A(n9378), .ZN(P1_U3550) );
  INV_X1 U10668 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9382) );
  AOI211_X1 U10669 ( .C1(n9381), .C2(n9648), .A(n9380), .B(n9379), .ZN(n9442)
         );
  MUX2_X1 U10670 ( .A(n9382), .B(n9442), .S(n9659), .Z(n9383) );
  OAI21_X1 U10671 ( .B1(n9446), .B2(n9384), .A(n9383), .ZN(P1_U3548) );
  NAND2_X1 U10672 ( .A1(n9386), .A2(n9385), .ZN(n9447) );
  MUX2_X1 U10673 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9447), .S(n9659), .Z(n9387) );
  AOI21_X1 U10674 ( .B1(n9414), .B2(n9449), .A(n9387), .ZN(n9388) );
  OAI21_X1 U10675 ( .B1(n9451), .B2(n9427), .A(n9388), .ZN(P1_U3547) );
  INV_X1 U10676 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9391) );
  AOI211_X1 U10677 ( .C1(n9430), .C2(n6269), .A(n9390), .B(n9389), .ZN(n9452)
         );
  MUX2_X1 U10678 ( .A(n9391), .B(n9452), .S(n9659), .Z(n9392) );
  OAI21_X1 U10679 ( .B1(n9455), .B2(n9427), .A(n9392), .ZN(P1_U3546) );
  NAND2_X1 U10680 ( .A1(n9394), .A2(n9393), .ZN(n9456) );
  MUX2_X1 U10681 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9456), .S(n9659), .Z(n9395) );
  AOI21_X1 U10682 ( .B1(n9414), .B2(n9458), .A(n9395), .ZN(n9396) );
  OAI21_X1 U10683 ( .B1(n9460), .B2(n9427), .A(n9396), .ZN(P1_U3545) );
  AOI21_X1 U10684 ( .B1(n9430), .B2(n9398), .A(n9397), .ZN(n9399) );
  OAI211_X1 U10685 ( .C1(n9401), .C2(n9433), .A(n9400), .B(n9399), .ZN(n9461)
         );
  MUX2_X1 U10686 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9461), .S(n9659), .Z(
        P1_U3544) );
  NAND2_X1 U10687 ( .A1(n9403), .A2(n9402), .ZN(n9462) );
  MUX2_X1 U10688 ( .A(n9462), .B(P1_REG1_REG_21__SCAN_IN), .S(n9656), .Z(n9404) );
  AOI21_X1 U10689 ( .B1(n9414), .B2(n9464), .A(n9404), .ZN(n9405) );
  OAI21_X1 U10690 ( .B1(n9466), .B2(n9427), .A(n9405), .ZN(P1_U3543) );
  AOI211_X1 U10691 ( .C1(n9430), .C2(n9408), .A(n9407), .B(n9406), .ZN(n9409)
         );
  OAI21_X1 U10692 ( .B1(n9410), .B2(n9433), .A(n9409), .ZN(n9467) );
  MUX2_X1 U10693 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9467), .S(n9659), .Z(
        P1_U3542) );
  NAND2_X1 U10694 ( .A1(n9412), .A2(n9411), .ZN(n9468) );
  MUX2_X1 U10695 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9468), .S(n9659), .Z(n9413) );
  AOI21_X1 U10696 ( .B1(n9414), .B2(n9470), .A(n9413), .ZN(n9415) );
  OAI21_X1 U10697 ( .B1(n9473), .B2(n9427), .A(n9415), .ZN(P1_U3541) );
  AOI21_X1 U10698 ( .B1(n9430), .B2(n9417), .A(n9416), .ZN(n9418) );
  OAI211_X1 U10699 ( .C1(n9420), .C2(n9433), .A(n9419), .B(n9418), .ZN(n9474)
         );
  MUX2_X1 U10700 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9474), .S(n9659), .Z(
        P1_U3540) );
  OAI211_X1 U10701 ( .C1(n9423), .C2(n9645), .A(n9422), .B(n9421), .ZN(n9424)
         );
  INV_X1 U10702 ( .A(n9424), .ZN(n9475) );
  MUX2_X1 U10703 ( .A(n9425), .B(n9475), .S(n9659), .Z(n9426) );
  OAI21_X1 U10704 ( .B1(n9479), .B2(n9427), .A(n9426), .ZN(P1_U3539) );
  AOI21_X1 U10705 ( .B1(n9430), .B2(n9429), .A(n9428), .ZN(n9431) );
  OAI211_X1 U10706 ( .C1(n9434), .C2(n9433), .A(n9432), .B(n9431), .ZN(n9481)
         );
  MUX2_X1 U10707 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9481), .S(n9659), .Z(
        P1_U3538) );
  MUX2_X1 U10708 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9435), .S(n9659), .Z(
        P1_U3522) );
  INV_X1 U10709 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9437) );
  MUX2_X1 U10710 ( .A(n9437), .B(n9436), .S(n9650), .Z(n9438) );
  OAI21_X1 U10711 ( .B1(n7902), .B2(n9445), .A(n9438), .ZN(P1_U3520) );
  INV_X1 U10712 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9440) );
  INV_X1 U10713 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9443) );
  MUX2_X1 U10714 ( .A(n9443), .B(n9442), .S(n9650), .Z(n9444) );
  OAI21_X1 U10715 ( .B1(n9446), .B2(n9445), .A(n9444), .ZN(P1_U3516) );
  MUX2_X1 U10716 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9447), .S(n9650), .Z(n9448) );
  AOI21_X1 U10717 ( .B1(n9471), .B2(n9449), .A(n9448), .ZN(n9450) );
  OAI21_X1 U10718 ( .B1(n9451), .B2(n9478), .A(n9450), .ZN(P1_U3515) );
  INV_X1 U10719 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9453) );
  MUX2_X1 U10720 ( .A(n9453), .B(n9452), .S(n9650), .Z(n9454) );
  OAI21_X1 U10721 ( .B1(n9455), .B2(n9478), .A(n9454), .ZN(P1_U3514) );
  MUX2_X1 U10722 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9456), .S(n9650), .Z(n9457) );
  AOI21_X1 U10723 ( .B1(n9471), .B2(n9458), .A(n9457), .ZN(n9459) );
  OAI21_X1 U10724 ( .B1(n9460), .B2(n9478), .A(n9459), .ZN(P1_U3513) );
  MUX2_X1 U10725 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9461), .S(n9480), .Z(
        P1_U3512) );
  MUX2_X1 U10726 ( .A(n9462), .B(P1_REG0_REG_21__SCAN_IN), .S(n6284), .Z(n9463) );
  AOI21_X1 U10727 ( .B1(n9471), .B2(n9464), .A(n9463), .ZN(n9465) );
  OAI21_X1 U10728 ( .B1(n9466), .B2(n9478), .A(n9465), .ZN(P1_U3511) );
  MUX2_X1 U10729 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9467), .S(n9480), .Z(
        P1_U3510) );
  MUX2_X1 U10730 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9468), .S(n9650), .Z(n9469) );
  AOI21_X1 U10731 ( .B1(n9471), .B2(n9470), .A(n9469), .ZN(n9472) );
  OAI21_X1 U10732 ( .B1(n9473), .B2(n9478), .A(n9472), .ZN(P1_U3509) );
  MUX2_X1 U10733 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9474), .S(n9480), .Z(
        P1_U3507) );
  INV_X1 U10734 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9476) );
  MUX2_X1 U10735 ( .A(n9476), .B(n9475), .S(n9480), .Z(n9477) );
  OAI21_X1 U10736 ( .B1(n9479), .B2(n9478), .A(n9477), .ZN(P1_U3504) );
  MUX2_X1 U10737 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9481), .S(n9480), .Z(
        P1_U3501) );
  MUX2_X1 U10738 ( .A(P1_D_REG_0__SCAN_IN), .B(n9482), .S(n9623), .Z(P1_U3439)
         );
  NOR4_X1 U10739 ( .A1(n9483), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n9484), .ZN(n9485) );
  AOI21_X1 U10740 ( .B1(n9486), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9485), .ZN(
        n9487) );
  OAI21_X1 U10741 ( .B1(n9489), .B2(n9488), .A(n9487), .ZN(P1_U3324) );
  OAI222_X1 U10742 ( .A1(n9493), .A2(n9492), .B1(n9491), .B2(P1_U3086), .C1(
        n10062), .C2(n9490), .ZN(P1_U3326) );
  INV_X1 U10743 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9505) );
  AOI211_X1 U10744 ( .C1(n9496), .C2(n9495), .A(n9540), .B(n9494), .ZN(n9501)
         );
  AOI211_X1 U10745 ( .C1(n9499), .C2(n9498), .A(n9607), .B(n9497), .ZN(n9500)
         );
  AOI211_X1 U10746 ( .C1(n9599), .C2(n9502), .A(n9501), .B(n9500), .ZN(n9504)
         );
  OAI211_X1 U10747 ( .C1(n9505), .C2(n9622), .A(n9504), .B(n9503), .ZN(
        P1_U3253) );
  XNOR2_X1 U10748 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  OAI21_X1 U10749 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n9507), .A(n9506), .ZN(
        n9508) );
  XNOR2_X1 U10750 ( .A(n9508), .B(n5674), .ZN(n9511) );
  AOI22_X1 U10751 ( .A1(n9586), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9509) );
  OAI21_X1 U10752 ( .B1(n9511), .B2(n9510), .A(n9509), .ZN(P1_U3243) );
  INV_X1 U10753 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9523) );
  AOI211_X1 U10754 ( .C1(n9514), .C2(n9513), .A(n9512), .B(n9607), .ZN(n9519)
         );
  AOI211_X1 U10755 ( .C1(n9517), .C2(n9516), .A(n9515), .B(n9540), .ZN(n9518)
         );
  AOI211_X1 U10756 ( .C1(n9599), .C2(n9520), .A(n9519), .B(n9518), .ZN(n9522)
         );
  OAI211_X1 U10757 ( .C1(n9523), .C2(n9622), .A(n9522), .B(n9521), .ZN(
        P1_U3254) );
  INV_X1 U10758 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9539) );
  INV_X1 U10759 ( .A(n9524), .ZN(n9535) );
  OAI21_X1 U10760 ( .B1(n9527), .B2(n9526), .A(n9525), .ZN(n9528) );
  NAND2_X1 U10761 ( .A1(n9602), .A2(n9528), .ZN(n9534) );
  OAI21_X1 U10762 ( .B1(n9531), .B2(n9530), .A(n9529), .ZN(n9532) );
  NAND2_X1 U10763 ( .A1(n9610), .A2(n9532), .ZN(n9533) );
  OAI211_X1 U10764 ( .C1(n9616), .C2(n9535), .A(n9534), .B(n9533), .ZN(n9536)
         );
  INV_X1 U10765 ( .A(n9536), .ZN(n9538) );
  OAI211_X1 U10766 ( .C1(n9539), .C2(n9622), .A(n9538), .B(n9537), .ZN(
        P1_U3255) );
  INV_X1 U10767 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9552) );
  AOI211_X1 U10768 ( .C1(n9543), .C2(n9542), .A(n9541), .B(n9540), .ZN(n9548)
         );
  AOI211_X1 U10769 ( .C1(n9546), .C2(n9545), .A(n9544), .B(n9607), .ZN(n9547)
         );
  AOI211_X1 U10770 ( .C1(n9599), .C2(n9549), .A(n9548), .B(n9547), .ZN(n9551)
         );
  OAI211_X1 U10771 ( .C1(n9552), .C2(n9622), .A(n9551), .B(n9550), .ZN(
        P1_U3256) );
  INV_X1 U10772 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9565) );
  OAI211_X1 U10773 ( .C1(n9555), .C2(n9554), .A(n9610), .B(n9553), .ZN(n9556)
         );
  INV_X1 U10774 ( .A(n9556), .ZN(n9561) );
  AOI211_X1 U10775 ( .C1(n9559), .C2(n9558), .A(n9557), .B(n9607), .ZN(n9560)
         );
  AOI211_X1 U10776 ( .C1(n9599), .C2(n9562), .A(n9561), .B(n9560), .ZN(n9564)
         );
  OAI211_X1 U10777 ( .C1(n9565), .C2(n9622), .A(n9564), .B(n9563), .ZN(
        P1_U3257) );
  INV_X1 U10778 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10016) );
  NAND2_X1 U10779 ( .A1(n9567), .A2(n9566), .ZN(n9570) );
  INV_X1 U10780 ( .A(n9568), .ZN(n9569) );
  NAND3_X1 U10781 ( .A1(n9610), .A2(n9570), .A3(n9569), .ZN(n9576) );
  AOI21_X1 U10782 ( .B1(n9573), .B2(n9572), .A(n9571), .ZN(n9574) );
  NAND2_X1 U10783 ( .A1(n9602), .A2(n9574), .ZN(n9575) );
  OAI211_X1 U10784 ( .C1(n9616), .C2(n9577), .A(n9576), .B(n9575), .ZN(n9578)
         );
  INV_X1 U10785 ( .A(n9578), .ZN(n9580) );
  OAI211_X1 U10786 ( .C1(n10016), .C2(n9622), .A(n9580), .B(n9579), .ZN(
        P1_U3258) );
  AOI211_X1 U10787 ( .C1(n9583), .C2(n9582), .A(n9581), .B(n9607), .ZN(n9584)
         );
  AOI211_X1 U10788 ( .C1(P1_ADDR_REG_16__SCAN_IN), .C2(n9586), .A(n9585), .B(
        n9584), .ZN(n9593) );
  OAI21_X1 U10789 ( .B1(n9589), .B2(n9588), .A(n9587), .ZN(n9591) );
  AOI22_X1 U10790 ( .A1(n9591), .A2(n9610), .B1(n9590), .B2(n9599), .ZN(n9592)
         );
  NAND2_X1 U10791 ( .A1(n9593), .A2(n9592), .ZN(P1_U3259) );
  INV_X1 U10792 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9606) );
  OAI21_X1 U10793 ( .B1(n9596), .B2(n9595), .A(n9594), .ZN(n9603) );
  XNOR2_X1 U10794 ( .A(n9598), .B(n9597), .ZN(n9601) );
  AOI222_X1 U10795 ( .A1(n9603), .A2(n9602), .B1(n9610), .B2(n9601), .C1(n9600), .C2(n9599), .ZN(n9605) );
  OAI211_X1 U10796 ( .C1(n9606), .C2(n9622), .A(n9605), .B(n9604), .ZN(
        P1_U3260) );
  AOI21_X1 U10797 ( .B1(n9609), .B2(n9608), .A(n9607), .ZN(n9619) );
  OAI211_X1 U10798 ( .C1(n9613), .C2(n9612), .A(n9611), .B(n9610), .ZN(n9614)
         );
  OAI21_X1 U10799 ( .B1(n9616), .B2(n9615), .A(n9614), .ZN(n9617) );
  AOI21_X1 U10800 ( .B1(n9619), .B2(n9618), .A(n9617), .ZN(n9621) );
  OAI211_X1 U10801 ( .C1(n9908), .C2(n9622), .A(n9621), .B(n9620), .ZN(
        P1_U3261) );
  AND2_X1 U10802 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9624), .ZN(P1_U3294) );
  AND2_X1 U10803 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9624), .ZN(P1_U3295) );
  AND2_X1 U10804 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9624), .ZN(P1_U3296) );
  AND2_X1 U10805 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9624), .ZN(P1_U3297) );
  AND2_X1 U10806 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9624), .ZN(P1_U3298) );
  AND2_X1 U10807 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9624), .ZN(P1_U3299) );
  AND2_X1 U10808 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9624), .ZN(P1_U3300) );
  AND2_X1 U10809 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9624), .ZN(P1_U3301) );
  AND2_X1 U10810 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9624), .ZN(P1_U3302) );
  AND2_X1 U10811 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9624), .ZN(P1_U3303) );
  INV_X1 U10812 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10054) );
  NOR2_X1 U10813 ( .A1(n9623), .A2(n10054), .ZN(P1_U3304) );
  AND2_X1 U10814 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9624), .ZN(P1_U3305) );
  AND2_X1 U10815 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9624), .ZN(P1_U3306) );
  AND2_X1 U10816 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9624), .ZN(P1_U3307) );
  AND2_X1 U10817 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9624), .ZN(P1_U3308) );
  AND2_X1 U10818 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9624), .ZN(P1_U3309) );
  AND2_X1 U10819 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9624), .ZN(P1_U3310) );
  AND2_X1 U10820 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9624), .ZN(P1_U3311) );
  AND2_X1 U10821 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9624), .ZN(P1_U3312) );
  AND2_X1 U10822 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9624), .ZN(P1_U3313) );
  AND2_X1 U10823 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9624), .ZN(P1_U3314) );
  AND2_X1 U10824 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9624), .ZN(P1_U3315) );
  AND2_X1 U10825 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9624), .ZN(P1_U3316) );
  AND2_X1 U10826 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9624), .ZN(P1_U3317) );
  AND2_X1 U10827 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9624), .ZN(P1_U3318) );
  AND2_X1 U10828 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9624), .ZN(P1_U3319) );
  AND2_X1 U10829 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9624), .ZN(P1_U3320) );
  INV_X1 U10830 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10003) );
  NOR2_X1 U10831 ( .A1(n9623), .A2(n10003), .ZN(P1_U3321) );
  AND2_X1 U10832 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9624), .ZN(P1_U3322) );
  AND2_X1 U10833 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9624), .ZN(P1_U3323) );
  OAI21_X1 U10834 ( .B1(n9626), .B2(n9645), .A(n9625), .ZN(n9628) );
  AOI211_X1 U10835 ( .C1(n9648), .C2(n9629), .A(n9628), .B(n9627), .ZN(n9651)
         );
  INV_X1 U10836 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9630) );
  AOI22_X1 U10837 ( .A1(n9650), .A2(n9651), .B1(n9630), .B2(n6284), .ZN(
        P1_U3465) );
  OAI21_X1 U10838 ( .B1(n9632), .B2(n9645), .A(n9631), .ZN(n9634) );
  AOI211_X1 U10839 ( .C1(n9648), .C2(n9635), .A(n9634), .B(n9633), .ZN(n9653)
         );
  INV_X1 U10840 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9636) );
  AOI22_X1 U10841 ( .A1(n9650), .A2(n9653), .B1(n9636), .B2(n6284), .ZN(
        P1_U3471) );
  OAI21_X1 U10842 ( .B1(n9638), .B2(n9645), .A(n9637), .ZN(n9640) );
  AOI211_X1 U10843 ( .C1(n9648), .C2(n9641), .A(n9640), .B(n9639), .ZN(n9655)
         );
  INV_X1 U10844 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9642) );
  AOI22_X1 U10845 ( .A1(n9650), .A2(n9655), .B1(n9642), .B2(n6284), .ZN(
        P1_U3480) );
  OAI211_X1 U10846 ( .C1(n9646), .C2(n9645), .A(n9644), .B(n9643), .ZN(n9647)
         );
  AOI21_X1 U10847 ( .B1(n9649), .B2(n9648), .A(n9647), .ZN(n9658) );
  INV_X1 U10848 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10070) );
  AOI22_X1 U10849 ( .A1(n9650), .A2(n9658), .B1(n10070), .B2(n6284), .ZN(
        P1_U3483) );
  AOI22_X1 U10850 ( .A1(n9659), .A2(n9651), .B1(n6365), .B2(n9656), .ZN(
        P1_U3526) );
  INV_X1 U10851 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9652) );
  AOI22_X1 U10852 ( .A1(n9659), .A2(n9653), .B1(n9652), .B2(n9656), .ZN(
        P1_U3528) );
  INV_X1 U10853 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9654) );
  AOI22_X1 U10854 ( .A1(n9659), .A2(n9655), .B1(n9654), .B2(n9656), .ZN(
        P1_U3531) );
  INV_X1 U10855 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9657) );
  AOI22_X1 U10856 ( .A1(n9659), .A2(n9658), .B1(n9657), .B2(n9656), .ZN(
        P1_U3532) );
  OAI21_X1 U10857 ( .B1(n9660), .B2(P2_REG2_REG_3__SCAN_IN), .A(n9694), .ZN(
        n9661) );
  INV_X1 U10858 ( .A(n9661), .ZN(n9669) );
  XNOR2_X1 U10859 ( .A(n9662), .B(n6714), .ZN(n9663) );
  OR2_X1 U10860 ( .A1(n9664), .A2(n9663), .ZN(n9668) );
  AOI21_X1 U10861 ( .B1(n9846), .B2(n9666), .A(n9665), .ZN(n9667) );
  OAI211_X1 U10862 ( .C1(n9860), .C2(n9669), .A(n9668), .B(n9667), .ZN(n9670)
         );
  INV_X1 U10863 ( .A(n9670), .ZN(n9678) );
  NAND2_X1 U10864 ( .A1(n9672), .A2(n9671), .ZN(n9674) );
  AOI21_X1 U10865 ( .B1(n9675), .B2(n9674), .A(n9673), .ZN(n9676) );
  AOI21_X1 U10866 ( .B1(n9845), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n9676), .ZN(
        n9677) );
  NAND2_X1 U10867 ( .A1(n9678), .A2(n9677), .ZN(P2_U3185) );
  INV_X1 U10868 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9703) );
  OAI21_X1 U10869 ( .B1(n9681), .B2(n9680), .A(n9679), .ZN(n9682) );
  NAND2_X1 U10870 ( .A1(n9856), .A2(n9682), .ZN(n9701) );
  INV_X1 U10871 ( .A(n9683), .ZN(n9686) );
  INV_X1 U10872 ( .A(n9684), .ZN(n9685) );
  AOI21_X1 U10873 ( .B1(n9846), .B2(n9686), .A(n9685), .ZN(n9700) );
  INV_X1 U10874 ( .A(n9687), .ZN(n9688) );
  XNOR2_X1 U10875 ( .A(n9689), .B(n9688), .ZN(n9690) );
  NAND2_X1 U10876 ( .A1(n9690), .A2(n9855), .ZN(n9699) );
  INV_X1 U10877 ( .A(n9691), .ZN(n9693) );
  NAND3_X1 U10878 ( .A1(n9694), .A2(n9693), .A3(n9692), .ZN(n9695) );
  AND2_X1 U10879 ( .A1(n9696), .A2(n9695), .ZN(n9697) );
  OR2_X1 U10880 ( .A1(n9860), .A2(n9697), .ZN(n9698) );
  AND4_X1 U10881 ( .A1(n9701), .A2(n9700), .A3(n9699), .A4(n9698), .ZN(n9702)
         );
  OAI21_X1 U10882 ( .B1(n9745), .B2(n9703), .A(n9702), .ZN(P2_U3186) );
  INV_X1 U10883 ( .A(n9704), .ZN(n9706) );
  NAND3_X1 U10884 ( .A1(n9707), .A2(n9706), .A3(n9705), .ZN(n9708) );
  AND2_X1 U10885 ( .A1(n9709), .A2(n9708), .ZN(n9719) );
  OAI21_X1 U10886 ( .B1(n9712), .B2(n9711), .A(n9710), .ZN(n9713) );
  NAND2_X1 U10887 ( .A1(n9856), .A2(n9713), .ZN(n9718) );
  INV_X1 U10888 ( .A(n9714), .ZN(n9716) );
  AOI21_X1 U10889 ( .B1(n9846), .B2(n9716), .A(n9715), .ZN(n9717) );
  OAI211_X1 U10890 ( .C1(n9719), .C2(n9860), .A(n9718), .B(n9717), .ZN(n9720)
         );
  INV_X1 U10891 ( .A(n9720), .ZN(n9726) );
  OAI21_X1 U10892 ( .B1(n9723), .B2(n9722), .A(n9721), .ZN(n9724) );
  AOI22_X1 U10893 ( .A1(n9724), .A2(n9855), .B1(n9845), .B2(
        P2_ADDR_REG_6__SCAN_IN), .ZN(n9725) );
  NAND2_X1 U10894 ( .A1(n9726), .A2(n9725), .ZN(P2_U3188) );
  AOI21_X1 U10895 ( .B1(n9729), .B2(n9728), .A(n9727), .ZN(n9737) );
  OAI21_X1 U10896 ( .B1(n9731), .B2(P2_REG1_REG_9__SCAN_IN), .A(n9730), .ZN(
        n9732) );
  NAND2_X1 U10897 ( .A1(n9856), .A2(n9732), .ZN(n9736) );
  AOI21_X1 U10898 ( .B1(n9846), .B2(n9734), .A(n9733), .ZN(n9735) );
  OAI211_X1 U10899 ( .C1(n9737), .C2(n9860), .A(n9736), .B(n9735), .ZN(n9738)
         );
  INV_X1 U10900 ( .A(n9738), .ZN(n9744) );
  OAI21_X1 U10901 ( .B1(n9741), .B2(n9740), .A(n9739), .ZN(n9742) );
  NAND2_X1 U10902 ( .A1(n9742), .A2(n9855), .ZN(n9743) );
  OAI211_X1 U10903 ( .C1(n10129), .C2(n9745), .A(n9744), .B(n9743), .ZN(
        P2_U3191) );
  AOI22_X1 U10904 ( .A1(n9746), .A2(n9846), .B1(n9845), .B2(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n9763) );
  OAI21_X1 U10905 ( .B1(n9749), .B2(n9748), .A(n9747), .ZN(n9754) );
  OAI21_X1 U10906 ( .B1(n9752), .B2(n9751), .A(n9750), .ZN(n9753) );
  AOI22_X1 U10907 ( .A1(n9754), .A2(n9856), .B1(n9855), .B2(n9753), .ZN(n9762)
         );
  INV_X1 U10908 ( .A(n9755), .ZN(n9761) );
  AOI21_X1 U10909 ( .B1(n9758), .B2(n9757), .A(n9756), .ZN(n9759) );
  OR2_X1 U10910 ( .A1(n9759), .A2(n9860), .ZN(n9760) );
  NAND4_X1 U10911 ( .A1(n9763), .A2(n9762), .A3(n9761), .A4(n9760), .ZN(
        P2_U3192) );
  AOI22_X1 U10912 ( .A1(n9845), .A2(P2_ADDR_REG_11__SCAN_IN), .B1(n9764), .B2(
        n9846), .ZN(n9777) );
  OAI21_X1 U10913 ( .B1(n9766), .B2(P2_REG1_REG_11__SCAN_IN), .A(n9765), .ZN(
        n9771) );
  OAI21_X1 U10914 ( .B1(n9769), .B2(n9768), .A(n9767), .ZN(n9770) );
  AOI22_X1 U10915 ( .A1(n9771), .A2(n9856), .B1(n9855), .B2(n9770), .ZN(n9776)
         );
  NAND2_X1 U10916 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9942) );
  AOI21_X1 U10917 ( .B1(n5277), .B2(n9773), .A(n9772), .ZN(n9774) );
  OR2_X1 U10918 ( .A1(n9860), .A2(n9774), .ZN(n9775) );
  NAND4_X1 U10919 ( .A1(n9777), .A2(n9776), .A3(n9942), .A4(n9775), .ZN(
        P2_U3193) );
  AOI22_X1 U10920 ( .A1(n9778), .A2(n9846), .B1(n9845), .B2(
        P2_ADDR_REG_12__SCAN_IN), .ZN(n9794) );
  OAI21_X1 U10921 ( .B1(n9781), .B2(n9780), .A(n9779), .ZN(n9786) );
  OAI21_X1 U10922 ( .B1(n9784), .B2(n9783), .A(n9782), .ZN(n9785) );
  AOI22_X1 U10923 ( .A1(n9786), .A2(n9856), .B1(n9855), .B2(n9785), .ZN(n9793)
         );
  INV_X1 U10924 ( .A(n9787), .ZN(n9792) );
  AOI21_X1 U10925 ( .B1(n4349), .B2(n9789), .A(n9788), .ZN(n9790) );
  OR2_X1 U10926 ( .A1(n9860), .A2(n9790), .ZN(n9791) );
  NAND4_X1 U10927 ( .A1(n9794), .A2(n9793), .A3(n9792), .A4(n9791), .ZN(
        P2_U3194) );
  AOI22_X1 U10928 ( .A1(n9795), .A2(n9846), .B1(n9845), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n9811) );
  OAI21_X1 U10929 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n9797), .A(n9796), .ZN(
        n9802) );
  OAI21_X1 U10930 ( .B1(n9800), .B2(n9799), .A(n9798), .ZN(n9801) );
  AOI22_X1 U10931 ( .A1(n9802), .A2(n9856), .B1(n9855), .B2(n9801), .ZN(n9810)
         );
  INV_X1 U10932 ( .A(n9803), .ZN(n9804) );
  NOR2_X1 U10933 ( .A1(n9804), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9806) );
  OAI21_X1 U10934 ( .B1(n9807), .B2(n9806), .A(n9805), .ZN(n9808) );
  NAND4_X1 U10935 ( .A1(n9811), .A2(n9810), .A3(n9809), .A4(n9808), .ZN(
        P2_U3195) );
  AOI22_X1 U10936 ( .A1(n9812), .A2(n9846), .B1(n9845), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n9829) );
  OAI21_X1 U10937 ( .B1(n9815), .B2(n9814), .A(n9813), .ZN(n9820) );
  OAI21_X1 U10938 ( .B1(n9818), .B2(n9817), .A(n9816), .ZN(n9819) );
  AOI22_X1 U10939 ( .A1(n9820), .A2(n9856), .B1(n9855), .B2(n9819), .ZN(n9828)
         );
  INV_X1 U10940 ( .A(n9821), .ZN(n9827) );
  AOI21_X1 U10941 ( .B1(n9824), .B2(n9823), .A(n9822), .ZN(n9825) );
  OR2_X1 U10942 ( .A1(n9825), .A2(n9860), .ZN(n9826) );
  NAND4_X1 U10943 ( .A1(n9829), .A2(n9828), .A3(n9827), .A4(n9826), .ZN(
        P2_U3196) );
  AOI22_X1 U10944 ( .A1(n9830), .A2(n9846), .B1(n9845), .B2(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n9844) );
  OAI21_X1 U10945 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n9832), .A(n9831), .ZN(
        n9837) );
  OAI21_X1 U10946 ( .B1(n9835), .B2(n9834), .A(n9833), .ZN(n9836) );
  AOI22_X1 U10947 ( .A1(n9837), .A2(n9856), .B1(n9855), .B2(n9836), .ZN(n9843)
         );
  AOI21_X1 U10948 ( .B1(n9839), .B2(n7525), .A(n9838), .ZN(n9840) );
  OR2_X1 U10949 ( .A1(n9860), .A2(n9840), .ZN(n9841) );
  NAND4_X1 U10950 ( .A1(n9844), .A2(n9843), .A3(n9842), .A4(n9841), .ZN(
        P2_U3197) );
  AOI22_X1 U10951 ( .A1(n9847), .A2(n9846), .B1(n9845), .B2(
        P2_ADDR_REG_16__SCAN_IN), .ZN(n9865) );
  OAI21_X1 U10952 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(n9857) );
  OAI21_X1 U10953 ( .B1(n9853), .B2(n9852), .A(n9851), .ZN(n9854) );
  AOI22_X1 U10954 ( .A1(n9857), .A2(n9856), .B1(n9855), .B2(n9854), .ZN(n9864)
         );
  NAND2_X1 U10955 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3151), .ZN(n9863) );
  AOI21_X1 U10956 ( .B1(n4379), .B2(n9859), .A(n9858), .ZN(n9861) );
  OR2_X1 U10957 ( .A1(n9861), .A2(n9860), .ZN(n9862) );
  NAND4_X1 U10958 ( .A1(n9865), .A2(n9864), .A3(n9863), .A4(n9862), .ZN(
        P2_U3198) );
  INV_X1 U10959 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9868) );
  OAI22_X1 U10960 ( .A1(n9869), .A2(n9868), .B1(n9867), .B2(n9866), .ZN(n9872)
         );
  INV_X1 U10961 ( .A(n9870), .ZN(n9871) );
  AOI211_X1 U10962 ( .C1(n9874), .C2(n9873), .A(n9872), .B(n9871), .ZN(n9875)
         );
  AOI22_X1 U10963 ( .A1(n9876), .A2(n6584), .B1(n9875), .B2(n8693), .ZN(
        P2_U3231) );
  INV_X1 U10964 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9877) );
  AOI22_X1 U10965 ( .A1(n9901), .A2(n9878), .B1(n9877), .B2(n9898), .ZN(
        P2_U3390) );
  AOI22_X1 U10966 ( .A1(n9901), .A2(n9879), .B1(n5098), .B2(n9898), .ZN(
        P2_U3393) );
  INV_X1 U10967 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9880) );
  AOI22_X1 U10968 ( .A1(n9901), .A2(n9881), .B1(n9880), .B2(n9898), .ZN(
        P2_U3396) );
  AOI22_X1 U10969 ( .A1(n9901), .A2(n9882), .B1(n5136), .B2(n9898), .ZN(
        P2_U3399) );
  INV_X1 U10970 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9883) );
  AOI22_X1 U10971 ( .A1(n9901), .A2(n9884), .B1(n9883), .B2(n9898), .ZN(
        P2_U3402) );
  INV_X1 U10972 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9885) );
  AOI22_X1 U10973 ( .A1(n9901), .A2(n9886), .B1(n9885), .B2(n9898), .ZN(
        P2_U3405) );
  INV_X1 U10974 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9887) );
  AOI22_X1 U10975 ( .A1(n9901), .A2(n9888), .B1(n9887), .B2(n9898), .ZN(
        P2_U3408) );
  INV_X1 U10976 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U10977 ( .A1(n9901), .A2(n9890), .B1(n9889), .B2(n9898), .ZN(
        P2_U3411) );
  INV_X1 U10978 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9962) );
  AOI22_X1 U10979 ( .A1(n9901), .A2(n9891), .B1(n9962), .B2(n9898), .ZN(
        P2_U3414) );
  INV_X1 U10980 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9892) );
  AOI22_X1 U10981 ( .A1(n9901), .A2(n9893), .B1(n9892), .B2(n9898), .ZN(
        P2_U3417) );
  INV_X1 U10982 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9894) );
  AOI22_X1 U10983 ( .A1(n9901), .A2(n9895), .B1(n9894), .B2(n9898), .ZN(
        P2_U3420) );
  INV_X1 U10984 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9896) );
  AOI22_X1 U10985 ( .A1(n9901), .A2(n9897), .B1(n9896), .B2(n9898), .ZN(
        P2_U3423) );
  INV_X1 U10986 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9899) );
  AOI22_X1 U10987 ( .A1(n9901), .A2(n9900), .B1(n9899), .B2(n9898), .ZN(
        P2_U3426) );
  INV_X1 U10988 ( .A(n9902), .ZN(n9903) );
  NAND2_X1 U10989 ( .A1(n9904), .A2(n9903), .ZN(n9905) );
  XNOR2_X1 U10990 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9905), .ZN(ADD_1068_U5) );
  XOR2_X1 U10991 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U10992 ( .B1(n9908), .B2(n9907), .A(n9906), .ZN(n9909) );
  XOR2_X1 U10993 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n9909), .Z(ADD_1068_U55) );
  OAI21_X1 U10994 ( .B1(n9912), .B2(n9911), .A(n9910), .ZN(ADD_1068_U56) );
  OAI21_X1 U10995 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(ADD_1068_U57) );
  OAI21_X1 U10996 ( .B1(n9918), .B2(n9917), .A(n9916), .ZN(ADD_1068_U58) );
  OAI21_X1 U10997 ( .B1(n9921), .B2(n9920), .A(n9919), .ZN(ADD_1068_U59) );
  OAI21_X1 U10998 ( .B1(n9924), .B2(n9923), .A(n9922), .ZN(ADD_1068_U60) );
  OAI21_X1 U10999 ( .B1(n9927), .B2(n9926), .A(n9925), .ZN(ADD_1068_U61) );
  NAND2_X1 U11000 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9928) );
  NAND2_X1 U11001 ( .A1(n9929), .A2(n9928), .ZN(n9931) );
  XNOR2_X1 U11002 ( .A(n9931), .B(n9930), .ZN(ADD_1068_U62) );
  INV_X1 U11003 ( .A(n9932), .ZN(n9934) );
  NOR2_X1 U11004 ( .A1(n9934), .A2(n9933), .ZN(n9935) );
  XNOR2_X1 U11005 ( .A(n9936), .B(n9935), .ZN(ADD_1068_U63) );
  OAI22_X1 U11006 ( .A1(n9938), .A2(n9937), .B1(n8306), .B2(n9944), .ZN(n9941)
         );
  XNOR2_X1 U11007 ( .A(n9939), .B(n4441), .ZN(n9940) );
  XNOR2_X1 U11008 ( .A(n9941), .B(n9940), .ZN(n9959) );
  INV_X1 U11009 ( .A(n9942), .ZN(n9943) );
  AOI21_X1 U11010 ( .B1(n9945), .B2(n9944), .A(n9943), .ZN(n9956) );
  INV_X1 U11011 ( .A(n9946), .ZN(n9947) );
  NAND2_X1 U11012 ( .A1(n9948), .A2(n9947), .ZN(n9955) );
  NAND2_X1 U11013 ( .A1(n9950), .A2(n9949), .ZN(n9954) );
  NAND2_X1 U11014 ( .A1(n9952), .A2(n9951), .ZN(n9953) );
  NAND4_X1 U11015 ( .A1(n9956), .A2(n9955), .A3(n9954), .A4(n9953), .ZN(n9957)
         );
  AOI21_X1 U11016 ( .B1(n9959), .B2(n9958), .A(n9957), .ZN(n9960) );
  INV_X1 U11017 ( .A(n9960), .ZN(n10121) );
  AOI22_X1 U11018 ( .A1(n9962), .A2(keyinput25), .B1(n5273), .B2(keyinput7), 
        .ZN(n9961) );
  OAI221_X1 U11019 ( .B1(n9962), .B2(keyinput25), .C1(n5273), .C2(keyinput7), 
        .A(n9961), .ZN(n9963) );
  INV_X1 U11020 ( .A(n9963), .ZN(n9979) );
  INV_X1 U11021 ( .A(keyinput44), .ZN(n9965) );
  AOI22_X1 U11022 ( .A1(n9966), .A2(keyinput40), .B1(P1_ADDR_REG_18__SCAN_IN), 
        .B2(n9965), .ZN(n9964) );
  OAI221_X1 U11023 ( .B1(n9966), .B2(keyinput40), .C1(n9965), .C2(
        P1_ADDR_REG_18__SCAN_IN), .A(n9964), .ZN(n9967) );
  INV_X1 U11024 ( .A(n9967), .ZN(n9978) );
  INV_X1 U11025 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9970) );
  AOI22_X1 U11026 ( .A1(n9970), .A2(keyinput2), .B1(n9969), .B2(keyinput20), 
        .ZN(n9968) );
  OAI221_X1 U11027 ( .B1(n9970), .B2(keyinput2), .C1(n9969), .C2(keyinput20), 
        .A(n9968), .ZN(n9973) );
  XNOR2_X1 U11028 ( .A(n9971), .B(keyinput18), .ZN(n9972) );
  NOR2_X1 U11029 ( .A1(n9973), .A2(n9972), .ZN(n9977) );
  INV_X1 U11030 ( .A(keyinput56), .ZN(n9975) );
  XNOR2_X1 U11031 ( .A(n9975), .B(n9974), .ZN(n9976) );
  AND4_X1 U11032 ( .A1(n9979), .A2(n9978), .A3(n9977), .A4(n9976), .ZN(n10119)
         );
  INV_X1 U11033 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9982) );
  AOI22_X1 U11034 ( .A1(n9982), .A2(keyinput6), .B1(keyinput62), .B2(n9981), 
        .ZN(n9980) );
  OAI221_X1 U11035 ( .B1(n9982), .B2(keyinput6), .C1(n9981), .C2(keyinput62), 
        .A(n9980), .ZN(n9993) );
  AOI22_X1 U11036 ( .A1(n6487), .A2(keyinput50), .B1(n9984), .B2(keyinput1), 
        .ZN(n9983) );
  OAI221_X1 U11037 ( .B1(n6487), .B2(keyinput50), .C1(n9984), .C2(keyinput1), 
        .A(n9983), .ZN(n9992) );
  AOI22_X1 U11038 ( .A1(n9987), .A2(keyinput52), .B1(n9986), .B2(keyinput26), 
        .ZN(n9985) );
  OAI221_X1 U11039 ( .B1(n9987), .B2(keyinput52), .C1(n9986), .C2(keyinput26), 
        .A(n9985), .ZN(n9991) );
  XNOR2_X1 U11040 ( .A(P2_REG1_REG_1__SCAN_IN), .B(keyinput4), .ZN(n9989) );
  XNOR2_X1 U11041 ( .A(P1_REG3_REG_9__SCAN_IN), .B(keyinput36), .ZN(n9988) );
  NAND2_X1 U11042 ( .A1(n9989), .A2(n9988), .ZN(n9990) );
  NOR4_X1 U11043 ( .A1(n9993), .A2(n9992), .A3(n9991), .A4(n9990), .ZN(n10118)
         );
  OAI22_X1 U11044 ( .A1(n9996), .A2(keyinput51), .B1(n9995), .B2(keyinput39), 
        .ZN(n9994) );
  AOI221_X1 U11045 ( .B1(n9996), .B2(keyinput51), .C1(keyinput39), .C2(n9995), 
        .A(n9994), .ZN(n10008) );
  INV_X1 U11046 ( .A(keyinput30), .ZN(n9998) );
  OAI22_X1 U11047 ( .A1(n5617), .A2(keyinput27), .B1(n9998), .B2(
        P2_ADDR_REG_1__SCAN_IN), .ZN(n9997) );
  AOI221_X1 U11048 ( .B1(n5617), .B2(keyinput27), .C1(P2_ADDR_REG_1__SCAN_IN), 
        .C2(n9998), .A(n9997), .ZN(n10007) );
  INV_X1 U11049 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10001) );
  INV_X1 U11050 ( .A(keyinput8), .ZN(n10000) );
  OAI22_X1 U11051 ( .A1(n10001), .A2(keyinput31), .B1(n10000), .B2(
        P1_ADDR_REG_8__SCAN_IN), .ZN(n9999) );
  AOI221_X1 U11052 ( .B1(n10001), .B2(keyinput31), .C1(P1_ADDR_REG_8__SCAN_IN), 
        .C2(n10000), .A(n9999), .ZN(n10006) );
  OAI22_X1 U11053 ( .A1(n10004), .A2(keyinput37), .B1(n10003), .B2(keyinput58), 
        .ZN(n10002) );
  AOI221_X1 U11054 ( .B1(n10004), .B2(keyinput37), .C1(keyinput58), .C2(n10003), .A(n10002), .ZN(n10005) );
  NAND4_X1 U11055 ( .A1(n10008), .A2(n10007), .A3(n10006), .A4(n10005), .ZN(
        n10085) );
  INV_X1 U11056 ( .A(keyinput12), .ZN(n10010) );
  OAI22_X1 U11057 ( .A1(n10011), .A2(keyinput61), .B1(n10010), .B2(
        P1_ADDR_REG_5__SCAN_IN), .ZN(n10009) );
  AOI221_X1 U11058 ( .B1(n10011), .B2(keyinput61), .C1(P1_ADDR_REG_5__SCAN_IN), 
        .C2(n10010), .A(n10009), .ZN(n10024) );
  INV_X1 U11059 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10013) );
  OAI22_X1 U11060 ( .A1(n9213), .A2(keyinput35), .B1(n10013), .B2(keyinput5), 
        .ZN(n10012) );
  AOI221_X1 U11061 ( .B1(n9213), .B2(keyinput35), .C1(keyinput5), .C2(n10013), 
        .A(n10012), .ZN(n10023) );
  INV_X1 U11062 ( .A(keyinput24), .ZN(n10015) );
  OAI22_X1 U11063 ( .A1(keyinput63), .A2(n10016), .B1(n10015), .B2(
        P2_ADDR_REG_4__SCAN_IN), .ZN(n10014) );
  AOI221_X1 U11064 ( .B1(n10016), .B2(keyinput63), .C1(n10015), .C2(
        P2_ADDR_REG_4__SCAN_IN), .A(n10014), .ZN(n10022) );
  XNOR2_X1 U11065 ( .A(n10017), .B(keyinput16), .ZN(n10020) );
  XNOR2_X1 U11066 ( .A(n10018), .B(keyinput34), .ZN(n10019) );
  NOR2_X1 U11067 ( .A1(n10020), .A2(n10019), .ZN(n10021) );
  NAND4_X1 U11068 ( .A1(n10024), .A2(n10023), .A3(n10022), .A4(n10021), .ZN(
        n10084) );
  AOI22_X1 U11069 ( .A1(n10027), .A2(keyinput49), .B1(keyinput59), .B2(n10026), 
        .ZN(n10025) );
  OAI221_X1 U11070 ( .B1(n10027), .B2(keyinput49), .C1(n10026), .C2(keyinput59), .A(n10025), .ZN(n10038) );
  AOI22_X1 U11071 ( .A1(n10029), .A2(keyinput32), .B1(n8683), .B2(keyinput14), 
        .ZN(n10028) );
  OAI221_X1 U11072 ( .B1(n10029), .B2(keyinput32), .C1(n8683), .C2(keyinput14), 
        .A(n10028), .ZN(n10037) );
  INV_X1 U11073 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10031) );
  AOI22_X1 U11074 ( .A1(n10032), .A2(keyinput21), .B1(keyinput41), .B2(n10031), 
        .ZN(n10030) );
  OAI221_X1 U11075 ( .B1(n10032), .B2(keyinput21), .C1(n10031), .C2(keyinput41), .A(n10030), .ZN(n10036) );
  XOR2_X1 U11076 ( .A(n7627), .B(keyinput55), .Z(n10034) );
  XNOR2_X1 U11077 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput47), .ZN(n10033) );
  NAND2_X1 U11078 ( .A1(n10034), .A2(n10033), .ZN(n10035) );
  NOR4_X1 U11079 ( .A1(n10038), .A2(n10037), .A3(n10036), .A4(n10035), .ZN(
        n10082) );
  INV_X1 U11080 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10041) );
  AOI22_X1 U11081 ( .A1(n10041), .A2(keyinput45), .B1(n10040), .B2(keyinput60), 
        .ZN(n10039) );
  OAI221_X1 U11082 ( .B1(n10041), .B2(keyinput45), .C1(n10040), .C2(keyinput60), .A(n10039), .ZN(n10050) );
  XNOR2_X1 U11083 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput38), .ZN(n10046) );
  XNOR2_X1 U11084 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput0), .ZN(n10045) );
  XNOR2_X1 U11085 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput10), .ZN(n10044)
         );
  XNOR2_X1 U11086 ( .A(keyinput3), .B(P1_REG0_REG_3__SCAN_IN), .ZN(n10043) );
  NAND4_X1 U11087 ( .A1(n10046), .A2(n10045), .A3(n10044), .A4(n10043), .ZN(
        n10049) );
  XNOR2_X1 U11088 ( .A(keyinput15), .B(n8705), .ZN(n10048) );
  XNOR2_X1 U11089 ( .A(keyinput48), .B(n5410), .ZN(n10047) );
  NOR4_X1 U11090 ( .A1(n10050), .A2(n10049), .A3(n10048), .A4(n10047), .ZN(
        n10081) );
  INV_X1 U11091 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10053) );
  AOI22_X1 U11092 ( .A1(n10053), .A2(keyinput46), .B1(n10052), .B2(keyinput11), 
        .ZN(n10051) );
  OAI221_X1 U11093 ( .B1(n10053), .B2(keyinput46), .C1(n10052), .C2(keyinput11), .A(n10051), .ZN(n10060) );
  XNOR2_X1 U11094 ( .A(n10054), .B(keyinput33), .ZN(n10059) );
  XNOR2_X1 U11095 ( .A(n10055), .B(keyinput57), .ZN(n10058) );
  XNOR2_X1 U11096 ( .A(n10056), .B(keyinput23), .ZN(n10057) );
  OR4_X1 U11097 ( .A1(n10060), .A2(n10059), .A3(n10058), .A4(n10057), .ZN(
        n10066) );
  AOI22_X1 U11098 ( .A1(n10062), .A2(keyinput19), .B1(keyinput9), .B2(n5665), 
        .ZN(n10061) );
  OAI221_X1 U11099 ( .B1(n10062), .B2(keyinput19), .C1(n5665), .C2(keyinput9), 
        .A(n10061), .ZN(n10065) );
  XNOR2_X1 U11100 ( .A(n10063), .B(keyinput29), .ZN(n10064) );
  NOR3_X1 U11101 ( .A1(n10066), .A2(n10065), .A3(n10064), .ZN(n10080) );
  AOI22_X1 U11102 ( .A1(n10068), .A2(keyinput17), .B1(keyinput53), .B2(n8774), 
        .ZN(n10067) );
  OAI221_X1 U11103 ( .B1(n10068), .B2(keyinput17), .C1(n8774), .C2(keyinput53), 
        .A(n10067), .ZN(n10078) );
  AOI22_X1 U11104 ( .A1(n10071), .A2(keyinput28), .B1(keyinput42), .B2(n10070), 
        .ZN(n10069) );
  OAI221_X1 U11105 ( .B1(n10071), .B2(keyinput28), .C1(n10070), .C2(keyinput42), .A(n10069), .ZN(n10077) );
  XNOR2_X1 U11106 ( .A(SI_23_), .B(keyinput13), .ZN(n10075) );
  XNOR2_X1 U11107 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput22), .ZN(n10074)
         );
  XNOR2_X1 U11108 ( .A(SI_1_), .B(keyinput43), .ZN(n10073) );
  XNOR2_X1 U11109 ( .A(keyinput54), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n10072) );
  NAND4_X1 U11110 ( .A1(n10075), .A2(n10074), .A3(n10073), .A4(n10072), .ZN(
        n10076) );
  NOR3_X1 U11111 ( .A1(n10078), .A2(n10077), .A3(n10076), .ZN(n10079) );
  NAND4_X1 U11112 ( .A1(n10082), .A2(n10081), .A3(n10080), .A4(n10079), .ZN(
        n10083) );
  NOR3_X1 U11113 ( .A1(n10085), .A2(n10084), .A3(n10083), .ZN(n10117) );
  NAND3_X1 U11114 ( .A1(keyinput55), .A2(keyinput21), .A3(keyinput41), .ZN(
        n10091) );
  NOR2_X1 U11115 ( .A1(keyinput10), .A2(keyinput3), .ZN(n10086) );
  NAND3_X1 U11116 ( .A1(keyinput38), .A2(keyinput48), .A3(n10086), .ZN(n10090)
         );
  NOR3_X1 U11117 ( .A1(keyinput14), .A2(keyinput49), .A3(keyinput59), .ZN(
        n10088) );
  NOR3_X1 U11118 ( .A1(keyinput45), .A2(keyinput60), .A3(keyinput15), .ZN(
        n10087) );
  NAND4_X1 U11119 ( .A1(keyinput32), .A2(n10088), .A3(keyinput0), .A4(n10087), 
        .ZN(n10089) );
  NOR4_X1 U11120 ( .A1(keyinput47), .A2(n10091), .A3(n10090), .A4(n10089), 
        .ZN(n10115) );
  NAND2_X1 U11121 ( .A1(keyinput19), .A2(keyinput9), .ZN(n10098) );
  NOR2_X1 U11122 ( .A1(keyinput28), .A2(keyinput42), .ZN(n10096) );
  NAND3_X1 U11123 ( .A1(keyinput23), .A2(keyinput46), .A3(keyinput11), .ZN(
        n10094) );
  INV_X1 U11124 ( .A(keyinput54), .ZN(n10092) );
  NAND3_X1 U11125 ( .A1(keyinput13), .A2(keyinput22), .A3(n10092), .ZN(n10093)
         );
  NOR4_X1 U11126 ( .A1(keyinput29), .A2(keyinput43), .A3(n10094), .A4(n10093), 
        .ZN(n10095) );
  NAND4_X1 U11127 ( .A1(keyinput17), .A2(keyinput53), .A3(n10096), .A4(n10095), 
        .ZN(n10097) );
  NOR4_X1 U11128 ( .A1(keyinput33), .A2(keyinput57), .A3(n10098), .A4(n10097), 
        .ZN(n10114) );
  NAND2_X1 U11129 ( .A1(keyinput61), .A2(keyinput35), .ZN(n10105) );
  NOR2_X1 U11130 ( .A1(keyinput27), .A2(keyinput51), .ZN(n10103) );
  NAND3_X1 U11131 ( .A1(keyinput63), .A2(keyinput16), .A3(keyinput34), .ZN(
        n10101) );
  INV_X1 U11132 ( .A(keyinput31), .ZN(n10099) );
  NAND3_X1 U11133 ( .A1(keyinput58), .A2(keyinput8), .A3(n10099), .ZN(n10100)
         );
  NOR4_X1 U11134 ( .A1(keyinput24), .A2(keyinput37), .A3(n10101), .A4(n10100), 
        .ZN(n10102) );
  NAND4_X1 U11135 ( .A1(keyinput30), .A2(keyinput39), .A3(n10103), .A4(n10102), 
        .ZN(n10104) );
  NOR4_X1 U11136 ( .A1(keyinput12), .A2(keyinput5), .A3(n10105), .A4(n10104), 
        .ZN(n10113) );
  NOR2_X1 U11137 ( .A1(keyinput2), .A2(keyinput44), .ZN(n10106) );
  NAND3_X1 U11138 ( .A1(keyinput20), .A2(keyinput40), .A3(n10106), .ZN(n10111)
         );
  NAND3_X1 U11139 ( .A1(keyinput7), .A2(keyinput18), .A3(keyinput56), .ZN(
        n10110) );
  NOR3_X1 U11140 ( .A1(keyinput50), .A2(keyinput1), .A3(keyinput52), .ZN(
        n10108) );
  NOR3_X1 U11141 ( .A1(keyinput36), .A2(keyinput4), .A3(keyinput6), .ZN(n10107) );
  NAND4_X1 U11142 ( .A1(keyinput26), .A2(n10108), .A3(keyinput62), .A4(n10107), 
        .ZN(n10109) );
  NOR4_X1 U11143 ( .A1(keyinput25), .A2(n10111), .A3(n10110), .A4(n10109), 
        .ZN(n10112) );
  NAND4_X1 U11144 ( .A1(n10115), .A2(n10114), .A3(n10113), .A4(n10112), .ZN(
        n10116) );
  NAND4_X1 U11145 ( .A1(n10119), .A2(n10118), .A3(n10117), .A4(n10116), .ZN(
        n10120) );
  XNOR2_X1 U11146 ( .A(n10121), .B(n10120), .ZN(P2_U3176) );
  XOR2_X1 U11147 ( .A(n10122), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1068_U50) );
  NOR2_X1 U11148 ( .A1(n10124), .A2(n10123), .ZN(n10126) );
  XNOR2_X1 U11149 ( .A(n10126), .B(n10125), .ZN(ADD_1068_U51) );
  AOI21_X1 U11150 ( .B1(n10129), .B2(n10128), .A(n10127), .ZN(ADD_1068_U47) );
  XOR2_X1 U11151 ( .A(n10130), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1068_U49) );
  XOR2_X1 U11152 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10131), .Z(ADD_1068_U48) );
  XOR2_X1 U11153 ( .A(n10133), .B(n10132), .Z(ADD_1068_U54) );
  XOR2_X1 U11154 ( .A(n10135), .B(n10134), .Z(ADD_1068_U53) );
  XNOR2_X1 U11155 ( .A(n10137), .B(n10136), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4854 ( .A(n5807), .Z(n6180) );
  CLKBUF_X1 U4861 ( .A(n6177), .Z(n4323) );
  CLKBUF_X1 U7387 ( .A(n5988), .Z(n4331) );
endmodule

