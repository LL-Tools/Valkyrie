

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938;

  INV_X1 U2374 ( .A(n2952), .ZN(n2803) );
  INV_X2 U2375 ( .A(n2905), .ZN(n2954) );
  INV_X1 U2376 ( .A(n2992), .ZN(n2976) );
  INV_X1 U2377 ( .A(n3909), .ZN(n2431) );
  AND2_X1 U2378 ( .A1(n3839), .A2(n3842), .ZN(n3813) );
  NAND2_X1 U2379 ( .A1(n3037), .A2(IR_REG_31__SCAN_IN), .ZN(n2329) );
  OAI211_X1 U2380 ( .C1(n2158), .C2(n4275), .A(n2675), .B(n2674), .ZN(n4018)
         );
  AND2_X1 U2381 ( .A1(n3180), .A2(n3890), .ZN(n4610) );
  AND2_X2 U2382 ( .A1(n2335), .A2(n4428), .ZN(n2363) );
  XNOR2_X1 U2383 ( .A(n2329), .B(n3038), .ZN(n2335) );
  NOR2_X2 U2384 ( .A1(n3560), .A2(n3559), .ZN(n3561) );
  NAND2_X2 U2385 ( .A1(n3833), .A2(n3836), .ZN(n3242) );
  INV_X4 U2386 ( .A(n2954), .ZN(n2988) );
  NAND4_X1 U2387 ( .A1(n2384), .A2(n2383), .A3(n2382), .A4(n2381), .ZN(n3911)
         );
  CLKBUF_X2 U2388 ( .A(n2346), .Z(n2438) );
  BUF_X4 U2389 ( .A(n2416), .Z(n2132) );
  NOR2_X1 U2390 ( .A1(n4307), .A2(n4306), .ZN(n4308) );
  AOI211_X1 U2391 ( .C1(n4230), .C2(n4007), .A(n3565), .B(n3564), .ZN(n4316)
         );
  NAND2_X1 U2392 ( .A1(n2857), .A2(n2856), .ZN(n3734) );
  OAI21_X1 U2393 ( .B1(n2186), .B2(n2185), .A(n2183), .ZN(n4005) );
  INV_X1 U2394 ( .A(n4027), .ZN(n2186) );
  AOI211_X1 U2395 ( .C1(n4247), .C2(n4250), .A(n4275), .B(n4249), .ZN(n4251)
         );
  NAND2_X1 U2396 ( .A1(n4107), .A2(n4106), .ZN(n4105) );
  NAND2_X1 U2397 ( .A1(n2642), .A2(n3854), .ZN(n3486) );
  NAND2_X1 U2398 ( .A1(n2641), .A2(n3847), .ZN(n3424) );
  NAND2_X1 U2399 ( .A1(n4220), .A2(n2524), .ZN(n4207) );
  NAND2_X1 U2400 ( .A1(n4222), .A2(n4221), .ZN(n4220) );
  NAND2_X1 U2401 ( .A1(n2638), .A2(n3844), .ZN(n3355) );
  INV_X1 U2402 ( .A(n2184), .ZN(n2183) );
  OAI21_X1 U2403 ( .B1(n2185), .B2(n2171), .A(n2617), .ZN(n2184) );
  NAND2_X1 U2404 ( .A1(n3256), .A2(n3838), .ZN(n3320) );
  NAND2_X1 U2405 ( .A1(n4007), .A2(n4006), .ZN(n4008) );
  NAND2_X1 U2406 ( .A1(n3257), .A2(n3815), .ZN(n3256) );
  AND2_X1 U2407 ( .A1(n2752), .A2(n2747), .ZN(n2295) );
  NAND2_X2 U2408 ( .A1(n3021), .A2(n4440), .ZN(n3738) );
  AND2_X1 U2409 ( .A1(n2639), .A2(n3848), .ZN(n3356) );
  AND2_X1 U2410 ( .A1(n3838), .A2(n3835), .ZN(n3815) );
  BUF_X1 U2411 ( .A(n2721), .Z(n2138) );
  OR2_X1 U2412 ( .A1(n3235), .A2(n3261), .ZN(n3838) );
  OR2_X1 U2413 ( .A1(n2730), .A2(n3250), .ZN(n3833) );
  NAND4_X1 U2414 ( .A1(n2395), .A2(n2394), .A3(n2393), .A4(n2392), .ZN(n3258)
         );
  NAND4_X1 U2415 ( .A1(n2425), .A2(n2424), .A3(n2423), .A4(n2422), .ZN(n3908)
         );
  NAND4_X1 U2416 ( .A1(n2367), .A2(n2366), .A3(n2365), .A4(n2364), .ZN(n3235)
         );
  OR2_X1 U2417 ( .A1(n2712), .A2(n3203), .ZN(n3832) );
  NAND4_X2 U2418 ( .A1(n2360), .A2(n2359), .A3(n2358), .A4(n2357), .ZN(n2730)
         );
  NAND4_X1 U2419 ( .A1(n2377), .A2(n2376), .A3(n2375), .A4(n2374), .ZN(n3910)
         );
  CLKBUF_X1 U2420 ( .A(n2139), .Z(n2670) );
  CLKBUF_X3 U2421 ( .A(n2438), .Z(n3756) );
  INV_X2 U2422 ( .A(n2418), .ZN(n2588) );
  MUX2_X1 U2423 ( .A(n3079), .B(n2361), .S(n2416), .Z(n3250) );
  NAND2_X2 U2424 ( .A1(n3012), .A2(n3215), .ZN(n2992) );
  INV_X1 U2425 ( .A(n2356), .ZN(n2418) );
  MUX2_X1 U2426 ( .A(n3076), .B(n2353), .S(n2416), .Z(n3203) );
  XNOR2_X1 U2427 ( .A(n2678), .B(n4881), .ZN(n3035) );
  NAND2_X1 U2428 ( .A1(n2677), .A2(IR_REG_31__SCAN_IN), .ZN(n2678) );
  AND2_X1 U2429 ( .A1(n2335), .A2(n2334), .ZN(n2356) );
  XNOR2_X1 U2430 ( .A(n2622), .B(IR_REG_22__SCAN_IN), .ZN(n4431) );
  XNOR2_X1 U2431 ( .A(n2332), .B(n2331), .ZN(n2334) );
  OR2_X1 U2432 ( .A1(n2676), .A2(n2679), .ZN(n2697) );
  OR2_X1 U2433 ( .A1(n2330), .A2(n2679), .ZN(n2332) );
  NOR2_X1 U2434 ( .A1(n2137), .A2(n2194), .ZN(n2330) );
  INV_X1 U2435 ( .A(n2194), .ZN(n2626) );
  NAND2_X1 U2436 ( .A1(n2157), .A2(n2262), .ZN(n2162) );
  NOR2_X1 U2437 ( .A1(n2257), .A2(IR_REG_18__SCAN_IN), .ZN(n2256) );
  NAND2_X1 U2438 ( .A1(n2297), .A2(n2258), .ZN(n2257) );
  AND2_X1 U2439 ( .A1(n2308), .A2(n2326), .ZN(n2297) );
  AND2_X1 U2440 ( .A1(n2306), .A2(n2327), .ZN(n2305) );
  AND2_X1 U2441 ( .A1(n4880), .A2(n4672), .ZN(n2306) );
  NOR2_X1 U2442 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2321)
         );
  INV_X1 U2443 ( .A(IR_REG_15__SCAN_IN), .ZN(n2510) );
  NOR2_X1 U2444 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2322)
         );
  NOR2_X1 U2445 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2323)
         );
  NOR2_X2 U2446 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n4890)
         );
  INV_X1 U2447 ( .A(IR_REG_16__SCAN_IN), .ZN(n4879) );
  INV_X1 U2448 ( .A(IR_REG_14__SCAN_IN), .ZN(n2326) );
  INV_X2 U2449 ( .A(IR_REG_3__SCAN_IN), .ZN(n2319) );
  INV_X1 U2450 ( .A(IR_REG_4__SCAN_IN), .ZN(n2398) );
  NOR2_X2 U2451 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2368)
         );
  NAND2_X1 U2452 ( .A1(n2653), .A2(n2136), .ZN(n2133) );
  AND2_X2 U2453 ( .A1(n2133), .A2(n2134), .ZN(n4083) );
  OR2_X1 U2454 ( .A1(n2135), .A2(n3867), .ZN(n2134) );
  INV_X1 U2455 ( .A(n3774), .ZN(n2135) );
  AND2_X1 U2456 ( .A1(n2652), .A2(n3774), .ZN(n2136) );
  OR2_X1 U2457 ( .A1(n4166), .A2(n3772), .ZN(n4142) );
  OR2_X1 U2458 ( .A1(n2164), .A2(n2162), .ZN(n2137) );
  OR2_X1 U2459 ( .A1(n2194), .A2(n2162), .ZN(n2343) );
  OAI21_X2 U2460 ( .B1(n3355), .B2(n2640), .A(n3848), .ZN(n3393) );
  NAND2_X1 U2461 ( .A1(n3245), .A2(n3833), .ZN(n3257) );
  NAND3_X2 U2462 ( .A1(n2195), .A2(n2256), .A3(n2148), .ZN(n2194) );
  AOI21_X1 U2463 ( .B1(n3197), .B2(n3821), .A(n2355), .ZN(n3240) );
  INV_X1 U2464 ( .A(n2334), .ZN(n4428) );
  NAND2_X1 U2465 ( .A1(n4427), .A2(n4428), .ZN(n2139) );
  NAND2_X1 U2466 ( .A1(n4427), .A2(n4428), .ZN(n2597) );
  OAI21_X2 U2467 ( .B1(n3320), .B2(n2632), .A(n3842), .ZN(n3335) );
  OAI21_X2 U2468 ( .B1(n3424), .B2(n3855), .A(n3852), .ZN(n3464) );
  NOR2_X1 U2469 ( .A1(n2335), .A2(n4428), .ZN(n2346) );
  INV_X1 U2470 ( .A(n2418), .ZN(n2140) );
  INV_X2 U2471 ( .A(n2418), .ZN(n2141) );
  NAND2_X1 U2472 ( .A1(n3588), .A2(n3583), .ZN(n2854) );
  OR2_X1 U2473 ( .A1(n2246), .A2(n3138), .ZN(n2245) );
  INV_X1 U2474 ( .A(n2404), .ZN(n2405) );
  NAND2_X1 U2475 ( .A1(n3890), .A2(n4432), .ZN(n3215) );
  INV_X1 U2476 ( .A(IR_REG_25__SCAN_IN), .ZN(n2681) );
  NAND3_X1 U2477 ( .A1(n4429), .A2(n3045), .A3(n4430), .ZN(n3028) );
  AND2_X1 U2478 ( .A1(n2284), .A2(n2283), .ZN(n3946) );
  NAND2_X1 U2479 ( .A1(n4435), .A2(REG1_REG_9__SCAN_IN), .ZN(n2283) );
  AND2_X1 U2480 ( .A1(n2220), .A2(n2219), .ZN(n4466) );
  INV_X1 U2481 ( .A(n4467), .ZN(n2219) );
  XNOR2_X1 U2482 ( .A(n3964), .B(n3963), .ZN(n4630) );
  OR2_X1 U2483 ( .A1(n2279), .A2(n3967), .ZN(n2205) );
  NAND2_X1 U2484 ( .A1(n2279), .A2(n2206), .ZN(n2203) );
  NOR2_X1 U2485 ( .A1(n2207), .A2(n4565), .ZN(n2206) );
  INV_X1 U2486 ( .A(n2278), .ZN(n2207) );
  NAND2_X1 U2487 ( .A1(n2281), .A2(n2280), .ZN(n2279) );
  INV_X1 U2488 ( .A(n4482), .ZN(n2280) );
  NOR2_X1 U2489 ( .A1(n2146), .A2(n2174), .ZN(n2289) );
  NAND2_X1 U2490 ( .A1(n2623), .A2(n2555), .ZN(n3985) );
  OR2_X1 U2491 ( .A1(n3939), .A2(n2168), .ZN(n2243) );
  INV_X1 U2492 ( .A(n3144), .ZN(n2216) );
  NOR2_X1 U2493 ( .A1(n2216), .A2(n2213), .ZN(n2212) );
  NAND2_X1 U2494 ( .A1(n2226), .A2(n2225), .ZN(n3968) );
  NAND2_X1 U2495 ( .A1(n4567), .A2(n4864), .ZN(n2225) );
  OR2_X1 U2496 ( .A1(n4479), .A2(n2317), .ZN(n2226) );
  INV_X1 U2497 ( .A(n4097), .ZN(n2927) );
  AND2_X1 U2498 ( .A1(n2149), .A2(n4214), .ZN(n2260) );
  NAND2_X1 U2499 ( .A1(n2637), .A2(n3361), .ZN(n2255) );
  INV_X1 U2500 ( .A(n4431), .ZN(n2672) );
  NOR2_X1 U2501 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2327)
         );
  INV_X1 U2502 ( .A(n3585), .ZN(n2844) );
  NAND2_X1 U2503 ( .A1(n3385), .A2(n3386), .ZN(n2294) );
  AND2_X1 U2504 ( .A1(n2292), .A2(n3724), .ZN(n2291) );
  INV_X1 U2505 ( .A(n3573), .ZN(n2292) );
  NAND2_X1 U2506 ( .A1(n3223), .A2(n3224), .ZN(n2296) );
  INV_X1 U2507 ( .A(n4432), .ZN(n3826) );
  NAND2_X1 U2508 ( .A1(n2363), .A2(REG1_REG_0__SCAN_IN), .ZN(n2336) );
  NAND3_X1 U2509 ( .A1(n2199), .A2(n3101), .A3(n2196), .ZN(n3102) );
  NAND2_X1 U2510 ( .A1(n2263), .A2(n2145), .ZN(n2199) );
  NAND2_X1 U2511 ( .A1(n2198), .A2(n2197), .ZN(n2196) );
  NAND2_X1 U2512 ( .A1(n3110), .A2(n3111), .ZN(n2246) );
  OR2_X1 U2513 ( .A1(n4450), .A2(n4451), .ZN(n2221) );
  NAND2_X1 U2514 ( .A1(n3957), .A2(n2173), .ZN(n3960) );
  OR2_X1 U2515 ( .A1(n4458), .A2(n3947), .ZN(n2220) );
  NAND2_X1 U2516 ( .A1(n4472), .A2(n3962), .ZN(n3964) );
  NAND2_X1 U2517 ( .A1(n4630), .A2(REG2_REG_12__SCAN_IN), .ZN(n4628) );
  OR2_X1 U2518 ( .A1(n4623), .A2(n3949), .ZN(n2281) );
  NAND2_X1 U2519 ( .A1(n4486), .A2(REG1_REG_13__SCAN_IN), .ZN(n2278) );
  NOR2_X1 U2520 ( .A1(n2209), .A2(n4491), .ZN(n2204) );
  OR2_X1 U2521 ( .A1(n4506), .A2(n4505), .ZN(n4503) );
  INV_X1 U2522 ( .A(n4440), .ZN(n3913) );
  NOR2_X1 U2523 ( .A1(n4564), .A2(n2240), .ZN(n2239) );
  INV_X1 U2524 ( .A(n3972), .ZN(n2240) );
  NAND2_X1 U2525 ( .A1(n2235), .A2(n3971), .ZN(n4500) );
  OAI211_X1 U2526 ( .C1(n2235), .C2(n2234), .A(n2231), .B(n2230), .ZN(n4513)
         );
  INV_X1 U2527 ( .A(n2237), .ZN(n2234) );
  AOI21_X1 U2528 ( .B1(n2237), .B2(n2233), .A(REG2_REG_16__SCAN_IN), .ZN(n2230) );
  NAND2_X1 U2529 ( .A1(n2235), .A2(n2232), .ZN(n2231) );
  AOI21_X1 U2530 ( .B1(n4124), .B2(n2572), .A(n2176), .ZN(n4107) );
  NAND2_X1 U2531 ( .A1(n4210), .A2(n2523), .ZN(n2524) );
  OR2_X1 U2532 ( .A1(n4253), .A2(n3593), .ZN(n2502) );
  OR2_X1 U2533 ( .A1(n3907), .A2(n3425), .ZN(n2189) );
  NAND2_X1 U2534 ( .A1(n2436), .A2(n2159), .ZN(n2191) );
  INV_X1 U2535 ( .A(n3403), .ZN(n2705) );
  AND2_X1 U2536 ( .A1(n2712), .A2(n2354), .ZN(n2355) );
  AND2_X1 U2537 ( .A1(n4440), .A2(n3050), .ZN(n4272) );
  NAND2_X1 U2538 ( .A1(n2628), .A2(n3985), .ZN(n4153) );
  INV_X1 U2539 ( .A(n2721), .ZN(n2629) );
  OR2_X1 U2540 ( .A1(n4440), .A2(n2985), .ZN(n4268) );
  NAND2_X1 U2541 ( .A1(n2686), .A2(n4429), .ZN(n3044) );
  NAND2_X1 U2542 ( .A1(n2343), .A2(n2342), .ZN(n3041) );
  AND2_X1 U2543 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2342)
         );
  NOR2_X1 U2544 ( .A1(n2499), .A2(n2257), .ZN(n2540) );
  OR3_X1 U2545 ( .A1(n2445), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2448) );
  NOR2_X1 U2546 ( .A1(n2448), .A2(IR_REG_9__SCAN_IN), .ZN(n2464) );
  INV_X1 U2547 ( .A(n2291), .ZN(n2290) );
  AND2_X1 U2548 ( .A1(n3006), .A2(n2987), .ZN(n3716) );
  AND2_X1 U2549 ( .A1(n3058), .A2(n3057), .ZN(n3075) );
  NOR2_X1 U2550 ( .A1(n4459), .A2(n4878), .ZN(n4458) );
  XNOR2_X1 U2551 ( .A(n3960), .B(n2282), .ZN(n4463) );
  NAND2_X1 U2552 ( .A1(n4463), .A2(REG2_REG_10__SCAN_IN), .ZN(n4462) );
  NAND2_X1 U2553 ( .A1(n4525), .A2(n2274), .ZN(n4534) );
  AOI21_X1 U2554 ( .B1(n4525), .B2(n2270), .A(n4622), .ZN(n2223) );
  NAND2_X1 U2555 ( .A1(n2249), .A2(n2248), .ZN(n3982) );
  OR2_X1 U2556 ( .A1(n2153), .A2(n3979), .ZN(n2248) );
  NAND2_X1 U2557 ( .A1(n4525), .A2(n2181), .ZN(n2264) );
  INV_X1 U2558 ( .A(n4529), .ZN(n4622) );
  INV_X1 U2559 ( .A(n3985), .ZN(n4434) );
  NAND2_X1 U2560 ( .A1(n3910), .A2(n3315), .ZN(n2403) );
  INV_X1 U2561 ( .A(n3199), .ZN(n3831) );
  INV_X1 U2562 ( .A(n2716), .ZN(n2952) );
  NOR2_X1 U2563 ( .A1(n2156), .A2(n2304), .ZN(n2303) );
  INV_X1 U2564 ( .A(n3659), .ZN(n2304) );
  INV_X1 U2565 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4897) );
  NOR2_X1 U2566 ( .A1(n4466), .A2(n2218), .ZN(n3948) );
  AND2_X1 U2567 ( .A1(n4569), .A2(REG1_REG_11__SCAN_IN), .ZN(n2218) );
  NOR2_X1 U2568 ( .A1(n2238), .A2(n2233), .ZN(n2232) );
  NAND2_X1 U2569 ( .A1(n2241), .A2(n3973), .ZN(n2238) );
  NOR2_X1 U2570 ( .A1(n2239), .A2(n2242), .ZN(n2237) );
  NAND2_X1 U2571 ( .A1(n4562), .A2(n2252), .ZN(n2251) );
  NAND2_X1 U2572 ( .A1(n3788), .A2(n2616), .ZN(n2185) );
  INV_X1 U2573 ( .A(n4132), .ZN(n2901) );
  INV_X1 U2574 ( .A(n3772), .ZN(n2652) );
  AND2_X1 U2575 ( .A1(n3501), .A2(n3858), .ZN(n3487) );
  NOR2_X1 U2576 ( .A1(n2386), .A2(n3292), .ZN(n2404) );
  INV_X1 U2577 ( .A(n2403), .ZN(n2386) );
  AND2_X1 U2578 ( .A1(n3050), .A2(n2698), .ZN(n3008) );
  INV_X1 U2579 ( .A(n4040), .ZN(n2961) );
  INV_X1 U2580 ( .A(IR_REG_28__SCAN_IN), .ZN(n2345) );
  INV_X1 U2581 ( .A(IR_REG_26__SCAN_IN), .ZN(n2262) );
  INV_X1 U2582 ( .A(IR_REG_20__SCAN_IN), .ZN(n2624) );
  INV_X1 U2583 ( .A(IR_REG_17__SCAN_IN), .ZN(n2258) );
  AOI21_X1 U2584 ( .B1(n2301), .B2(n3518), .A(n2300), .ZN(n2299) );
  AND2_X1 U2585 ( .A1(n2132), .A2(DATAI_25_), .ZN(n2706) );
  AND2_X1 U2586 ( .A1(n3599), .A2(n3600), .ZN(n3598) );
  INV_X1 U2587 ( .A(n2952), .ZN(n2989) );
  INV_X1 U2588 ( .A(n2313), .ZN(n2301) );
  AND2_X1 U2589 ( .A1(n3636), .A2(n3666), .ZN(n3715) );
  AND2_X1 U2590 ( .A1(n2983), .A2(n3213), .ZN(n3006) );
  NAND2_X1 U2591 ( .A1(n2854), .A2(n2855), .ZN(n3733) );
  INV_X1 U2592 ( .A(IR_REG_19__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U2593 ( .A1(n2554), .A2(n2553), .ZN(n2623) );
  NAND2_X1 U2594 ( .A1(n2228), .A2(n2227), .ZN(n3921) );
  OR2_X1 U2595 ( .A1(n3079), .A2(n3071), .ZN(n2228) );
  NAND2_X1 U2596 ( .A1(n3079), .A2(n3071), .ZN(n2227) );
  AOI21_X1 U2597 ( .B1(n3923), .B2(n3922), .A(n3921), .ZN(n3920) );
  NAND2_X1 U2598 ( .A1(n2263), .A2(n3080), .ZN(n2198) );
  OR2_X1 U2599 ( .A1(n3939), .A2(n2247), .ZN(n2244) );
  NAND2_X1 U2600 ( .A1(n2243), .A2(n2245), .ZN(n3137) );
  AND3_X1 U2601 ( .A1(n2243), .A2(n2245), .A3(n2177), .ZN(n3127) );
  NAND2_X1 U2602 ( .A1(n2214), .A2(n2211), .ZN(n3120) );
  INV_X1 U2603 ( .A(n2215), .ZN(n2214) );
  OAI21_X1 U2604 ( .B1(n3103), .B2(n2216), .A(n3105), .ZN(n2215) );
  INV_X1 U2605 ( .A(n3164), .ZN(n2285) );
  NAND2_X1 U2606 ( .A1(n2221), .A2(n2154), .ZN(n2286) );
  AOI21_X1 U2607 ( .B1(n3149), .B2(REG2_REG_7__SCAN_IN), .A(n3148), .ZN(n3151)
         );
  NOR2_X1 U2608 ( .A1(n4624), .A2(n4774), .ZN(n4623) );
  INV_X1 U2609 ( .A(IR_REG_6__SCAN_IN), .ZN(n4894) );
  XNOR2_X1 U2610 ( .A(n3968), .B(n3967), .ZN(n4493) );
  INV_X1 U2611 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3590) );
  AND2_X1 U2612 ( .A1(n4503), .A2(n3951), .ZN(n3952) );
  NAND2_X1 U2613 ( .A1(n4562), .A2(n4354), .ZN(n2274) );
  NAND2_X1 U2614 ( .A1(n4522), .A2(n2251), .ZN(n4536) );
  INV_X1 U2615 ( .A(n4535), .ZN(n2250) );
  NOR2_X1 U2616 ( .A1(n4533), .A2(n2271), .ZN(n2270) );
  INV_X1 U2617 ( .A(n2274), .ZN(n2271) );
  AND2_X1 U2618 ( .A1(n2664), .A2(n2665), .ZN(n3796) );
  OR3_X1 U2619 ( .A1(n2595), .A2(n3651), .A3(n3682), .ZN(n2605) );
  AND2_X1 U2620 ( .A1(n4116), .A2(n2927), .ZN(n2586) );
  AND4_X1 U2621 ( .A1(n2601), .A2(n2600), .A3(n2599), .A4(n2598), .ZN(n4069)
         );
  NAND2_X1 U2622 ( .A1(n4105), .A2(n2579), .ZN(n4082) );
  NAND2_X1 U2623 ( .A1(n4128), .A2(n4108), .ZN(n2579) );
  NOR2_X1 U2624 ( .A1(n2573), .A2(n3706), .ZN(n2580) );
  NOR2_X1 U2625 ( .A1(n4157), .A2(n2901), .ZN(n2261) );
  AND2_X1 U2626 ( .A1(n4149), .A2(n4180), .ZN(n2556) );
  AND2_X1 U2627 ( .A1(n2546), .A2(REG3_REG_19__SCAN_IN), .ZN(n2558) );
  NOR2_X1 U2628 ( .A1(n2534), .A2(n4886), .ZN(n2546) );
  AND2_X1 U2629 ( .A1(n4231), .A2(n3672), .ZN(n2531) );
  AOI21_X1 U2630 ( .B1(n4239), .B2(n2513), .A(n2175), .ZN(n4222) );
  INV_X1 U2631 ( .A(n4240), .ZN(n4245) );
  INV_X1 U2632 ( .A(n4250), .ZN(n2650) );
  NOR2_X1 U2633 ( .A1(n2493), .A2(n3590), .ZN(n2503) );
  AND2_X1 U2634 ( .A1(n3904), .A2(n4277), .ZN(n2491) );
  AND2_X1 U2635 ( .A1(n3862), .A2(n3800), .ZN(n4264) );
  INV_X1 U2636 ( .A(n3801), .ZN(n3508) );
  OR2_X1 U2637 ( .A1(n2471), .A2(n2470), .ZN(n2483) );
  INV_X1 U2638 ( .A(n3490), .ZN(n3496) );
  AND2_X1 U2639 ( .A1(n2450), .A2(REG3_REG_10__SCAN_IN), .ZN(n2457) );
  AND2_X1 U2640 ( .A1(n3854), .A2(n3857), .ZN(n3806) );
  INV_X1 U2641 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3155) );
  AND2_X1 U2642 ( .A1(n3851), .A2(n3847), .ZN(n3805) );
  AND2_X1 U2643 ( .A1(n3845), .A2(n3841), .ZN(n3804) );
  OAI211_X1 U2644 ( .C1(n2362), .C2(n2193), .A(n2192), .B(n2371), .ZN(n3290)
         );
  AND2_X1 U2645 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2387) );
  AND2_X1 U2646 ( .A1(n3327), .A2(n3250), .ZN(n2259) );
  INV_X1 U2647 ( .A(n4272), .ZN(n4234) );
  INV_X1 U2648 ( .A(n4268), .ZN(n4230) );
  NOR2_X1 U2649 ( .A1(n3270), .A2(n3269), .ZN(n3268) );
  NAND2_X1 U2650 ( .A1(n3195), .A2(n3250), .ZN(n3270) );
  INV_X1 U2651 ( .A(n4299), .ZN(n4267) );
  INV_X1 U2652 ( .A(n4153), .ZN(n4265) );
  AND2_X1 U2653 ( .A1(n2672), .A2(n3826), .ZN(n3180) );
  INV_X1 U2654 ( .A(n3018), .ZN(n4006) );
  AND2_X1 U2655 ( .A1(n3180), .A2(n4433), .ZN(n4299) );
  OR2_X1 U2656 ( .A1(n4076), .A2(n2706), .ZN(n2314) );
  NAND2_X1 U2657 ( .A1(n4073), .A2(n4074), .ZN(n4076) );
  INV_X1 U2658 ( .A(n2261), .ZN(n4131) );
  AND2_X1 U2659 ( .A1(n4241), .A2(n2150), .ZN(n4181) );
  NAND2_X1 U2660 ( .A1(n4241), .A2(n2260), .ZN(n4213) );
  NOR2_X1 U2661 ( .A1(n4279), .A2(n3593), .ZN(n4241) );
  INV_X1 U2662 ( .A(n4266), .ZN(n4277) );
  OR2_X1 U2663 ( .A1(n3509), .A2(n4277), .ZN(n4279) );
  NOR2_X1 U2664 ( .A1(n3495), .A2(n3496), .ZN(n3511) );
  OR2_X1 U2665 ( .A1(n3471), .A2(n3470), .ZN(n3495) );
  INV_X1 U2666 ( .A(n4610), .ZN(n4600) );
  NAND2_X1 U2667 ( .A1(n4153), .A2(n4605), .ZN(n4602) );
  NOR2_X1 U2668 ( .A1(n2255), .A2(n3419), .ZN(n2254) );
  INV_X1 U2669 ( .A(n4602), .ZN(n4591) );
  AND2_X1 U2670 ( .A1(n4548), .A2(n2672), .ZN(n4583) );
  INV_X1 U2671 ( .A(IR_REG_29__SCAN_IN), .ZN(n2331) );
  XNOR2_X1 U2672 ( .A(n2682), .B(n2681), .ZN(n2699) );
  AND2_X1 U2673 ( .A1(n2626), .A2(n2305), .ZN(n2680) );
  INV_X1 U2674 ( .A(IR_REG_23__SCAN_IN), .ZN(n2696) );
  INV_X1 U2675 ( .A(IR_REG_24__SCAN_IN), .ZN(n4881) );
  XNOR2_X1 U2676 ( .A(n2697), .B(n2696), .ZN(n3051) );
  XNOR2_X1 U2677 ( .A(n2625), .B(n2624), .ZN(n3890) );
  NAND2_X1 U2678 ( .A1(n2623), .A2(IR_REG_31__SCAN_IN), .ZN(n2625) );
  INV_X1 U2679 ( .A(IR_REG_13__SCAN_IN), .ZN(n2325) );
  XNOR2_X1 U2680 ( .A(n2229), .B(n4844), .ZN(n3079) );
  NAND2_X1 U2681 ( .A1(n2352), .A2(IR_REG_31__SCAN_IN), .ZN(n2229) );
  NAND2_X1 U2682 ( .A1(n2293), .A2(n3724), .ZN(n3574) );
  INV_X1 U2683 ( .A(n3548), .ZN(n3593) );
  INV_X1 U2684 ( .A(n3438), .ZN(n2808) );
  INV_X1 U2685 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4898) );
  INV_X1 U2686 ( .A(n2706), .ZN(n4055) );
  INV_X1 U2687 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3682) );
  INV_X1 U2688 ( .A(n3232), .ZN(n2752) );
  NAND2_X1 U2689 ( .A1(n2132), .A2(DATAI_20_), .ZN(n4155) );
  INV_X1 U2690 ( .A(n3740), .ZN(n3719) );
  NAND3_X1 U2691 ( .A1(n3015), .A2(n3173), .A3(n3898), .ZN(n3743) );
  OAI211_X1 U2692 ( .C1(n3575), .C2(n2670), .A(n2615), .B(n2614), .ZN(n3178)
         );
  INV_X1 U2693 ( .A(n4069), .ZN(n4036) );
  OR2_X1 U2694 ( .A1(n2139), .A2(n3087), .ZN(n2351) );
  OR2_X1 U2695 ( .A1(n2597), .A2(n2333), .ZN(n2339) );
  NAND2_X1 U2696 ( .A1(n2217), .A2(n3103), .ZN(n3143) );
  NAND2_X1 U2697 ( .A1(n3938), .A2(REG1_REG_4__SCAN_IN), .ZN(n2217) );
  NAND2_X1 U2698 ( .A1(n3143), .A2(n3144), .ZN(n3142) );
  NAND2_X1 U2699 ( .A1(n2154), .A2(n2222), .ZN(n4450) );
  NAND2_X1 U2700 ( .A1(n3162), .A2(n4571), .ZN(n2222) );
  INV_X1 U2701 ( .A(n2221), .ZN(n4449) );
  XNOR2_X1 U2702 ( .A(n3946), .B(n2282), .ZN(n4459) );
  NAND2_X1 U2703 ( .A1(n4462), .A2(n3961), .ZN(n4473) );
  INV_X1 U2704 ( .A(n2220), .ZN(n4468) );
  NAND2_X1 U2705 ( .A1(n4628), .A2(n3966), .ZN(n4479) );
  INV_X1 U2706 ( .A(n2279), .ZN(n4481) );
  INV_X1 U2707 ( .A(n2281), .ZN(n4483) );
  AND2_X1 U2708 ( .A1(n2210), .A2(n2144), .ZN(n4506) );
  AND2_X1 U2709 ( .A1(n2279), .A2(n2278), .ZN(n3950) );
  XNOR2_X1 U2710 ( .A(n3952), .B(n3973), .ZN(n4516) );
  OAI211_X1 U2711 ( .C1(n4500), .C2(n3973), .A(n2241), .B(n2236), .ZN(n4514)
         );
  NAND2_X1 U2712 ( .A1(n4500), .A2(n2239), .ZN(n2236) );
  AND2_X1 U2713 ( .A1(n3075), .A2(n3059), .ZN(n4529) );
  NAND2_X1 U2714 ( .A1(n4539), .A2(REG1_REG_18__SCAN_IN), .ZN(n2273) );
  OAI21_X1 U2715 ( .B1(n2272), .B2(n2267), .A(n2266), .ZN(n2265) );
  NAND2_X1 U2716 ( .A1(n2272), .A2(n2273), .ZN(n2266) );
  NOR2_X1 U2717 ( .A1(n2270), .A2(n2268), .ZN(n2267) );
  INV_X1 U2718 ( .A(n2273), .ZN(n2268) );
  NAND2_X1 U2719 ( .A1(n2261), .A2(n4119), .ZN(n4333) );
  AND2_X1 U2720 ( .A1(n4556), .A2(n3296), .ZN(n4019) );
  AND2_X1 U2721 ( .A1(n2188), .A2(n2187), .ZN(n3430) );
  NAND2_X1 U2722 ( .A1(n3365), .A2(n2437), .ZN(n2187) );
  INV_X1 U2723 ( .A(n2436), .ZN(n2188) );
  INV_X1 U2724 ( .A(n4445), .ZN(n4282) );
  OR2_X1 U2725 ( .A1(n3053), .A2(n3016), .ZN(n4242) );
  AND2_X1 U2726 ( .A1(n4204), .A2(n4610), .ZN(n4445) );
  AND2_X1 U2727 ( .A1(n3890), .A2(n4434), .ZN(n4548) );
  INV_X1 U2728 ( .A(n4242), .ZN(n4552) );
  INV_X2 U2729 ( .A(n4619), .ZN(n4621) );
  INV_X1 U2730 ( .A(n3035), .ZN(n3045) );
  INV_X1 U2731 ( .A(n4560), .ZN(n3046) );
  INV_X1 U2732 ( .A(IR_REG_30__SCAN_IN), .ZN(n3038) );
  XNOR2_X1 U2733 ( .A(n2671), .B(IR_REG_28__SCAN_IN), .ZN(n4440) );
  XNOR2_X1 U2734 ( .A(n2685), .B(IR_REG_26__SCAN_IN), .ZN(n4429) );
  INV_X1 U2735 ( .A(n2699), .ZN(n4430) );
  NAND2_X1 U2736 ( .A1(n2160), .A2(IR_REG_31__SCAN_IN), .ZN(n2622) );
  XNOR2_X1 U2737 ( .A(n2627), .B(IR_REG_21__SCAN_IN), .ZN(n4432) );
  XNOR2_X1 U2738 ( .A(n2478), .B(IR_REG_11__SCAN_IN), .ZN(n4569) );
  NOR2_X1 U2739 ( .A1(n2449), .A2(n2464), .ZN(n4435) );
  NAND2_X1 U2740 ( .A1(n2352), .A2(n2275), .ZN(n3076) );
  INV_X1 U2741 ( .A(n2276), .ZN(n2275) );
  OAI21_X1 U2742 ( .B1(IR_REG_31__SCAN_IN), .B2(IR_REG_1__SCAN_IN), .A(n2277), 
        .ZN(n2276) );
  INV_X2 U2743 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  AOI21_X1 U2744 ( .B1(n2289), .B2(n2290), .A(n2165), .ZN(n2287) );
  AOI21_X1 U2745 ( .B1(n2224), .B2(n2223), .A(n4543), .ZN(n4546) );
  NAND2_X1 U2746 ( .A1(n4534), .A2(n4533), .ZN(n2224) );
  NAND2_X1 U2747 ( .A1(n3954), .A2(n2273), .ZN(n2269) );
  MUX2_X1 U2748 ( .A(n4789), .B(n4310), .S(n4621), .Z(n4314) );
  OR2_X1 U2749 ( .A1(n2314), .A2(n2151), .ZN(n2142) );
  AND2_X1 U2750 ( .A1(n4241), .A2(n2149), .ZN(n2143) );
  AOI21_X1 U2751 ( .B1(n2186), .B2(n2171), .A(n2611), .ZN(n3566) );
  OR2_X1 U2752 ( .A1(n3950), .A2(n3967), .ZN(n2144) );
  AND3_X1 U2753 ( .A1(n4438), .A2(REG1_REG_3__SCAN_IN), .A3(n3080), .ZN(n2145)
         );
  NAND2_X1 U2754 ( .A1(n2195), .A2(n2256), .ZN(n2552) );
  INV_X1 U2755 ( .A(n3203), .ZN(n2354) );
  NAND2_X1 U2756 ( .A1(n3001), .A2(n3000), .ZN(n2146) );
  AND2_X1 U2757 ( .A1(n2808), .A2(n2802), .ZN(n2147) );
  AND2_X1 U2758 ( .A1(n2553), .A2(n2624), .ZN(n2148) );
  AND2_X2 U2759 ( .A1(n3028), .A2(n2711), .ZN(n2905) );
  INV_X1 U2760 ( .A(n3959), .ZN(n2282) );
  INV_X1 U2761 ( .A(n4228), .ZN(n2523) );
  AND2_X1 U2762 ( .A1(n4245), .A2(n4228), .ZN(n2149) );
  AND2_X1 U2763 ( .A1(n2260), .A2(n4191), .ZN(n2150) );
  INV_X1 U2764 ( .A(n4285), .ZN(n4556) );
  OR2_X1 U2765 ( .A1(n2961), .A2(n2973), .ZN(n2151) );
  OR3_X1 U2766 ( .A1(n2151), .A2(n4006), .A3(n4014), .ZN(n2152) );
  INV_X1 U2767 ( .A(n3971), .ZN(n2233) );
  AND2_X1 U2768 ( .A1(n2251), .A2(n2250), .ZN(n2153) );
  OR2_X1 U2769 ( .A1(n3162), .A2(n4571), .ZN(n2154) );
  NOR2_X1 U2770 ( .A1(n3479), .A2(n2318), .ZN(n2155) );
  OR2_X1 U2771 ( .A1(n2312), .A2(n2920), .ZN(n2156) );
  AND2_X1 U2772 ( .A1(n2305), .A2(n2681), .ZN(n2157) );
  XOR2_X1 U2773 ( .A(n4004), .B(n3993), .Z(n2158) );
  NAND2_X1 U2774 ( .A1(n3907), .A2(n3425), .ZN(n2159) );
  AOI21_X1 U2775 ( .B1(n4165), .B2(n2557), .A(n2556), .ZN(n4140) );
  AOI21_X1 U2776 ( .B1(n4082), .B2(n2587), .A(n2586), .ZN(n4063) );
  NAND2_X1 U2777 ( .A1(n2626), .A2(n4880), .ZN(n2160) );
  NAND2_X1 U2778 ( .A1(n4225), .A2(n3765), .ZN(n4166) );
  INV_X1 U2779 ( .A(n3419), .ZN(n3404) );
  INV_X1 U2780 ( .A(n3196), .ZN(n3182) );
  MUX2_X1 U2781 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2416), .Z(n3196) );
  AND2_X1 U2782 ( .A1(n2288), .A2(n2287), .ZN(n2161) );
  AND2_X1 U2783 ( .A1(n4522), .A2(n2153), .ZN(n2163) );
  NAND2_X1 U2784 ( .A1(n2626), .A2(n2157), .ZN(n2684) );
  NAND2_X1 U2785 ( .A1(n2328), .A2(n2345), .ZN(n2164) );
  INV_X1 U2786 ( .A(IR_REG_18__SCAN_IN), .ZN(n2541) );
  NOR2_X1 U2787 ( .A1(n2314), .A2(n2152), .ZN(n4287) );
  NAND2_X1 U2788 ( .A1(n3026), .A2(n3025), .ZN(n2165) );
  NOR2_X1 U2789 ( .A1(n2314), .A2(n2961), .ZN(n3567) );
  AND2_X1 U2790 ( .A1(n2293), .A2(n2291), .ZN(n2166) );
  AND2_X1 U2791 ( .A1(n4500), .A2(n3972), .ZN(n2167) );
  OR2_X1 U2792 ( .A1(n3138), .A2(n2247), .ZN(n2168) );
  INV_X1 U2793 ( .A(n2370), .ZN(n2193) );
  OR2_X1 U2794 ( .A1(n2156), .A2(n2907), .ZN(n2169) );
  INV_X1 U2795 ( .A(IR_REG_31__SCAN_IN), .ZN(n2679) );
  INV_X1 U2796 ( .A(n3534), .ZN(n2300) );
  XOR2_X1 U2797 ( .A(n3900), .B(n4011), .Z(n2170) );
  NAND2_X1 U2798 ( .A1(n3901), .A2(n2961), .ZN(n2171) );
  NOR2_X1 U2799 ( .A1(n4333), .A2(n2927), .ZN(n4073) );
  AND2_X1 U2800 ( .A1(n4181), .A2(n4180), .ZN(n4154) );
  NAND2_X1 U2801 ( .A1(n2838), .A2(n2837), .ZN(n3584) );
  NAND2_X1 U2802 ( .A1(n2294), .A2(n2802), .ZN(n3437) );
  NAND2_X1 U2803 ( .A1(n2489), .A2(n2325), .ZN(n2499) );
  NAND2_X1 U2804 ( .A1(n2195), .A2(n2297), .ZN(n2529) );
  NAND2_X1 U2805 ( .A1(n2195), .A2(n2326), .ZN(n2509) );
  INV_X1 U2806 ( .A(n4128), .ZN(n3642) );
  NAND2_X1 U2807 ( .A1(n4241), .A2(n4245), .ZN(n2172) );
  NOR3_X1 U2808 ( .A1(n2314), .A2(n4006), .A3(n2151), .ZN(n4012) );
  OR2_X1 U2809 ( .A1(n3958), .A2(n3433), .ZN(n2173) );
  AND2_X1 U2810 ( .A1(n2291), .A2(n3725), .ZN(n2174) );
  AND2_X1 U2811 ( .A1(n4235), .A2(n4245), .ZN(n2175) );
  NOR2_X1 U2812 ( .A1(n4147), .A2(n2901), .ZN(n2176) );
  INV_X1 U2813 ( .A(n3788), .ZN(n2611) );
  INV_X1 U2814 ( .A(n4214), .ZN(n3672) );
  NAND2_X1 U2815 ( .A1(n4437), .A2(REG2_REG_5__SCAN_IN), .ZN(n2177) );
  INV_X1 U2816 ( .A(n4176), .ZN(n2544) );
  NOR2_X1 U2817 ( .A1(n3340), .A2(n3315), .ZN(n3287) );
  NOR2_X1 U2818 ( .A1(n3340), .A2(n2255), .ZN(n3362) );
  AOI21_X1 U2819 ( .B1(n2469), .B2(n2155), .A(n2468), .ZN(n3507) );
  INV_X1 U2820 ( .A(IR_REG_10__SCAN_IN), .ZN(n2463) );
  NAND2_X1 U2821 ( .A1(n2416), .A2(DATAI_27_), .ZN(n3576) );
  NAND2_X1 U2822 ( .A1(n3240), .A2(n3242), .ZN(n3241) );
  NAND2_X1 U2823 ( .A1(n2296), .A2(n2747), .ZN(n3231) );
  INV_X1 U2824 ( .A(n4119), .ZN(n4108) );
  NAND2_X1 U2825 ( .A1(n2132), .A2(DATAI_22_), .ZN(n4119) );
  NAND2_X1 U2826 ( .A1(n2781), .A2(n2780), .ZN(n2178) );
  NAND4_X1 U2827 ( .A1(n2411), .A2(n2410), .A3(n2409), .A4(n2408), .ZN(n3909)
         );
  AND2_X1 U2828 ( .A1(n3203), .A2(n3182), .ZN(n3195) );
  AND2_X2 U2829 ( .A1(n2703), .A2(n3211), .ZN(n4613) );
  INV_X1 U2830 ( .A(n4613), .ZN(n4611) );
  INV_X1 U2831 ( .A(n4565), .ZN(n3967) );
  INV_X1 U2832 ( .A(n2209), .ZN(n2208) );
  NOR2_X1 U2833 ( .A1(n2278), .A2(n3967), .ZN(n2209) );
  INV_X1 U2834 ( .A(n2242), .ZN(n2241) );
  NOR2_X1 U2835 ( .A1(n3973), .A2(n3972), .ZN(n2242) );
  AND2_X1 U2836 ( .A1(n4524), .A2(n3978), .ZN(n2179) );
  AND2_X1 U2837 ( .A1(n2244), .A2(n2246), .ZN(n2180) );
  INV_X1 U2838 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2213) );
  NAND2_X1 U2839 ( .A1(n2330), .A2(n2331), .ZN(n3037) );
  AND2_X1 U2840 ( .A1(n2272), .A2(n2270), .ZN(n2181) );
  INV_X1 U2841 ( .A(n3954), .ZN(n2272) );
  AND2_X1 U2842 ( .A1(n4438), .A2(n3080), .ZN(n2182) );
  INV_X1 U2843 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2252) );
  INV_X1 U2844 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2200) );
  NAND3_X1 U2845 ( .A1(n2191), .A2(n2190), .A3(n2189), .ZN(n3469) );
  NAND3_X1 U2846 ( .A1(n3365), .A2(n2437), .A3(n2159), .ZN(n2190) );
  AOI21_X2 U2847 ( .B1(n4207), .B2(n2532), .A(n2531), .ZN(n4189) );
  NAND3_X1 U2848 ( .A1(n3240), .A2(n3242), .A3(n2370), .ZN(n2192) );
  NAND2_X1 U2849 ( .A1(n3241), .A2(n2362), .ZN(n3264) );
  INV_X1 U2850 ( .A(n2343), .ZN(n2341) );
  INV_X2 U2851 ( .A(n2499), .ZN(n2195) );
  NAND2_X1 U2852 ( .A1(n2198), .A2(n3081), .ZN(n2202) );
  NOR2_X1 U2853 ( .A1(n4438), .A2(n2200), .ZN(n2197) );
  NAND2_X1 U2854 ( .A1(n2182), .A2(n2263), .ZN(n2201) );
  NAND2_X1 U2855 ( .A1(n2202), .A2(n2201), .ZN(n3099) );
  NAND2_X1 U2856 ( .A1(n2263), .A2(n3080), .ZN(n3100) );
  NAND3_X1 U2857 ( .A1(n2205), .A2(n2208), .A3(n2203), .ZN(n4490) );
  NAND3_X1 U2858 ( .A1(n2205), .A2(n2204), .A3(n2203), .ZN(n2210) );
  INV_X1 U2859 ( .A(n2210), .ZN(n4489) );
  NAND2_X1 U2860 ( .A1(n3938), .A2(n2212), .ZN(n2211) );
  INV_X1 U2861 ( .A(n4502), .ZN(n2235) );
  INV_X1 U2862 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2247) );
  NAND2_X1 U2863 ( .A1(n4523), .A2(n2179), .ZN(n2249) );
  NAND2_X1 U2864 ( .A1(n4523), .A2(n4524), .ZN(n4522) );
  INV_X1 U2865 ( .A(n3340), .ZN(n2253) );
  NAND2_X1 U2866 ( .A1(n2253), .A2(n2254), .ZN(n3403) );
  INV_X1 U2867 ( .A(n3326), .ZN(n2704) );
  NAND3_X1 U2868 ( .A1(n3261), .A2(n3195), .A3(n2259), .ZN(n3326) );
  NAND2_X1 U2869 ( .A1(n3927), .A2(n3926), .ZN(n2263) );
  OAI211_X1 U2870 ( .C1(n4525), .C2(n2269), .A(n2265), .B(n2264), .ZN(n3989)
         );
  NAND3_X1 U2871 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .A3(
        IR_REG_0__SCAN_IN), .ZN(n2277) );
  INV_X1 U2872 ( .A(n2286), .ZN(n3165) );
  INV_X1 U2873 ( .A(n2284), .ZN(n3945) );
  NAND2_X1 U2874 ( .A1(n2286), .A2(n2285), .ZN(n2284) );
  NAND3_X1 U2875 ( .A1(n2838), .A2(n2837), .A3(n2844), .ZN(n3588) );
  NAND2_X1 U2876 ( .A1(n2968), .A2(n2289), .ZN(n2288) );
  NAND2_X1 U2877 ( .A1(n2968), .A2(n2967), .ZN(n2293) );
  NAND2_X1 U2878 ( .A1(n2294), .A2(n2147), .ZN(n3439) );
  NAND2_X1 U2879 ( .A1(n2296), .A2(n2295), .ZN(n3233) );
  AND2_X1 U2880 ( .A1(n2341), .A2(n2328), .ZN(n2344) );
  OAI21_X1 U2881 ( .B1(n3517), .B2(n2301), .A(n3518), .ZN(n3537) );
  NAND2_X1 U2882 ( .A1(n2298), .A2(n2299), .ZN(n2835) );
  NAND2_X1 U2883 ( .A1(n3517), .A2(n3518), .ZN(n2298) );
  NAND2_X1 U2884 ( .A1(n2302), .A2(n2169), .ZN(n2926) );
  NAND3_X1 U2885 ( .A1(n2867), .A2(n3734), .A3(n2303), .ZN(n2302) );
  INV_X1 U2886 ( .A(n2926), .ZN(n3701) );
  NAND3_X1 U2887 ( .A1(n2867), .A2(n3734), .A3(n3659), .ZN(n3607) );
  AND2_X1 U2888 ( .A1(n2626), .A2(n2306), .ZN(n2676) );
  NAND2_X1 U2889 ( .A1(n2705), .A2(n3431), .ZN(n3471) );
  NAND2_X1 U2890 ( .A1(n4154), .A2(n4155), .ZN(n4157) );
  NAND2_X1 U2891 ( .A1(n2704), .A2(n2633), .ZN(n3340) );
  NAND2_X1 U2892 ( .A1(n2401), .A2(n2400), .ZN(n3365) );
  AND2_X1 U2893 ( .A1(n2138), .A2(n3196), .ZN(n3197) );
  INV_X1 U2894 ( .A(n3537), .ZN(n2836) );
  INV_X1 U2895 ( .A(n3561), .ZN(n3562) );
  NOR2_X2 U2896 ( .A1(n3561), .A2(n3750), .ZN(n3993) );
  INV_X1 U2897 ( .A(n2335), .ZN(n4427) );
  AOI21_X2 U2898 ( .B1(n4140), .B2(n2565), .A(n2564), .ZN(n4124) );
  INV_X1 U2899 ( .A(n4629), .ZN(n4537) );
  AND2_X1 U2900 ( .A1(n2709), .A2(n2708), .ZN(n2307) );
  INV_X1 U2901 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2419) );
  AND2_X1 U2902 ( .A1(n4879), .A2(n2510), .ZN(n2308) );
  AND2_X1 U2903 ( .A1(n2328), .A2(n2679), .ZN(n2309) );
  OR2_X1 U2904 ( .A1(n3028), .A2(n4877), .ZN(n2310) );
  INV_X1 U2905 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2470) );
  INV_X2 U2906 ( .A(IR_REG_2__SCAN_IN), .ZN(n4844) );
  INV_X1 U2907 ( .A(n4191), .ZN(n4196) );
  INV_X1 U2908 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U2909 ( .A1(n3291), .A2(n2403), .ZN(n2311) );
  NOR2_X1 U2910 ( .A1(n2915), .A2(n3631), .ZN(n2312) );
  NAND2_X1 U2911 ( .A1(n2826), .A2(n2827), .ZN(n2313) );
  NOR2_X1 U2912 ( .A1(n3703), .A2(n2948), .ZN(n2315) );
  NOR2_X1 U2913 ( .A1(n2942), .A2(n3675), .ZN(n2316) );
  AND2_X1 U2914 ( .A1(n4486), .A2(REG2_REG_13__SCAN_IN), .ZN(n2317) );
  NOR2_X1 U2915 ( .A1(n3905), .A2(n3496), .ZN(n2318) );
  AND2_X1 U2916 ( .A1(n4143), .A2(n2658), .ZN(n3867) );
  NOR2_X1 U2917 ( .A1(n3908), .A2(n3419), .ZN(n2432) );
  INV_X1 U2918 ( .A(n2430), .ZN(n2435) );
  INV_X1 U2919 ( .A(IR_REG_27__SCAN_IN), .ZN(n2328) );
  INV_X1 U2920 ( .A(n3703), .ZN(n2925) );
  INV_X1 U2921 ( .A(n3633), .ZN(n2920) );
  INV_X1 U2922 ( .A(n3965), .ZN(n3963) );
  INV_X1 U2923 ( .A(n4275), .ZN(n3995) );
  AND2_X1 U2924 ( .A1(n3366), .A2(n2430), .ZN(n2437) );
  NAND2_X1 U2925 ( .A1(n2631), .A2(n3814), .ZN(n3245) );
  XNOR2_X1 U2926 ( .A(n2715), .B(n2992), .ZN(n2728) );
  NAND2_X1 U2927 ( .A1(n2926), .A2(n2315), .ZN(n2950) );
  OR2_X1 U2928 ( .A1(n2914), .A2(n2913), .ZN(n3688) );
  INV_X1 U2929 ( .A(n3006), .ZN(n3020) );
  OR2_X1 U2930 ( .A1(n3751), .A2(n3992), .ZN(n4004) );
  AND2_X1 U2931 ( .A1(n3902), .A2(n4146), .ZN(n2564) );
  NAND2_X1 U2932 ( .A1(n2544), .A2(n4191), .ZN(n2545) );
  NAND2_X1 U2933 ( .A1(n2416), .A2(DATAI_28_), .ZN(n3018) );
  AND2_X1 U2934 ( .A1(n4431), .A2(n4432), .ZN(n3050) );
  OR2_X1 U2935 ( .A1(n2483), .A2(n4897), .ZN(n2493) );
  OR2_X1 U2936 ( .A1(n3690), .A2(n3688), .ZN(n3631) );
  AND2_X1 U2937 ( .A1(n3667), .A2(n2866), .ZN(n3659) );
  NAND2_X1 U2938 ( .A1(n2950), .A2(n2949), .ZN(n3678) );
  INV_X1 U2939 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3706) );
  XNOR2_X1 U2940 ( .A(n2733), .B(n2976), .ZN(n2738) );
  INV_X1 U2941 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4920) );
  NOR2_X1 U2942 ( .A1(n2605), .A2(n4920), .ZN(n2612) );
  OR2_X1 U2943 ( .A1(n2597), .A2(n3300), .ZN(n2360) );
  AOI22_X1 U2944 ( .A1(n3129), .A2(REG2_REG_6__SCAN_IN), .B1(n4436), .B2(n3128), .ZN(n3131) );
  NAND2_X1 U2945 ( .A1(n4540), .A2(n4539), .ZN(n4541) );
  INV_X1 U2946 ( .A(n4011), .ZN(n4014) );
  AOI21_X1 U2947 ( .B1(n4263), .B2(n2492), .A(n2491), .ZN(n3545) );
  NAND2_X1 U2948 ( .A1(n4583), .A2(n3826), .ZN(n3016) );
  OR2_X1 U2949 ( .A1(n4613), .A2(n2707), .ZN(n2708) );
  NAND2_X1 U2950 ( .A1(n2132), .A2(DATAI_24_), .ZN(n4074) );
  INV_X1 U2951 ( .A(n3523), .ZN(n3510) );
  AND2_X1 U2952 ( .A1(n2667), .A2(n2666), .ZN(n4275) );
  INV_X1 U2953 ( .A(n4583), .ZN(n4605) );
  NAND2_X1 U2954 ( .A1(n3028), .A2(n4560), .ZN(n3053) );
  AND2_X1 U2955 ( .A1(n2416), .A2(n3052), .ZN(n3058) );
  OR2_X1 U2956 ( .A1(n2420), .A2(n2419), .ZN(n2439) );
  OR2_X1 U2957 ( .A1(n2566), .A2(n4898), .ZN(n2573) );
  OR2_X1 U2958 ( .A1(n2515), .A2(n2514), .ZN(n2534) );
  NOR2_X1 U2959 ( .A1(n2439), .A2(n3155), .ZN(n2450) );
  OR2_X1 U2960 ( .A1(n2618), .A2(n4904), .ZN(n3990) );
  OR2_X1 U2961 ( .A1(n2597), .A2(n3342), .ZN(n2381) );
  AND2_X1 U2962 ( .A1(n3075), .A2(n3913), .ZN(n4540) );
  AND2_X1 U2963 ( .A1(n3075), .A2(n3894), .ZN(n4629) );
  AND2_X1 U2964 ( .A1(n4556), .A2(n3985), .ZN(n4204) );
  OR2_X1 U2965 ( .A1(n3290), .A2(n3813), .ZN(n3333) );
  NAND2_X1 U2966 ( .A1(n3214), .A2(n4242), .ZN(n4236) );
  AND2_X1 U2967 ( .A1(n4621), .A2(n4610), .ZN(n4311) );
  NAND2_X1 U2968 ( .A1(n2132), .A2(DATAI_26_), .ZN(n4040) );
  NAND2_X1 U2969 ( .A1(n2132), .A2(DATAI_23_), .ZN(n4097) );
  INV_X1 U2970 ( .A(n3618), .ZN(n4180) );
  OR2_X1 U2971 ( .A1(n3369), .A2(n3356), .ZN(n4595) );
  AND2_X1 U2972 ( .A1(n4613), .A2(n4610), .ZN(n3459) );
  OAI22_X1 U2973 ( .A1(n3044), .A2(D_REG_0__SCAN_IN), .B1(n3045), .B2(n4429), 
        .ZN(n3211) );
  NOR2_X2 U2974 ( .A1(n3058), .A2(n3054), .ZN(n4627) );
  INV_X1 U2975 ( .A(n3743), .ZN(n3722) );
  INV_X1 U2976 ( .A(n3716), .ZN(n3746) );
  OAI211_X1 U2977 ( .C1(n3728), .C2(n2670), .A(n2610), .B(n2609), .ZN(n3901)
         );
  OR2_X1 U2978 ( .A1(n3028), .A2(n3046), .ZN(n3912) );
  INV_X1 U2979 ( .A(n4569), .ZN(n4477) );
  INV_X1 U2980 ( .A(n4540), .ZN(n4633) );
  INV_X1 U2981 ( .A(n4627), .ZN(n4547) );
  AND2_X1 U2982 ( .A1(n3402), .A2(n3401), .ZN(n3447) );
  INV_X1 U2983 ( .A(n4019), .ZN(n4257) );
  INV_X1 U2984 ( .A(n4311), .ZN(n4376) );
  OR2_X1 U2985 ( .A1(n3185), .A2(n3211), .ZN(n4619) );
  INV_X1 U2986 ( .A(n3459), .ZN(n4425) );
  AND2_X1 U2987 ( .A1(n4577), .A2(n4576), .ZN(n4614) );
  INV_X1 U2988 ( .A(n4558), .ZN(n4559) );
  NAND2_X1 U2989 ( .A1(n3174), .A2(n3044), .ZN(n4558) );
  AND2_X1 U2990 ( .A1(n3051), .A2(STATE_REG_SCAN_IN), .ZN(n4560) );
  AND2_X1 U2991 ( .A1(n2512), .A2(n2521), .ZN(n4509) );
  INV_X2 U2992 ( .A(n3912), .ZN(U4043) );
  AND3_X2 U2993 ( .A1(n2398), .A2(n2319), .A3(n4844), .ZN(n2320) );
  NAND2_X1 U2994 ( .A1(n2320), .A2(n2368), .ZN(n2378) );
  NAND4_X1 U2995 ( .A1(n4890), .A2(n2323), .A3(n2322), .A4(n2321), .ZN(n2324)
         );
  NOR2_X2 U2996 ( .A1(n2378), .A2(n2324), .ZN(n2489) );
  NAND2_X1 U2997 ( .A1(n2438), .A2(REG2_REG_0__SCAN_IN), .ZN(n2340) );
  INV_X1 U2998 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2333) );
  NAND2_X1 U2999 ( .A1(n2356), .A2(REG0_REG_0__SCAN_IN), .ZN(n2337) );
  AND2_X1 U3000 ( .A1(n2337), .A2(n2336), .ZN(n2338) );
  NAND3_X1 U3001 ( .A1(n2340), .A2(n2339), .A3(n2338), .ZN(n2721) );
  NOR2_X1 U3002 ( .A1(n2344), .A2(n2309), .ZN(n3042) );
  MUX2_X2 U3003 ( .A(n3041), .B(n3042), .S(n2345), .Z(n2416) );
  INV_X1 U3004 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3087) );
  NAND2_X1 U3005 ( .A1(n2346), .A2(REG2_REG_1__SCAN_IN), .ZN(n2349) );
  NAND2_X1 U3006 ( .A1(n2363), .A2(REG1_REG_1__SCAN_IN), .ZN(n2348) );
  NAND2_X1 U3007 ( .A1(n2356), .A2(REG0_REG_1__SCAN_IN), .ZN(n2347) );
  AND3_X1 U3008 ( .A1(n2349), .A2(n2348), .A3(n2347), .ZN(n2350) );
  NAND2_X2 U3009 ( .A1(n2351), .A2(n2350), .ZN(n2712) );
  INV_X1 U3010 ( .A(n2368), .ZN(n2352) );
  INV_X1 U3011 ( .A(DATAI_1_), .ZN(n2353) );
  NAND2_X1 U3012 ( .A1(n2712), .A2(n3203), .ZN(n3829) );
  NAND2_X2 U3013 ( .A1(n3832), .A2(n3829), .ZN(n3821) );
  INV_X1 U3014 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3300) );
  NAND2_X1 U3015 ( .A1(n2140), .A2(REG0_REG_2__SCAN_IN), .ZN(n2359) );
  NAND2_X1 U3016 ( .A1(n2363), .A2(REG1_REG_2__SCAN_IN), .ZN(n2358) );
  NAND2_X1 U3017 ( .A1(n2438), .A2(REG2_REG_2__SCAN_IN), .ZN(n2357) );
  INV_X1 U3018 ( .A(DATAI_2_), .ZN(n2361) );
  NAND2_X1 U3019 ( .A1(n2730), .A2(n3250), .ZN(n3836) );
  INV_X1 U3020 ( .A(n3250), .ZN(n3191) );
  OR2_X1 U3021 ( .A1(n2730), .A2(n3191), .ZN(n2362) );
  NAND2_X1 U3022 ( .A1(n2588), .A2(REG0_REG_3__SCAN_IN), .ZN(n2367) );
  NAND2_X1 U3023 ( .A1(n2438), .A2(REG2_REG_3__SCAN_IN), .ZN(n2366) );
  NAND2_X1 U3024 ( .A1(n3755), .A2(REG1_REG_3__SCAN_IN), .ZN(n2365) );
  OR2_X1 U3025 ( .A1(n2597), .A2(REG3_REG_3__SCAN_IN), .ZN(n2364) );
  NAND2_X1 U3026 ( .A1(n2368), .A2(n4844), .ZN(n2369) );
  NAND2_X1 U3027 ( .A1(n2369), .A2(IR_REG_31__SCAN_IN), .ZN(n2396) );
  XNOR2_X1 U3028 ( .A(n2396), .B(IR_REG_3__SCAN_IN), .ZN(n4438) );
  MUX2_X1 U3029 ( .A(n4438), .B(DATAI_3_), .S(n2416), .Z(n3269) );
  NAND2_X1 U3030 ( .A1(n3235), .A2(n3269), .ZN(n2370) );
  OR2_X1 U3031 ( .A1(n3235), .A2(n3269), .ZN(n2371) );
  INV_X1 U3032 ( .A(n3290), .ZN(n2401) );
  NAND2_X1 U3033 ( .A1(n3755), .A2(REG1_REG_6__SCAN_IN), .ZN(n2377) );
  NAND2_X1 U3034 ( .A1(n2588), .A2(REG0_REG_6__SCAN_IN), .ZN(n2376) );
  NAND2_X1 U3035 ( .A1(n2438), .A2(REG2_REG_6__SCAN_IN), .ZN(n2375) );
  NAND2_X1 U3036 ( .A1(n2387), .A2(REG3_REG_5__SCAN_IN), .ZN(n2380) );
  INV_X1 U3037 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2372) );
  AND2_X1 U3038 ( .A1(n2380), .A2(n2372), .ZN(n2373) );
  NOR2_X1 U3039 ( .A1(n2380), .A2(n2372), .ZN(n2406) );
  OR2_X1 U3040 ( .A1(n2373), .A2(n2406), .ZN(n3318) );
  OR2_X1 U3041 ( .A1(n2597), .A2(n3318), .ZN(n2374) );
  NOR2_X1 U3042 ( .A1(n2378), .A2(IR_REG_5__SCAN_IN), .ZN(n2412) );
  OR2_X1 U3043 ( .A1(n2412), .A2(n2679), .ZN(n2379) );
  XNOR2_X1 U3044 ( .A(n2379), .B(IR_REG_6__SCAN_IN), .ZN(n4436) );
  MUX2_X1 U3045 ( .A(n4436), .B(DATAI_6_), .S(n2132), .Z(n3315) );
  NAND2_X1 U3046 ( .A1(n2588), .A2(REG0_REG_5__SCAN_IN), .ZN(n2384) );
  NAND2_X1 U3047 ( .A1(n2438), .A2(REG2_REG_5__SCAN_IN), .ZN(n2383) );
  NAND2_X1 U3048 ( .A1(n3755), .A2(REG1_REG_5__SCAN_IN), .ZN(n2382) );
  OAI21_X1 U3049 ( .B1(n2387), .B2(REG3_REG_5__SCAN_IN), .A(n2380), .ZN(n3342)
         );
  NAND2_X1 U3050 ( .A1(n2378), .A2(IR_REG_31__SCAN_IN), .ZN(n2385) );
  XNOR2_X1 U3051 ( .A(n2385), .B(IR_REG_5__SCAN_IN), .ZN(n4437) );
  MUX2_X1 U3052 ( .A(n4437), .B(DATAI_5_), .S(n2132), .Z(n3341) );
  OR2_X1 U3053 ( .A1(n3911), .A2(n3341), .ZN(n3292) );
  INV_X1 U3054 ( .A(n2387), .ZN(n2391) );
  INV_X1 U3055 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2389) );
  INV_X1 U3056 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2388) );
  NAND2_X1 U3057 ( .A1(n2389), .A2(n2388), .ZN(n2390) );
  NAND2_X1 U3058 ( .A1(n2391), .A2(n2390), .ZN(n3328) );
  OR2_X1 U3059 ( .A1(n2597), .A2(n3328), .ZN(n2395) );
  NAND2_X1 U3060 ( .A1(n2588), .A2(REG0_REG_4__SCAN_IN), .ZN(n2394) );
  NAND2_X1 U3061 ( .A1(n2438), .A2(REG2_REG_4__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U3062 ( .A1(n3755), .A2(REG1_REG_4__SCAN_IN), .ZN(n2392) );
  NAND2_X1 U3063 ( .A1(n2396), .A2(n2319), .ZN(n2397) );
  NAND2_X1 U3064 ( .A1(n2397), .A2(IR_REG_31__SCAN_IN), .ZN(n2399) );
  XNOR2_X1 U3065 ( .A(n2399), .B(n2398), .ZN(n3935) );
  INV_X1 U3066 ( .A(DATAI_4_), .ZN(n3030) );
  MUX2_X1 U3067 ( .A(n3935), .B(n3030), .S(n2132), .Z(n3327) );
  OR2_X1 U3068 ( .A1(n3258), .A2(n3327), .ZN(n3839) );
  NAND2_X1 U3069 ( .A1(n3258), .A2(n3327), .ZN(n3842) );
  NOR2_X1 U3070 ( .A1(n2404), .A2(n3813), .ZN(n2400) );
  INV_X1 U3071 ( .A(n3327), .ZN(n3237) );
  NAND2_X1 U3072 ( .A1(n3258), .A2(n3237), .ZN(n3332) );
  NAND2_X1 U3073 ( .A1(n3911), .A2(n3341), .ZN(n2402) );
  AND2_X1 U3074 ( .A1(n3332), .A2(n2402), .ZN(n3291) );
  NAND2_X1 U3075 ( .A1(n2311), .A2(n2405), .ZN(n3366) );
  NAND2_X1 U3076 ( .A1(n2406), .A2(REG3_REG_7__SCAN_IN), .ZN(n2420) );
  OR2_X1 U3077 ( .A1(n2406), .A2(REG3_REG_7__SCAN_IN), .ZN(n2407) );
  NAND2_X1 U3078 ( .A1(n2420), .A2(n2407), .ZN(n3384) );
  OR2_X1 U3079 ( .A1(n2597), .A2(n3384), .ZN(n2411) );
  NAND2_X1 U3080 ( .A1(n2141), .A2(REG0_REG_7__SCAN_IN), .ZN(n2410) );
  NAND2_X1 U3081 ( .A1(n3755), .A2(REG1_REG_7__SCAN_IN), .ZN(n2409) );
  NAND2_X1 U3082 ( .A1(n2438), .A2(REG2_REG_7__SCAN_IN), .ZN(n2408) );
  NAND2_X1 U3083 ( .A1(n2412), .A2(n4894), .ZN(n2445) );
  NAND2_X1 U3084 ( .A1(n2445), .A2(IR_REG_31__SCAN_IN), .ZN(n2414) );
  INV_X1 U3085 ( .A(IR_REG_7__SCAN_IN), .ZN(n2413) );
  NAND2_X1 U3086 ( .A1(n2414), .A2(n2413), .ZN(n2426) );
  OR2_X1 U3087 ( .A1(n2414), .A2(n2413), .ZN(n2415) );
  NAND2_X1 U3088 ( .A1(n2426), .A2(n2415), .ZN(n3159) );
  INV_X1 U3089 ( .A(DATAI_7_), .ZN(n2417) );
  MUX2_X1 U3090 ( .A(n3159), .B(n2417), .S(n2132), .Z(n3361) );
  INV_X1 U3091 ( .A(n3361), .ZN(n3381) );
  NAND2_X1 U3092 ( .A1(n3909), .A2(n3381), .ZN(n3399) );
  NAND2_X1 U3093 ( .A1(n2588), .A2(REG0_REG_8__SCAN_IN), .ZN(n2425) );
  NAND2_X1 U3094 ( .A1(n2438), .A2(REG2_REG_8__SCAN_IN), .ZN(n2424) );
  NAND2_X1 U3095 ( .A1(n2420), .A2(n2419), .ZN(n2421) );
  NAND2_X1 U3096 ( .A1(n2439), .A2(n2421), .ZN(n3422) );
  OR2_X1 U3097 ( .A1(n2597), .A2(n3422), .ZN(n2423) );
  NAND2_X1 U3098 ( .A1(n3755), .A2(REG1_REG_8__SCAN_IN), .ZN(n2422) );
  NAND2_X1 U3099 ( .A1(n2426), .A2(IR_REG_31__SCAN_IN), .ZN(n2427) );
  XNOR2_X1 U3100 ( .A(n2427), .B(n4671), .ZN(n4571) );
  INV_X1 U3101 ( .A(n4571), .ZN(n3150) );
  MUX2_X1 U3102 ( .A(n3150), .B(DATAI_8_), .S(n2132), .Z(n3419) );
  NAND2_X1 U3103 ( .A1(n3908), .A2(n3419), .ZN(n2428) );
  AND2_X1 U3104 ( .A1(n3399), .A2(n2428), .ZN(n2429) );
  OR2_X1 U3105 ( .A1(n2429), .A2(n2432), .ZN(n2430) );
  NAND2_X1 U3106 ( .A1(n2431), .A2(n3381), .ZN(n2639) );
  NAND2_X1 U3107 ( .A1(n3909), .A2(n3361), .ZN(n3848) );
  NOR2_X1 U3108 ( .A1(n3356), .A2(n2432), .ZN(n2433) );
  OR2_X1 U3109 ( .A1(n3910), .A2(n3315), .ZN(n3367) );
  AND2_X1 U3110 ( .A1(n2433), .A2(n3367), .ZN(n2434) );
  NOR2_X1 U3111 ( .A1(n2435), .A2(n2434), .ZN(n2436) );
  NAND2_X1 U3112 ( .A1(n3755), .A2(REG1_REG_9__SCAN_IN), .ZN(n2444) );
  NAND2_X1 U3113 ( .A1(n2588), .A2(REG0_REG_9__SCAN_IN), .ZN(n2443) );
  NAND2_X1 U3114 ( .A1(n3756), .A2(REG2_REG_9__SCAN_IN), .ZN(n2442) );
  AND2_X1 U3115 ( .A1(n2439), .A2(n3155), .ZN(n2440) );
  OR2_X1 U3116 ( .A1(n2440), .A2(n2450), .ZN(n3432) );
  OR2_X1 U3117 ( .A1(n2597), .A2(n3432), .ZN(n2441) );
  NAND4_X1 U3118 ( .A1(n2444), .A2(n2443), .A3(n2442), .A4(n2441), .ZN(n3907)
         );
  NAND2_X1 U3119 ( .A1(n2448), .A2(IR_REG_31__SCAN_IN), .ZN(n2446) );
  MUX2_X1 U3120 ( .A(IR_REG_31__SCAN_IN), .B(n2446), .S(IR_REG_9__SCAN_IN), 
        .Z(n2447) );
  INV_X1 U3121 ( .A(n2447), .ZN(n2449) );
  MUX2_X1 U3122 ( .A(n4435), .B(DATAI_9_), .S(n2132), .Z(n3425) );
  INV_X1 U3123 ( .A(n3469), .ZN(n2469) );
  NAND2_X1 U3124 ( .A1(n2588), .A2(REG0_REG_10__SCAN_IN), .ZN(n2455) );
  NAND2_X1 U3125 ( .A1(n3756), .A2(REG2_REG_10__SCAN_IN), .ZN(n2454) );
  NAND2_X1 U3126 ( .A1(n3755), .A2(REG1_REG_10__SCAN_IN), .ZN(n2453) );
  NOR2_X1 U3127 ( .A1(n2450), .A2(REG3_REG_10__SCAN_IN), .ZN(n2451) );
  OR2_X1 U3128 ( .A1(n2457), .A2(n2451), .ZN(n3473) );
  OR2_X1 U3129 ( .A1(n2597), .A2(n3473), .ZN(n2452) );
  NAND4_X1 U3130 ( .A1(n2455), .A2(n2454), .A3(n2453), .A4(n2452), .ZN(n3906)
         );
  OR2_X1 U3131 ( .A1(n2464), .A2(n2679), .ZN(n2456) );
  XNOR2_X1 U3132 ( .A(n2456), .B(IR_REG_10__SCAN_IN), .ZN(n3959) );
  MUX2_X1 U3133 ( .A(n3959), .B(DATAI_10_), .S(n2132), .Z(n3470) );
  NOR2_X1 U3134 ( .A1(n3906), .A2(n3470), .ZN(n3479) );
  NAND2_X1 U3135 ( .A1(n2588), .A2(REG0_REG_11__SCAN_IN), .ZN(n2462) );
  NAND2_X1 U3136 ( .A1(n3756), .A2(REG2_REG_11__SCAN_IN), .ZN(n2461) );
  BUF_X4 U3137 ( .A(n2363), .Z(n3755) );
  NAND2_X1 U3138 ( .A1(n3755), .A2(REG1_REG_11__SCAN_IN), .ZN(n2460) );
  NAND2_X1 U3139 ( .A1(n2457), .A2(REG3_REG_11__SCAN_IN), .ZN(n2471) );
  OR2_X1 U3140 ( .A1(n2457), .A2(REG3_REG_11__SCAN_IN), .ZN(n2458) );
  NAND2_X1 U3141 ( .A1(n2471), .A2(n2458), .ZN(n3497) );
  OR2_X1 U3142 ( .A1(n2139), .A2(n3497), .ZN(n2459) );
  NAND4_X1 U3143 ( .A1(n2462), .A2(n2461), .A3(n2460), .A4(n2459), .ZN(n3905)
         );
  NAND2_X1 U3144 ( .A1(n2464), .A2(n2463), .ZN(n2465) );
  NAND2_X1 U3145 ( .A1(n2465), .A2(IR_REG_31__SCAN_IN), .ZN(n2478) );
  INV_X1 U3146 ( .A(DATAI_11_), .ZN(n2466) );
  MUX2_X1 U3147 ( .A(n4477), .B(n2466), .S(n2132), .Z(n3490) );
  OR2_X1 U31480 ( .A1(n3905), .A2(n3490), .ZN(n3501) );
  NAND2_X1 U31490 ( .A1(n3905), .A2(n3490), .ZN(n3858) );
  INV_X1 U3150 ( .A(n3487), .ZN(n2467) );
  NAND2_X1 U3151 ( .A1(n3906), .A2(n3470), .ZN(n3481) );
  AND2_X1 U3152 ( .A1(n2467), .A2(n3481), .ZN(n3480) );
  NOR2_X1 U3153 ( .A1(n2318), .A2(n3480), .ZN(n2468) );
  NAND2_X1 U3154 ( .A1(n3755), .A2(REG1_REG_12__SCAN_IN), .ZN(n2476) );
  NAND2_X1 U3155 ( .A1(n2588), .A2(REG0_REG_12__SCAN_IN), .ZN(n2475) );
  NAND2_X1 U3156 ( .A1(n3756), .A2(REG2_REG_12__SCAN_IN), .ZN(n2474) );
  NAND2_X1 U3157 ( .A1(n2471), .A2(n2470), .ZN(n2472) );
  NAND2_X1 U3158 ( .A1(n2483), .A2(n2472), .ZN(n3526) );
  OR2_X1 U3159 ( .A1(n2139), .A2(n3526), .ZN(n2473) );
  NAND4_X1 U3160 ( .A1(n2476), .A2(n2475), .A3(n2474), .A4(n2473), .ZN(n4271)
         );
  INV_X1 U3161 ( .A(IR_REG_11__SCAN_IN), .ZN(n2477) );
  NAND2_X1 U3162 ( .A1(n2478), .A2(n2477), .ZN(n2479) );
  NAND2_X1 U3163 ( .A1(n2479), .A2(IR_REG_31__SCAN_IN), .ZN(n2480) );
  XNOR2_X1 U3164 ( .A(n2480), .B(IR_REG_12__SCAN_IN), .ZN(n3965) );
  MUX2_X1 U3165 ( .A(n3965), .B(DATAI_12_), .S(n2132), .Z(n3523) );
  NAND2_X1 U3166 ( .A1(n4271), .A2(n3523), .ZN(n2482) );
  NOR2_X1 U3167 ( .A1(n4271), .A2(n3523), .ZN(n2481) );
  AOI21_X1 U3168 ( .B1(n3507), .B2(n2482), .A(n2481), .ZN(n4263) );
  NAND2_X1 U3169 ( .A1(n3755), .A2(REG1_REG_13__SCAN_IN), .ZN(n2488) );
  NAND2_X1 U3170 ( .A1(n2588), .A2(REG0_REG_13__SCAN_IN), .ZN(n2487) );
  NAND2_X1 U3171 ( .A1(n3756), .A2(REG2_REG_13__SCAN_IN), .ZN(n2486) );
  NAND2_X1 U3172 ( .A1(n2483), .A2(n4897), .ZN(n2484) );
  NAND2_X1 U3173 ( .A1(n2493), .A2(n2484), .ZN(n3538) );
  OR2_X1 U3174 ( .A1(n2670), .A2(n3538), .ZN(n2485) );
  NAND4_X1 U3175 ( .A1(n2488), .A2(n2487), .A3(n2486), .A4(n2485), .ZN(n3904)
         );
  INV_X1 U3176 ( .A(n3904), .ZN(n3591) );
  OR2_X1 U3177 ( .A1(n2489), .A2(n2679), .ZN(n2490) );
  XNOR2_X1 U3178 ( .A(n2490), .B(IR_REG_13__SCAN_IN), .ZN(n4486) );
  INV_X1 U3179 ( .A(n4486), .ZN(n4567) );
  INV_X1 U3180 ( .A(DATAI_13_), .ZN(n4640) );
  MUX2_X1 U3181 ( .A(n4567), .B(n4640), .S(n2132), .Z(n4266) );
  NAND2_X1 U3182 ( .A1(n3591), .A2(n4266), .ZN(n2492) );
  NAND2_X1 U3183 ( .A1(n2588), .A2(REG0_REG_14__SCAN_IN), .ZN(n2498) );
  NAND2_X1 U3184 ( .A1(n3756), .A2(REG2_REG_14__SCAN_IN), .ZN(n2497) );
  NAND2_X1 U3185 ( .A1(n3755), .A2(REG1_REG_14__SCAN_IN), .ZN(n2496) );
  AND2_X1 U3186 ( .A1(n2493), .A2(n3590), .ZN(n2494) );
  OR2_X1 U3187 ( .A1(n2494), .A2(n2503), .ZN(n3596) );
  OR2_X1 U3188 ( .A1(n2670), .A2(n3596), .ZN(n2495) );
  NAND4_X1 U3189 ( .A1(n2498), .A2(n2497), .A3(n2496), .A4(n2495), .ZN(n4253)
         );
  NAND2_X1 U3190 ( .A1(n2499), .A2(IR_REG_31__SCAN_IN), .ZN(n2500) );
  XNOR2_X1 U3191 ( .A(n2500), .B(IR_REG_14__SCAN_IN), .ZN(n4565) );
  INV_X1 U3192 ( .A(DATAI_14_), .ZN(n2501) );
  MUX2_X1 U3193 ( .A(n3967), .B(n2501), .S(n2132), .Z(n3548) );
  OR2_X1 U3194 ( .A1(n4253), .A2(n3548), .ZN(n3764) );
  NAND2_X1 U3195 ( .A1(n4253), .A2(n3548), .ZN(n3771) );
  NAND2_X1 U3196 ( .A1(n3764), .A2(n3771), .ZN(n3544) );
  NAND2_X1 U3197 ( .A1(n3545), .A2(n3544), .ZN(n3543) );
  NAND2_X1 U3198 ( .A1(n3543), .A2(n2502), .ZN(n4239) );
  NAND2_X1 U3199 ( .A1(n3755), .A2(REG1_REG_15__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U3200 ( .A1(n2588), .A2(REG0_REG_15__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U3201 ( .A1(n3756), .A2(REG2_REG_15__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U3202 ( .A1(n2503), .A2(REG3_REG_15__SCAN_IN), .ZN(n2515) );
  OR2_X1 U3203 ( .A1(n2503), .A2(REG3_REG_15__SCAN_IN), .ZN(n2504) );
  NAND2_X1 U3204 ( .A1(n2515), .A2(n2504), .ZN(n4243) );
  OR2_X1 U3205 ( .A1(n2670), .A2(n4243), .ZN(n2505) );
  NAND4_X1 U3206 ( .A1(n2508), .A2(n2507), .A3(n2506), .A4(n2505), .ZN(n3903)
         );
  NAND2_X1 U3207 ( .A1(n2509), .A2(IR_REG_31__SCAN_IN), .ZN(n2511) );
  OR2_X1 U3208 ( .A1(n2511), .A2(n2510), .ZN(n2512) );
  NAND2_X1 U3209 ( .A1(n2511), .A2(n2510), .ZN(n2521) );
  MUX2_X1 U32100 ( .A(n4509), .B(DATAI_15_), .S(n2132), .Z(n4240) );
  NAND2_X1 U32110 ( .A1(n3903), .A2(n4240), .ZN(n2513) );
  INV_X1 U32120 ( .A(n3903), .ZN(n4235) );
  NAND2_X1 U32130 ( .A1(n3755), .A2(REG1_REG_16__SCAN_IN), .ZN(n2520) );
  NAND2_X1 U32140 ( .A1(n2588), .A2(REG0_REG_16__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U32150 ( .A1(n3756), .A2(REG2_REG_16__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U32160 ( .A1(n2515), .A2(n2514), .ZN(n2516) );
  NAND2_X1 U32170 ( .A1(n2534), .A2(n2516), .ZN(n4223) );
  OR2_X1 U32180 ( .A1(n2670), .A2(n4223), .ZN(n2517) );
  NAND4_X1 U32190 ( .A1(n2520), .A2(n2519), .A3(n2518), .A4(n2517), .ZN(n4210)
         );
  NAND2_X1 U32200 ( .A1(n2521), .A2(IR_REG_31__SCAN_IN), .ZN(n2522) );
  XNOR2_X1 U32210 ( .A(n2522), .B(n4879), .ZN(n4564) );
  INV_X1 U32220 ( .A(DATAI_16_), .ZN(n4563) );
  MUX2_X1 U32230 ( .A(n4564), .B(n4563), .S(n2132), .Z(n4228) );
  OR2_X1 U32240 ( .A1(n4210), .A2(n4228), .ZN(n3866) );
  NAND2_X1 U32250 ( .A1(n4210), .A2(n4228), .ZN(n3765) );
  NAND2_X1 U32260 ( .A1(n3866), .A2(n3765), .ZN(n4221) );
  INV_X1 U32270 ( .A(n4210), .ZN(n4246) );
  NAND2_X1 U32280 ( .A1(n2588), .A2(REG0_REG_17__SCAN_IN), .ZN(n2528) );
  NAND2_X1 U32290 ( .A1(n3756), .A2(REG2_REG_17__SCAN_IN), .ZN(n2527) );
  NAND2_X1 U32300 ( .A1(n3755), .A2(REG1_REG_17__SCAN_IN), .ZN(n2526) );
  INV_X1 U32310 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4664) );
  XNOR2_X1 U32320 ( .A(n2534), .B(n4664), .ZN(n4215) );
  OR2_X1 U32330 ( .A1(n2670), .A2(n4215), .ZN(n2525) );
  NAND4_X1 U32340 ( .A1(n2528), .A2(n2527), .A3(n2526), .A4(n2525), .ZN(n4231)
         );
  INV_X1 U32350 ( .A(n4231), .ZN(n4199) );
  NAND2_X1 U32360 ( .A1(n2529), .A2(IR_REG_31__SCAN_IN), .ZN(n2530) );
  XNOR2_X1 U32370 ( .A(n2530), .B(IR_REG_17__SCAN_IN), .ZN(n3975) );
  INV_X1 U32380 ( .A(n3975), .ZN(n4562) );
  INV_X1 U32390 ( .A(DATAI_17_), .ZN(n4561) );
  MUX2_X1 U32400 ( .A(n4562), .B(n4561), .S(n2132), .Z(n4214) );
  NAND2_X1 U32410 ( .A1(n4199), .A2(n4214), .ZN(n2532) );
  NAND2_X1 U32420 ( .A1(n2141), .A2(REG0_REG_18__SCAN_IN), .ZN(n2539) );
  NAND2_X1 U32430 ( .A1(n3756), .A2(REG2_REG_18__SCAN_IN), .ZN(n2538) );
  NAND2_X1 U32440 ( .A1(n3755), .A2(REG1_REG_18__SCAN_IN), .ZN(n2537) );
  INV_X1 U32450 ( .A(n2534), .ZN(n2533) );
  AOI21_X1 U32460 ( .B1(n2533), .B2(REG3_REG_17__SCAN_IN), .A(
        REG3_REG_18__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U32470 ( .A1(REG3_REG_18__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .ZN(
        n4886) );
  OR2_X1 U32480 ( .A1(n2535), .A2(n2546), .ZN(n4193) );
  OR2_X1 U32490 ( .A1(n2670), .A2(n4193), .ZN(n2536) );
  NAND4_X1 U32500 ( .A1(n2539), .A2(n2538), .A3(n2537), .A4(n2536), .ZN(n4176)
         );
  OR2_X1 U32510 ( .A1(n2540), .A2(n2679), .ZN(n2542) );
  XNOR2_X1 U32520 ( .A(n2542), .B(n2541), .ZN(n3976) );
  INV_X1 U32530 ( .A(DATAI_18_), .ZN(n2543) );
  MUX2_X1 U32540 ( .A(n3976), .B(n2543), .S(n2132), .Z(n4191) );
  OR2_X1 U32550 ( .A1(n4176), .A2(n4191), .ZN(n4169) );
  NAND2_X1 U32560 ( .A1(n4176), .A2(n4191), .ZN(n4170) );
  NAND2_X1 U32570 ( .A1(n4169), .A2(n4170), .ZN(n4188) );
  NAND2_X1 U32580 ( .A1(n4189), .A2(n4188), .ZN(n4187) );
  NAND2_X1 U32590 ( .A1(n4187), .A2(n2545), .ZN(n4165) );
  NAND2_X1 U32600 ( .A1(n3755), .A2(REG1_REG_19__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U32610 ( .A1(n2141), .A2(REG0_REG_19__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U32620 ( .A1(n3756), .A2(REG2_REG_19__SCAN_IN), .ZN(n2549) );
  NOR2_X1 U32630 ( .A1(n2546), .A2(REG3_REG_19__SCAN_IN), .ZN(n2547) );
  OR2_X1 U32640 ( .A1(n2558), .A2(n2547), .ZN(n4182) );
  OR2_X1 U32650 ( .A1(n2670), .A2(n4182), .ZN(n2548) );
  NAND4_X1 U32660 ( .A1(n2551), .A2(n2550), .A3(n2549), .A4(n2548), .ZN(n4197)
         );
  NAND2_X1 U32670 ( .A1(n2552), .A2(IR_REG_31__SCAN_IN), .ZN(n2554) );
  OR2_X1 U32680 ( .A1(n2554), .A2(n2553), .ZN(n2555) );
  MUX2_X1 U32690 ( .A(n4434), .B(DATAI_19_), .S(n2132), .Z(n3618) );
  NAND2_X1 U32700 ( .A1(n4197), .A2(n3618), .ZN(n2557) );
  INV_X1 U32710 ( .A(n4197), .ZN(n4149) );
  NAND2_X1 U32720 ( .A1(n3755), .A2(REG1_REG_20__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U32730 ( .A1(n2141), .A2(REG0_REG_20__SCAN_IN), .ZN(n2562) );
  NAND2_X1 U32740 ( .A1(n3756), .A2(REG2_REG_20__SCAN_IN), .ZN(n2561) );
  NAND2_X1 U32750 ( .A1(n2558), .A2(REG3_REG_20__SCAN_IN), .ZN(n2566) );
  OR2_X1 U32760 ( .A1(n2558), .A2(REG3_REG_20__SCAN_IN), .ZN(n2559) );
  NAND2_X1 U32770 ( .A1(n2566), .A2(n2559), .ZN(n4158) );
  OR2_X1 U32780 ( .A1(n2670), .A2(n4158), .ZN(n2560) );
  NAND4_X1 U32790 ( .A1(n2563), .A2(n2562), .A3(n2561), .A4(n2560), .ZN(n3902)
         );
  INV_X1 U32800 ( .A(n3902), .ZN(n4174) );
  NAND2_X1 U32810 ( .A1(n4174), .A2(n4155), .ZN(n2565) );
  INV_X1 U32820 ( .A(n4155), .ZN(n4146) );
  NAND2_X1 U32830 ( .A1(n3755), .A2(REG1_REG_21__SCAN_IN), .ZN(n2571) );
  NAND2_X1 U32840 ( .A1(n2141), .A2(REG0_REG_21__SCAN_IN), .ZN(n2570) );
  NAND2_X1 U32850 ( .A1(n3756), .A2(REG2_REG_21__SCAN_IN), .ZN(n2569) );
  NAND2_X1 U32860 ( .A1(n2566), .A2(n4898), .ZN(n2567) );
  NAND2_X1 U32870 ( .A1(n2573), .A2(n2567), .ZN(n4134) );
  OR2_X1 U32880 ( .A1(n2670), .A2(n4134), .ZN(n2568) );
  NAND4_X1 U32890 ( .A1(n2571), .A2(n2570), .A3(n2569), .A4(n2568), .ZN(n4147)
         );
  NAND2_X1 U32900 ( .A1(n2132), .A2(DATAI_21_), .ZN(n4132) );
  NAND2_X1 U32910 ( .A1(n4147), .A2(n2901), .ZN(n2572) );
  NAND2_X1 U32920 ( .A1(n2588), .A2(REG0_REG_22__SCAN_IN), .ZN(n2578) );
  NAND2_X1 U32930 ( .A1(n3756), .A2(REG2_REG_22__SCAN_IN), .ZN(n2577) );
  NAND2_X1 U32940 ( .A1(n3755), .A2(REG1_REG_22__SCAN_IN), .ZN(n2576) );
  AND2_X1 U32950 ( .A1(n2573), .A2(n3706), .ZN(n2574) );
  OR2_X1 U32960 ( .A1(n2574), .A2(n2580), .ZN(n4109) );
  OR2_X1 U32970 ( .A1(n2670), .A2(n4109), .ZN(n2575) );
  NAND4_X1 U32980 ( .A1(n2578), .A2(n2577), .A3(n2576), .A4(n2575), .ZN(n4128)
         );
  NAND2_X1 U32990 ( .A1(n3642), .A2(n4108), .ZN(n4088) );
  NAND2_X1 U33000 ( .A1(n4128), .A2(n4119), .ZN(n2660) );
  NAND2_X1 U33010 ( .A1(n4088), .A2(n2660), .ZN(n4106) );
  NAND2_X1 U33020 ( .A1(n3755), .A2(REG1_REG_23__SCAN_IN), .ZN(n2585) );
  NAND2_X1 U33030 ( .A1(n2141), .A2(REG0_REG_23__SCAN_IN), .ZN(n2584) );
  NAND2_X1 U33040 ( .A1(n3756), .A2(REG2_REG_23__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U33050 ( .A1(n2580), .A2(REG3_REG_23__SCAN_IN), .ZN(n2595) );
  OR2_X1 U33060 ( .A1(n2580), .A2(REG3_REG_23__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U33070 ( .A1(n2595), .A2(n2581), .ZN(n4099) );
  OR2_X1 U33080 ( .A1(n2670), .A2(n4099), .ZN(n2582) );
  NAND4_X1 U33090 ( .A1(n2585), .A2(n2584), .A3(n2583), .A4(n2582), .ZN(n4116)
         );
  INV_X1 U33100 ( .A(n4116), .ZN(n3705) );
  NAND2_X1 U33110 ( .A1(n3705), .A2(n4097), .ZN(n2587) );
  NAND2_X1 U33120 ( .A1(n3755), .A2(REG1_REG_24__SCAN_IN), .ZN(n2592) );
  NAND2_X1 U33130 ( .A1(n2141), .A2(REG0_REG_24__SCAN_IN), .ZN(n2591) );
  NAND2_X1 U33140 ( .A1(n3756), .A2(REG2_REG_24__SCAN_IN), .ZN(n2590) );
  XNOR2_X1 U33150 ( .A(n2595), .B(n3682), .ZN(n3681) );
  OR2_X1 U33160 ( .A1(n2670), .A2(n3681), .ZN(n2589) );
  NAND4_X1 U33170 ( .A1(n2592), .A2(n2591), .A3(n2590), .A4(n2589), .ZN(n4092)
         );
  INV_X1 U33180 ( .A(n4074), .ZN(n2934) );
  NAND2_X1 U33190 ( .A1(n4092), .A2(n2934), .ZN(n2594) );
  NOR2_X1 U33200 ( .A1(n4092), .A2(n2934), .ZN(n2593) );
  AOI21_X1 U33210 ( .B1(n4063), .B2(n2594), .A(n2593), .ZN(n4047) );
  NAND2_X1 U33220 ( .A1(n2588), .A2(REG0_REG_25__SCAN_IN), .ZN(n2601) );
  NAND2_X1 U33230 ( .A1(n3756), .A2(REG2_REG_25__SCAN_IN), .ZN(n2600) );
  NAND2_X1 U33240 ( .A1(n3755), .A2(REG1_REG_25__SCAN_IN), .ZN(n2599) );
  INV_X1 U33250 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3651) );
  OAI21_X1 U33260 ( .B1(n2595), .B2(n3682), .A(n3651), .ZN(n2596) );
  NAND2_X1 U33270 ( .A1(n2596), .A2(n2605), .ZN(n4057) );
  OR2_X1 U33280 ( .A1(n4057), .A2(n2670), .ZN(n2598) );
  NAND2_X1 U33290 ( .A1(n4069), .A2(n4055), .ZN(n2602) );
  NAND2_X1 U33300 ( .A1(n4047), .A2(n2602), .ZN(n2604) );
  NAND2_X1 U33310 ( .A1(n4036), .A2(n2706), .ZN(n2603) );
  NAND2_X1 U33320 ( .A1(n2604), .A2(n2603), .ZN(n4027) );
  AND2_X1 U33330 ( .A1(n2605), .A2(n4920), .ZN(n2606) );
  OR2_X1 U33340 ( .A1(n2606), .A2(n2612), .ZN(n3728) );
  NAND2_X1 U33350 ( .A1(n2141), .A2(REG0_REG_26__SCAN_IN), .ZN(n2608) );
  NAND2_X1 U33360 ( .A1(n3756), .A2(REG2_REG_26__SCAN_IN), .ZN(n2607) );
  AND2_X1 U33370 ( .A1(n2608), .A2(n2607), .ZN(n2610) );
  NAND2_X1 U33380 ( .A1(n3755), .A2(REG1_REG_26__SCAN_IN), .ZN(n2609) );
  OR2_X1 U33390 ( .A1(n3901), .A2(n2961), .ZN(n3788) );
  NAND2_X1 U33400 ( .A1(n2612), .A2(REG3_REG_27__SCAN_IN), .ZN(n2618) );
  OR2_X1 U33410 ( .A1(n2612), .A2(REG3_REG_27__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U33420 ( .A1(n2618), .A2(n2613), .ZN(n3575) );
  AOI22_X1 U33430 ( .A1(n2141), .A2(REG0_REG_27__SCAN_IN), .B1(n3755), .B2(
        REG1_REG_27__SCAN_IN), .ZN(n2615) );
  NAND2_X1 U33440 ( .A1(n3756), .A2(REG2_REG_27__SCAN_IN), .ZN(n2614) );
  INV_X1 U33450 ( .A(n3178), .ZN(n4034) );
  NAND2_X1 U33460 ( .A1(n4034), .A2(n3576), .ZN(n2616) );
  INV_X1 U33470 ( .A(n3576), .ZN(n2973) );
  NAND2_X1 U33480 ( .A1(n3178), .A2(n2973), .ZN(n2617) );
  INV_X1 U33490 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4904) );
  NAND2_X1 U33500 ( .A1(n2618), .A2(n4904), .ZN(n2619) );
  NAND2_X1 U33510 ( .A1(n3990), .A2(n2619), .ZN(n4022) );
  AOI22_X1 U33520 ( .A1(n2141), .A2(REG0_REG_28__SCAN_IN), .B1(n3755), .B2(
        REG1_REG_28__SCAN_IN), .ZN(n2621) );
  NAND2_X1 U3353 ( .A1(n3756), .A2(REG2_REG_28__SCAN_IN), .ZN(n2620) );
  OAI211_X1 U33540 ( .C1(n4022), .C2(n2670), .A(n2621), .B(n2620), .ZN(n4007)
         );
  OR2_X1 U3355 ( .A1(n4007), .A2(n3018), .ZN(n3991) );
  INV_X1 U3356 ( .A(n3991), .ZN(n3751) );
  AND2_X1 U3357 ( .A1(n4007), .A2(n3018), .ZN(n3992) );
  INV_X1 U3358 ( .A(n4004), .ZN(n3797) );
  XNOR2_X1 U3359 ( .A(n4005), .B(n3797), .ZN(n4020) );
  NAND2_X1 U3360 ( .A1(n2194), .A2(IR_REG_31__SCAN_IN), .ZN(n2627) );
  XNOR2_X1 U3361 ( .A(n4431), .B(n3215), .ZN(n2628) );
  NAND2_X1 U3362 ( .A1(n2629), .A2(n3196), .ZN(n3199) );
  INV_X1 U3363 ( .A(n3821), .ZN(n2630) );
  NAND2_X1 U3364 ( .A1(n3831), .A2(n2630), .ZN(n3243) );
  NAND2_X1 U3365 ( .A1(n3243), .A2(n3832), .ZN(n2631) );
  INV_X1 U3366 ( .A(n3242), .ZN(n3814) );
  INV_X1 U3367 ( .A(n3269), .ZN(n3261) );
  NAND2_X1 U3368 ( .A1(n3235), .A2(n3261), .ZN(n3835) );
  INV_X1 U3369 ( .A(n3839), .ZN(n2632) );
  INV_X1 U3370 ( .A(n3341), .ZN(n2633) );
  OR2_X1 U3371 ( .A1(n3911), .A2(n2633), .ZN(n3845) );
  NAND2_X1 U3372 ( .A1(n3335), .A2(n3845), .ZN(n2634) );
  NAND2_X1 U3373 ( .A1(n3911), .A2(n2633), .ZN(n3841) );
  NAND2_X1 U3374 ( .A1(n2634), .A2(n3841), .ZN(n3283) );
  INV_X1 U3375 ( .A(n3283), .ZN(n2636) );
  INV_X1 U3376 ( .A(n3315), .ZN(n2637) );
  AND2_X1 U3377 ( .A1(n3910), .A2(n2637), .ZN(n3846) );
  INV_X1 U3378 ( .A(n3846), .ZN(n2635) );
  NAND2_X1 U3379 ( .A1(n2636), .A2(n2635), .ZN(n2638) );
  OR2_X1 U3380 ( .A1(n3910), .A2(n2637), .ZN(n3844) );
  INV_X1 U3381 ( .A(n2639), .ZN(n2640) );
  OR2_X1 U3382 ( .A1(n3908), .A2(n3404), .ZN(n3851) );
  NAND2_X1 U3383 ( .A1(n3393), .A2(n3851), .ZN(n2641) );
  NAND2_X1 U3384 ( .A1(n3908), .A2(n3404), .ZN(n3847) );
  INV_X1 U3385 ( .A(n3425), .ZN(n3431) );
  AND2_X1 U3386 ( .A1(n3907), .A2(n3431), .ZN(n3855) );
  OR2_X1 U3387 ( .A1(n3907), .A2(n3431), .ZN(n3852) );
  INV_X1 U3388 ( .A(n3470), .ZN(n3465) );
  NAND2_X1 U3389 ( .A1(n3906), .A2(n3465), .ZN(n3857) );
  NAND2_X1 U3390 ( .A1(n3464), .A2(n3857), .ZN(n2642) );
  OR2_X1 U3391 ( .A1(n3906), .A2(n3465), .ZN(n3854) );
  NAND2_X1 U3392 ( .A1(n4271), .A2(n3510), .ZN(n4258) );
  NAND2_X1 U3393 ( .A1(n3904), .A2(n4266), .ZN(n3800) );
  NAND2_X1 U3394 ( .A1(n4258), .A2(n3800), .ZN(n2645) );
  INV_X1 U3395 ( .A(n3858), .ZN(n2643) );
  NOR2_X1 U3396 ( .A1(n2645), .A2(n2643), .ZN(n2644) );
  NAND2_X1 U3397 ( .A1(n3486), .A2(n2644), .ZN(n2648) );
  INV_X1 U3398 ( .A(n2645), .ZN(n3859) );
  OR2_X1 U3399 ( .A1(n4271), .A2(n3510), .ZN(n4260) );
  NAND2_X1 U3400 ( .A1(n3501), .A2(n4260), .ZN(n2646) );
  NAND2_X1 U3401 ( .A1(n3859), .A2(n2646), .ZN(n3863) );
  OR2_X1 U3402 ( .A1(n3904), .A2(n4266), .ZN(n3862) );
  AND2_X1 U3403 ( .A1(n3863), .A2(n3862), .ZN(n2647) );
  NAND2_X1 U3404 ( .A1(n2648), .A2(n2647), .ZN(n3546) );
  INV_X1 U3405 ( .A(n3544), .ZN(n3812) );
  NAND2_X1 U3406 ( .A1(n3546), .A2(n3812), .ZN(n2649) );
  NAND2_X1 U3407 ( .A1(n2649), .A2(n3764), .ZN(n4247) );
  INV_X1 U3408 ( .A(n4247), .ZN(n2651) );
  OR2_X1 U3409 ( .A1(n3903), .A2(n4245), .ZN(n3767) );
  NAND2_X1 U3410 ( .A1(n3903), .A2(n4245), .ZN(n3770) );
  NAND2_X1 U3411 ( .A1(n3767), .A2(n3770), .ZN(n4250) );
  NAND2_X1 U3412 ( .A1(n2651), .A2(n2650), .ZN(n4248) );
  NAND2_X1 U3413 ( .A1(n4248), .A2(n3770), .ZN(n4227) );
  INV_X1 U3414 ( .A(n4221), .ZN(n4226) );
  NAND2_X1 U3415 ( .A1(n4227), .A2(n4226), .ZN(n4225) );
  INV_X1 U3416 ( .A(n4166), .ZN(n2653) );
  NAND2_X1 U3417 ( .A1(n4197), .A2(n4180), .ZN(n3792) );
  NAND2_X1 U3418 ( .A1(n4170), .A2(n3792), .ZN(n2654) );
  AND2_X1 U3419 ( .A1(n4231), .A2(n4214), .ZN(n4168) );
  OR2_X1 U3420 ( .A1(n2654), .A2(n4168), .ZN(n3772) );
  INV_X1 U3421 ( .A(n2654), .ZN(n2657) );
  OR2_X1 U3422 ( .A1(n4231), .A2(n4214), .ZN(n4167) );
  NAND2_X1 U3423 ( .A1(n4169), .A2(n4167), .ZN(n2656) );
  OR2_X1 U3424 ( .A1(n4197), .A2(n4180), .ZN(n3793) );
  INV_X1 U3425 ( .A(n3793), .ZN(n2655) );
  AOI21_X1 U3426 ( .B1(n2657), .B2(n2656), .A(n2655), .ZN(n4143) );
  OR2_X1 U3427 ( .A1(n3902), .A2(n4155), .ZN(n2658) );
  NAND2_X1 U3428 ( .A1(n3902), .A2(n4155), .ZN(n3774) );
  INV_X1 U3429 ( .A(n4088), .ZN(n2659) );
  NOR2_X1 U3430 ( .A1(n4147), .A2(n4132), .ZN(n4085) );
  NOR2_X1 U3431 ( .A1(n2659), .A2(n4085), .ZN(n3874) );
  AND2_X1 U3432 ( .A1(n4147), .A2(n4132), .ZN(n4084) );
  NAND2_X1 U3433 ( .A1(n4088), .A2(n4084), .ZN(n2661) );
  NAND2_X1 U3434 ( .A1(n4116), .A2(n4097), .ZN(n3799) );
  AND2_X1 U3435 ( .A1(n2660), .A2(n3799), .ZN(n3878) );
  NAND2_X1 U3436 ( .A1(n2661), .A2(n3878), .ZN(n3777) );
  AOI21_X1 U3437 ( .B1(n4083), .B2(n3874), .A(n3777), .ZN(n4066) );
  OR2_X1 U3438 ( .A1(n4116), .A2(n4097), .ZN(n4064) );
  OR2_X1 U3439 ( .A1(n4092), .A2(n4074), .ZN(n3798) );
  NAND2_X1 U3440 ( .A1(n4064), .A2(n3798), .ZN(n3876) );
  OR2_X2 U3441 ( .A1(n4066), .A2(n3876), .ZN(n4028) );
  NAND2_X1 U3442 ( .A1(n4069), .A2(n2706), .ZN(n4029) );
  OAI21_X1 U3443 ( .B1(n3901), .B2(n4040), .A(n4029), .ZN(n3875) );
  NAND2_X1 U3444 ( .A1(n4036), .A2(n4055), .ZN(n3791) );
  NAND2_X1 U3445 ( .A1(n4092), .A2(n4074), .ZN(n4048) );
  AND2_X1 U3446 ( .A1(n3791), .A2(n4048), .ZN(n4031) );
  OR2_X1 U3447 ( .A1(n4031), .A2(n3875), .ZN(n2662) );
  NAND2_X1 U3448 ( .A1(n3901), .A2(n4040), .ZN(n3761) );
  NAND2_X1 U3449 ( .A1(n2662), .A2(n3761), .ZN(n3881) );
  INV_X1 U3450 ( .A(n3881), .ZN(n2663) );
  OAI21_X2 U3451 ( .B1(n4028), .B2(n3875), .A(n2663), .ZN(n3560) );
  AND2_X1 U3452 ( .A1(n3178), .A2(n3576), .ZN(n3883) );
  INV_X1 U3453 ( .A(n3883), .ZN(n2664) );
  OR2_X1 U3454 ( .A1(n3178), .A2(n3576), .ZN(n2665) );
  INV_X1 U3455 ( .A(n3796), .ZN(n3559) );
  INV_X1 U3456 ( .A(n2665), .ZN(n3750) );
  NAND2_X1 U3457 ( .A1(n4431), .A2(n4434), .ZN(n2667) );
  INV_X1 U34580 ( .A(n3890), .ZN(n4433) );
  NAND2_X1 U34590 ( .A1(n4433), .A2(n4432), .ZN(n2666) );
  AOI22_X1 U3460 ( .A1(n3756), .A2(REG2_REG_29__SCAN_IN), .B1(n3755), .B2(
        REG1_REG_29__SCAN_IN), .ZN(n2669) );
  NAND2_X1 U3461 ( .A1(n2588), .A2(REG0_REG_29__SCAN_IN), .ZN(n2668) );
  OAI211_X1 U3462 ( .C1(n3990), .C2(n2670), .A(n2669), .B(n2668), .ZN(n3900)
         );
  OR2_X1 U3463 ( .A1(n2344), .A2(n2679), .ZN(n2671) );
  INV_X1 U3464 ( .A(n3050), .ZN(n2985) );
  NOR2_X1 U3465 ( .A1(n3018), .A2(n4267), .ZN(n2673) );
  AOI21_X1 U3466 ( .B1(n3900), .B2(n4230), .A(n2673), .ZN(n2675) );
  NAND2_X1 U34670 ( .A1(n3178), .A2(n4272), .ZN(n2674) );
  AOI21_X1 U3468 ( .B1(n4020), .B2(n4602), .A(n4018), .ZN(n4310) );
  NAND2_X1 U34690 ( .A1(n2697), .A2(n2696), .ZN(n2677) );
  OR2_X1 U3470 ( .A1(n2680), .A2(n2679), .ZN(n2682) );
  NAND2_X1 U34710 ( .A1(n3035), .A2(n2699), .ZN(n2683) );
  MUX2_X1 U3472 ( .A(n3035), .B(n2683), .S(B_REG_SCAN_IN), .Z(n2686) );
  NAND2_X1 U34730 ( .A1(n2684), .A2(IR_REG_31__SCAN_IN), .ZN(n2685) );
  INV_X1 U3474 ( .A(n3044), .ZN(n2982) );
  NOR3_X1 U34750 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .ZN(n2688) );
  NOR4_X1 U3476 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2687) );
  INV_X1 U34770 ( .A(D_REG_4__SCAN_IN), .ZN(n4689) );
  INV_X1 U3478 ( .A(D_REG_6__SCAN_IN), .ZN(n4688) );
  NAND4_X1 U34790 ( .A1(n2688), .A2(n2687), .A3(n4689), .A4(n4688), .ZN(n4928)
         );
  OR4_X1 U3480 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n2694) );
  NOR4_X1 U34810 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2692) );
  NOR4_X1 U3482 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2691) );
  NOR4_X1 U34830 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n2690) );
  NOR4_X1 U3484 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2689) );
  NAND4_X1 U34850 ( .A1(n2692), .A2(n2691), .A3(n2690), .A4(n2689), .ZN(n2693)
         );
  NOR4_X1 U3486 ( .A1(D_REG_25__SCAN_IN), .A2(n4928), .A3(n2694), .A4(n2693), 
        .ZN(n2979) );
  INV_X1 U34870 ( .A(n2979), .ZN(n2695) );
  NAND2_X1 U3488 ( .A1(n2982), .A2(n2695), .ZN(n2702) );
  NAND2_X1 U34890 ( .A1(n3890), .A2(n3985), .ZN(n2698) );
  NOR2_X1 U3490 ( .A1(n3053), .A2(n3008), .ZN(n3212) );
  INV_X1 U34910 ( .A(n4429), .ZN(n2700) );
  NAND2_X1 U3492 ( .A1(n2700), .A2(n2699), .ZN(n2980) );
  OAI21_X1 U34930 ( .B1(n3044), .B2(D_REG_1__SCAN_IN), .A(n2980), .ZN(n2701)
         );
  NAND4_X1 U3494 ( .A1(n2702), .A2(n3212), .A3(n2701), .A4(n3016), .ZN(n3185)
         );
  INV_X1 U34950 ( .A(n3185), .ZN(n2703) );
  OR2_X1 U3496 ( .A1(n4310), .A2(n4611), .ZN(n2710) );
  NAND2_X1 U34970 ( .A1(n3511), .A2(n3510), .ZN(n3509) );
  INV_X1 U3498 ( .A(n4012), .ZN(n4013) );
  AOI21_X1 U34990 ( .B1(n4006), .B2(n2142), .A(n4012), .ZN(n4312) );
  NAND2_X1 U3500 ( .A1(n4312), .A2(n3459), .ZN(n2709) );
  INV_X1 U35010 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2707) );
  NAND2_X1 U3502 ( .A1(n2710), .A2(n2307), .ZN(U3514) );
  INV_X1 U35030 ( .A(n3215), .ZN(n2711) );
  NAND2_X1 U3504 ( .A1(n2712), .A2(n2905), .ZN(n2714) );
  AND2_X1 U35050 ( .A1(n3028), .A2(n3215), .ZN(n2716) );
  NAND2_X1 U35060 ( .A1(n2354), .A2(n2803), .ZN(n2713) );
  NAND2_X1 U35070 ( .A1(n2714), .A2(n2713), .ZN(n2715) );
  NAND2_X1 U35080 ( .A1(n4431), .A2(n3985), .ZN(n3012) );
  NAND2_X1 U35090 ( .A1(n2716), .A2(n4600), .ZN(n2955) );
  NOR2_X1 U35100 ( .A1(n3203), .A2(n2954), .ZN(n2717) );
  AOI21_X1 U35110 ( .B1(n2712), .B2(n2994), .A(n2717), .ZN(n2726) );
  XNOR2_X1 U35120 ( .A(n2728), .B(n2726), .ZN(n3621) );
  NAND2_X1 U35130 ( .A1(n2138), .A2(n2905), .ZN(n2719) );
  NAND2_X1 U35140 ( .A1(n3196), .A2(n2803), .ZN(n2718) );
  NAND2_X1 U35150 ( .A1(n2719), .A2(n2718), .ZN(n2724) );
  INV_X1 U35160 ( .A(n2724), .ZN(n2720) );
  INV_X1 U35170 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4877) );
  NAND2_X1 U35180 ( .A1(n2720), .A2(n2310), .ZN(n3171) );
  INV_X2 U35190 ( .A(n2955), .ZN(n2994) );
  NAND2_X1 U35200 ( .A1(n2138), .A2(n2994), .ZN(n2723) );
  INV_X1 U35210 ( .A(n3028), .ZN(n3011) );
  AOI22_X1 U35220 ( .A1(n3196), .A2(n2905), .B1(IR_REG_0__SCAN_IN), .B2(n3011), 
        .ZN(n2722) );
  NAND2_X1 U35230 ( .A1(n2723), .A2(n2722), .ZN(n3170) );
  NAND2_X1 U35240 ( .A1(n3171), .A2(n3170), .ZN(n3169) );
  OR2_X1 U35250 ( .A1(n2724), .A2(n2992), .ZN(n2725) );
  NAND2_X1 U35260 ( .A1(n3169), .A2(n2725), .ZN(n3623) );
  NAND2_X1 U35270 ( .A1(n3621), .A2(n3623), .ZN(n3622) );
  INV_X1 U35280 ( .A(n2726), .ZN(n2727) );
  NAND2_X1 U35290 ( .A1(n2728), .A2(n2727), .ZN(n2729) );
  NAND2_X1 U35300 ( .A1(n3622), .A2(n2729), .ZN(n3187) );
  INV_X1 U35310 ( .A(n3187), .ZN(n2736) );
  NAND2_X1 U35320 ( .A1(n2730), .A2(n2905), .ZN(n2732) );
  NAND2_X1 U35330 ( .A1(n3191), .A2(n2803), .ZN(n2731) );
  NAND2_X1 U35340 ( .A1(n2732), .A2(n2731), .ZN(n2733) );
  NOR2_X1 U35350 ( .A1(n3250), .A2(n2954), .ZN(n2734) );
  AOI21_X1 U35360 ( .B1(n2730), .B2(n2994), .A(n2734), .ZN(n2737) );
  XNOR2_X1 U35370 ( .A(n2738), .B(n2737), .ZN(n3190) );
  INV_X1 U35380 ( .A(n3190), .ZN(n2735) );
  NAND2_X1 U35390 ( .A1(n2736), .A2(n2735), .ZN(n3188) );
  NAND2_X1 U35400 ( .A1(n2738), .A2(n2737), .ZN(n2739) );
  NAND2_X1 U35410 ( .A1(n3188), .A2(n2739), .ZN(n3223) );
  NAND2_X1 U35420 ( .A1(n3235), .A2(n2905), .ZN(n2741) );
  NAND2_X1 U35430 ( .A1(n3269), .A2(n2803), .ZN(n2740) );
  NAND2_X1 U35440 ( .A1(n2741), .A2(n2740), .ZN(n2742) );
  XNOR2_X1 U35450 ( .A(n2742), .B(n2992), .ZN(n2744) );
  AND2_X1 U35460 ( .A1(n3269), .A2(n2988), .ZN(n2743) );
  AOI21_X1 U35470 ( .B1(n3235), .B2(n2994), .A(n2743), .ZN(n2745) );
  XNOR2_X1 U35480 ( .A(n2744), .B(n2745), .ZN(n3224) );
  INV_X1 U35490 ( .A(n2744), .ZN(n2746) );
  NAND2_X1 U35500 ( .A1(n2746), .A2(n2745), .ZN(n2747) );
  NAND2_X1 U35510 ( .A1(n3258), .A2(n2905), .ZN(n2749) );
  NAND2_X1 U35520 ( .A1(n3237), .A2(n2803), .ZN(n2748) );
  NAND2_X1 U35530 ( .A1(n2749), .A2(n2748), .ZN(n2750) );
  XNOR2_X1 U35540 ( .A(n2750), .B(n2976), .ZN(n2753) );
  NOR2_X1 U35550 ( .A1(n3327), .A2(n2954), .ZN(n2751) );
  AOI21_X1 U35560 ( .B1(n3258), .B2(n2994), .A(n2751), .ZN(n2754) );
  XNOR2_X1 U35570 ( .A(n2753), .B(n2754), .ZN(n3232) );
  INV_X1 U35580 ( .A(n2753), .ZN(n2756) );
  INV_X1 U35590 ( .A(n2754), .ZN(n2755) );
  NAND2_X1 U35600 ( .A1(n2756), .A2(n2755), .ZN(n2757) );
  NAND2_X1 U35610 ( .A1(n3233), .A2(n2757), .ZN(n3278) );
  NAND2_X1 U35620 ( .A1(n3911), .A2(n2905), .ZN(n2759) );
  NAND2_X1 U35630 ( .A1(n3341), .A2(n2803), .ZN(n2758) );
  NAND2_X1 U35640 ( .A1(n2759), .A2(n2758), .ZN(n2760) );
  XNOR2_X1 U35650 ( .A(n2760), .B(n2992), .ZN(n2764) );
  AND2_X1 U35660 ( .A1(n3341), .A2(n2988), .ZN(n2761) );
  AOI21_X1 U35670 ( .B1(n3911), .B2(n2994), .A(n2761), .ZN(n2762) );
  XNOR2_X1 U35680 ( .A(n2764), .B(n2762), .ZN(n3277) );
  NAND2_X1 U35690 ( .A1(n3278), .A2(n3277), .ZN(n3276) );
  INV_X1 U35700 ( .A(n2762), .ZN(n2763) );
  NAND2_X1 U35710 ( .A1(n2764), .A2(n2763), .ZN(n2765) );
  NAND2_X1 U35720 ( .A1(n3276), .A2(n2765), .ZN(n3310) );
  NAND2_X1 U35730 ( .A1(n3910), .A2(n2994), .ZN(n2767) );
  NAND2_X1 U35740 ( .A1(n3315), .A2(n2905), .ZN(n2766) );
  NAND2_X1 U35750 ( .A1(n2767), .A2(n2766), .ZN(n3307) );
  NAND2_X1 U35760 ( .A1(n3310), .A2(n3307), .ZN(n3375) );
  NAND2_X1 U35770 ( .A1(n3908), .A2(n2905), .ZN(n2769) );
  NAND2_X1 U35780 ( .A1(n3419), .A2(n2803), .ZN(n2768) );
  NAND2_X1 U35790 ( .A1(n2769), .A2(n2768), .ZN(n2770) );
  XNOR2_X1 U35800 ( .A(n2770), .B(n2992), .ZN(n2781) );
  INV_X1 U35810 ( .A(n2781), .ZN(n2774) );
  NAND2_X1 U3582 ( .A1(n3908), .A2(n2994), .ZN(n2772) );
  NAND2_X1 U3583 ( .A1(n3419), .A2(n2905), .ZN(n2771) );
  NAND2_X1 U3584 ( .A1(n2772), .A2(n2771), .ZN(n2780) );
  INV_X1 U3585 ( .A(n2780), .ZN(n2773) );
  NAND2_X1 U3586 ( .A1(n2774), .A2(n2773), .ZN(n3414) );
  INV_X1 U3587 ( .A(n3414), .ZN(n2783) );
  NAND2_X1 U3588 ( .A1(n3909), .A2(n2988), .ZN(n2776) );
  NAND2_X1 U3589 ( .A1(n3381), .A2(n2989), .ZN(n2775) );
  NAND2_X1 U3590 ( .A1(n2776), .A2(n2775), .ZN(n2777) );
  XNOR2_X1 U3591 ( .A(n2777), .B(n2992), .ZN(n2790) );
  NOR2_X1 U3592 ( .A1(n3361), .A2(n2954), .ZN(n2778) );
  AOI21_X1 U3593 ( .B1(n3909), .B2(n2994), .A(n2778), .ZN(n2789) );
  INV_X1 U3594 ( .A(n2789), .ZN(n2779) );
  NAND2_X1 U3595 ( .A1(n2790), .A2(n2779), .ZN(n3412) );
  AND2_X1 U3596 ( .A1(n3412), .A2(n2178), .ZN(n2782) );
  OR2_X1 U3597 ( .A1(n2783), .A2(n2782), .ZN(n2788) );
  AND2_X1 U3598 ( .A1(n3375), .A2(n2788), .ZN(n2787) );
  NAND2_X1 U3599 ( .A1(n3910), .A2(n2988), .ZN(n2785) );
  NAND2_X1 U3600 ( .A1(n3315), .A2(n2803), .ZN(n2784) );
  NAND2_X1 U3601 ( .A1(n2785), .A2(n2784), .ZN(n2786) );
  XNOR2_X1 U3602 ( .A(n2786), .B(n2992), .ZN(n3308) );
  OAI21_X1 U3603 ( .B1(n3310), .B2(n3307), .A(n3308), .ZN(n3376) );
  NAND2_X1 U3604 ( .A1(n2787), .A2(n3376), .ZN(n2794) );
  INV_X1 U3605 ( .A(n2788), .ZN(n2792) );
  XNOR2_X1 U3606 ( .A(n2790), .B(n2789), .ZN(n3410) );
  AND2_X1 U3607 ( .A1(n3410), .A2(n3414), .ZN(n2791) );
  OR2_X1 U3608 ( .A1(n2792), .A2(n2791), .ZN(n2793) );
  NAND2_X1 U3609 ( .A1(n2794), .A2(n2793), .ZN(n3385) );
  NAND2_X1 U3610 ( .A1(n3907), .A2(n2905), .ZN(n2796) );
  NAND2_X1 U3611 ( .A1(n3425), .A2(n2803), .ZN(n2795) );
  NAND2_X1 U3612 ( .A1(n2796), .A2(n2795), .ZN(n2797) );
  XNOR2_X1 U3613 ( .A(n2797), .B(n2992), .ZN(n2799) );
  AND2_X1 U3614 ( .A1(n3425), .A2(n2988), .ZN(n2798) );
  AOI21_X1 U3615 ( .B1(n3907), .B2(n2994), .A(n2798), .ZN(n2800) );
  XNOR2_X1 U3616 ( .A(n2799), .B(n2800), .ZN(n3386) );
  INV_X1 U3617 ( .A(n2799), .ZN(n2801) );
  NAND2_X1 U3618 ( .A1(n2801), .A2(n2800), .ZN(n2802) );
  NAND2_X1 U3619 ( .A1(n3906), .A2(n2988), .ZN(n2805) );
  NAND2_X1 U3620 ( .A1(n3470), .A2(n2803), .ZN(n2804) );
  NAND2_X1 U3621 ( .A1(n2805), .A2(n2804), .ZN(n2806) );
  XNOR2_X1 U3622 ( .A(n2806), .B(n2976), .ZN(n2809) );
  AND2_X1 U3623 ( .A1(n3470), .A2(n2988), .ZN(n2807) );
  AOI21_X1 U3624 ( .B1(n3906), .B2(n2994), .A(n2807), .ZN(n2810) );
  XNOR2_X1 U3625 ( .A(n2809), .B(n2810), .ZN(n3438) );
  INV_X1 U3626 ( .A(n2809), .ZN(n2812) );
  INV_X1 U3627 ( .A(n2810), .ZN(n2811) );
  NAND2_X1 U3628 ( .A1(n2812), .A2(n2811), .ZN(n2813) );
  NAND2_X1 U3629 ( .A1(n3439), .A2(n2813), .ZN(n3453) );
  NAND2_X1 U3630 ( .A1(n3905), .A2(n2994), .ZN(n2815) );
  NAND2_X1 U3631 ( .A1(n3496), .A2(n2988), .ZN(n2814) );
  NAND2_X1 U3632 ( .A1(n2815), .A2(n2814), .ZN(n3451) );
  NAND2_X1 U3633 ( .A1(n3905), .A2(n2988), .ZN(n2817) );
  NAND2_X1 U3634 ( .A1(n3496), .A2(n2989), .ZN(n2816) );
  NAND2_X1 U3635 ( .A1(n2817), .A2(n2816), .ZN(n2818) );
  XNOR2_X1 U3636 ( .A(n2818), .B(n2992), .ZN(n3450) );
  OAI21_X1 U3637 ( .B1(n3453), .B2(n3451), .A(n3450), .ZN(n2820) );
  NAND2_X1 U3638 ( .A1(n3453), .A2(n3451), .ZN(n2819) );
  NAND2_X1 U3639 ( .A1(n2820), .A2(n2819), .ZN(n3517) );
  NAND2_X1 U3640 ( .A1(n4271), .A2(n2988), .ZN(n2822) );
  NAND2_X1 U3641 ( .A1(n3523), .A2(n2989), .ZN(n2821) );
  NAND2_X1 U3642 ( .A1(n2822), .A2(n2821), .ZN(n2823) );
  XNOR2_X1 U3643 ( .A(n2823), .B(n2992), .ZN(n2826) );
  NAND2_X1 U3644 ( .A1(n4271), .A2(n2994), .ZN(n2825) );
  NAND2_X1 U3645 ( .A1(n3523), .A2(n2988), .ZN(n2824) );
  NAND2_X1 U3646 ( .A1(n2825), .A2(n2824), .ZN(n2827) );
  INV_X1 U3647 ( .A(n2826), .ZN(n2829) );
  INV_X1 U3648 ( .A(n2827), .ZN(n2828) );
  NAND2_X1 U3649 ( .A1(n2829), .A2(n2828), .ZN(n3518) );
  NAND2_X1 U3650 ( .A1(n3904), .A2(n2988), .ZN(n2831) );
  NAND2_X1 U3651 ( .A1(n4277), .A2(n2989), .ZN(n2830) );
  NAND2_X1 U3652 ( .A1(n2831), .A2(n2830), .ZN(n2832) );
  XNOR2_X1 U3653 ( .A(n2832), .B(n2976), .ZN(n3534) );
  NAND2_X1 U3654 ( .A1(n3904), .A2(n2994), .ZN(n2834) );
  NAND2_X1 U3655 ( .A1(n4277), .A2(n2988), .ZN(n2833) );
  NAND2_X1 U3656 ( .A1(n2834), .A2(n2833), .ZN(n3535) );
  NAND2_X1 U3657 ( .A1(n2835), .A2(n3535), .ZN(n2838) );
  NAND2_X1 U3658 ( .A1(n2836), .A2(n2300), .ZN(n2837) );
  NAND2_X1 U3659 ( .A1(n4253), .A2(n2988), .ZN(n2840) );
  NAND2_X1 U3660 ( .A1(n3593), .A2(n2989), .ZN(n2839) );
  NAND2_X1 U3661 ( .A1(n2840), .A2(n2839), .ZN(n2841) );
  XNOR2_X1 U3662 ( .A(n2841), .B(n2992), .ZN(n2845) );
  NAND2_X1 U3663 ( .A1(n4253), .A2(n2994), .ZN(n2843) );
  NAND2_X1 U3664 ( .A1(n3593), .A2(n2988), .ZN(n2842) );
  NAND2_X1 U3665 ( .A1(n2843), .A2(n2842), .ZN(n2846) );
  AND2_X1 U3666 ( .A1(n2845), .A2(n2846), .ZN(n3585) );
  INV_X1 U3667 ( .A(n2845), .ZN(n2848) );
  INV_X1 U3668 ( .A(n2846), .ZN(n2847) );
  NAND2_X1 U3669 ( .A1(n2848), .A2(n2847), .ZN(n3583) );
  NAND2_X1 U3670 ( .A1(n3903), .A2(n2988), .ZN(n2850) );
  NAND2_X1 U3671 ( .A1(n4240), .A2(n2989), .ZN(n2849) );
  NAND2_X1 U3672 ( .A1(n2850), .A2(n2849), .ZN(n2851) );
  XNOR2_X1 U3673 ( .A(n2851), .B(n2976), .ZN(n2855) );
  NAND2_X1 U3674 ( .A1(n3903), .A2(n2994), .ZN(n2853) );
  NAND2_X1 U3675 ( .A1(n4240), .A2(n2988), .ZN(n2852) );
  NAND2_X1 U3676 ( .A1(n2853), .A2(n2852), .ZN(n3736) );
  NAND2_X1 U3677 ( .A1(n3733), .A2(n3736), .ZN(n2867) );
  INV_X1 U3678 ( .A(n2854), .ZN(n2857) );
  INV_X1 U3679 ( .A(n2855), .ZN(n2856) );
  NAND2_X1 U3680 ( .A1(n4210), .A2(n2988), .ZN(n2859) );
  NAND2_X1 U3681 ( .A1(n2523), .A2(n2989), .ZN(n2858) );
  NAND2_X1 U3682 ( .A1(n2859), .A2(n2858), .ZN(n2860) );
  XNOR2_X1 U3683 ( .A(n2860), .B(n2976), .ZN(n2862) );
  NOR2_X1 U3684 ( .A1(n4228), .A2(n2954), .ZN(n2861) );
  AOI21_X1 U3685 ( .B1(n4210), .B2(n2994), .A(n2861), .ZN(n2863) );
  NAND2_X1 U3686 ( .A1(n2862), .A2(n2863), .ZN(n3667) );
  INV_X1 U3687 ( .A(n2862), .ZN(n2865) );
  INV_X1 U3688 ( .A(n2863), .ZN(n2864) );
  NAND2_X1 U3689 ( .A1(n2865), .A2(n2864), .ZN(n2866) );
  NAND2_X1 U3690 ( .A1(n4231), .A2(n2988), .ZN(n2869) );
  NAND2_X1 U3691 ( .A1(n3672), .A2(n2989), .ZN(n2868) );
  NAND2_X1 U3692 ( .A1(n2869), .A2(n2868), .ZN(n2870) );
  XNOR2_X1 U3693 ( .A(n2870), .B(n2992), .ZN(n2910) );
  INV_X1 U3694 ( .A(n2910), .ZN(n2874) );
  NAND2_X1 U3695 ( .A1(n4231), .A2(n2994), .ZN(n2872) );
  NAND2_X1 U3696 ( .A1(n3672), .A2(n2988), .ZN(n2871) );
  NAND2_X1 U3697 ( .A1(n2872), .A2(n2871), .ZN(n2909) );
  INV_X1 U3698 ( .A(n2909), .ZN(n2873) );
  NAND2_X1 U3699 ( .A1(n2874), .A2(n2873), .ZN(n3665) );
  AND2_X1 U3700 ( .A1(n3667), .A2(n3665), .ZN(n3608) );
  NAND2_X1 U3701 ( .A1(n3902), .A2(n2988), .ZN(n2876) );
  NAND2_X1 U3702 ( .A1(n4146), .A2(n2989), .ZN(n2875) );
  NAND2_X1 U3703 ( .A1(n2876), .A2(n2875), .ZN(n2877) );
  XNOR2_X1 U3704 ( .A(n2877), .B(n2992), .ZN(n2897) );
  NAND2_X1 U3705 ( .A1(n3902), .A2(n2994), .ZN(n2879) );
  OR2_X1 U3706 ( .A1(n4155), .A2(n2954), .ZN(n2878) );
  NAND2_X1 U3707 ( .A1(n2879), .A2(n2878), .ZN(n2898) );
  NAND2_X1 U3708 ( .A1(n2897), .A2(n2898), .ZN(n3694) );
  INV_X1 U3709 ( .A(n3694), .ZN(n2896) );
  NAND2_X1 U3710 ( .A1(n4197), .A2(n2988), .ZN(n2881) );
  NAND2_X1 U3711 ( .A1(n3618), .A2(n2989), .ZN(n2880) );
  NAND2_X1 U3712 ( .A1(n2881), .A2(n2880), .ZN(n2882) );
  XNOR2_X1 U3713 ( .A(n2882), .B(n2992), .ZN(n2891) );
  NAND2_X1 U3714 ( .A1(n4197), .A2(n2994), .ZN(n2884) );
  NAND2_X1 U3715 ( .A1(n3618), .A2(n2988), .ZN(n2883) );
  NAND2_X1 U3716 ( .A1(n2884), .A2(n2883), .ZN(n2892) );
  NAND2_X1 U3717 ( .A1(n2891), .A2(n2892), .ZN(n3613) );
  NAND2_X1 U3718 ( .A1(n4176), .A2(n2994), .ZN(n2886) );
  NAND2_X1 U3719 ( .A1(n4196), .A2(n2988), .ZN(n2885) );
  NAND2_X1 U3720 ( .A1(n2886), .A2(n2885), .ZN(n3609) );
  INV_X1 U3721 ( .A(n3609), .ZN(n3712) );
  NAND2_X1 U3722 ( .A1(n4176), .A2(n2988), .ZN(n2888) );
  NAND2_X1 U3723 ( .A1(n4196), .A2(n2989), .ZN(n2887) );
  NAND2_X1 U3724 ( .A1(n2888), .A2(n2887), .ZN(n2889) );
  XNOR2_X1 U3725 ( .A(n2889), .B(n2992), .ZN(n3713) );
  INV_X1 U3726 ( .A(n3713), .ZN(n2890) );
  NAND3_X1 U3727 ( .A1(n3613), .A2(n3712), .A3(n2890), .ZN(n2895) );
  INV_X1 U3728 ( .A(n2891), .ZN(n2894) );
  INV_X1 U3729 ( .A(n2892), .ZN(n2893) );
  NAND2_X1 U3730 ( .A1(n2894), .A2(n2893), .ZN(n3612) );
  AND2_X1 U3731 ( .A1(n2895), .A2(n3612), .ZN(n3637) );
  OR2_X1 U3732 ( .A1(n2896), .A2(n3637), .ZN(n2908) );
  AND2_X1 U3733 ( .A1(n3608), .A2(n2908), .ZN(n3687) );
  INV_X1 U3734 ( .A(n2897), .ZN(n2900) );
  INV_X1 U3735 ( .A(n2898), .ZN(n2899) );
  NAND2_X1 U3736 ( .A1(n2900), .A2(n2899), .ZN(n3693) );
  AND2_X1 U3737 ( .A1(n3687), .A2(n3693), .ZN(n3630) );
  NAND2_X1 U3738 ( .A1(n4147), .A2(n2988), .ZN(n2903) );
  NAND2_X1 U3739 ( .A1(n2901), .A2(n2989), .ZN(n2902) );
  NAND2_X1 U3740 ( .A1(n2903), .A2(n2902), .ZN(n2904) );
  XNOR2_X1 U3741 ( .A(n2904), .B(n2976), .ZN(n2916) );
  NOR2_X1 U3742 ( .A1(n4132), .A2(n2954), .ZN(n2906) );
  AOI21_X1 U3743 ( .B1(n4147), .B2(n2994), .A(n2906), .ZN(n2917) );
  AND2_X1 U3744 ( .A1(n2916), .A2(n2917), .ZN(n2915) );
  INV_X1 U3745 ( .A(n2915), .ZN(n3634) );
  AND2_X1 U3746 ( .A1(n3630), .A2(n3634), .ZN(n2907) );
  INV_X1 U3747 ( .A(n3693), .ZN(n3690) );
  INV_X1 U3748 ( .A(n2908), .ZN(n2914) );
  NAND2_X1 U3749 ( .A1(n2910), .A2(n2909), .ZN(n3666) );
  NAND2_X1 U3750 ( .A1(n3713), .A2(n3609), .ZN(n2911) );
  AND2_X1 U3751 ( .A1(n3613), .A2(n2911), .ZN(n2912) );
  AND2_X1 U3752 ( .A1(n3666), .A2(n2912), .ZN(n3635) );
  AND2_X1 U3753 ( .A1(n3635), .A2(n3694), .ZN(n2913) );
  INV_X1 U3754 ( .A(n2916), .ZN(n2919) );
  INV_X1 U3755 ( .A(n2917), .ZN(n2918) );
  NAND2_X1 U3756 ( .A1(n2919), .A2(n2918), .ZN(n3633) );
  NAND2_X1 U3757 ( .A1(n4128), .A2(n2988), .ZN(n2922) );
  NAND2_X1 U3758 ( .A1(n4108), .A2(n2989), .ZN(n2921) );
  NAND2_X1 U3759 ( .A1(n2922), .A2(n2921), .ZN(n2923) );
  XNOR2_X1 U3760 ( .A(n2923), .B(n2976), .ZN(n2933) );
  NOR2_X1 U3761 ( .A1(n4119), .A2(n2954), .ZN(n2924) );
  AOI21_X1 U3762 ( .B1(n4128), .B2(n2994), .A(n2924), .ZN(n2932) );
  XNOR2_X1 U3763 ( .A(n2933), .B(n2932), .ZN(n3703) );
  NAND2_X1 U3764 ( .A1(n2926), .A2(n2925), .ZN(n3597) );
  NAND2_X1 U3765 ( .A1(n4116), .A2(n2988), .ZN(n2929) );
  NAND2_X1 U3766 ( .A1(n2927), .A2(n2989), .ZN(n2928) );
  NAND2_X1 U3767 ( .A1(n2929), .A2(n2928), .ZN(n2930) );
  XNOR2_X1 U3768 ( .A(n2930), .B(n2992), .ZN(n2940) );
  NOR2_X1 U3769 ( .A1(n4097), .A2(n2954), .ZN(n2931) );
  AOI21_X1 U3770 ( .B1(n4116), .B2(n2994), .A(n2931), .ZN(n2938) );
  XNOR2_X1 U3771 ( .A(n2940), .B(n2938), .ZN(n3599) );
  NAND2_X1 U3772 ( .A1(n2933), .A2(n2932), .ZN(n3600) );
  NAND2_X1 U3773 ( .A1(n4092), .A2(n2988), .ZN(n2936) );
  NAND2_X1 U3774 ( .A1(n2934), .A2(n2989), .ZN(n2935) );
  NAND2_X1 U3775 ( .A1(n2936), .A2(n2935), .ZN(n2937) );
  XNOR2_X1 U3776 ( .A(n2937), .B(n2992), .ZN(n3680) );
  AND2_X1 U3777 ( .A1(n3598), .A2(n3680), .ZN(n2943) );
  INV_X1 U3778 ( .A(n3680), .ZN(n2942) );
  INV_X1 U3779 ( .A(n2938), .ZN(n2939) );
  NAND2_X1 U3780 ( .A1(n2940), .A2(n2939), .ZN(n2944) );
  NOR2_X1 U3781 ( .A1(n4074), .A2(n2954), .ZN(n2941) );
  AOI21_X1 U3782 ( .B1(n4092), .B2(n2994), .A(n2941), .ZN(n2945) );
  AND2_X1 U3783 ( .A1(n2944), .A2(n2945), .ZN(n3675) );
  AOI21_X1 U3784 ( .B1(n3597), .B2(n2943), .A(n2316), .ZN(n2951) );
  NOR2_X1 U3785 ( .A1(n2945), .A2(n2944), .ZN(n2948) );
  INV_X1 U3786 ( .A(n2945), .ZN(n2946) );
  AND2_X1 U3787 ( .A1(n3598), .A2(n2946), .ZN(n2947) );
  OR2_X1 U3788 ( .A1(n2948), .A2(n2947), .ZN(n2949) );
  NAND2_X1 U3789 ( .A1(n2951), .A2(n3678), .ZN(n3649) );
  OAI22_X1 U3790 ( .A1(n4069), .A2(n2954), .B1(n4055), .B2(n2952), .ZN(n2953)
         );
  XNOR2_X1 U3791 ( .A(n2953), .B(n2976), .ZN(n2957) );
  OAI22_X1 U3792 ( .A1(n4069), .A2(n2955), .B1(n4055), .B2(n2954), .ZN(n2958)
         );
  INV_X1 U3793 ( .A(n2958), .ZN(n2956) );
  NAND2_X1 U3794 ( .A1(n2957), .A2(n2956), .ZN(n3647) );
  NAND2_X1 U3795 ( .A1(n3649), .A2(n3647), .ZN(n2960) );
  INV_X1 U3796 ( .A(n2957), .ZN(n2959) );
  NAND2_X1 U3797 ( .A1(n2959), .A2(n2958), .ZN(n3648) );
  NAND2_X1 U3798 ( .A1(n2960), .A2(n3648), .ZN(n3723) );
  INV_X1 U3799 ( .A(n3723), .ZN(n2968) );
  NAND2_X1 U3800 ( .A1(n3901), .A2(n2988), .ZN(n2963) );
  NAND2_X1 U3801 ( .A1(n2961), .A2(n2989), .ZN(n2962) );
  NAND2_X1 U3802 ( .A1(n2963), .A2(n2962), .ZN(n2964) );
  XNOR2_X1 U3803 ( .A(n2964), .B(n2992), .ZN(n2969) );
  NAND2_X1 U3804 ( .A1(n3901), .A2(n2994), .ZN(n2966) );
  OR2_X1 U3805 ( .A1(n4040), .A2(n2954), .ZN(n2965) );
  NAND2_X1 U3806 ( .A1(n2966), .A2(n2965), .ZN(n2970) );
  AND2_X1 U3807 ( .A1(n2969), .A2(n2970), .ZN(n3725) );
  INV_X1 U3808 ( .A(n3725), .ZN(n2967) );
  INV_X1 U3809 ( .A(n2969), .ZN(n2972) );
  INV_X1 U3810 ( .A(n2970), .ZN(n2971) );
  NAND2_X1 U3811 ( .A1(n2972), .A2(n2971), .ZN(n3724) );
  NAND2_X1 U3812 ( .A1(n3178), .A2(n2988), .ZN(n2975) );
  NAND2_X1 U3813 ( .A1(n2973), .A2(n2989), .ZN(n2974) );
  NAND2_X1 U3814 ( .A1(n2975), .A2(n2974), .ZN(n2977) );
  XNOR2_X1 U3815 ( .A(n2977), .B(n2976), .ZN(n2999) );
  NOR2_X1 U3816 ( .A1(n3576), .A2(n2954), .ZN(n2978) );
  AOI21_X1 U3817 ( .B1(n3178), .B2(n2994), .A(n2978), .ZN(n2998) );
  XNOR2_X1 U3818 ( .A(n2999), .B(n2998), .ZN(n3573) );
  INV_X1 U3819 ( .A(n3211), .ZN(n2983) );
  NAND2_X1 U3820 ( .A1(n2979), .A2(D_REG_1__SCAN_IN), .ZN(n2981) );
  INV_X1 U3821 ( .A(n2980), .ZN(n3049) );
  AOI21_X1 U3822 ( .B1(n2982), .B2(n2981), .A(n3049), .ZN(n3213) );
  NAND2_X1 U3823 ( .A1(n3180), .A2(n4434), .ZN(n2984) );
  NAND2_X1 U3824 ( .A1(n2985), .A2(n2984), .ZN(n2986) );
  OR2_X1 U3825 ( .A1(n2986), .A2(n4299), .ZN(n3005) );
  NOR2_X1 U3826 ( .A1(n3053), .A2(n3005), .ZN(n2987) );
  NAND2_X1 U3827 ( .A1(n4007), .A2(n2988), .ZN(n2991) );
  NAND2_X1 U3828 ( .A1(n4006), .A2(n2989), .ZN(n2990) );
  NAND2_X1 U3829 ( .A1(n2991), .A2(n2990), .ZN(n2993) );
  XNOR2_X1 U3830 ( .A(n2993), .B(n2992), .ZN(n2997) );
  NAND2_X1 U3831 ( .A1(n4007), .A2(n2994), .ZN(n2995) );
  OAI21_X1 U3832 ( .B1(n2954), .B2(n3018), .A(n2995), .ZN(n2996) );
  XNOR2_X1 U3833 ( .A(n2997), .B(n2996), .ZN(n3004) );
  NAND3_X1 U3834 ( .A1(n2166), .A2(n3716), .A3(n3004), .ZN(n3027) );
  INV_X1 U3835 ( .A(n3004), .ZN(n3001) );
  OR2_X1 U3836 ( .A1(n2999), .A2(n2998), .ZN(n3002) );
  AND2_X1 U3837 ( .A1(n3002), .A2(n3716), .ZN(n3000) );
  INV_X1 U3838 ( .A(n3002), .ZN(n3003) );
  NAND3_X1 U3839 ( .A1(n3004), .A2(n3716), .A3(n3003), .ZN(n3026) );
  INV_X1 U3840 ( .A(n4022), .ZN(n3024) );
  INV_X1 U3841 ( .A(n3005), .ZN(n3007) );
  OAI21_X1 U3842 ( .B1(n4299), .B2(n3007), .A(n3020), .ZN(n3010) );
  INV_X1 U3843 ( .A(n3008), .ZN(n3009) );
  NAND2_X1 U3844 ( .A1(n3010), .A2(n3009), .ZN(n3172) );
  OAI21_X1 U3845 ( .B1(n3172), .B2(n3011), .A(STATE_REG_SCAN_IN), .ZN(n3015)
         );
  INV_X1 U3846 ( .A(n3012), .ZN(n3013) );
  NAND3_X1 U3847 ( .A1(n2988), .A2(n4560), .A3(n3013), .ZN(n3019) );
  INV_X1 U3848 ( .A(n3019), .ZN(n3895) );
  NAND2_X1 U3849 ( .A1(n3020), .A2(n3895), .ZN(n3173) );
  INV_X1 U3850 ( .A(n3051), .ZN(n3014) );
  NAND2_X1 U3851 ( .A1(n3014), .A2(STATE_REG_SCAN_IN), .ZN(n3898) );
  NOR3_X1 U3852 ( .A1(n3020), .A2(n4267), .A3(n3053), .ZN(n3017) );
  NOR2_X2 U3853 ( .A1(n3017), .A2(n4552), .ZN(n3740) );
  OAI22_X1 U3854 ( .A1(n3740), .A2(n3018), .B1(STATE_REG_SCAN_IN), .B2(n4904), 
        .ZN(n3023) );
  INV_X1 U3855 ( .A(n3900), .ZN(n3748) );
  NOR2_X1 U3856 ( .A1(n3020), .A2(n3019), .ZN(n3021) );
  NAND2_X2 U3857 ( .A1(n3021), .A2(n3913), .ZN(n3737) );
  OAI22_X1 U3858 ( .A1(n3748), .A2(n3737), .B1(n4034), .B2(n3738), .ZN(n3022)
         );
  AOI211_X1 U3859 ( .C1(n3024), .C2(n3743), .A(n3023), .B(n3022), .ZN(n3025)
         );
  NAND2_X1 U3860 ( .A1(n3027), .A2(n2161), .ZN(U3217) );
  MUX2_X1 U3861 ( .A(n3076), .B(n2353), .S(U3149), .Z(n3029) );
  INV_X1 U3862 ( .A(n3029), .ZN(U3351) );
  MUX2_X1 U3863 ( .A(n3030), .B(n3935), .S(STATE_REG_SCAN_IN), .Z(n3031) );
  INV_X1 U3864 ( .A(n3031), .ZN(U3348) );
  MUX2_X1 U3865 ( .A(n3159), .B(n2417), .S(U3149), .Z(n3032) );
  INV_X1 U3866 ( .A(n3032), .ZN(U3345) );
  INV_X1 U3867 ( .A(n3976), .ZN(n4539) );
  NAND2_X1 U3868 ( .A1(n4539), .A2(STATE_REG_SCAN_IN), .ZN(n3033) );
  OAI21_X1 U3869 ( .B1(STATE_REG_SCAN_IN), .B2(n2543), .A(n3033), .ZN(U3334)
         );
  INV_X1 U3870 ( .A(DATAI_24_), .ZN(n3034) );
  MUX2_X1 U3871 ( .A(n3035), .B(n3034), .S(U3149), .Z(n3036) );
  INV_X1 U3872 ( .A(n3036), .ZN(U3328) );
  NAND3_X1 U3873 ( .A1(n3038), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3040) );
  INV_X1 U3874 ( .A(DATAI_31_), .ZN(n3039) );
  OAI22_X1 U3875 ( .A1(n3037), .A2(n3040), .B1(STATE_REG_SCAN_IN), .B2(n3039), 
        .ZN(U3321) );
  INV_X1 U3876 ( .A(DATAI_27_), .ZN(n4635) );
  AND2_X1 U3877 ( .A1(n3042), .A2(n3041), .ZN(n3997) );
  NAND2_X1 U3878 ( .A1(n3997), .A2(STATE_REG_SCAN_IN), .ZN(n3043) );
  OAI21_X1 U3879 ( .B1(STATE_REG_SCAN_IN), .B2(n4635), .A(n3043), .ZN(U3325)
         );
  INV_X1 U3880 ( .A(n3053), .ZN(n3174) );
  INV_X1 U3881 ( .A(D_REG_0__SCAN_IN), .ZN(n3048) );
  NOR3_X1 U3882 ( .A1(n3046), .A2(n3045), .A3(n4429), .ZN(n3047) );
  AOI21_X1 U3883 ( .B1(n4558), .B2(n3048), .A(n3047), .ZN(U3458) );
  INV_X1 U3884 ( .A(D_REG_1__SCAN_IN), .ZN(n4693) );
  AOI22_X1 U3885 ( .A1(n4558), .A2(n4693), .B1(n3049), .B2(n4560), .ZN(U3459)
         );
  NAND2_X1 U3886 ( .A1(n3051), .A2(n3050), .ZN(n3052) );
  NAND2_X1 U3887 ( .A1(n3053), .A2(n3898), .ZN(n3057) );
  INV_X1 U3888 ( .A(n3057), .ZN(n3054) );
  NOR2_X1 U3889 ( .A1(n4627), .A2(U4043), .ZN(U3148) );
  INV_X1 U3890 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3055) );
  AOI21_X1 U3891 ( .B1(n3997), .B2(n3055), .A(n3913), .ZN(n3918) );
  OAI21_X1 U3892 ( .B1(REG1_REG_0__SCAN_IN), .B2(n3997), .A(n3918), .ZN(n3056)
         );
  MUX2_X1 U3893 ( .A(n3056), .B(n3918), .S(IR_REG_0__SCAN_IN), .Z(n3063) );
  INV_X1 U3894 ( .A(n3075), .ZN(n3062) );
  AOI22_X1 U3895 ( .A1(n4627), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n3061) );
  INV_X1 U3896 ( .A(n3997), .ZN(n3059) );
  NAND3_X1 U3897 ( .A1(n4529), .A2(IR_REG_0__SCAN_IN), .A3(n4877), .ZN(n3060)
         );
  OAI211_X1 U3898 ( .C1(n3063), .C2(n3062), .A(n3061), .B(n3060), .ZN(U3240)
         );
  INV_X1 U3899 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n4911) );
  NAND2_X1 U3900 ( .A1(n3258), .A2(U4043), .ZN(n3064) );
  OAI21_X1 U3901 ( .B1(U4043), .B2(n4911), .A(n3064), .ZN(U3554) );
  INV_X1 U3902 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4820) );
  NAND2_X1 U3903 ( .A1(n2138), .A2(U4043), .ZN(n3065) );
  OAI21_X1 U3904 ( .B1(U4043), .B2(n4820), .A(n3065), .ZN(U3550) );
  INV_X1 U3905 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n4912) );
  NAND2_X1 U3906 ( .A1(n2712), .A2(U4043), .ZN(n3066) );
  OAI21_X1 U3907 ( .B1(U4043), .B2(n4912), .A(n3066), .ZN(U3551) );
  INV_X1 U3908 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4833) );
  NAND2_X1 U3909 ( .A1(n4116), .A2(U4043), .ZN(n3067) );
  OAI21_X1 U3910 ( .B1(U4043), .B2(n4833), .A(n3067), .ZN(U3573) );
  INV_X1 U3911 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4839) );
  NAND2_X1 U3912 ( .A1(n4092), .A2(U4043), .ZN(n3068) );
  OAI21_X1 U3913 ( .B1(U4043), .B2(n4839), .A(n3068), .ZN(U3574) );
  NOR2_X1 U3914 ( .A1(STATE_REG_SCAN_IN), .A2(n2389), .ZN(n3228) );
  INV_X1 U3915 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4915) );
  AND2_X1 U3916 ( .A1(n4440), .A2(n3997), .ZN(n3894) );
  INV_X1 U3917 ( .A(n3079), .ZN(n4439) );
  INV_X1 U3918 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3069) );
  MUX2_X1 U3919 ( .A(n3069), .B(REG2_REG_1__SCAN_IN), .S(n3076), .Z(n3091) );
  AND2_X1 U3920 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3070)
         );
  NAND2_X1 U3921 ( .A1(n3091), .A2(n3070), .ZN(n3923) );
  INV_X1 U3922 ( .A(n3076), .ZN(n3090) );
  NAND2_X1 U3923 ( .A1(n3090), .A2(REG2_REG_1__SCAN_IN), .ZN(n3922) );
  INV_X1 U3924 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3071) );
  AOI21_X1 U3925 ( .B1(REG2_REG_2__SCAN_IN), .B2(n4439), .A(n3920), .ZN(n3106)
         );
  XNOR2_X1 U3926 ( .A(n3106), .B(n4438), .ZN(n3108) );
  XOR2_X1 U3927 ( .A(REG2_REG_3__SCAN_IN), .B(n3108), .Z(n3072) );
  NAND2_X1 U3928 ( .A1(n4629), .A2(n3072), .ZN(n3073) );
  OAI21_X1 U3929 ( .B1(n4915), .B2(n4547), .A(n3073), .ZN(n3074) );
  NOR2_X1 U3930 ( .A1(n3228), .A2(n3074), .ZN(n3084) );
  XNOR2_X1 U3931 ( .A(n3076), .B(REG1_REG_1__SCAN_IN), .ZN(n3086) );
  AND2_X1 U3932 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3085)
         );
  NAND2_X1 U3933 ( .A1(n3086), .A2(n3085), .ZN(n3078) );
  NAND2_X1 U3934 ( .A1(n3090), .A2(REG1_REG_1__SCAN_IN), .ZN(n3077) );
  NAND2_X1 U3935 ( .A1(n3078), .A2(n3077), .ZN(n3927) );
  XNOR2_X1 U3936 ( .A(n3079), .B(REG1_REG_2__SCAN_IN), .ZN(n3926) );
  NAND2_X1 U3937 ( .A1(n4439), .A2(REG1_REG_2__SCAN_IN), .ZN(n3080) );
  INV_X1 U3938 ( .A(n4438), .ZN(n3081) );
  XOR2_X1 U3939 ( .A(n3099), .B(REG1_REG_3__SCAN_IN), .Z(n3082) );
  AOI22_X1 U3940 ( .A1(n4438), .A2(n4540), .B1(n4529), .B2(n3082), .ZN(n3083)
         );
  NAND2_X1 U3941 ( .A1(n3084), .A2(n3083), .ZN(U3243) );
  XNOR2_X1 U3942 ( .A(n3086), .B(n3085), .ZN(n3094) );
  INV_X1 U3943 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n3088) );
  OAI22_X1 U3944 ( .A1(n4547), .A2(n3088), .B1(STATE_REG_SCAN_IN), .B2(n3087), 
        .ZN(n3089) );
  AOI21_X1 U3945 ( .B1(n3090), .B2(n4540), .A(n3089), .ZN(n3093) );
  NAND2_X1 U3946 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3914) );
  OAI211_X1 U3947 ( .C1(n3070), .C2(n3091), .A(n4629), .B(n3923), .ZN(n3092)
         );
  OAI211_X1 U3948 ( .C1(n4622), .C2(n3094), .A(n3093), .B(n3092), .ZN(U3241)
         );
  INV_X1 U3949 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4828) );
  NAND2_X1 U3950 ( .A1(n4231), .A2(U4043), .ZN(n3095) );
  OAI21_X1 U3951 ( .B1(U4043), .B2(n4828), .A(n3095), .ZN(U3567) );
  INV_X1 U3952 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n4831) );
  NAND2_X1 U3953 ( .A1(n4176), .A2(U4043), .ZN(n3096) );
  OAI21_X1 U3954 ( .B1(U4043), .B2(n4831), .A(n3096), .ZN(U3568) );
  INV_X1 U3955 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4826) );
  NAND2_X1 U3956 ( .A1(n3235), .A2(U4043), .ZN(n3097) );
  OAI21_X1 U3957 ( .B1(U4043), .B2(n4826), .A(n3097), .ZN(U3553) );
  INV_X1 U3958 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4919) );
  NAND2_X1 U3959 ( .A1(n4147), .A2(U4043), .ZN(n3098) );
  OAI21_X1 U3960 ( .B1(U4043), .B2(n4919), .A(n3098), .ZN(U3571) );
  NAND2_X1 U3961 ( .A1(n3100), .A2(n4438), .ZN(n3101) );
  XNOR2_X1 U3962 ( .A(n3102), .B(n3935), .ZN(n3938) );
  INV_X1 U3963 ( .A(n3935), .ZN(n3111) );
  NAND2_X1 U3964 ( .A1(n3102), .A2(n3111), .ZN(n3103) );
  INV_X1 U3965 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3104) );
  MUX2_X1 U3966 ( .A(REG1_REG_5__SCAN_IN), .B(n3104), .S(n4437), .Z(n3144) );
  NAND2_X1 U3967 ( .A1(n4437), .A2(REG1_REG_5__SCAN_IN), .ZN(n3105) );
  INV_X1 U3968 ( .A(n4436), .ZN(n3114) );
  XNOR2_X1 U3969 ( .A(n3120), .B(n3114), .ZN(n3122) );
  XNOR2_X1 U3970 ( .A(n3122), .B(REG1_REG_6__SCAN_IN), .ZN(n3118) );
  INV_X1 U3971 ( .A(n3106), .ZN(n3107) );
  AOI22_X1 U3972 ( .A1(n3108), .A2(REG2_REG_3__SCAN_IN), .B1(n4438), .B2(n3107), .ZN(n3109) );
  XNOR2_X1 U3973 ( .A(n3109), .B(n3935), .ZN(n3939) );
  INV_X1 U3974 ( .A(n3109), .ZN(n3110) );
  INV_X1 U3975 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3112) );
  MUX2_X1 U3976 ( .A(n3112), .B(REG2_REG_5__SCAN_IN), .S(n4437), .Z(n3138) );
  XNOR2_X1 U3977 ( .A(n3127), .B(n4436), .ZN(n3129) );
  INV_X1 U3978 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3289) );
  XNOR2_X1 U3979 ( .A(n3129), .B(n3289), .ZN(n3116) );
  NOR2_X1 U3980 ( .A1(STATE_REG_SCAN_IN), .A2(n2372), .ZN(n3314) );
  AOI21_X1 U3981 ( .B1(n4627), .B2(ADDR_REG_6__SCAN_IN), .A(n3314), .ZN(n3113)
         );
  OAI21_X1 U3982 ( .B1(n4633), .B2(n3114), .A(n3113), .ZN(n3115) );
  AOI21_X1 U3983 ( .B1(n3116), .B2(n4629), .A(n3115), .ZN(n3117) );
  OAI21_X1 U3984 ( .B1(n3118), .B2(n4622), .A(n3117), .ZN(U3246) );
  INV_X1 U3985 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U3986 ( .A1(n4128), .A2(U4043), .ZN(n3119) );
  OAI21_X1 U3987 ( .B1(U4043), .B2(n4918), .A(n3119), .ZN(U3572) );
  AND2_X1 U3988 ( .A1(n3120), .A2(n4436), .ZN(n3121) );
  AOI21_X1 U3989 ( .B1(n3122), .B2(REG1_REG_6__SCAN_IN), .A(n3121), .ZN(n3157)
         );
  MUX2_X1 U3990 ( .A(REG1_REG_7__SCAN_IN), .B(n3158), .S(n3159), .Z(n3123) );
  XNOR2_X1 U3991 ( .A(n3157), .B(n3123), .ZN(n3135) );
  INV_X1 U3992 ( .A(n3159), .ZN(n3149) );
  INV_X1 U3993 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n3126) );
  INV_X1 U3994 ( .A(REG3_REG_7__SCAN_IN), .ZN(n3124) );
  NOR2_X1 U3995 ( .A1(STATE_REG_SCAN_IN), .A2(n3124), .ZN(n3380) );
  INV_X1 U3996 ( .A(n3380), .ZN(n3125) );
  OAI21_X1 U3997 ( .B1(n4547), .B2(n3126), .A(n3125), .ZN(n3133) );
  INV_X1 U3998 ( .A(n3127), .ZN(n3128) );
  INV_X1 U3999 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3364) );
  MUX2_X1 U4000 ( .A(REG2_REG_7__SCAN_IN), .B(n3364), .S(n3159), .Z(n3130) );
  NOR2_X1 U4001 ( .A1(n3131), .A2(n3130), .ZN(n3148) );
  AOI211_X1 U4002 ( .C1(n3131), .C2(n3130), .A(n4537), .B(n3148), .ZN(n3132)
         );
  AOI211_X1 U4003 ( .C1(n4540), .C2(n3149), .A(n3133), .B(n3132), .ZN(n3134)
         );
  OAI21_X1 U4004 ( .B1(n4622), .B2(n3135), .A(n3134), .ZN(U3247) );
  INV_X1 U4005 ( .A(n4437), .ZN(n3147) );
  INV_X1 U4006 ( .A(REG3_REG_5__SCAN_IN), .ZN(n3136) );
  NOR2_X1 U4007 ( .A1(STATE_REG_SCAN_IN), .A2(n3136), .ZN(n3280) );
  INV_X1 U4008 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4816) );
  AOI211_X1 U4009 ( .C1(n2180), .C2(n3138), .A(n3137), .B(n4537), .ZN(n3139)
         );
  INV_X1 U4010 ( .A(n3139), .ZN(n3140) );
  OAI21_X1 U4011 ( .B1(n4547), .B2(n4816), .A(n3140), .ZN(n3141) );
  NOR2_X1 U4012 ( .A1(n3280), .A2(n3141), .ZN(n3146) );
  OAI211_X1 U4013 ( .C1(n3144), .C2(n3143), .A(n4529), .B(n3142), .ZN(n3145)
         );
  OAI211_X1 U4014 ( .C1(n4633), .C2(n3147), .A(n3146), .B(n3145), .ZN(U3245)
         );
  INV_X1 U4015 ( .A(n4435), .ZN(n3958) );
  OR2_X1 U4016 ( .A1(n3151), .A2(n4571), .ZN(n3152) );
  XNOR2_X1 U4017 ( .A(n3151), .B(n3150), .ZN(n4455) );
  NAND2_X1 U4018 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4455), .ZN(n4454) );
  NAND2_X1 U4019 ( .A1(n3152), .A2(n4454), .ZN(n3154) );
  INV_X1 U4020 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3433) );
  MUX2_X1 U4021 ( .A(REG2_REG_9__SCAN_IN), .B(n3433), .S(n4435), .Z(n3153) );
  NAND2_X1 U4022 ( .A1(n3154), .A2(n3153), .ZN(n3957) );
  OAI211_X1 U4023 ( .C1(n3154), .C2(n3153), .A(n3957), .B(n4629), .ZN(n3168)
         );
  NOR2_X1 U4024 ( .A1(STATE_REG_SCAN_IN), .A2(n3155), .ZN(n3390) );
  INV_X1 U4025 ( .A(REG1_REG_7__SCAN_IN), .ZN(n3158) );
  OR2_X1 U4026 ( .A1(n3159), .A2(n3158), .ZN(n3156) );
  NAND2_X1 U4027 ( .A1(n3157), .A2(n3156), .ZN(n3161) );
  NAND2_X1 U4028 ( .A1(n3159), .A2(n3158), .ZN(n3160) );
  NAND2_X1 U4029 ( .A1(n3161), .A2(n3160), .ZN(n3162) );
  INV_X1 U4030 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4451) );
  INV_X1 U4031 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3163) );
  MUX2_X1 U4032 ( .A(n3163), .B(REG1_REG_9__SCAN_IN), .S(n4435), .Z(n3164) );
  AOI211_X1 U4033 ( .C1(n3165), .C2(n3164), .A(n3945), .B(n4622), .ZN(n3166)
         );
  AOI211_X1 U4034 ( .C1(n4627), .C2(ADDR_REG_9__SCAN_IN), .A(n3390), .B(n3166), 
        .ZN(n3167) );
  OAI211_X1 U4035 ( .C1(n4633), .C2(n3958), .A(n3168), .B(n3167), .ZN(U3249)
         );
  OAI21_X1 U4036 ( .B1(n3171), .B2(n3170), .A(n3169), .ZN(n3916) );
  INV_X1 U4037 ( .A(n3172), .ZN(n3175) );
  NAND3_X1 U4038 ( .A1(n3175), .A2(n3174), .A3(n3173), .ZN(n3626) );
  INV_X1 U4039 ( .A(n2712), .ZN(n3184) );
  OAI22_X1 U4040 ( .A1(n3740), .A2(n3182), .B1(n3184), .B2(n3737), .ZN(n3176)
         );
  AOI21_X1 U4041 ( .B1(REG3_REG_0__SCAN_IN), .B2(n3626), .A(n3176), .ZN(n3177)
         );
  OAI21_X1 U4042 ( .B1(n3746), .B2(n3916), .A(n3177), .ZN(U3229) );
  INV_X1 U40430 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4917) );
  NAND2_X1 U4044 ( .A1(n3178), .A2(U4043), .ZN(n3179) );
  OAI21_X1 U4045 ( .B1(U4043), .B2(n4917), .A(n3179), .ZN(U3577) );
  NAND2_X1 U4046 ( .A1(n2138), .A2(n3182), .ZN(n3830) );
  NAND2_X1 U4047 ( .A1(n3199), .A2(n3830), .ZN(n4554) );
  INV_X1 U4048 ( .A(n3180), .ZN(n3181) );
  NOR2_X1 U4049 ( .A1(n3182), .A2(n3181), .ZN(n4551) );
  OAI21_X1 U4050 ( .B1(n4265), .B2(n3995), .A(n4554), .ZN(n3183) );
  OAI21_X1 U4051 ( .B1(n3184), .B2(n4268), .A(n3183), .ZN(n4549) );
  AOI211_X1 U4052 ( .C1(n4583), .C2(n4554), .A(n4551), .B(n4549), .ZN(n4572)
         );
  NAND2_X1 U4053 ( .A1(n4619), .A2(REG1_REG_0__SCAN_IN), .ZN(n3186) );
  OAI21_X1 U4054 ( .B1(n4572), .B2(n4619), .A(n3186), .ZN(U3518) );
  INV_X1 U4055 ( .A(n3188), .ZN(n3189) );
  AOI21_X1 U4056 ( .B1(n3190), .B2(n3187), .A(n3189), .ZN(n3194) );
  INV_X1 U4057 ( .A(n3738), .ZN(n3624) );
  AOI22_X1 U4058 ( .A1(n3719), .A2(n3191), .B1(n3624), .B2(n2712), .ZN(n3193)
         );
  INV_X1 U4059 ( .A(n3737), .ZN(n3625) );
  AOI22_X1 U4060 ( .A1(n3626), .A2(REG3_REG_2__SCAN_IN), .B1(n3625), .B2(n3235), .ZN(n3192) );
  OAI211_X1 U4061 ( .C1(n3194), .C2(n3746), .A(n3193), .B(n3192), .ZN(U3234)
         );
  AOI21_X1 U4062 ( .B1(n3196), .B2(n2354), .A(n3195), .ZN(n3219) );
  INV_X1 U4063 ( .A(n3197), .ZN(n3198) );
  XNOR2_X1 U4064 ( .A(n3821), .B(n3198), .ZN(n3206) );
  INV_X1 U4065 ( .A(n3206), .ZN(n3222) );
  NOR2_X1 U4066 ( .A1(n3222), .A2(n4605), .ZN(n3209) );
  NAND2_X1 U4067 ( .A1(n3821), .A2(n3199), .ZN(n3200) );
  NAND2_X1 U4068 ( .A1(n3243), .A2(n3200), .ZN(n3205) );
  NAND2_X1 U4069 ( .A1(n2138), .A2(n4272), .ZN(n3202) );
  NAND2_X1 U4070 ( .A1(n2730), .A2(n4230), .ZN(n3201) );
  OAI211_X1 U4071 ( .C1(n4267), .C2(n3203), .A(n3202), .B(n3201), .ZN(n3204)
         );
  AOI21_X1 U4072 ( .B1(n3205), .B2(n3995), .A(n3204), .ZN(n3208) );
  NAND2_X1 U4073 ( .A1(n3206), .A2(n4265), .ZN(n3207) );
  NAND2_X1 U4074 ( .A1(n3208), .A2(n3207), .ZN(n3217) );
  AOI211_X1 U4075 ( .C1(n4610), .C2(n3219), .A(n3209), .B(n3217), .ZN(n4573)
         );
  NAND2_X1 U4076 ( .A1(n4619), .A2(REG1_REG_1__SCAN_IN), .ZN(n3210) );
  OAI21_X1 U4077 ( .B1(n4573), .B2(n4619), .A(n3210), .ZN(U3519) );
  NAND3_X1 U4078 ( .A1(n3213), .A2(n3212), .A3(n3211), .ZN(n3214) );
  INV_X2 U4079 ( .A(n4236), .ZN(n4285) );
  OR2_X1 U4080 ( .A1(n3215), .A2(n3985), .ZN(n3295) );
  INV_X1 U4081 ( .A(n3295), .ZN(n3216) );
  NAND2_X1 U4082 ( .A1(n4556), .A2(n3216), .ZN(n4164) );
  MUX2_X1 U4083 ( .A(REG2_REG_1__SCAN_IN), .B(n3217), .S(n4556), .Z(n3218) );
  INV_X1 U4084 ( .A(n3218), .ZN(n3221) );
  AOI22_X1 U4085 ( .A1(n3219), .A2(n4445), .B1(REG3_REG_1__SCAN_IN), .B2(n4552), .ZN(n3220) );
  OAI211_X1 U4086 ( .C1(n3222), .C2(n4164), .A(n3221), .B(n3220), .ZN(U3289)
         );
  XNOR2_X1 U4087 ( .A(n3223), .B(n3224), .ZN(n3225) );
  NAND2_X1 U4088 ( .A1(n3225), .A2(n3716), .ZN(n3230) );
  INV_X1 U4089 ( .A(n2730), .ZN(n3226) );
  INV_X1 U4090 ( .A(n3258), .ZN(n3337) );
  OAI22_X1 U4091 ( .A1(n3226), .A2(n3738), .B1(n3337), .B2(n3737), .ZN(n3227)
         );
  AOI211_X1 U4092 ( .C1(n3269), .C2(n3719), .A(n3228), .B(n3227), .ZN(n3229)
         );
  OAI211_X1 U4093 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3722), .A(n3230), .B(n3229), 
        .ZN(U3215) );
  AOI21_X1 U4094 ( .B1(n3231), .B2(n3232), .A(n3746), .ZN(n3234) );
  NAND2_X1 U4095 ( .A1(n3234), .A2(n3233), .ZN(n3239) );
  AND2_X1 U4096 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3937) );
  INV_X1 U4097 ( .A(n3911), .ZN(n3312) );
  INV_X1 U4098 ( .A(n3235), .ZN(n3321) );
  OAI22_X1 U4099 ( .A1(n3312), .A2(n3737), .B1(n3321), .B2(n3738), .ZN(n3236)
         );
  AOI211_X1 U4100 ( .C1(n3237), .C2(n3719), .A(n3937), .B(n3236), .ZN(n3238)
         );
  OAI211_X1 U4101 ( .C1(n3722), .C2(n3328), .A(n3239), .B(n3238), .ZN(U3227)
         );
  OAI21_X1 U4102 ( .B1(n3240), .B2(n3242), .A(n3241), .ZN(n3305) );
  INV_X1 U4103 ( .A(n3305), .ZN(n3249) );
  OAI22_X1 U4104 ( .A1(n3321), .A2(n4268), .B1(n3250), .B2(n4267), .ZN(n3247)
         );
  NAND3_X1 U4105 ( .A1(n3243), .A2(n3242), .A3(n3832), .ZN(n3244) );
  AOI21_X1 U4106 ( .B1(n3245), .B2(n3244), .A(n4275), .ZN(n3246) );
  AOI211_X1 U4107 ( .C1(n4272), .C2(n2712), .A(n3247), .B(n3246), .ZN(n3248)
         );
  OAI21_X1 U4108 ( .B1(n3249), .B2(n4153), .A(n3248), .ZN(n3302) );
  AOI21_X1 U4109 ( .B1(n4583), .B2(n3305), .A(n3302), .ZN(n3255) );
  OAI21_X1 U4110 ( .B1(n3195), .B2(n3250), .A(n3270), .ZN(n3301) );
  INV_X1 U4111 ( .A(n3301), .ZN(n3253) );
  AOI22_X1 U4112 ( .A1(n3253), .A2(n4311), .B1(REG1_REG_2__SCAN_IN), .B2(n4619), .ZN(n3251) );
  OAI21_X1 U4113 ( .B1(n3255), .B2(n4619), .A(n3251), .ZN(U3520) );
  INV_X1 U4114 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4737) );
  NOR2_X1 U4115 ( .A1(n4613), .A2(n4737), .ZN(n3252) );
  AOI21_X1 U4116 ( .B1(n3253), .B2(n3459), .A(n3252), .ZN(n3254) );
  OAI21_X1 U4117 ( .B1(n3255), .B2(n4611), .A(n3254), .ZN(U3471) );
  OAI21_X1 U4118 ( .B1(n3815), .B2(n3257), .A(n3256), .ZN(n3263) );
  NAND2_X1 U4119 ( .A1(n2730), .A2(n4272), .ZN(n3260) );
  NAND2_X1 U4120 ( .A1(n3258), .A2(n4230), .ZN(n3259) );
  OAI211_X1 U4121 ( .C1(n4267), .C2(n3261), .A(n3260), .B(n3259), .ZN(n3262)
         );
  AOI21_X1 U4122 ( .B1(n3263), .B2(n3995), .A(n3262), .ZN(n3267) );
  INV_X1 U4123 ( .A(n3815), .ZN(n3265) );
  XNOR2_X1 U4124 ( .A(n3264), .B(n3265), .ZN(n4575) );
  NAND2_X1 U4125 ( .A1(n4575), .A2(n4265), .ZN(n3266) );
  AND2_X1 U4126 ( .A1(n3267), .A2(n3266), .ZN(n4577) );
  INV_X1 U4127 ( .A(n4164), .ZN(n4553) );
  AND2_X1 U4128 ( .A1(n3270), .A2(n3269), .ZN(n3271) );
  NOR2_X1 U4129 ( .A1(n3268), .A2(n3271), .ZN(n4574) );
  INV_X1 U4130 ( .A(n4574), .ZN(n3273) );
  AOI22_X1 U4131 ( .A1(n4285), .A2(REG2_REG_3__SCAN_IN), .B1(n4552), .B2(n2389), .ZN(n3272) );
  OAI21_X1 U4132 ( .B1(n3273), .B2(n4282), .A(n3272), .ZN(n3274) );
  AOI21_X1 U4133 ( .B1(n4575), .B2(n4553), .A(n3274), .ZN(n3275) );
  OAI21_X1 U4134 ( .B1(n4577), .B2(n4285), .A(n3275), .ZN(U3287) );
  OAI211_X1 U4135 ( .C1(n3278), .C2(n3277), .A(n3276), .B(n3716), .ZN(n3282)
         );
  INV_X1 U4136 ( .A(n3910), .ZN(n3378) );
  OAI22_X1 U4137 ( .A1(n3337), .A2(n3738), .B1(n3378), .B2(n3737), .ZN(n3279)
         );
  AOI211_X1 U4138 ( .C1(n3341), .C2(n3719), .A(n3280), .B(n3279), .ZN(n3281)
         );
  OAI211_X1 U4139 ( .C1(n3722), .C2(n3342), .A(n3282), .B(n3281), .ZN(U3224)
         );
  NAND2_X1 U4140 ( .A1(n2635), .A2(n3844), .ZN(n3819) );
  XNOR2_X1 U4141 ( .A(n3283), .B(n3819), .ZN(n3286) );
  AOI22_X1 U4142 ( .A1(n3909), .A2(n4230), .B1(n4299), .B2(n3315), .ZN(n3284)
         );
  OAI21_X1 U4143 ( .B1(n3312), .B2(n4234), .A(n3284), .ZN(n3285) );
  AOI21_X1 U4144 ( .B1(n3286), .B2(n3995), .A(n3285), .ZN(n3346) );
  AND2_X1 U4145 ( .A1(n3340), .A2(n3315), .ZN(n3288) );
  NOR2_X1 U4146 ( .A1(n3287), .A2(n3288), .ZN(n3352) );
  OAI22_X1 U4147 ( .A1(n4556), .A2(n3289), .B1(n3318), .B2(n4242), .ZN(n3298)
         );
  NAND2_X1 U4148 ( .A1(n3333), .A2(n3291), .ZN(n3293) );
  AND2_X1 U4149 ( .A1(n3293), .A2(n3292), .ZN(n3294) );
  XNOR2_X1 U4150 ( .A(n3294), .B(n3819), .ZN(n3347) );
  NAND2_X1 U4151 ( .A1(n4153), .A2(n3295), .ZN(n3296) );
  NOR2_X1 U4152 ( .A1(n3347), .A2(n4257), .ZN(n3297) );
  AOI211_X1 U4153 ( .C1(n3352), .C2(n4445), .A(n3298), .B(n3297), .ZN(n3299)
         );
  OAI21_X1 U4154 ( .B1(n4285), .B2(n3346), .A(n3299), .ZN(U3284) );
  OAI22_X1 U4155 ( .A1(n4282), .A2(n3301), .B1(n3300), .B2(n4242), .ZN(n3304)
         );
  MUX2_X1 U4156 ( .A(REG2_REG_2__SCAN_IN), .B(n3302), .S(n4556), .Z(n3303) );
  AOI211_X1 U4157 ( .C1(n4553), .C2(n3305), .A(n3304), .B(n3303), .ZN(n3306)
         );
  INV_X1 U4158 ( .A(n3306), .ZN(U3288) );
  XNOR2_X1 U4159 ( .A(n3308), .B(n3307), .ZN(n3309) );
  XNOR2_X1 U4160 ( .A(n3310), .B(n3309), .ZN(n3311) );
  NAND2_X1 U4161 ( .A1(n3311), .A2(n3716), .ZN(n3317) );
  OAI22_X1 U4162 ( .A1(n3312), .A2(n3738), .B1(n2431), .B2(n3737), .ZN(n3313)
         );
  AOI211_X1 U4163 ( .C1(n3315), .C2(n3719), .A(n3314), .B(n3313), .ZN(n3316)
         );
  OAI211_X1 U4164 ( .C1(n3722), .C2(n3318), .A(n3317), .B(n3316), .ZN(U3236)
         );
  NAND2_X1 U4165 ( .A1(n3290), .A2(n3813), .ZN(n3319) );
  NAND2_X1 U4166 ( .A1(n3333), .A2(n3319), .ZN(n4579) );
  XOR2_X1 U4167 ( .A(n3813), .B(n3320), .Z(n3325) );
  OAI22_X1 U4168 ( .A1(n3321), .A2(n4234), .B1(n3327), .B2(n4267), .ZN(n3323)
         );
  NOR2_X1 U4169 ( .A1(n4579), .A2(n4153), .ZN(n3322) );
  AOI211_X1 U4170 ( .C1(n4230), .C2(n3911), .A(n3323), .B(n3322), .ZN(n3324)
         );
  OAI21_X1 U4171 ( .B1(n4275), .B2(n3325), .A(n3324), .ZN(n4581) );
  OAI211_X1 U4172 ( .C1(n3268), .C2(n3327), .A(n3326), .B(n4610), .ZN(n4580)
         );
  OAI22_X1 U4173 ( .A1(n4580), .A2(n4434), .B1(n4242), .B2(n3328), .ZN(n3329)
         );
  OAI21_X1 U4174 ( .B1(n4581), .B2(n3329), .A(n4236), .ZN(n3331) );
  NAND2_X1 U4175 ( .A1(n4285), .A2(REG2_REG_4__SCAN_IN), .ZN(n3330) );
  OAI211_X1 U4176 ( .C1(n4579), .C2(n4164), .A(n3331), .B(n3330), .ZN(U3286)
         );
  NAND2_X1 U4177 ( .A1(n3333), .A2(n3332), .ZN(n3334) );
  XOR2_X1 U4178 ( .A(n3804), .B(n3334), .Z(n4586) );
  XOR2_X1 U4179 ( .A(n3335), .B(n3804), .Z(n3339) );
  AOI22_X1 U4180 ( .A1(n3910), .A2(n4230), .B1(n4299), .B2(n3341), .ZN(n3336)
         );
  OAI21_X1 U4181 ( .B1(n3337), .B2(n4234), .A(n3336), .ZN(n3338) );
  AOI21_X1 U4182 ( .B1(n3339), .B2(n3995), .A(n3338), .ZN(n4587) );
  MUX2_X1 U4183 ( .A(n4587), .B(n3112), .S(n4285), .Z(n3345) );
  AOI21_X1 U4184 ( .B1(n3341), .B2(n3326), .A(n2253), .ZN(n4590) );
  INV_X1 U4185 ( .A(n3342), .ZN(n3343) );
  AOI22_X1 U4186 ( .A1(n4590), .A2(n4445), .B1(n3343), .B2(n4552), .ZN(n3344)
         );
  OAI211_X1 U4187 ( .C1(n4257), .C2(n4586), .A(n3345), .B(n3344), .ZN(U3285)
         );
  INV_X1 U4188 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3350) );
  OAI21_X1 U4189 ( .B1(n4591), .B2(n3347), .A(n3346), .ZN(n3351) );
  NAND2_X1 U4190 ( .A1(n3351), .A2(n4621), .ZN(n3349) );
  NAND2_X1 U4191 ( .A1(n3352), .A2(n4311), .ZN(n3348) );
  OAI211_X1 U4192 ( .C1(n4621), .C2(n3350), .A(n3349), .B(n3348), .ZN(U3524)
         );
  INV_X1 U4193 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4861) );
  NAND2_X1 U4194 ( .A1(n3351), .A2(n4613), .ZN(n3354) );
  NAND2_X1 U4195 ( .A1(n3352), .A2(n3459), .ZN(n3353) );
  OAI211_X1 U4196 ( .C1(n4613), .C2(n4861), .A(n3354), .B(n3353), .ZN(U3479)
         );
  XNOR2_X1 U4197 ( .A(n3355), .B(n3356), .ZN(n3357) );
  NAND2_X1 U4198 ( .A1(n3357), .A2(n3995), .ZN(n3360) );
  NOR2_X1 U4199 ( .A1(n3361), .A2(n4267), .ZN(n3358) );
  AOI21_X1 U4200 ( .B1(n3908), .B2(n4230), .A(n3358), .ZN(n3359) );
  OAI211_X1 U4201 ( .C1(n3378), .C2(n4234), .A(n3360), .B(n3359), .ZN(n4593)
         );
  INV_X1 U4202 ( .A(n4593), .ZN(n3374) );
  OAI21_X1 U4203 ( .B1(n3287), .B2(n3361), .A(n4610), .ZN(n3363) );
  NOR2_X1 U4204 ( .A1(n3363), .A2(n3362), .ZN(n4594) );
  OAI22_X1 U4205 ( .A1(n4556), .A2(n3364), .B1(n3384), .B2(n4242), .ZN(n3372)
         );
  NAND2_X1 U4206 ( .A1(n3365), .A2(n3366), .ZN(n3368) );
  NAND2_X1 U4207 ( .A1(n3368), .A2(n3367), .ZN(n3369) );
  INV_X1 U4208 ( .A(n4595), .ZN(n3370) );
  AND2_X1 U4209 ( .A1(n3369), .A2(n3356), .ZN(n4592) );
  NOR3_X1 U4210 ( .A1(n3370), .A2(n4592), .A3(n4257), .ZN(n3371) );
  AOI211_X1 U4211 ( .C1(n4204), .C2(n4594), .A(n3372), .B(n3371), .ZN(n3373)
         );
  OAI21_X1 U4212 ( .B1(n4285), .B2(n3374), .A(n3373), .ZN(U3283) );
  NAND2_X1 U4213 ( .A1(n3376), .A2(n3375), .ZN(n3411) );
  XOR2_X1 U4214 ( .A(n3410), .B(n3411), .Z(n3377) );
  NAND2_X1 U4215 ( .A1(n3377), .A2(n3716), .ZN(n3383) );
  INV_X1 U4216 ( .A(n3908), .ZN(n3427) );
  OAI22_X1 U4217 ( .A1(n3427), .A2(n3737), .B1(n3378), .B2(n3738), .ZN(n3379)
         );
  AOI211_X1 U4218 ( .C1(n3381), .C2(n3719), .A(n3380), .B(n3379), .ZN(n3382)
         );
  OAI211_X1 U4219 ( .C1(n3722), .C2(n3384), .A(n3383), .B(n3382), .ZN(U3210)
         );
  XNOR2_X1 U4220 ( .A(n3385), .B(n3386), .ZN(n3387) );
  NAND2_X1 U4221 ( .A1(n3387), .A2(n3716), .ZN(n3392) );
  INV_X1 U4222 ( .A(n3906), .ZN(n3388) );
  OAI22_X1 U4223 ( .A1(n3427), .A2(n3738), .B1(n3388), .B2(n3737), .ZN(n3389)
         );
  AOI211_X1 U4224 ( .C1(n3425), .C2(n3719), .A(n3390), .B(n3389), .ZN(n3391)
         );
  OAI211_X1 U4225 ( .C1(n3722), .C2(n3432), .A(n3392), .B(n3391), .ZN(U3228)
         );
  INV_X1 U4226 ( .A(n3805), .ZN(n3394) );
  XNOR2_X1 U4227 ( .A(n3393), .B(n3394), .ZN(n3398) );
  NAND2_X1 U4228 ( .A1(n3909), .A2(n4272), .ZN(n3396) );
  NAND2_X1 U4229 ( .A1(n3907), .A2(n4230), .ZN(n3395) );
  OAI211_X1 U4230 ( .C1(n4267), .C2(n3404), .A(n3396), .B(n3395), .ZN(n3397)
         );
  AOI21_X1 U4231 ( .B1(n3398), .B2(n3995), .A(n3397), .ZN(n3402) );
  NAND2_X1 U4232 ( .A1(n4595), .A2(n3399), .ZN(n3400) );
  XNOR2_X1 U4233 ( .A(n3400), .B(n3805), .ZN(n3445) );
  NAND2_X1 U4234 ( .A1(n3445), .A2(n4265), .ZN(n3401) );
  OR2_X1 U4235 ( .A1(n3362), .A2(n3404), .ZN(n3405) );
  NAND2_X1 U4236 ( .A1(n3403), .A2(n3405), .ZN(n3463) );
  NOR2_X1 U4237 ( .A1(n3463), .A2(n4282), .ZN(n3408) );
  INV_X1 U4238 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3406) );
  OAI22_X1 U4239 ( .A1(n4556), .A2(n3406), .B1(n3422), .B2(n4242), .ZN(n3407)
         );
  AOI211_X1 U4240 ( .C1(n3445), .C2(n4553), .A(n3408), .B(n3407), .ZN(n3409)
         );
  OAI21_X1 U4241 ( .B1(n3447), .B2(n4285), .A(n3409), .ZN(U3282) );
  NAND2_X1 U4242 ( .A1(n3411), .A2(n3410), .ZN(n3413) );
  NAND2_X1 U4243 ( .A1(n3413), .A2(n3412), .ZN(n3416) );
  NAND2_X1 U4244 ( .A1(n2178), .A2(n3414), .ZN(n3415) );
  XNOR2_X1 U4245 ( .A(n3416), .B(n3415), .ZN(n3417) );
  NAND2_X1 U4246 ( .A1(n3417), .A2(n3716), .ZN(n3421) );
  NOR2_X1 U4247 ( .A1(STATE_REG_SCAN_IN), .A2(n2419), .ZN(n4452) );
  INV_X1 U4248 ( .A(n3907), .ZN(n3441) );
  OAI22_X1 U4249 ( .A1(n2431), .A2(n3738), .B1(n3441), .B2(n3737), .ZN(n3418)
         );
  AOI211_X1 U4250 ( .C1(n3419), .C2(n3719), .A(n4452), .B(n3418), .ZN(n3420)
         );
  OAI211_X1 U4251 ( .C1(n3722), .C2(n3422), .A(n3421), .B(n3420), .ZN(U3218)
         );
  INV_X1 U4252 ( .A(n3855), .ZN(n3423) );
  AND2_X1 U4253 ( .A1(n3423), .A2(n3852), .ZN(n3807) );
  XOR2_X1 U4254 ( .A(n3807), .B(n3424), .Z(n3429) );
  AOI22_X1 U4255 ( .A1(n3906), .A2(n4230), .B1(n4299), .B2(n3425), .ZN(n3426)
         );
  OAI21_X1 U4256 ( .B1(n3427), .B2(n4234), .A(n3426), .ZN(n3428) );
  AOI21_X1 U4257 ( .B1(n3429), .B2(n3995), .A(n3428), .ZN(n4598) );
  XNOR2_X1 U4258 ( .A(n3430), .B(n3807), .ZN(n4603) );
  OAI21_X1 U4259 ( .B1(n2705), .B2(n3431), .A(n3471), .ZN(n4599) );
  NOR2_X1 U4260 ( .A1(n4599), .A2(n4282), .ZN(n3435) );
  OAI22_X1 U4261 ( .A1(n4556), .A2(n3433), .B1(n3432), .B2(n4242), .ZN(n3434)
         );
  AOI211_X1 U4262 ( .C1(n4603), .C2(n4019), .A(n3435), .B(n3434), .ZN(n3436)
         );
  OAI21_X1 U4263 ( .B1(n4598), .B2(n4285), .A(n3436), .ZN(U3281) );
  AOI21_X1 U4264 ( .B1(n3437), .B2(n3438), .A(n3746), .ZN(n3440) );
  NAND2_X1 U4265 ( .A1(n3440), .A2(n3439), .ZN(n3444) );
  AND2_X1 U4266 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n4461) );
  INV_X1 U4267 ( .A(n3905), .ZN(n3521) );
  OAI22_X1 U4268 ( .A1(n3441), .A2(n3738), .B1(n3521), .B2(n3737), .ZN(n3442)
         );
  AOI211_X1 U4269 ( .C1(n3470), .C2(n3719), .A(n4461), .B(n3442), .ZN(n3443)
         );
  OAI211_X1 U4270 ( .C1(n3722), .C2(n3473), .A(n3444), .B(n3443), .ZN(U3214)
         );
  NAND2_X1 U4271 ( .A1(n3445), .A2(n4583), .ZN(n3446) );
  NAND2_X1 U4272 ( .A1(n3447), .A2(n3446), .ZN(n3460) );
  MUX2_X1 U4273 ( .A(REG1_REG_8__SCAN_IN), .B(n3460), .S(n4621), .Z(n3448) );
  INV_X1 U4274 ( .A(n3448), .ZN(n3449) );
  OAI21_X1 U4275 ( .B1(n3463), .B2(n4376), .A(n3449), .ZN(U3526) );
  XOR2_X1 U4276 ( .A(n3451), .B(n3450), .Z(n3452) );
  XNOR2_X1 U4277 ( .A(n3453), .B(n3452), .ZN(n3458) );
  INV_X1 U4278 ( .A(n3497), .ZN(n3456) );
  AOI22_X1 U4279 ( .A1(n3625), .A2(n4271), .B1(n3624), .B2(n3906), .ZN(n3454)
         );
  NAND2_X1 U4280 ( .A1(REG3_REG_11__SCAN_IN), .A2(U3149), .ZN(n4469) );
  OAI211_X1 U4281 ( .C1(n3740), .C2(n3490), .A(n3454), .B(n4469), .ZN(n3455)
         );
  AOI21_X1 U4282 ( .B1(n3456), .B2(n3743), .A(n3455), .ZN(n3457) );
  OAI21_X1 U4283 ( .B1(n3458), .B2(n3746), .A(n3457), .ZN(U3233) );
  INV_X1 U4284 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4739) );
  INV_X1 U4285 ( .A(n3460), .ZN(n3461) );
  MUX2_X1 U4286 ( .A(n4739), .B(n3461), .S(n4613), .Z(n3462) );
  OAI21_X1 U4287 ( .B1(n3463), .B2(n4425), .A(n3462), .ZN(U3483) );
  XOR2_X1 U4288 ( .A(n3806), .B(n3464), .Z(n3468) );
  OAI22_X1 U4289 ( .A1(n3521), .A2(n4268), .B1(n4267), .B2(n3465), .ZN(n3466)
         );
  AOI21_X1 U4290 ( .B1(n4272), .B2(n3907), .A(n3466), .ZN(n3467) );
  OAI21_X1 U4291 ( .B1(n3468), .B2(n4275), .A(n3467), .ZN(n3527) );
  INV_X1 U4292 ( .A(n3527), .ZN(n3478) );
  XOR2_X1 U4293 ( .A(n3469), .B(n3806), .Z(n3528) );
  NAND2_X1 U4294 ( .A1(n3471), .A2(n3470), .ZN(n3472) );
  NAND2_X1 U4295 ( .A1(n3495), .A2(n3472), .ZN(n3533) );
  NOR2_X1 U4296 ( .A1(n3533), .A2(n4282), .ZN(n3476) );
  INV_X1 U4297 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3474) );
  OAI22_X1 U4298 ( .A1(n4236), .A2(n3474), .B1(n3473), .B2(n4242), .ZN(n3475)
         );
  AOI211_X1 U4299 ( .C1(n3528), .C2(n4019), .A(n3476), .B(n3475), .ZN(n3477)
         );
  OAI21_X1 U4300 ( .B1(n3478), .B2(n4285), .A(n3477), .ZN(U3280) );
  OR2_X1 U4301 ( .A1(n3469), .A2(n3479), .ZN(n3482) );
  NAND2_X1 U4302 ( .A1(n3482), .A2(n3480), .ZN(n3485) );
  NAND2_X1 U4303 ( .A1(n3482), .A2(n3481), .ZN(n3483) );
  NAND2_X1 U4304 ( .A1(n3483), .A2(n3487), .ZN(n3484) );
  NAND2_X1 U4305 ( .A1(n3485), .A2(n3484), .ZN(n3492) );
  INV_X1 U4306 ( .A(n3492), .ZN(n4606) );
  XNOR2_X1 U4307 ( .A(n3486), .B(n2467), .ZN(n3494) );
  NAND2_X1 U4308 ( .A1(n3906), .A2(n4272), .ZN(n3489) );
  NAND2_X1 U4309 ( .A1(n4271), .A2(n4230), .ZN(n3488) );
  OAI211_X1 U4310 ( .C1(n4267), .C2(n3490), .A(n3489), .B(n3488), .ZN(n3491)
         );
  AOI21_X1 U4311 ( .B1(n3492), .B2(n4265), .A(n3491), .ZN(n3493) );
  OAI21_X1 U4312 ( .B1(n4275), .B2(n3494), .A(n3493), .ZN(n4607) );
  NAND2_X1 U4313 ( .A1(n4607), .A2(n4236), .ZN(n3500) );
  AOI21_X1 U4314 ( .B1(n3496), .B2(n3495), .A(n3511), .ZN(n4609) );
  OAI22_X1 U4315 ( .A1(n4556), .A2(n3956), .B1(n3497), .B2(n4242), .ZN(n3498)
         );
  AOI21_X1 U4316 ( .B1(n4609), .B2(n4445), .A(n3498), .ZN(n3499) );
  OAI211_X1 U4317 ( .C1(n4606), .C2(n4164), .A(n3500), .B(n3499), .ZN(U3279)
         );
  INV_X1 U4318 ( .A(n3501), .ZN(n3502) );
  AOI21_X1 U4319 ( .B1(n3486), .B2(n3858), .A(n3502), .ZN(n4261) );
  AND2_X1 U4320 ( .A1(n4260), .A2(n4258), .ZN(n3801) );
  XNOR2_X1 U4321 ( .A(n4261), .B(n3508), .ZN(n3506) );
  NAND2_X1 U4322 ( .A1(n3905), .A2(n4272), .ZN(n3504) );
  NAND2_X1 U4323 ( .A1(n3904), .A2(n4230), .ZN(n3503) );
  OAI211_X1 U4324 ( .C1(n4267), .C2(n3510), .A(n3504), .B(n3503), .ZN(n3505)
         );
  AOI21_X1 U4325 ( .B1(n3506), .B2(n3995), .A(n3505), .ZN(n4373) );
  XNOR2_X1 U4326 ( .A(n3507), .B(n3508), .ZN(n4371) );
  OR2_X1 U4327 ( .A1(n3511), .A2(n3510), .ZN(n3512) );
  NAND2_X1 U4328 ( .A1(n3509), .A2(n3512), .ZN(n4426) );
  NOR2_X1 U4329 ( .A1(n4426), .A2(n4282), .ZN(n3515) );
  INV_X1 U4330 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3513) );
  OAI22_X1 U4331 ( .A1(n4236), .A2(n3513), .B1(n3526), .B2(n4242), .ZN(n3514)
         );
  AOI211_X1 U4332 ( .C1(n4371), .C2(n4019), .A(n3515), .B(n3514), .ZN(n3516)
         );
  OAI21_X1 U4333 ( .B1(n4373), .B2(n4285), .A(n3516), .ZN(U3278) );
  NAND2_X1 U4334 ( .A1(n2313), .A2(n3518), .ZN(n3519) );
  XNOR2_X1 U4335 ( .A(n3517), .B(n3519), .ZN(n3520) );
  NAND2_X1 U4336 ( .A1(n3520), .A2(n3716), .ZN(n3525) );
  NOR2_X1 U4337 ( .A1(STATE_REG_SCAN_IN), .A2(n2470), .ZN(n4625) );
  OAI22_X1 U4338 ( .A1(n3521), .A2(n3738), .B1(n3591), .B2(n3737), .ZN(n3522)
         );
  AOI211_X1 U4339 ( .C1(n3523), .C2(n3719), .A(n4625), .B(n3522), .ZN(n3524)
         );
  OAI211_X1 U4340 ( .C1(n3722), .C2(n3526), .A(n3525), .B(n3524), .ZN(U3221)
         );
  INV_X1 U4341 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3529) );
  AOI21_X1 U4342 ( .B1(n4602), .B2(n3528), .A(n3527), .ZN(n3531) );
  MUX2_X1 U4343 ( .A(n3529), .B(n3531), .S(n4613), .Z(n3530) );
  OAI21_X1 U4344 ( .B1(n3533), .B2(n4425), .A(n3530), .ZN(U3487) );
  INV_X1 U4345 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4878) );
  MUX2_X1 U4346 ( .A(n4878), .B(n3531), .S(n4621), .Z(n3532) );
  OAI21_X1 U4347 ( .B1(n3533), .B2(n4376), .A(n3532), .ZN(U3528) );
  XOR2_X1 U4348 ( .A(n3535), .B(n3534), .Z(n3536) );
  XNOR2_X1 U4349 ( .A(n3537), .B(n3536), .ZN(n3542) );
  INV_X1 U4350 ( .A(n3538), .ZN(n4280) );
  AOI22_X1 U4351 ( .A1(n3624), .A2(n4271), .B1(n3625), .B2(n4253), .ZN(n3539)
         );
  NAND2_X1 U4352 ( .A1(REG3_REG_13__SCAN_IN), .A2(U3149), .ZN(n4487) );
  OAI211_X1 U4353 ( .C1(n3740), .C2(n4266), .A(n3539), .B(n4487), .ZN(n3540)
         );
  AOI21_X1 U4354 ( .B1(n4280), .B2(n3743), .A(n3540), .ZN(n3541) );
  OAI21_X1 U4355 ( .B1(n3542), .B2(n3746), .A(n3541), .ZN(U3231) );
  OAI21_X1 U4356 ( .B1(n3545), .B2(n3544), .A(n3543), .ZN(n4365) );
  INV_X1 U4357 ( .A(n4365), .ZN(n3558) );
  XNOR2_X1 U4358 ( .A(n3546), .B(n3812), .ZN(n3547) );
  NAND2_X1 U4359 ( .A1(n3547), .A2(n3995), .ZN(n3551) );
  NOR2_X1 U4360 ( .A1(n3548), .A2(n4267), .ZN(n3549) );
  AOI21_X1 U4361 ( .B1(n3903), .B2(n4230), .A(n3549), .ZN(n3550) );
  OAI211_X1 U4362 ( .C1(n3591), .C2(n4234), .A(n3551), .B(n3550), .ZN(n4364)
         );
  INV_X1 U4363 ( .A(n4241), .ZN(n3553) );
  NAND2_X1 U4364 ( .A1(n4279), .A2(n3593), .ZN(n3552) );
  NAND2_X1 U4365 ( .A1(n3553), .A2(n3552), .ZN(n4418) );
  INV_X1 U4366 ( .A(n3596), .ZN(n3554) );
  AOI22_X1 U4367 ( .A1(n4285), .A2(REG2_REG_14__SCAN_IN), .B1(n3554), .B2(
        n4552), .ZN(n3555) );
  OAI21_X1 U4368 ( .B1(n4418), .B2(n4282), .A(n3555), .ZN(n3556) );
  AOI21_X1 U4369 ( .B1(n4364), .B2(n4236), .A(n3556), .ZN(n3557) );
  OAI21_X1 U4370 ( .B1(n3558), .B2(n4257), .A(n3557), .ZN(U3276) );
  INV_X1 U4371 ( .A(n3901), .ZN(n4051) );
  OAI22_X1 U4372 ( .A1(n4051), .A2(n4234), .B1(n3576), .B2(n4267), .ZN(n3565)
         );
  NAND2_X1 U4373 ( .A1(n3560), .A2(n3559), .ZN(n3563) );
  AOI21_X1 U4374 ( .B1(n3563), .B2(n3562), .A(n4275), .ZN(n3564) );
  XNOR2_X1 U4375 ( .A(n3566), .B(n3796), .ZN(n4315) );
  NAND2_X1 U4376 ( .A1(n4315), .A2(n4019), .ZN(n3572) );
  OAI21_X1 U4377 ( .B1(n3567), .B2(n3576), .A(n2142), .ZN(n4318) );
  INV_X1 U4378 ( .A(n4318), .ZN(n3570) );
  INV_X1 U4379 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3568) );
  OAI22_X1 U4380 ( .A1(n3575), .A2(n4242), .B1(n3568), .B2(n4236), .ZN(n3569)
         );
  AOI21_X1 U4381 ( .B1(n3570), .B2(n4445), .A(n3569), .ZN(n3571) );
  OAI211_X1 U4382 ( .C1(n4316), .C2(n4285), .A(n3572), .B(n3571), .ZN(U3263)
         );
  XNOR2_X1 U4383 ( .A(n3574), .B(n3573), .ZN(n3582) );
  INV_X1 U4384 ( .A(n3575), .ZN(n3580) );
  OAI22_X1 U4385 ( .A1(n3740), .A2(n3576), .B1(STATE_REG_SCAN_IN), .B2(n4891), 
        .ZN(n3579) );
  INV_X1 U4386 ( .A(n4007), .ZN(n3577) );
  OAI22_X1 U4387 ( .A1(n3577), .A2(n3737), .B1(n4051), .B2(n3738), .ZN(n3578)
         );
  AOI211_X1 U4388 ( .C1(n3580), .C2(n3743), .A(n3579), .B(n3578), .ZN(n3581)
         );
  OAI21_X1 U4389 ( .B1(n3582), .B2(n3746), .A(n3581), .ZN(U3211) );
  INV_X1 U4390 ( .A(n3583), .ZN(n3587) );
  OAI21_X1 U4391 ( .B1(n3587), .B2(n3585), .A(n3584), .ZN(n3586) );
  OAI21_X1 U4392 ( .B1(n3588), .B2(n3587), .A(n3586), .ZN(n3589) );
  NAND2_X1 U4393 ( .A1(n3589), .A2(n3716), .ZN(n3595) );
  NOR2_X1 U4394 ( .A1(STATE_REG_SCAN_IN), .A2(n3590), .ZN(n4497) );
  OAI22_X1 U4395 ( .A1(n4235), .A2(n3737), .B1(n3591), .B2(n3738), .ZN(n3592)
         );
  AOI211_X1 U4396 ( .C1(n3593), .C2(n3719), .A(n4497), .B(n3592), .ZN(n3594)
         );
  OAI211_X1 U4397 ( .C1(n3722), .C2(n3596), .A(n3595), .B(n3594), .ZN(U3212)
         );
  NAND2_X1 U4398 ( .A1(n3597), .A2(n3598), .ZN(n3676) );
  NAND2_X1 U4399 ( .A1(n3676), .A2(n3716), .ZN(n3606) );
  AOI21_X1 U4400 ( .B1(n3597), .B2(n3600), .A(n3599), .ZN(n3605) );
  INV_X1 U4401 ( .A(n4099), .ZN(n3603) );
  INV_X1 U4402 ( .A(n4092), .ZN(n3652) );
  OAI22_X1 U4403 ( .A1(n3642), .A2(n3738), .B1(n3652), .B2(n3737), .ZN(n3602)
         );
  INV_X1 U4404 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4653) );
  OAI22_X1 U4405 ( .A1(n3740), .A2(n4097), .B1(STATE_REG_SCAN_IN), .B2(n4653), 
        .ZN(n3601) );
  AOI211_X1 U4406 ( .C1(n3603), .C2(n3743), .A(n3602), .B(n3601), .ZN(n3604)
         );
  OAI21_X1 U4407 ( .B1(n3606), .B2(n3605), .A(n3604), .ZN(U3213) );
  NAND2_X1 U4408 ( .A1(n3607), .A2(n3608), .ZN(n3636) );
  INV_X1 U4409 ( .A(n3715), .ZN(n3610) );
  OAI21_X1 U4410 ( .B1(n3610), .B2(n3609), .A(n3713), .ZN(n3611) );
  OAI21_X1 U4411 ( .B1(n3712), .B2(n3715), .A(n3611), .ZN(n3615) );
  NAND2_X1 U4412 ( .A1(n3613), .A2(n3612), .ZN(n3614) );
  XNOR2_X1 U4413 ( .A(n3615), .B(n3614), .ZN(n3616) );
  NAND2_X1 U4414 ( .A1(n3616), .A2(n3716), .ZN(n3620) );
  AND2_X1 U4415 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3983) );
  OAI22_X1 U4416 ( .A1(n2544), .A2(n3738), .B1(n4174), .B2(n3737), .ZN(n3617)
         );
  AOI211_X1 U4417 ( .C1(n3618), .C2(n3719), .A(n3983), .B(n3617), .ZN(n3619)
         );
  OAI211_X1 U4418 ( .C1(n3722), .C2(n4182), .A(n3620), .B(n3619), .ZN(U3216)
         );
  OAI211_X1 U4419 ( .C1(n3621), .C2(n3623), .A(n3622), .B(n3716), .ZN(n3629)
         );
  AOI22_X1 U4420 ( .A1(n3719), .A2(n2354), .B1(n3624), .B2(n2138), .ZN(n3628)
         );
  AOI22_X1 U4421 ( .A1(n3626), .A2(REG3_REG_1__SCAN_IN), .B1(n3625), .B2(n2730), .ZN(n3627) );
  NAND3_X1 U4422 ( .A1(n3629), .A2(n3628), .A3(n3627), .ZN(U3219) );
  NAND2_X1 U4423 ( .A1(n3607), .A2(n3630), .ZN(n3632) );
  AND2_X1 U4424 ( .A1(n3632), .A2(n3631), .ZN(n3641) );
  NAND2_X1 U4425 ( .A1(n3634), .A2(n3633), .ZN(n3640) );
  NAND2_X1 U4426 ( .A1(n3636), .A2(n3635), .ZN(n3638) );
  NAND2_X1 U4427 ( .A1(n3638), .A2(n3637), .ZN(n3692) );
  OAI211_X1 U4428 ( .C1(n3692), .C2(n3690), .A(n3694), .B(n3640), .ZN(n3639)
         );
  OAI211_X1 U4429 ( .C1(n3641), .C2(n3640), .A(n3716), .B(n3639), .ZN(n3646)
         );
  OAI22_X1 U4430 ( .A1(n3740), .A2(n4132), .B1(STATE_REG_SCAN_IN), .B2(n4898), 
        .ZN(n3644) );
  OAI22_X1 U4431 ( .A1(n4174), .A2(n3738), .B1(n3642), .B2(n3737), .ZN(n3643)
         );
  NOR2_X1 U4432 ( .A1(n3644), .A2(n3643), .ZN(n3645) );
  OAI211_X1 U4433 ( .C1(n3722), .C2(n4134), .A(n3646), .B(n3645), .ZN(U3220)
         );
  NAND2_X1 U4434 ( .A1(n3648), .A2(n3647), .ZN(n3650) );
  XOR2_X1 U4435 ( .A(n3650), .B(n3649), .Z(n3657) );
  INV_X1 U4436 ( .A(n4057), .ZN(n3655) );
  OAI22_X1 U4437 ( .A1(n3740), .A2(n4055), .B1(STATE_REG_SCAN_IN), .B2(n3651), 
        .ZN(n3654) );
  OAI22_X1 U4438 ( .A1(n4051), .A2(n3737), .B1(n3652), .B2(n3738), .ZN(n3653)
         );
  AOI211_X1 U4439 ( .C1(n3655), .C2(n3743), .A(n3654), .B(n3653), .ZN(n3656)
         );
  OAI21_X1 U4440 ( .B1(n3657), .B2(n3746), .A(n3656), .ZN(U3222) );
  INV_X1 U4441 ( .A(n3734), .ZN(n3658) );
  OAI21_X1 U4442 ( .B1(n3658), .B2(n3736), .A(n3733), .ZN(n3660) );
  XNOR2_X1 U4443 ( .A(n3660), .B(n3659), .ZN(n3661) );
  NAND2_X1 U4444 ( .A1(n3661), .A2(n3716), .ZN(n3664) );
  NOR2_X1 U4445 ( .A1(STATE_REG_SCAN_IN), .A2(n2514), .ZN(n4512) );
  OAI22_X1 U4446 ( .A1(n4199), .A2(n3737), .B1(n4235), .B2(n3738), .ZN(n3662)
         );
  AOI211_X1 U4447 ( .C1(n2523), .C2(n3719), .A(n4512), .B(n3662), .ZN(n3663)
         );
  OAI211_X1 U4448 ( .C1(n3722), .C2(n4223), .A(n3664), .B(n3663), .ZN(U3223)
         );
  NAND2_X1 U4449 ( .A1(n3666), .A2(n3665), .ZN(n3669) );
  NAND2_X1 U4450 ( .A1(n3607), .A2(n3667), .ZN(n3668) );
  XOR2_X1 U4451 ( .A(n3669), .B(n3668), .Z(n3670) );
  NAND2_X1 U4452 ( .A1(n3670), .A2(n3716), .ZN(n3674) );
  NOR2_X1 U4453 ( .A1(STATE_REG_SCAN_IN), .A2(n4664), .ZN(n4521) );
  OAI22_X1 U4454 ( .A1(n4246), .A2(n3738), .B1(n2544), .B2(n3737), .ZN(n3671)
         );
  AOI211_X1 U4455 ( .C1(n3672), .C2(n3719), .A(n4521), .B(n3671), .ZN(n3673)
         );
  OAI211_X1 U4456 ( .C1(n3722), .C2(n4215), .A(n3674), .B(n3673), .ZN(U3225)
         );
  NAND2_X1 U4457 ( .A1(n3676), .A2(n3675), .ZN(n3677) );
  NAND2_X1 U4458 ( .A1(n3678), .A2(n3677), .ZN(n3679) );
  XOR2_X1 U4459 ( .A(n3680), .B(n3679), .Z(n3686) );
  INV_X1 U4460 ( .A(n3681), .ZN(n4077) );
  OAI22_X1 U4461 ( .A1(n3705), .A2(n3738), .B1(n4069), .B2(n3737), .ZN(n3684)
         );
  OAI22_X1 U4462 ( .A1(n3740), .A2(n4074), .B1(STATE_REG_SCAN_IN), .B2(n3682), 
        .ZN(n3683) );
  AOI211_X1 U4463 ( .C1(n4077), .C2(n3743), .A(n3684), .B(n3683), .ZN(n3685)
         );
  OAI21_X1 U4464 ( .B1(n3686), .B2(n3746), .A(n3685), .ZN(U3226) );
  NAND2_X1 U4465 ( .A1(n3607), .A2(n3687), .ZN(n3689) );
  NAND2_X1 U4466 ( .A1(n3689), .A2(n3688), .ZN(n3691) );
  NOR2_X1 U4467 ( .A1(n3691), .A2(n3690), .ZN(n3696) );
  AOI21_X1 U4468 ( .B1(n3694), .B2(n3693), .A(n3692), .ZN(n3695) );
  OAI21_X1 U4469 ( .B1(n3696), .B2(n3695), .A(n3716), .ZN(n3700) );
  INV_X1 U4470 ( .A(n4147), .ZN(n3704) );
  OAI22_X1 U4471 ( .A1(n4149), .A2(n3738), .B1(n3704), .B2(n3737), .ZN(n3698)
         );
  NOR2_X1 U4472 ( .A1(n3740), .A2(n4155), .ZN(n3697) );
  AOI211_X1 U4473 ( .C1(REG3_REG_20__SCAN_IN), .C2(U3149), .A(n3698), .B(n3697), .ZN(n3699) );
  OAI211_X1 U4474 ( .C1(n3722), .C2(n4158), .A(n3700), .B(n3699), .ZN(U3230)
         );
  INV_X1 U4475 ( .A(n3597), .ZN(n3702) );
  AOI21_X1 U4476 ( .B1(n3703), .B2(n3701), .A(n3702), .ZN(n3711) );
  INV_X1 U4477 ( .A(n4109), .ZN(n3709) );
  OAI22_X1 U4478 ( .A1(n3705), .A2(n3737), .B1(n3704), .B2(n3738), .ZN(n3708)
         );
  OAI22_X1 U4479 ( .A1(n3740), .A2(n4119), .B1(STATE_REG_SCAN_IN), .B2(n3706), 
        .ZN(n3707) );
  AOI211_X1 U4480 ( .C1(n3709), .C2(n3743), .A(n3708), .B(n3707), .ZN(n3710)
         );
  OAI21_X1 U4481 ( .B1(n3711), .B2(n3746), .A(n3710), .ZN(U3232) );
  XNOR2_X1 U4482 ( .A(n3713), .B(n3712), .ZN(n3714) );
  XNOR2_X1 U4483 ( .A(n3715), .B(n3714), .ZN(n3717) );
  NAND2_X1 U4484 ( .A1(n3717), .A2(n3716), .ZN(n3721) );
  INV_X1 U4485 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4842) );
  NOR2_X1 U4486 ( .A1(STATE_REG_SCAN_IN), .A2(n4842), .ZN(n4544) );
  OAI22_X1 U4487 ( .A1(n4149), .A2(n3737), .B1(n4199), .B2(n3738), .ZN(n3718)
         );
  AOI211_X1 U4488 ( .C1(n4196), .C2(n3719), .A(n4544), .B(n3718), .ZN(n3720)
         );
  OAI211_X1 U4489 ( .C1(n3722), .C2(n4193), .A(n3721), .B(n3720), .ZN(U3235)
         );
  INV_X1 U4490 ( .A(n3724), .ZN(n3726) );
  NOR2_X1 U4491 ( .A1(n3726), .A2(n3725), .ZN(n3727) );
  XNOR2_X1 U4492 ( .A(n3723), .B(n3727), .ZN(n3732) );
  INV_X1 U4493 ( .A(n3728), .ZN(n4042) );
  OAI22_X1 U4494 ( .A1(n3740), .A2(n4040), .B1(STATE_REG_SCAN_IN), .B2(n4920), 
        .ZN(n3730) );
  OAI22_X1 U4495 ( .A1(n4034), .A2(n3737), .B1(n4069), .B2(n3738), .ZN(n3729)
         );
  AOI211_X1 U4496 ( .C1(n4042), .C2(n3743), .A(n3730), .B(n3729), .ZN(n3731)
         );
  OAI21_X1 U4497 ( .B1(n3732), .B2(n3746), .A(n3731), .ZN(U3237) );
  NAND2_X1 U4498 ( .A1(n3734), .A2(n3733), .ZN(n3735) );
  XOR2_X1 U4499 ( .A(n3736), .B(n3735), .Z(n3747) );
  INV_X1 U4500 ( .A(n4243), .ZN(n3744) );
  INV_X1 U4501 ( .A(n4253), .ZN(n4269) );
  OAI22_X1 U4502 ( .A1(n4269), .A2(n3738), .B1(n4246), .B2(n3737), .ZN(n3742)
         );
  INV_X1 U4503 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3739) );
  OAI22_X1 U4504 ( .A1(n3740), .A2(n4245), .B1(STATE_REG_SCAN_IN), .B2(n3739), 
        .ZN(n3741) );
  AOI211_X1 U4505 ( .C1(n3744), .C2(n3743), .A(n3742), .B(n3741), .ZN(n3745)
         );
  OAI21_X1 U4506 ( .B1(n3747), .B2(n3746), .A(n3745), .ZN(U3238) );
  NAND2_X1 U4507 ( .A1(n2416), .A2(DATAI_29_), .ZN(n4011) );
  NOR2_X1 U4508 ( .A1(n3748), .A2(n4014), .ZN(n3749) );
  NOR2_X1 U4509 ( .A1(n3749), .A2(n3992), .ZN(n3879) );
  OR2_X1 U4510 ( .A1(n3751), .A2(n3750), .ZN(n3762) );
  NOR2_X1 U4511 ( .A1(n3900), .A2(n4011), .ZN(n3763) );
  NAND2_X1 U4512 ( .A1(n3755), .A2(REG1_REG_31__SCAN_IN), .ZN(n3754) );
  NAND2_X1 U4513 ( .A1(n3756), .A2(REG2_REG_31__SCAN_IN), .ZN(n3753) );
  NAND2_X1 U4514 ( .A1(n2141), .A2(REG0_REG_31__SCAN_IN), .ZN(n3752) );
  NAND3_X1 U4515 ( .A1(n3754), .A2(n3753), .A3(n3752), .ZN(n4291) );
  NAND2_X1 U4516 ( .A1(n2132), .A2(DATAI_31_), .ZN(n4289) );
  NAND2_X1 U4517 ( .A1(n4291), .A2(n4289), .ZN(n3885) );
  NAND2_X1 U4518 ( .A1(n3755), .A2(REG1_REG_30__SCAN_IN), .ZN(n3759) );
  NAND2_X1 U4519 ( .A1(n3756), .A2(REG2_REG_30__SCAN_IN), .ZN(n3758) );
  NAND2_X1 U4520 ( .A1(n2141), .A2(REG0_REG_30__SCAN_IN), .ZN(n3757) );
  NAND3_X1 U4521 ( .A1(n3759), .A2(n3758), .A3(n3757), .ZN(n3998) );
  NAND2_X1 U4522 ( .A1(n2132), .A2(DATAI_30_), .ZN(n4288) );
  OR2_X1 U4523 ( .A1(n3998), .A2(n4288), .ZN(n3760) );
  NAND2_X1 U4524 ( .A1(n3885), .A2(n3760), .ZN(n3820) );
  AOI211_X1 U4525 ( .C1(n3879), .C2(n3762), .A(n3763), .B(n3820), .ZN(n3884)
         );
  NAND3_X1 U4526 ( .A1(n3796), .A2(n3879), .A3(n3761), .ZN(n3782) );
  NOR4_X1 U4527 ( .A1(n3763), .A2(n3875), .A3(n3762), .A4(n3820), .ZN(n3781)
         );
  INV_X1 U4528 ( .A(n3866), .ZN(n3768) );
  NAND2_X1 U4529 ( .A1(n3764), .A2(n3767), .ZN(n3861) );
  NOR3_X1 U4530 ( .A1(n3546), .A2(n3768), .A3(n3861), .ZN(n3766) );
  INV_X1 U4531 ( .A(n3765), .ZN(n3868) );
  OAI21_X1 U4532 ( .B1(n3766), .B2(n3868), .A(n3867), .ZN(n3776) );
  INV_X1 U4533 ( .A(n3767), .ZN(n3769) );
  AOI211_X1 U4534 ( .C1(n3771), .C2(n3770), .A(n3769), .B(n3768), .ZN(n3773)
         );
  OAI21_X1 U4535 ( .B1(n3773), .B2(n3772), .A(n3867), .ZN(n3775) );
  AND2_X1 U4536 ( .A1(n3775), .A2(n3774), .ZN(n3871) );
  NAND2_X1 U4537 ( .A1(n3776), .A2(n3871), .ZN(n3778) );
  AOI21_X1 U4538 ( .B1(n3874), .B2(n3778), .A(n3777), .ZN(n3779) );
  OAI21_X1 U4539 ( .B1(n3779), .B2(n3876), .A(n4031), .ZN(n3780) );
  AOI22_X1 U4540 ( .A1(n3884), .A2(n3782), .B1(n3781), .B2(n3780), .ZN(n3787)
         );
  NOR2_X1 U4541 ( .A1(n4291), .A2(n4288), .ZN(n3786) );
  INV_X1 U4542 ( .A(n3998), .ZN(n3783) );
  INV_X1 U4543 ( .A(n4288), .ZN(n4300) );
  NOR2_X1 U4544 ( .A1(n3783), .A2(n4300), .ZN(n3789) );
  INV_X1 U4545 ( .A(n4291), .ZN(n3784) );
  NOR2_X1 U4546 ( .A1(n3789), .A2(n3784), .ZN(n3785) );
  OAI22_X1 U4547 ( .A1(n3787), .A2(n3786), .B1(n3785), .B2(n4289), .ZN(n3828)
         );
  NAND2_X1 U4548 ( .A1(n2171), .A2(n3788), .ZN(n4032) );
  NOR2_X1 U4549 ( .A1(n4291), .A2(n4289), .ZN(n3790) );
  NOR2_X1 U4550 ( .A1(n3790), .A2(n3789), .ZN(n3887) );
  AND2_X1 U4551 ( .A1(n4032), .A2(n3887), .ZN(n3795) );
  NAND2_X1 U4552 ( .A1(n3791), .A2(n4029), .ZN(n4050) );
  NAND2_X1 U4553 ( .A1(n3793), .A2(n3792), .ZN(n4173) );
  NOR2_X1 U4554 ( .A1(n4050), .A2(n4173), .ZN(n3794) );
  NAND4_X1 U4555 ( .A1(n3797), .A2(n3796), .A3(n3795), .A4(n3794), .ZN(n3811)
         );
  XNOR2_X1 U4556 ( .A(n3902), .B(n4155), .ZN(n4141) );
  INV_X1 U4557 ( .A(n4141), .ZN(n4144) );
  NAND2_X1 U4558 ( .A1(n2170), .A2(n4144), .ZN(n3810) );
  NAND2_X1 U4559 ( .A1(n3798), .A2(n4048), .ZN(n4068) );
  INV_X1 U4560 ( .A(n4068), .ZN(n3803) );
  NAND2_X1 U4561 ( .A1(n4064), .A2(n3799), .ZN(n4089) );
  INV_X1 U4562 ( .A(n4089), .ZN(n3802) );
  NAND4_X1 U4563 ( .A1(n3803), .A2(n3802), .A3(n4264), .A4(n3801), .ZN(n3809)
         );
  NAND4_X1 U4564 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3808)
         );
  NOR4_X1 U4565 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n3825)
         );
  INV_X1 U4566 ( .A(n4188), .ZN(n4194) );
  NAND4_X1 U4567 ( .A1(n3813), .A2(n3356), .A3(n4194), .A4(n3812), .ZN(n3817)
         );
  NAND2_X1 U4568 ( .A1(n3815), .A2(n3814), .ZN(n3816) );
  OR2_X1 U4569 ( .A1(n4085), .A2(n4084), .ZN(n4125) );
  NOR4_X1 U4570 ( .A1(n3817), .A2(n3816), .A3(n4125), .A4(n4250), .ZN(n3824)
         );
  INV_X1 U4571 ( .A(n4168), .ZN(n3818) );
  NAND2_X1 U4572 ( .A1(n3818), .A2(n4167), .ZN(n4208) );
  NOR4_X1 U4573 ( .A1(n4208), .A2(n3819), .A3(n4106), .A4(n4221), .ZN(n3823)
         );
  NOR4_X1 U4574 ( .A1(n2467), .A2(n3821), .A3(n4554), .A4(n3820), .ZN(n3822)
         );
  NAND4_X1 U4575 ( .A1(n3825), .A2(n3824), .A3(n3823), .A4(n3822), .ZN(n3827)
         );
  MUX2_X1 U4576 ( .A(n3828), .B(n3827), .S(n3826), .Z(n3892) );
  OAI211_X1 U4577 ( .C1(n3831), .C2(n4432), .A(n3830), .B(n3829), .ZN(n3834)
         );
  NAND3_X1 U4578 ( .A1(n3834), .A2(n3833), .A3(n3832), .ZN(n3837) );
  NAND3_X1 U4579 ( .A1(n3837), .A2(n3836), .A3(n3835), .ZN(n3840) );
  NAND3_X1 U4580 ( .A1(n3840), .A2(n3839), .A3(n3838), .ZN(n3843) );
  AND4_X1 U4581 ( .A1(n3843), .A2(n3842), .A3(n2635), .A4(n3841), .ZN(n3850)
         );
  OAI211_X1 U4582 ( .C1(n3846), .C2(n3845), .A(n3356), .B(n3844), .ZN(n3849)
         );
  OAI211_X1 U4583 ( .C1(n3850), .C2(n3849), .A(n3848), .B(n3847), .ZN(n3853)
         );
  AND3_X1 U4584 ( .A1(n3853), .A2(n3852), .A3(n3851), .ZN(n3856) );
  OAI21_X1 U4585 ( .B1(n3856), .B2(n3855), .A(n3854), .ZN(n3860) );
  NAND4_X1 U4586 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3865)
         );
  INV_X1 U4587 ( .A(n3861), .ZN(n3864) );
  AND4_X1 U4588 ( .A1(n3865), .A2(n3864), .A3(n3863), .A4(n3862), .ZN(n3869)
         );
  OAI211_X1 U4589 ( .C1(n3869), .C2(n3868), .A(n3867), .B(n3866), .ZN(n3872)
         );
  INV_X1 U4590 ( .A(n4084), .ZN(n3870) );
  NAND3_X1 U4591 ( .A1(n3872), .A2(n3871), .A3(n3870), .ZN(n3873) );
  NAND2_X1 U4592 ( .A1(n3874), .A2(n3873), .ZN(n3877) );
  AOI211_X1 U4593 ( .C1(n3878), .C2(n3877), .A(n3876), .B(n3875), .ZN(n3882)
         );
  INV_X1 U4594 ( .A(n3879), .ZN(n3880) );
  NOR4_X1 U4595 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3889)
         );
  INV_X1 U4596 ( .A(n3884), .ZN(n3888) );
  INV_X1 U4597 ( .A(n3885), .ZN(n3886) );
  OAI22_X1 U4598 ( .A1(n3889), .A2(n3888), .B1(n3887), .B2(n3886), .ZN(n3891)
         );
  MUX2_X1 U4599 ( .A(n3892), .B(n3891), .S(n3890), .Z(n3893) );
  XNOR2_X1 U4600 ( .A(n3893), .B(n3985), .ZN(n3899) );
  NAND2_X1 U4601 ( .A1(n3895), .A2(n3894), .ZN(n3896) );
  OAI211_X1 U4602 ( .C1(n4431), .C2(n3898), .A(n3896), .B(B_REG_SCAN_IN), .ZN(
        n3897) );
  OAI21_X1 U4603 ( .B1(n3899), .B2(n3898), .A(n3897), .ZN(U3239) );
  MUX2_X1 U4604 ( .A(DATAO_REG_31__SCAN_IN), .B(n4291), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4605 ( .A(DATAO_REG_30__SCAN_IN), .B(n3998), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4606 ( .A(n3900), .B(DATAO_REG_29__SCAN_IN), .S(n3912), .Z(U3579)
         );
  MUX2_X1 U4607 ( .A(n4007), .B(DATAO_REG_28__SCAN_IN), .S(n3912), .Z(U3578)
         );
  MUX2_X1 U4608 ( .A(n3901), .B(DATAO_REG_26__SCAN_IN), .S(n3912), .Z(U3576)
         );
  MUX2_X1 U4609 ( .A(n4036), .B(DATAO_REG_25__SCAN_IN), .S(n3912), .Z(U3575)
         );
  MUX2_X1 U4610 ( .A(n3902), .B(DATAO_REG_20__SCAN_IN), .S(n3912), .Z(U3570)
         );
  MUX2_X1 U4611 ( .A(n4197), .B(DATAO_REG_19__SCAN_IN), .S(n3912), .Z(U3569)
         );
  MUX2_X1 U4612 ( .A(n4210), .B(DATAO_REG_16__SCAN_IN), .S(n3912), .Z(U3566)
         );
  MUX2_X1 U4613 ( .A(n3903), .B(DATAO_REG_15__SCAN_IN), .S(n3912), .Z(U3565)
         );
  MUX2_X1 U4614 ( .A(n4253), .B(DATAO_REG_14__SCAN_IN), .S(n3912), .Z(U3564)
         );
  MUX2_X1 U4615 ( .A(n3904), .B(DATAO_REG_13__SCAN_IN), .S(n3912), .Z(U3563)
         );
  MUX2_X1 U4616 ( .A(n4271), .B(DATAO_REG_12__SCAN_IN), .S(n3912), .Z(U3562)
         );
  MUX2_X1 U4617 ( .A(n3905), .B(DATAO_REG_11__SCAN_IN), .S(n3912), .Z(U3561)
         );
  MUX2_X1 U4618 ( .A(n3906), .B(DATAO_REG_10__SCAN_IN), .S(n3912), .Z(U3560)
         );
  MUX2_X1 U4619 ( .A(n3907), .B(DATAO_REG_9__SCAN_IN), .S(n3912), .Z(U3559) );
  MUX2_X1 U4620 ( .A(n3908), .B(DATAO_REG_8__SCAN_IN), .S(n3912), .Z(U3558) );
  MUX2_X1 U4621 ( .A(n3909), .B(DATAO_REG_7__SCAN_IN), .S(n3912), .Z(U3557) );
  MUX2_X1 U4622 ( .A(n3910), .B(DATAO_REG_6__SCAN_IN), .S(n3912), .Z(U3556) );
  MUX2_X1 U4623 ( .A(n3911), .B(DATAO_REG_5__SCAN_IN), .S(n3912), .Z(U3555) );
  MUX2_X1 U4624 ( .A(n2730), .B(DATAO_REG_2__SCAN_IN), .S(n3912), .Z(U3552) );
  AOI21_X1 U4625 ( .B1(n3997), .B2(n3914), .A(n3913), .ZN(n3915) );
  OAI21_X1 U4626 ( .B1(n3916), .B2(n3997), .A(n3915), .ZN(n3917) );
  OAI211_X1 U4627 ( .C1(IR_REG_0__SCAN_IN), .C2(n3918), .A(n3917), .B(U4043), 
        .ZN(n3944) );
  NOR2_X1 U4628 ( .A1(STATE_REG_SCAN_IN), .A2(n3300), .ZN(n3919) );
  AOI21_X1 U4629 ( .B1(n4627), .B2(ADDR_REG_2__SCAN_IN), .A(n3919), .ZN(n3934)
         );
  INV_X1 U4630 ( .A(n3920), .ZN(n3925) );
  NAND3_X1 U4631 ( .A1(n3923), .A2(n3922), .A3(n3921), .ZN(n3924) );
  NAND3_X1 U4632 ( .A1(n4629), .A2(n3925), .A3(n3924), .ZN(n3931) );
  INV_X1 U4633 ( .A(n3926), .ZN(n3928) );
  XNOR2_X1 U4634 ( .A(n3928), .B(n3927), .ZN(n3929) );
  NAND2_X1 U4635 ( .A1(n4529), .A2(n3929), .ZN(n3930) );
  AND2_X1 U4636 ( .A1(n3931), .A2(n3930), .ZN(n3933) );
  NAND2_X1 U4637 ( .A1(n4540), .A2(n4439), .ZN(n3932) );
  NAND4_X1 U4638 ( .A1(n3944), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(U3242)
         );
  NOR2_X1 U4639 ( .A1(n4633), .A2(n3935), .ZN(n3936) );
  AOI211_X1 U4640 ( .C1(n4627), .C2(ADDR_REG_4__SCAN_IN), .A(n3937), .B(n3936), 
        .ZN(n3943) );
  XOR2_X1 U4641 ( .A(n3938), .B(REG1_REG_4__SCAN_IN), .Z(n3941) );
  XNOR2_X1 U4642 ( .A(n3939), .B(REG2_REG_4__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4643 ( .A1(n4529), .A2(n3941), .B1(n4629), .B2(n3940), .ZN(n3942)
         );
  NAND3_X1 U4644 ( .A1(n3944), .A2(n3943), .A3(n3942), .ZN(U3244) );
  INV_X1 U4645 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4354) );
  AOI22_X1 U4646 ( .A1(n3975), .A2(REG1_REG_17__SCAN_IN), .B1(n4354), .B2(
        n4562), .ZN(n4527) );
  NOR2_X1 U4647 ( .A1(n3946), .A2(n2282), .ZN(n3947) );
  INV_X1 U4648 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4887) );
  AOI22_X1 U4649 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4477), .B1(n4569), .B2(
        n4887), .ZN(n4467) );
  NOR2_X1 U4650 ( .A1(n3948), .A2(n3963), .ZN(n3949) );
  INV_X1 U4651 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4774) );
  XNOR2_X1 U4652 ( .A(n3948), .B(n3963), .ZN(n4624) );
  INV_X1 U4653 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4369) );
  AOI22_X1 U4654 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4567), .B1(n4486), .B2(
        n4369), .ZN(n4482) );
  INV_X1 U4655 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4491) );
  XNOR2_X1 U4656 ( .A(n4509), .B(REG1_REG_15__SCAN_IN), .ZN(n4505) );
  NAND2_X1 U4657 ( .A1(n4509), .A2(REG1_REG_15__SCAN_IN), .ZN(n3951) );
  NAND2_X1 U4658 ( .A1(n3952), .A2(n4564), .ZN(n3953) );
  INV_X1 U4659 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4773) );
  NAND2_X1 U4660 ( .A1(n4516), .A2(n4773), .ZN(n4515) );
  NAND2_X1 U4661 ( .A1(n3953), .A2(n4515), .ZN(n4526) );
  NAND2_X1 U4662 ( .A1(n4527), .A2(n4526), .ZN(n4525) );
  XOR2_X1 U4663 ( .A(REG1_REG_18__SCAN_IN), .B(n3976), .Z(n4533) );
  XNOR2_X1 U4664 ( .A(n4434), .B(REG1_REG_19__SCAN_IN), .ZN(n3954) );
  NOR2_X1 U4665 ( .A1(n3975), .A2(REG2_REG_17__SCAN_IN), .ZN(n3955) );
  AOI21_X1 U4666 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3975), .A(n3955), .ZN(n4524) );
  INV_X1 U4667 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4668 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4569), .B1(n4477), .B2(
        n3956), .ZN(n4474) );
  NAND2_X1 U4669 ( .A1(n3959), .A2(n3960), .ZN(n3961) );
  NAND2_X1 U4670 ( .A1(n4474), .A2(n4473), .ZN(n4472) );
  NAND2_X1 U4671 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4569), .ZN(n3962) );
  NAND2_X1 U4672 ( .A1(n3965), .A2(n3964), .ZN(n3966) );
  NOR2_X1 U4673 ( .A1(n3967), .A2(n3968), .ZN(n3969) );
  INV_X1 U4674 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4494) );
  NOR2_X1 U4675 ( .A1(n4494), .A2(n4493), .ZN(n4492) );
  NOR2_X1 U4676 ( .A1(n3969), .A2(n4492), .ZN(n4502) );
  INV_X1 U4677 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4244) );
  NAND2_X1 U4678 ( .A1(n4509), .A2(n4244), .ZN(n3970) );
  OAI21_X1 U4679 ( .B1(n4509), .B2(n4244), .A(n3970), .ZN(n3971) );
  NAND2_X1 U4680 ( .A1(n4509), .A2(REG2_REG_15__SCAN_IN), .ZN(n3972) );
  NAND2_X1 U4681 ( .A1(n2167), .A2(n4564), .ZN(n3974) );
  INV_X1 U4682 ( .A(n4564), .ZN(n3973) );
  INV_X1 U4683 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4794) );
  NAND2_X1 U4684 ( .A1(n3974), .A2(n4513), .ZN(n4523) );
  NAND2_X1 U4685 ( .A1(n4539), .A2(REG2_REG_18__SCAN_IN), .ZN(n3978) );
  NAND2_X1 U4686 ( .A1(n3976), .A2(n4804), .ZN(n3977) );
  NAND2_X1 U4687 ( .A1(n3978), .A2(n3977), .ZN(n4535) );
  INV_X1 U4688 ( .A(n3978), .ZN(n3979) );
  INV_X1 U4689 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3980) );
  MUX2_X1 U4690 ( .A(n3980), .B(REG2_REG_19__SCAN_IN), .S(n3985), .Z(n3981) );
  XNOR2_X1 U4691 ( .A(n3982), .B(n3981), .ZN(n3987) );
  AOI21_X1 U4692 ( .B1(n4627), .B2(ADDR_REG_19__SCAN_IN), .A(n3983), .ZN(n3984) );
  OAI21_X1 U4693 ( .B1(n4633), .B2(n3985), .A(n3984), .ZN(n3986) );
  AOI21_X1 U4694 ( .B1(n3987), .B2(n4629), .A(n3986), .ZN(n3988) );
  OAI21_X1 U4695 ( .B1(n3989), .B2(n4622), .A(n3988), .ZN(U3259) );
  INV_X1 U4696 ( .A(n3990), .ZN(n4003) );
  OAI21_X1 U4697 ( .B1(n3993), .B2(n3992), .A(n3991), .ZN(n3994) );
  XNOR2_X1 U4698 ( .A(n3994), .B(n2170), .ZN(n3996) );
  NAND2_X1 U4699 ( .A1(n3996), .A2(n3995), .ZN(n4002) );
  NAND2_X1 U4700 ( .A1(n4007), .A2(n4272), .ZN(n4000) );
  AOI21_X1 U4701 ( .B1(n3997), .B2(B_REG_SCAN_IN), .A(n4268), .ZN(n4290) );
  AOI22_X1 U4702 ( .A1(n3998), .A2(n4290), .B1(n4014), .B2(n4299), .ZN(n3999)
         );
  AND2_X1 U4703 ( .A1(n4000), .A2(n3999), .ZN(n4001) );
  NAND2_X1 U4704 ( .A1(n4002), .A2(n4001), .ZN(n4307) );
  AOI21_X1 U4705 ( .B1(n4003), .B2(n4552), .A(n4307), .ZN(n4017) );
  NAND2_X1 U4706 ( .A1(n4005), .A2(n4004), .ZN(n4009) );
  NAND2_X1 U4707 ( .A1(n4009), .A2(n4008), .ZN(n4010) );
  XNOR2_X1 U4708 ( .A(n4010), .B(n2170), .ZN(n4303) );
  NAND2_X1 U4709 ( .A1(n4303), .A2(n4019), .ZN(n4016) );
  AOI21_X1 U4710 ( .B1(n4014), .B2(n4013), .A(n4287), .ZN(n4304) );
  AOI22_X1 U4711 ( .A1(n4304), .A2(n4445), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4285), .ZN(n4015) );
  OAI211_X1 U4712 ( .C1(n4285), .C2(n4017), .A(n4016), .B(n4015), .ZN(U3354)
         );
  INV_X1 U4713 ( .A(n4018), .ZN(n4026) );
  NAND2_X1 U4714 ( .A1(n4020), .A2(n4019), .ZN(n4025) );
  INV_X1 U4715 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4021) );
  OAI22_X1 U4716 ( .A1(n4022), .A2(n4242), .B1(n4021), .B2(n4236), .ZN(n4023)
         );
  AOI21_X1 U4717 ( .B1(n4312), .B2(n4445), .A(n4023), .ZN(n4024) );
  OAI211_X1 U4718 ( .C1(n4026), .C2(n4285), .A(n4025), .B(n4024), .ZN(U3262)
         );
  XNOR2_X1 U4719 ( .A(n4027), .B(n4032), .ZN(n4320) );
  INV_X1 U4720 ( .A(n4320), .ZN(n4046) );
  INV_X1 U4721 ( .A(n4029), .ZN(n4030) );
  AOI21_X1 U4722 ( .B1(n4028), .B2(n4031), .A(n4030), .ZN(n4033) );
  XNOR2_X1 U4723 ( .A(n4033), .B(n4032), .ZN(n4038) );
  OAI22_X1 U4724 ( .A1(n4034), .A2(n4268), .B1(n4267), .B2(n4040), .ZN(n4035)
         );
  AOI21_X1 U4725 ( .B1(n4272), .B2(n4036), .A(n4035), .ZN(n4037) );
  OAI21_X1 U4726 ( .B1(n4038), .B2(n4275), .A(n4037), .ZN(n4319) );
  INV_X1 U4727 ( .A(n2314), .ZN(n4041) );
  INV_X1 U4728 ( .A(n3567), .ZN(n4039) );
  OAI21_X1 U4729 ( .B1(n4041), .B2(n4040), .A(n4039), .ZN(n4386) );
  AOI22_X1 U4730 ( .A1(n4042), .A2(n4552), .B1(n4285), .B2(
        REG2_REG_26__SCAN_IN), .ZN(n4043) );
  OAI21_X1 U4731 ( .B1(n4386), .B2(n4282), .A(n4043), .ZN(n4044) );
  AOI21_X1 U4732 ( .B1(n4319), .B2(n4236), .A(n4044), .ZN(n4045) );
  OAI21_X1 U4733 ( .B1(n4046), .B2(n4257), .A(n4045), .ZN(U3264) );
  XOR2_X1 U4734 ( .A(n4050), .B(n4047), .Z(n4324) );
  INV_X1 U4735 ( .A(n4324), .ZN(n4062) );
  NAND2_X1 U4736 ( .A1(n4028), .A2(n4048), .ZN(n4049) );
  XOR2_X1 U4737 ( .A(n4050), .B(n4049), .Z(n4054) );
  OAI22_X1 U4738 ( .A1(n4051), .A2(n4268), .B1(n4267), .B2(n4055), .ZN(n4052)
         );
  AOI21_X1 U4739 ( .B1(n4272), .B2(n4092), .A(n4052), .ZN(n4053) );
  OAI21_X1 U4740 ( .B1(n4054), .B2(n4275), .A(n4053), .ZN(n4323) );
  INV_X1 U4741 ( .A(n4076), .ZN(n4056) );
  OAI21_X1 U4742 ( .B1(n4056), .B2(n4055), .A(n2314), .ZN(n4389) );
  NOR2_X1 U4743 ( .A1(n4389), .A2(n4282), .ZN(n4060) );
  INV_X1 U4744 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4058) );
  OAI22_X1 U4745 ( .A1(n4236), .A2(n4058), .B1(n4057), .B2(n4242), .ZN(n4059)
         );
  AOI211_X1 U4746 ( .C1(n4323), .C2(n4236), .A(n4060), .B(n4059), .ZN(n4061)
         );
  OAI21_X1 U4747 ( .B1(n4062), .B2(n4257), .A(n4061), .ZN(U3265) );
  XNOR2_X1 U4748 ( .A(n4063), .B(n4068), .ZN(n4327) );
  INV_X1 U4749 ( .A(n4327), .ZN(n4081) );
  INV_X1 U4750 ( .A(n4064), .ZN(n4065) );
  NOR2_X1 U4751 ( .A1(n4066), .A2(n4065), .ZN(n4067) );
  XOR2_X1 U4752 ( .A(n4068), .B(n4067), .Z(n4072) );
  OAI22_X1 U4753 ( .A1(n4069), .A2(n4268), .B1(n4267), .B2(n4074), .ZN(n4070)
         );
  AOI21_X1 U4754 ( .B1(n4272), .B2(n4116), .A(n4070), .ZN(n4071) );
  OAI21_X1 U4755 ( .B1(n4072), .B2(n4275), .A(n4071), .ZN(n4326) );
  OR2_X1 U4756 ( .A1(n4073), .A2(n4074), .ZN(n4075) );
  NAND2_X1 U4757 ( .A1(n4076), .A2(n4075), .ZN(n4392) );
  AOI22_X1 U4758 ( .A1(n4285), .A2(REG2_REG_24__SCAN_IN), .B1(n4077), .B2(
        n4552), .ZN(n4078) );
  OAI21_X1 U4759 ( .B1(n4392), .B2(n4282), .A(n4078), .ZN(n4079) );
  AOI21_X1 U4760 ( .B1(n4326), .B2(n4236), .A(n4079), .ZN(n4080) );
  OAI21_X1 U4761 ( .B1(n4081), .B2(n4257), .A(n4080), .ZN(U3266) );
  XOR2_X1 U4762 ( .A(n4089), .B(n4082), .Z(n4330) );
  INV_X1 U4763 ( .A(n4330), .ZN(n4104) );
  OR2_X1 U4764 ( .A1(n4083), .A2(n4084), .ZN(n4087) );
  INV_X1 U4765 ( .A(n4085), .ZN(n4086) );
  NAND2_X1 U4766 ( .A1(n4087), .A2(n4086), .ZN(n4114) );
  INV_X1 U4767 ( .A(n4106), .ZN(n4115) );
  NAND2_X1 U4768 ( .A1(n4114), .A2(n4115), .ZN(n4113) );
  NAND2_X1 U4769 ( .A1(n4113), .A2(n4088), .ZN(n4090) );
  XNOR2_X1 U4770 ( .A(n4090), .B(n4089), .ZN(n4095) );
  NOR2_X1 U4771 ( .A1(n4097), .A2(n4267), .ZN(n4091) );
  AOI21_X1 U4772 ( .B1(n4092), .B2(n4230), .A(n4091), .ZN(n4094) );
  NAND2_X1 U4773 ( .A1(n4128), .A2(n4272), .ZN(n4093) );
  OAI211_X1 U4774 ( .C1(n4095), .C2(n4275), .A(n4094), .B(n4093), .ZN(n4329)
         );
  INV_X1 U4775 ( .A(n4333), .ZN(n4098) );
  INV_X1 U4776 ( .A(n4073), .ZN(n4096) );
  OAI21_X1 U4777 ( .B1(n4098), .B2(n4097), .A(n4096), .ZN(n4396) );
  NOR2_X1 U4778 ( .A1(n4396), .A2(n4282), .ZN(n4102) );
  INV_X1 U4779 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4100) );
  OAI22_X1 U4780 ( .A1(n4236), .A2(n4100), .B1(n4099), .B2(n4242), .ZN(n4101)
         );
  AOI211_X1 U4781 ( .C1(n4329), .C2(n4236), .A(n4102), .B(n4101), .ZN(n4103)
         );
  OAI21_X1 U4782 ( .B1(n4104), .B2(n4257), .A(n4103), .ZN(U3267) );
  OAI21_X1 U4783 ( .B1(n4107), .B2(n4106), .A(n4105), .ZN(n4336) );
  NAND2_X1 U4784 ( .A1(n4131), .A2(n4108), .ZN(n4332) );
  AND2_X1 U4785 ( .A1(n4332), .A2(n4445), .ZN(n4112) );
  INV_X1 U4786 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4110) );
  OAI22_X1 U4787 ( .A1(n4556), .A2(n4110), .B1(n4109), .B2(n4242), .ZN(n4111)
         );
  AOI21_X1 U4788 ( .B1(n4112), .B2(n4333), .A(n4111), .ZN(n4123) );
  OAI21_X1 U4789 ( .B1(n4115), .B2(n4114), .A(n4113), .ZN(n4121) );
  NAND2_X1 U4790 ( .A1(n4147), .A2(n4272), .ZN(n4118) );
  NAND2_X1 U4791 ( .A1(n4116), .A2(n4230), .ZN(n4117) );
  OAI211_X1 U4792 ( .C1(n4267), .C2(n4119), .A(n4118), .B(n4117), .ZN(n4120)
         );
  AOI21_X1 U4793 ( .B1(n4121), .B2(n3995), .A(n4120), .ZN(n4335) );
  OR2_X1 U4794 ( .A1(n4335), .A2(n4285), .ZN(n4122) );
  OAI211_X1 U4795 ( .C1(n4336), .C2(n4257), .A(n4123), .B(n4122), .ZN(U3268)
         );
  XNOR2_X1 U4796 ( .A(n4124), .B(n4125), .ZN(n4338) );
  INV_X1 U4797 ( .A(n4338), .ZN(n4139) );
  XNOR2_X1 U4798 ( .A(n4083), .B(n4125), .ZN(n4126) );
  NAND2_X1 U4799 ( .A1(n4126), .A2(n3995), .ZN(n4130) );
  NOR2_X1 U4800 ( .A1(n4132), .A2(n4267), .ZN(n4127) );
  AOI21_X1 U4801 ( .B1(n4128), .B2(n4230), .A(n4127), .ZN(n4129) );
  OAI211_X1 U4802 ( .C1(n4174), .C2(n4234), .A(n4130), .B(n4129), .ZN(n4337)
         );
  INV_X1 U4803 ( .A(n4157), .ZN(n4133) );
  OAI21_X1 U4804 ( .B1(n4133), .B2(n4132), .A(n4131), .ZN(n4401) );
  NOR2_X1 U4805 ( .A1(n4401), .A2(n4282), .ZN(n4137) );
  INV_X1 U4806 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4135) );
  OAI22_X1 U4807 ( .A1(n4236), .A2(n4135), .B1(n4134), .B2(n4242), .ZN(n4136)
         );
  AOI211_X1 U4808 ( .C1(n4337), .C2(n4236), .A(n4137), .B(n4136), .ZN(n4138)
         );
  OAI21_X1 U4809 ( .B1(n4139), .B2(n4257), .A(n4138), .ZN(U3269) );
  XNOR2_X1 U4810 ( .A(n4140), .B(n4141), .ZN(n4341) );
  NAND2_X1 U4811 ( .A1(n4142), .A2(n4143), .ZN(n4145) );
  XNOR2_X1 U4812 ( .A(n4145), .B(n4144), .ZN(n4151) );
  AOI22_X1 U4813 ( .A1(n4147), .A2(n4230), .B1(n4299), .B2(n4146), .ZN(n4148)
         );
  OAI21_X1 U4814 ( .B1(n4149), .B2(n4234), .A(n4148), .ZN(n4150) );
  AOI21_X1 U4815 ( .B1(n4151), .B2(n3995), .A(n4150), .ZN(n4152) );
  OAI21_X1 U4816 ( .B1(n4341), .B2(n4153), .A(n4152), .ZN(n4342) );
  NAND2_X1 U4817 ( .A1(n4342), .A2(n4236), .ZN(n4163) );
  OR2_X1 U4818 ( .A1(n4154), .A2(n4155), .ZN(n4156) );
  NAND2_X1 U4819 ( .A1(n4157), .A2(n4156), .ZN(n4404) );
  INV_X1 U4820 ( .A(n4404), .ZN(n4161) );
  INV_X1 U4821 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4159) );
  OAI22_X1 U4822 ( .A1(n4236), .A2(n4159), .B1(n4158), .B2(n4242), .ZN(n4160)
         );
  AOI21_X1 U4823 ( .B1(n4161), .B2(n4445), .A(n4160), .ZN(n4162) );
  OAI211_X1 U4824 ( .C1(n4341), .C2(n4164), .A(n4163), .B(n4162), .ZN(U3270)
         );
  XNOR2_X1 U4825 ( .A(n4165), .B(n4173), .ZN(n4346) );
  INV_X1 U4826 ( .A(n4346), .ZN(n4186) );
  OAI21_X1 U4827 ( .B1(n4166), .B2(n4168), .A(n4167), .ZN(n4195) );
  INV_X1 U4828 ( .A(n4169), .ZN(n4171) );
  OAI21_X1 U4829 ( .B1(n4195), .B2(n4171), .A(n4170), .ZN(n4172) );
  XOR2_X1 U4830 ( .A(n4173), .B(n4172), .Z(n4178) );
  OAI22_X1 U4831 ( .A1(n4174), .A2(n4268), .B1(n4267), .B2(n4180), .ZN(n4175)
         );
  AOI21_X1 U4832 ( .B1(n4272), .B2(n4176), .A(n4175), .ZN(n4177) );
  OAI21_X1 U4833 ( .B1(n4178), .B2(n4275), .A(n4177), .ZN(n4345) );
  INV_X1 U4834 ( .A(n4154), .ZN(n4179) );
  OAI21_X1 U4835 ( .B1(n4181), .B2(n4180), .A(n4179), .ZN(n4408) );
  NOR2_X1 U4836 ( .A1(n4408), .A2(n4282), .ZN(n4184) );
  OAI22_X1 U4837 ( .A1(n4556), .A2(n3980), .B1(n4182), .B2(n4242), .ZN(n4183)
         );
  AOI211_X1 U4838 ( .C1(n4345), .C2(n4236), .A(n4184), .B(n4183), .ZN(n4185)
         );
  OAI21_X1 U4839 ( .B1(n4186), .B2(n4257), .A(n4185), .ZN(U3271) );
  OAI21_X1 U4840 ( .B1(n4189), .B2(n4188), .A(n4187), .ZN(n4190) );
  INV_X1 U4841 ( .A(n4190), .ZN(n4351) );
  XNOR2_X1 U4842 ( .A(n4213), .B(n4191), .ZN(n4192) );
  NAND2_X1 U4843 ( .A1(n4192), .A2(n4610), .ZN(n4349) );
  INV_X1 U4844 ( .A(n4349), .ZN(n4205) );
  OAI22_X1 U4845 ( .A1(n4556), .A2(n4804), .B1(n4193), .B2(n4242), .ZN(n4203)
         );
  XNOR2_X1 U4846 ( .A(n4195), .B(n4194), .ZN(n4201) );
  AOI22_X1 U4847 ( .A1(n4197), .A2(n4230), .B1(n4196), .B2(n4299), .ZN(n4198)
         );
  OAI21_X1 U4848 ( .B1(n4199), .B2(n4234), .A(n4198), .ZN(n4200) );
  AOI21_X1 U4849 ( .B1(n4201), .B2(n3995), .A(n4200), .ZN(n4350) );
  NOR2_X1 U4850 ( .A1(n4350), .A2(n4285), .ZN(n4202) );
  AOI211_X1 U4851 ( .C1(n4205), .C2(n4204), .A(n4203), .B(n4202), .ZN(n4206)
         );
  OAI21_X1 U4852 ( .B1(n4351), .B2(n4257), .A(n4206), .ZN(U3272) );
  XOR2_X1 U4853 ( .A(n4208), .B(n4207), .Z(n4353) );
  INV_X1 U4854 ( .A(n4353), .ZN(n4219) );
  XOR2_X1 U4855 ( .A(n4208), .B(n4166), .Z(n4212) );
  OAI22_X1 U4856 ( .A1(n2544), .A2(n4268), .B1(n4267), .B2(n4214), .ZN(n4209)
         );
  AOI21_X1 U4857 ( .B1(n4272), .B2(n4210), .A(n4209), .ZN(n4211) );
  OAI21_X1 U4858 ( .B1(n4212), .B2(n4275), .A(n4211), .ZN(n4352) );
  OAI21_X1 U4859 ( .B1(n2143), .B2(n4214), .A(n4213), .ZN(n4413) );
  NOR2_X1 U4860 ( .A1(n4413), .A2(n4282), .ZN(n4217) );
  OAI22_X1 U4861 ( .A1(n4236), .A2(n2252), .B1(n4215), .B2(n4242), .ZN(n4216)
         );
  AOI211_X1 U4862 ( .C1(n4352), .C2(n4236), .A(n4217), .B(n4216), .ZN(n4218)
         );
  OAI21_X1 U4863 ( .B1(n4219), .B2(n4257), .A(n4218), .ZN(U3273) );
  OAI21_X1 U4864 ( .B1(n4222), .B2(n4221), .A(n4220), .ZN(n4359) );
  AOI21_X1 U4865 ( .B1(n2523), .B2(n2172), .A(n2143), .ZN(n4357) );
  OAI22_X1 U4866 ( .A1(n4556), .A2(n4794), .B1(n4223), .B2(n4242), .ZN(n4224)
         );
  AOI21_X1 U4867 ( .B1(n4357), .B2(n4445), .A(n4224), .ZN(n4238) );
  OAI211_X1 U4868 ( .C1(n4227), .C2(n4226), .A(n4225), .B(n3995), .ZN(n4233)
         );
  NOR2_X1 U4869 ( .A1(n4228), .A2(n4267), .ZN(n4229) );
  AOI21_X1 U4870 ( .B1(n4231), .B2(n4230), .A(n4229), .ZN(n4232) );
  OAI211_X1 U4871 ( .C1(n4235), .C2(n4234), .A(n4233), .B(n4232), .ZN(n4356)
         );
  NAND2_X1 U4872 ( .A1(n4356), .A2(n4236), .ZN(n4237) );
  OAI211_X1 U4873 ( .C1(n4359), .C2(n4257), .A(n4238), .B(n4237), .ZN(U3274)
         );
  XOR2_X1 U4874 ( .A(n4250), .B(n4239), .Z(n4363) );
  XNOR2_X1 U4875 ( .A(n4241), .B(n4240), .ZN(n4360) );
  OAI22_X1 U4876 ( .A1(n4236), .A2(n4244), .B1(n4243), .B2(n4242), .ZN(n4255)
         );
  OAI22_X1 U4877 ( .A1(n4246), .A2(n4268), .B1(n4267), .B2(n4245), .ZN(n4252)
         );
  INV_X1 U4878 ( .A(n4248), .ZN(n4249) );
  AOI211_X1 U4879 ( .C1(n4272), .C2(n4253), .A(n4252), .B(n4251), .ZN(n4362)
         );
  NOR2_X1 U4880 ( .A1(n4362), .A2(n4285), .ZN(n4254) );
  AOI211_X1 U4881 ( .C1(n4445), .C2(n4360), .A(n4255), .B(n4254), .ZN(n4256)
         );
  OAI21_X1 U4882 ( .B1(n4363), .B2(n4257), .A(n4256), .ZN(U3275) );
  INV_X1 U4883 ( .A(n4258), .ZN(n4259) );
  AOI21_X1 U4884 ( .B1(n4261), .B2(n4260), .A(n4259), .ZN(n4262) );
  XOR2_X1 U4885 ( .A(n4264), .B(n4262), .Z(n4276) );
  XNOR2_X1 U4886 ( .A(n4263), .B(n4264), .ZN(n4368) );
  NAND2_X1 U4887 ( .A1(n4368), .A2(n4265), .ZN(n4274) );
  OAI22_X1 U4888 ( .A1(n4269), .A2(n4268), .B1(n4267), .B2(n4266), .ZN(n4270)
         );
  AOI21_X1 U4889 ( .B1(n4272), .B2(n4271), .A(n4270), .ZN(n4273) );
  OAI211_X1 U4890 ( .C1(n4276), .C2(n4275), .A(n4274), .B(n4273), .ZN(n4367)
         );
  INV_X1 U4891 ( .A(n4367), .ZN(n4286) );
  NAND2_X1 U4892 ( .A1(n3509), .A2(n4277), .ZN(n4278) );
  NAND2_X1 U4893 ( .A1(n4279), .A2(n4278), .ZN(n4421) );
  AOI22_X1 U4894 ( .A1(n4285), .A2(REG2_REG_13__SCAN_IN), .B1(n4280), .B2(
        n4552), .ZN(n4281) );
  OAI21_X1 U4895 ( .B1(n4421), .B2(n4282), .A(n4281), .ZN(n4283) );
  AOI21_X1 U4896 ( .B1(n4368), .B2(n4553), .A(n4283), .ZN(n4284) );
  OAI21_X1 U4897 ( .B1(n4286), .B2(n4285), .A(n4284), .ZN(U3277) );
  NAND2_X1 U4898 ( .A1(n4287), .A2(n4288), .ZN(n4295) );
  XNOR2_X1 U4899 ( .A(n4295), .B(n4289), .ZN(n4442) );
  INV_X1 U4900 ( .A(n4442), .ZN(n4378) );
  INV_X1 U4901 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4293) );
  INV_X1 U4902 ( .A(n4289), .ZN(n4292) );
  AND2_X1 U4903 ( .A1(n4291), .A2(n4290), .ZN(n4298) );
  AOI21_X1 U4904 ( .B1(n4292), .B2(n4299), .A(n4298), .ZN(n4444) );
  MUX2_X1 U4905 ( .A(n4293), .B(n4444), .S(n4621), .Z(n4294) );
  OAI21_X1 U4906 ( .B1(n4378), .B2(n4376), .A(n4294), .ZN(U3549) );
  INV_X1 U4907 ( .A(n4287), .ZN(n4297) );
  INV_X1 U4908 ( .A(n4295), .ZN(n4296) );
  AOI21_X1 U4909 ( .B1(n4300), .B2(n4297), .A(n4296), .ZN(n4446) );
  INV_X1 U4910 ( .A(n4446), .ZN(n4380) );
  INV_X1 U4911 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4301) );
  AOI21_X1 U4912 ( .B1(n4300), .B2(n4299), .A(n4298), .ZN(n4448) );
  MUX2_X1 U4913 ( .A(n4301), .B(n4448), .S(n4621), .Z(n4302) );
  OAI21_X1 U4914 ( .B1(n4380), .B2(n4376), .A(n4302), .ZN(U3548) );
  NAND2_X1 U4915 ( .A1(n4303), .A2(n4602), .ZN(n4309) );
  INV_X1 U4916 ( .A(n4304), .ZN(n4305) );
  NOR2_X1 U4917 ( .A1(n4305), .A2(n4600), .ZN(n4306) );
  NAND2_X1 U4918 ( .A1(n4309), .A2(n4308), .ZN(n4381) );
  MUX2_X1 U4919 ( .A(REG1_REG_29__SCAN_IN), .B(n4381), .S(n4621), .Z(U3547) );
  INV_X1 U4920 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4789) );
  NAND2_X1 U4921 ( .A1(n4312), .A2(n4311), .ZN(n4313) );
  NAND2_X1 U4922 ( .A1(n4314), .A2(n4313), .ZN(U3546) );
  NAND2_X1 U4923 ( .A1(n4315), .A2(n4602), .ZN(n4317) );
  OAI211_X1 U4924 ( .C1(n4600), .C2(n4318), .A(n4317), .B(n4316), .ZN(n4382)
         );
  MUX2_X1 U4925 ( .A(REG1_REG_27__SCAN_IN), .B(n4382), .S(n4621), .Z(U3545) );
  INV_X1 U4926 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4321) );
  AOI21_X1 U4927 ( .B1(n4320), .B2(n4602), .A(n4319), .ZN(n4383) );
  MUX2_X1 U4928 ( .A(n4321), .B(n4383), .S(n4621), .Z(n4322) );
  OAI21_X1 U4929 ( .B1(n4376), .B2(n4386), .A(n4322), .ZN(U3544) );
  INV_X1 U4930 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4782) );
  AOI21_X1 U4931 ( .B1(n4324), .B2(n4602), .A(n4323), .ZN(n4387) );
  MUX2_X1 U4932 ( .A(n4782), .B(n4387), .S(n4621), .Z(n4325) );
  OAI21_X1 U4933 ( .B1(n4376), .B2(n4389), .A(n4325), .ZN(U3543) );
  INV_X1 U4934 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4779) );
  AOI21_X1 U4935 ( .B1(n4327), .B2(n4602), .A(n4326), .ZN(n4390) );
  MUX2_X1 U4936 ( .A(n4779), .B(n4390), .S(n4621), .Z(n4328) );
  OAI21_X1 U4937 ( .B1(n4376), .B2(n4392), .A(n4328), .ZN(U3542) );
  INV_X1 U4938 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4870) );
  AOI21_X1 U4939 ( .B1(n4330), .B2(n4602), .A(n4329), .ZN(n4393) );
  MUX2_X1 U4940 ( .A(n4870), .B(n4393), .S(n4621), .Z(n4331) );
  OAI21_X1 U4941 ( .B1(n4376), .B2(n4396), .A(n4331), .ZN(U3541) );
  NAND3_X1 U4942 ( .A1(n4333), .A2(n4610), .A3(n4332), .ZN(n4334) );
  OAI211_X1 U4943 ( .C1(n4336), .C2(n4591), .A(n4335), .B(n4334), .ZN(n4397)
         );
  MUX2_X1 U4944 ( .A(REG1_REG_22__SCAN_IN), .B(n4397), .S(n4621), .Z(U3540) );
  INV_X1 U4945 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4339) );
  AOI21_X1 U4946 ( .B1(n4338), .B2(n4602), .A(n4337), .ZN(n4398) );
  MUX2_X1 U4947 ( .A(n4339), .B(n4398), .S(n4621), .Z(n4340) );
  OAI21_X1 U4948 ( .B1(n4376), .B2(n4401), .A(n4340), .ZN(U3539) );
  INV_X1 U4949 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4776) );
  INV_X1 U4950 ( .A(n4341), .ZN(n4343) );
  AOI21_X1 U4951 ( .B1(n4583), .B2(n4343), .A(n4342), .ZN(n4402) );
  MUX2_X1 U4952 ( .A(n4776), .B(n4402), .S(n4621), .Z(n4344) );
  OAI21_X1 U4953 ( .B1(n4376), .B2(n4404), .A(n4344), .ZN(U3538) );
  INV_X1 U4954 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4347) );
  AOI21_X1 U4955 ( .B1(n4346), .B2(n4602), .A(n4345), .ZN(n4405) );
  MUX2_X1 U4956 ( .A(n4347), .B(n4405), .S(n4621), .Z(n4348) );
  OAI21_X1 U4957 ( .B1(n4376), .B2(n4408), .A(n4348), .ZN(U3537) );
  OAI211_X1 U4958 ( .C1(n4351), .C2(n4591), .A(n4350), .B(n4349), .ZN(n4409)
         );
  MUX2_X1 U4959 ( .A(REG1_REG_18__SCAN_IN), .B(n4409), .S(n4621), .Z(U3536) );
  AOI21_X1 U4960 ( .B1(n4353), .B2(n4602), .A(n4352), .ZN(n4410) );
  MUX2_X1 U4961 ( .A(n4354), .B(n4410), .S(n4621), .Z(n4355) );
  OAI21_X1 U4962 ( .B1(n4376), .B2(n4413), .A(n4355), .ZN(U3535) );
  AOI21_X1 U4963 ( .B1(n4610), .B2(n4357), .A(n4356), .ZN(n4358) );
  OAI21_X1 U4964 ( .B1(n4359), .B2(n4591), .A(n4358), .ZN(n4414) );
  MUX2_X1 U4965 ( .A(REG1_REG_16__SCAN_IN), .B(n4414), .S(n4621), .Z(U3534) );
  NAND2_X1 U4966 ( .A1(n4360), .A2(n4610), .ZN(n4361) );
  OAI211_X1 U4967 ( .C1(n4591), .C2(n4363), .A(n4362), .B(n4361), .ZN(n4415)
         );
  MUX2_X1 U4968 ( .A(REG1_REG_15__SCAN_IN), .B(n4415), .S(n4621), .Z(U3533) );
  AOI21_X1 U4969 ( .B1(n4365), .B2(n4602), .A(n4364), .ZN(n4416) );
  MUX2_X1 U4970 ( .A(n4491), .B(n4416), .S(n4621), .Z(n4366) );
  OAI21_X1 U4971 ( .B1(n4376), .B2(n4418), .A(n4366), .ZN(U3532) );
  AOI21_X1 U4972 ( .B1(n4583), .B2(n4368), .A(n4367), .ZN(n4419) );
  MUX2_X1 U4973 ( .A(n4369), .B(n4419), .S(n4621), .Z(n4370) );
  OAI21_X1 U4974 ( .B1(n4376), .B2(n4421), .A(n4370), .ZN(U3531) );
  NAND2_X1 U4975 ( .A1(n4371), .A2(n4602), .ZN(n4372) );
  NAND2_X1 U4976 ( .A1(n4373), .A2(n4372), .ZN(n4422) );
  MUX2_X1 U4977 ( .A(REG1_REG_12__SCAN_IN), .B(n4422), .S(n4621), .Z(n4374) );
  INV_X1 U4978 ( .A(n4374), .ZN(n4375) );
  OAI21_X1 U4979 ( .B1(n4376), .B2(n4426), .A(n4375), .ZN(U3530) );
  INV_X1 U4980 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4866) );
  MUX2_X1 U4981 ( .A(n4866), .B(n4444), .S(n4613), .Z(n4377) );
  OAI21_X1 U4982 ( .B1(n4378), .B2(n4425), .A(n4377), .ZN(U3517) );
  INV_X1 U4983 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4868) );
  MUX2_X1 U4984 ( .A(n4868), .B(n4448), .S(n4613), .Z(n4379) );
  OAI21_X1 U4985 ( .B1(n4380), .B2(n4425), .A(n4379), .ZN(U3516) );
  MUX2_X1 U4986 ( .A(REG0_REG_29__SCAN_IN), .B(n4381), .S(n4613), .Z(U3515) );
  MUX2_X1 U4987 ( .A(REG0_REG_27__SCAN_IN), .B(n4382), .S(n4613), .Z(U3513) );
  INV_X1 U4988 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4384) );
  MUX2_X1 U4989 ( .A(n4384), .B(n4383), .S(n4613), .Z(n4385) );
  OAI21_X1 U4990 ( .B1(n4386), .B2(n4425), .A(n4385), .ZN(U3512) );
  INV_X1 U4991 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4867) );
  MUX2_X1 U4992 ( .A(n4867), .B(n4387), .S(n4613), .Z(n4388) );
  OAI21_X1 U4993 ( .B1(n4389), .B2(n4425), .A(n4388), .ZN(U3511) );
  INV_X1 U4994 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4869) );
  MUX2_X1 U4995 ( .A(n4869), .B(n4390), .S(n4613), .Z(n4391) );
  OAI21_X1 U4996 ( .B1(n4392), .B2(n4425), .A(n4391), .ZN(U3510) );
  INV_X1 U4997 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4394) );
  MUX2_X1 U4998 ( .A(n4394), .B(n4393), .S(n4613), .Z(n4395) );
  OAI21_X1 U4999 ( .B1(n4396), .B2(n4425), .A(n4395), .ZN(U3509) );
  MUX2_X1 U5000 ( .A(REG0_REG_22__SCAN_IN), .B(n4397), .S(n4613), .Z(U3508) );
  INV_X1 U5001 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4399) );
  MUX2_X1 U5002 ( .A(n4399), .B(n4398), .S(n4613), .Z(n4400) );
  OAI21_X1 U5003 ( .B1(n4401), .B2(n4425), .A(n4400), .ZN(U3507) );
  INV_X1 U5004 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4755) );
  MUX2_X1 U5005 ( .A(n4755), .B(n4402), .S(n4613), .Z(n4403) );
  OAI21_X1 U5006 ( .B1(n4404), .B2(n4425), .A(n4403), .ZN(U3506) );
  INV_X1 U5007 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4406) );
  MUX2_X1 U5008 ( .A(n4406), .B(n4405), .S(n4613), .Z(n4407) );
  OAI21_X1 U5009 ( .B1(n4408), .B2(n4425), .A(n4407), .ZN(U3505) );
  MUX2_X1 U5010 ( .A(REG0_REG_18__SCAN_IN), .B(n4409), .S(n4613), .Z(U3503) );
  INV_X1 U5011 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4411) );
  MUX2_X1 U5012 ( .A(n4411), .B(n4410), .S(n4613), .Z(n4412) );
  OAI21_X1 U5013 ( .B1(n4413), .B2(n4425), .A(n4412), .ZN(U3501) );
  MUX2_X1 U5014 ( .A(REG0_REG_16__SCAN_IN), .B(n4414), .S(n4613), .Z(U3499) );
  MUX2_X1 U5015 ( .A(REG0_REG_15__SCAN_IN), .B(n4415), .S(n4613), .Z(U3497) );
  INV_X1 U5016 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4752) );
  MUX2_X1 U5017 ( .A(n4752), .B(n4416), .S(n4613), .Z(n4417) );
  OAI21_X1 U5018 ( .B1(n4418), .B2(n4425), .A(n4417), .ZN(U3495) );
  INV_X1 U5019 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4741) );
  MUX2_X1 U5020 ( .A(n4741), .B(n4419), .S(n4613), .Z(n4420) );
  OAI21_X1 U5021 ( .B1(n4421), .B2(n4425), .A(n4420), .ZN(U3493) );
  MUX2_X1 U5022 ( .A(REG0_REG_12__SCAN_IN), .B(n4422), .S(n4613), .Z(n4423) );
  INV_X1 U5023 ( .A(n4423), .ZN(n4424) );
  OAI21_X1 U5024 ( .B1(n4426), .B2(n4425), .A(n4424), .ZN(U3491) );
  MUX2_X1 U5025 ( .A(DATAI_30_), .B(n4427), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U5026 ( .A(DATAI_29_), .B(n4428), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U5027 ( .A(n4429), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5028 ( .A(n4430), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5029 ( .A(n4431), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5030 ( .A(n4432), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5031 ( .A(DATAI_20_), .B(n4433), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5032 ( .A(n4434), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5033 ( .A(n4509), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U5034 ( .A(n4435), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5035 ( .A(n4436), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5036 ( .A(n4437), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5037 ( .A(DATAI_3_), .B(n4438), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5038 ( .A(n4439), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5039 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  OAI22_X1 U5040 ( .A1(U3149), .A2(n4440), .B1(DATAI_28_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4441) );
  INV_X1 U5041 ( .A(n4441), .ZN(U3324) );
  AOI22_X1 U5042 ( .A1(n4442), .A2(n4445), .B1(n4285), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4443) );
  OAI21_X1 U5043 ( .B1(n4285), .B2(n4444), .A(n4443), .ZN(U3260) );
  AOI22_X1 U5044 ( .A1(n4446), .A2(n4445), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4285), .ZN(n4447) );
  OAI21_X1 U5045 ( .B1(n4285), .B2(n4448), .A(n4447), .ZN(U3261) );
  AOI211_X1 U5046 ( .C1(n4451), .C2(n4450), .A(n4449), .B(n4622), .ZN(n4453)
         );
  AOI211_X1 U5047 ( .C1(n4627), .C2(ADDR_REG_8__SCAN_IN), .A(n4453), .B(n4452), 
        .ZN(n4457) );
  OAI211_X1 U5048 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4455), .A(n4629), .B(n4454), 
        .ZN(n4456) );
  OAI211_X1 U5049 ( .C1(n4633), .C2(n4571), .A(n4457), .B(n4456), .ZN(U3248)
         );
  AOI211_X1 U5050 ( .C1(n4878), .C2(n4459), .A(n4458), .B(n4622), .ZN(n4460)
         );
  AOI211_X1 U5051 ( .C1(n4627), .C2(ADDR_REG_10__SCAN_IN), .A(n4461), .B(n4460), .ZN(n4465) );
  OAI211_X1 U5052 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4463), .A(n4629), .B(n4462), .ZN(n4464) );
  OAI211_X1 U5053 ( .C1(n4633), .C2(n2282), .A(n4465), .B(n4464), .ZN(U3250)
         );
  AOI211_X1 U5054 ( .C1(n4468), .C2(n4467), .A(n4466), .B(n4622), .ZN(n4471)
         );
  INV_X1 U5055 ( .A(n4469), .ZN(n4470) );
  AOI211_X1 U5056 ( .C1(n4627), .C2(ADDR_REG_11__SCAN_IN), .A(n4471), .B(n4470), .ZN(n4476) );
  OAI211_X1 U5057 ( .C1(n4474), .C2(n4473), .A(n4629), .B(n4472), .ZN(n4475)
         );
  OAI211_X1 U5058 ( .C1(n4633), .C2(n4477), .A(n4476), .B(n4475), .ZN(U3251)
         );
  INV_X1 U5059 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4916) );
  INV_X1 U5060 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4864) );
  AOI22_X1 U5061 ( .A1(REG2_REG_13__SCAN_IN), .A2(n4486), .B1(n4567), .B2(
        n4864), .ZN(n4480) );
  OAI21_X1 U5062 ( .B1(n4480), .B2(n4479), .A(n4629), .ZN(n4478) );
  AOI21_X1 U5063 ( .B1(n4480), .B2(n4479), .A(n4478), .ZN(n4485) );
  AOI211_X1 U5064 ( .C1(n4483), .C2(n4482), .A(n4481), .B(n4622), .ZN(n4484)
         );
  AOI211_X1 U5065 ( .C1(n4540), .C2(n4486), .A(n4485), .B(n4484), .ZN(n4488)
         );
  OAI211_X1 U5066 ( .C1(n4547), .C2(n4916), .A(n4488), .B(n4487), .ZN(U3253)
         );
  INV_X1 U5067 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4808) );
  AOI211_X1 U5068 ( .C1(n4491), .C2(n4490), .A(n4489), .B(n4622), .ZN(n4496)
         );
  AOI211_X1 U5069 ( .C1(n4494), .C2(n4493), .A(n4492), .B(n4537), .ZN(n4495)
         );
  AOI211_X1 U5070 ( .C1(n4540), .C2(n4565), .A(n4496), .B(n4495), .ZN(n4499)
         );
  INV_X1 U5071 ( .A(n4497), .ZN(n4498) );
  OAI211_X1 U5072 ( .C1(n4547), .C2(n4808), .A(n4499), .B(n4498), .ZN(U3254)
         );
  AOI22_X1 U5073 ( .A1(ADDR_REG_15__SCAN_IN), .A2(n4627), .B1(
        REG3_REG_15__SCAN_IN), .B2(U3149), .ZN(n4511) );
  INV_X1 U5074 ( .A(n4500), .ZN(n4501) );
  AOI211_X1 U5075 ( .C1(n4502), .C2(n2233), .A(n4537), .B(n4501), .ZN(n4508)
         );
  INV_X1 U5076 ( .A(n4503), .ZN(n4504) );
  AOI211_X1 U5077 ( .C1(n4506), .C2(n4505), .A(n4622), .B(n4504), .ZN(n4507)
         );
  AOI211_X1 U5078 ( .C1(n4540), .C2(n4509), .A(n4508), .B(n4507), .ZN(n4510)
         );
  NAND2_X1 U5079 ( .A1(n4511), .A2(n4510), .ZN(U3255) );
  AOI21_X1 U5080 ( .B1(n4627), .B2(ADDR_REG_16__SCAN_IN), .A(n4512), .ZN(n4520) );
  OAI21_X1 U5081 ( .B1(n4514), .B2(n4794), .A(n4513), .ZN(n4518) );
  OAI21_X1 U5082 ( .B1(n4516), .B2(n4773), .A(n4515), .ZN(n4517) );
  AOI22_X1 U5083 ( .A1(n4629), .A2(n4518), .B1(n4529), .B2(n4517), .ZN(n4519)
         );
  OAI211_X1 U5084 ( .C1(n4564), .C2(n4633), .A(n4520), .B(n4519), .ZN(U3256)
         );
  AOI21_X1 U5085 ( .B1(n4627), .B2(ADDR_REG_17__SCAN_IN), .A(n4521), .ZN(n4532) );
  OAI21_X1 U5086 ( .B1(n4524), .B2(n4523), .A(n4522), .ZN(n4530) );
  OAI21_X1 U5087 ( .B1(n4527), .B2(n4526), .A(n4525), .ZN(n4528) );
  AOI22_X1 U5088 ( .A1(n4629), .A2(n4530), .B1(n4529), .B2(n4528), .ZN(n4531)
         );
  OAI211_X1 U5089 ( .C1(n4562), .C2(n4633), .A(n4532), .B(n4531), .ZN(U3257)
         );
  INV_X1 U5090 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n4863) );
  NAND2_X1 U5091 ( .A1(n4536), .A2(n4535), .ZN(n4538) );
  NAND2_X1 U5092 ( .A1(n4538), .A2(n4629), .ZN(n4542) );
  OAI21_X1 U5093 ( .B1(n4542), .B2(n2163), .A(n4541), .ZN(n4543) );
  INV_X1 U5094 ( .A(n4544), .ZN(n4545) );
  OAI211_X1 U5095 ( .C1(n4547), .C2(n4863), .A(n4546), .B(n4545), .ZN(U3258)
         );
  INV_X1 U5096 ( .A(n4548), .ZN(n4550) );
  AOI21_X1 U5097 ( .B1(n4551), .B2(n4550), .A(n4549), .ZN(n4557) );
  AOI22_X1 U5098 ( .A1(n4554), .A2(n4553), .B1(REG3_REG_0__SCAN_IN), .B2(n4552), .ZN(n4555) );
  OAI221_X1 U5099 ( .B1(n4285), .B2(n4557), .C1(n4556), .C2(n3055), .A(n4555), 
        .ZN(U3290) );
  INV_X1 U5100 ( .A(D_REG_31__SCAN_IN), .ZN(n4728) );
  NOR2_X1 U5101 ( .A1(n4559), .A2(n4728), .ZN(U3291) );
  INV_X1 U5102 ( .A(D_REG_30__SCAN_IN), .ZN(n4727) );
  NOR2_X1 U5103 ( .A1(n4559), .A2(n4727), .ZN(U3292) );
  AND2_X1 U5104 ( .A1(D_REG_29__SCAN_IN), .A2(n4558), .ZN(U3293) );
  INV_X1 U5105 ( .A(D_REG_28__SCAN_IN), .ZN(n4725) );
  NOR2_X1 U5106 ( .A1(n4559), .A2(n4725), .ZN(U3294) );
  AND2_X1 U5107 ( .A1(D_REG_27__SCAN_IN), .A2(n4558), .ZN(U3295) );
  INV_X1 U5108 ( .A(D_REG_26__SCAN_IN), .ZN(n4724) );
  NOR2_X1 U5109 ( .A1(n4559), .A2(n4724), .ZN(U3296) );
  AND2_X1 U5110 ( .A1(D_REG_25__SCAN_IN), .A2(n4558), .ZN(U3297) );
  INV_X1 U5111 ( .A(D_REG_24__SCAN_IN), .ZN(n4721) );
  NOR2_X1 U5112 ( .A1(n4559), .A2(n4721), .ZN(U3298) );
  AND2_X1 U5113 ( .A1(D_REG_23__SCAN_IN), .A2(n4558), .ZN(U3299) );
  INV_X1 U5114 ( .A(D_REG_22__SCAN_IN), .ZN(n4722) );
  NOR2_X1 U5115 ( .A1(n4559), .A2(n4722), .ZN(U3300) );
  INV_X1 U5116 ( .A(D_REG_21__SCAN_IN), .ZN(n4719) );
  NOR2_X1 U5117 ( .A1(n4559), .A2(n4719), .ZN(U3301) );
  INV_X1 U5118 ( .A(D_REG_20__SCAN_IN), .ZN(n4718) );
  NOR2_X1 U5119 ( .A1(n4559), .A2(n4718), .ZN(U3302) );
  INV_X1 U5120 ( .A(D_REG_19__SCAN_IN), .ZN(n4712) );
  NOR2_X1 U5121 ( .A1(n4559), .A2(n4712), .ZN(U3303) );
  INV_X1 U5122 ( .A(D_REG_18__SCAN_IN), .ZN(n4711) );
  NOR2_X1 U5123 ( .A1(n4559), .A2(n4711), .ZN(U3304) );
  INV_X1 U5124 ( .A(D_REG_17__SCAN_IN), .ZN(n4708) );
  NOR2_X1 U5125 ( .A1(n4559), .A2(n4708), .ZN(U3305) );
  AND2_X1 U5126 ( .A1(D_REG_16__SCAN_IN), .A2(n4558), .ZN(U3306) );
  AND2_X1 U5127 ( .A1(D_REG_15__SCAN_IN), .A2(n4558), .ZN(U3307) );
  INV_X1 U5128 ( .A(D_REG_14__SCAN_IN), .ZN(n4709) );
  NOR2_X1 U5129 ( .A1(n4559), .A2(n4709), .ZN(U3308) );
  AND2_X1 U5130 ( .A1(D_REG_13__SCAN_IN), .A2(n4558), .ZN(U3309) );
  AND2_X1 U5131 ( .A1(D_REG_12__SCAN_IN), .A2(n4558), .ZN(U3310) );
  INV_X1 U5132 ( .A(D_REG_11__SCAN_IN), .ZN(n4706) );
  NOR2_X1 U5133 ( .A1(n4559), .A2(n4706), .ZN(U3311) );
  INV_X1 U5134 ( .A(D_REG_10__SCAN_IN), .ZN(n4705) );
  NOR2_X1 U5135 ( .A1(n4559), .A2(n4705), .ZN(U3312) );
  AND2_X1 U5136 ( .A1(D_REG_9__SCAN_IN), .A2(n4558), .ZN(U3313) );
  INV_X1 U5137 ( .A(D_REG_8__SCAN_IN), .ZN(n4703) );
  NOR2_X1 U5138 ( .A1(n4559), .A2(n4703), .ZN(U3314) );
  INV_X1 U5139 ( .A(D_REG_7__SCAN_IN), .ZN(n4702) );
  NOR2_X1 U5140 ( .A1(n4559), .A2(n4702), .ZN(U3315) );
  NOR2_X1 U5141 ( .A1(n4559), .A2(n4688), .ZN(U3316) );
  AND2_X1 U5142 ( .A1(D_REG_5__SCAN_IN), .A2(n4558), .ZN(U3317) );
  NOR2_X1 U5143 ( .A1(n4559), .A2(n4689), .ZN(U3318) );
  INV_X1 U5144 ( .A(D_REG_3__SCAN_IN), .ZN(n4691) );
  NOR2_X1 U5145 ( .A1(n4559), .A2(n4691), .ZN(U3319) );
  INV_X1 U5146 ( .A(D_REG_2__SCAN_IN), .ZN(n4692) );
  NOR2_X1 U5147 ( .A1(n4559), .A2(n4692), .ZN(U3320) );
  INV_X1 U5148 ( .A(DATAI_23_), .ZN(n4638) );
  AOI21_X1 U5149 ( .B1(U3149), .B2(n4638), .A(n4560), .ZN(U3329) );
  AOI22_X1 U5150 ( .A1(STATE_REG_SCAN_IN), .A2(n4562), .B1(n4561), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5151 ( .A1(STATE_REG_SCAN_IN), .A2(n4564), .B1(n4563), .B2(U3149), 
        .ZN(U3336) );
  OAI22_X1 U5152 ( .A1(U3149), .A2(n4565), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4566) );
  INV_X1 U5153 ( .A(n4566), .ZN(U3338) );
  AOI22_X1 U5154 ( .A1(STATE_REG_SCAN_IN), .A2(n4567), .B1(n4640), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5155 ( .A(DATAI_12_), .ZN(n4568) );
  AOI22_X1 U5156 ( .A1(STATE_REG_SCAN_IN), .A2(n3963), .B1(n4568), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5157 ( .A1(U3149), .A2(n4569), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4570) );
  INV_X1 U5158 ( .A(n4570), .ZN(U3341) );
  INV_X1 U5159 ( .A(DATAI_10_), .ZN(n4644) );
  AOI22_X1 U5160 ( .A1(STATE_REG_SCAN_IN), .A2(n2282), .B1(n4644), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5161 ( .A(DATAI_8_), .ZN(n4650) );
  AOI22_X1 U5162 ( .A1(STATE_REG_SCAN_IN), .A2(n4571), .B1(n4650), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5163 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4862) );
  AOI22_X1 U5164 ( .A1(n4613), .A2(n4572), .B1(n4862), .B2(n4611), .ZN(U3467)
         );
  INV_X1 U5165 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4734) );
  AOI22_X1 U5166 ( .A1(n4613), .A2(n4573), .B1(n4734), .B2(n4611), .ZN(U3469)
         );
  AOI22_X1 U5167 ( .A1(n4575), .A2(n4583), .B1(n4610), .B2(n4574), .ZN(n4576)
         );
  INV_X1 U5168 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4578) );
  AOI22_X1 U5169 ( .A1(n4613), .A2(n4614), .B1(n4578), .B2(n4611), .ZN(U3473)
         );
  INV_X1 U5170 ( .A(n4579), .ZN(n4584) );
  INV_X1 U5171 ( .A(n4580), .ZN(n4582) );
  AOI211_X1 U5172 ( .C1(n4584), .C2(n4583), .A(n4582), .B(n4581), .ZN(n4615)
         );
  INV_X1 U5173 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4585) );
  AOI22_X1 U5174 ( .A1(n4613), .A2(n4615), .B1(n4585), .B2(n4611), .ZN(U3475)
         );
  NOR2_X1 U5175 ( .A1(n4586), .A2(n4591), .ZN(n4589) );
  INV_X1 U5176 ( .A(n4587), .ZN(n4588) );
  AOI211_X1 U5177 ( .C1(n4610), .C2(n4590), .A(n4589), .B(n4588), .ZN(n4616)
         );
  INV_X1 U5178 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4736) );
  AOI22_X1 U5179 ( .A1(n4613), .A2(n4616), .B1(n4736), .B2(n4611), .ZN(U3477)
         );
  NOR2_X1 U5180 ( .A1(n4592), .A2(n4591), .ZN(n4596) );
  AOI211_X1 U5181 ( .C1(n4596), .C2(n4595), .A(n4594), .B(n4593), .ZN(n4617)
         );
  INV_X1 U5182 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4597) );
  AOI22_X1 U5183 ( .A1(n4613), .A2(n4617), .B1(n4597), .B2(n4611), .ZN(U3481)
         );
  OAI21_X1 U5184 ( .B1(n4600), .B2(n4599), .A(n4598), .ZN(n4601) );
  AOI21_X1 U5185 ( .B1(n4603), .B2(n4602), .A(n4601), .ZN(n4618) );
  INV_X1 U5186 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4604) );
  AOI22_X1 U5187 ( .A1(n4613), .A2(n4618), .B1(n4604), .B2(n4611), .ZN(U3485)
         );
  NOR2_X1 U5188 ( .A1(n4606), .A2(n4605), .ZN(n4608) );
  AOI211_X1 U5189 ( .C1(n4610), .C2(n4609), .A(n4608), .B(n4607), .ZN(n4620)
         );
  INV_X1 U5190 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4612) );
  AOI22_X1 U5191 ( .A1(n4613), .A2(n4620), .B1(n4612), .B2(n4611), .ZN(U3489)
         );
  AOI22_X1 U5192 ( .A1(n4621), .A2(n4614), .B1(n2200), .B2(n4619), .ZN(U3521)
         );
  AOI22_X1 U5193 ( .A1(n4621), .A2(n4615), .B1(n2213), .B2(n4619), .ZN(U3522)
         );
  AOI22_X1 U5194 ( .A1(n4621), .A2(n4616), .B1(n3104), .B2(n4619), .ZN(U3523)
         );
  AOI22_X1 U5195 ( .A1(n4621), .A2(n4617), .B1(n3158), .B2(n4619), .ZN(U3525)
         );
  AOI22_X1 U5196 ( .A1(n4621), .A2(n4618), .B1(n3163), .B2(n4619), .ZN(U3527)
         );
  AOI22_X1 U5197 ( .A1(n4621), .A2(n4620), .B1(n4887), .B2(n4619), .ZN(U3529)
         );
  AOI211_X1 U5198 ( .C1(n4774), .C2(n4624), .A(n4623), .B(n4622), .ZN(n4626)
         );
  AOI211_X1 U5199 ( .C1(n4627), .C2(ADDR_REG_12__SCAN_IN), .A(n4626), .B(n4625), .ZN(n4632) );
  OAI211_X1 U5200 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4630), .A(n4629), .B(n4628), .ZN(n4631) );
  OAI211_X1 U5201 ( .C1(n4633), .C2(n3963), .A(n4632), .B(n4631), .ZN(n4860)
         );
  INV_X1 U5202 ( .A(DATAI_30_), .ZN(n4910) );
  AOI22_X1 U5203 ( .A1(n4635), .A2(keyinput108), .B1(keyinput106), .B2(n4910), 
        .ZN(n4634) );
  OAI221_X1 U5204 ( .B1(n4635), .B2(keyinput108), .C1(n4910), .C2(keyinput106), 
        .A(n4634), .ZN(n4648) );
  INV_X1 U5205 ( .A(DATAI_22_), .ZN(n4637) );
  AOI22_X1 U5206 ( .A1(n4638), .A2(keyinput97), .B1(keyinput112), .B2(n4637), 
        .ZN(n4636) );
  OAI221_X1 U5207 ( .B1(n4638), .B2(keyinput97), .C1(n4637), .C2(keyinput112), 
        .A(n4636), .ZN(n4647) );
  INV_X1 U5208 ( .A(DATAI_19_), .ZN(n4641) );
  AOI22_X1 U5209 ( .A1(n4641), .A2(keyinput37), .B1(keyinput64), .B2(n4640), 
        .ZN(n4639) );
  OAI221_X1 U5210 ( .B1(n4641), .B2(keyinput37), .C1(n4640), .C2(keyinput64), 
        .A(n4639), .ZN(n4646) );
  INV_X1 U5211 ( .A(DATAI_9_), .ZN(n4643) );
  AOI22_X1 U5212 ( .A1(n4644), .A2(keyinput99), .B1(keyinput0), .B2(n4643), 
        .ZN(n4642) );
  OAI221_X1 U5213 ( .B1(n4644), .B2(keyinput99), .C1(n4643), .C2(keyinput0), 
        .A(n4642), .ZN(n4645) );
  NOR4_X1 U5214 ( .A1(n4648), .A2(n4647), .A3(n4646), .A4(n4645), .ZN(n4686)
         );
  INV_X1 U5215 ( .A(DATAI_6_), .ZN(n4651) );
  AOI22_X1 U5216 ( .A1(n4651), .A2(keyinput125), .B1(n4650), .B2(keyinput52), 
        .ZN(n4649) );
  OAI221_X1 U5217 ( .B1(n4651), .B2(keyinput125), .C1(n4650), .C2(keyinput52), 
        .A(n4649), .ZN(n4660) );
  AOI22_X1 U5218 ( .A1(n4904), .A2(keyinput89), .B1(keyinput79), .B2(n4653), 
        .ZN(n4652) );
  OAI221_X1 U5219 ( .B1(n4904), .B2(keyinput89), .C1(n4653), .C2(keyinput79), 
        .A(n4652), .ZN(n4659) );
  INV_X1 U5220 ( .A(DATAI_0_), .ZN(n4903) );
  XOR2_X1 U5221 ( .A(n4903), .B(keyinput24), .Z(n4657) );
  XNOR2_X1 U5222 ( .A(keyinput123), .B(DATAI_5_), .ZN(n4656) );
  XNOR2_X1 U5223 ( .A(DATAI_4_), .B(keyinput96), .ZN(n4655) );
  XNOR2_X1 U5224 ( .A(DATAI_3_), .B(keyinput71), .ZN(n4654) );
  NAND4_X1 U5225 ( .A1(n4657), .A2(n4656), .A3(n4655), .A4(n4654), .ZN(n4658)
         );
  NOR3_X1 U5226 ( .A1(n4660), .A2(n4659), .A3(n4658), .ZN(n4685) );
  AOI22_X1 U5227 ( .A1(n2470), .A2(keyinput2), .B1(n2514), .B2(keyinput110), 
        .ZN(n4661) );
  OAI221_X1 U5228 ( .B1(n2470), .B2(keyinput2), .C1(n2514), .C2(keyinput110), 
        .A(n4661), .ZN(n4670) );
  AOI22_X1 U5229 ( .A1(n2419), .A2(keyinput115), .B1(n4898), .B2(keyinput7), 
        .ZN(n4662) );
  OAI221_X1 U5230 ( .B1(n2419), .B2(keyinput115), .C1(n4898), .C2(keyinput7), 
        .A(n4662), .ZN(n4669) );
  AOI22_X1 U5231 ( .A1(n4897), .A2(keyinput92), .B1(n4664), .B2(keyinput111), 
        .ZN(n4663) );
  OAI221_X1 U5232 ( .B1(n4897), .B2(keyinput92), .C1(n4664), .C2(keyinput111), 
        .A(n4663), .ZN(n4668) );
  XOR2_X1 U5233 ( .A(n2319), .B(keyinput14), .Z(n4666) );
  XNOR2_X1 U5234 ( .A(IR_REG_1__SCAN_IN), .B(keyinput33), .ZN(n4665) );
  NAND2_X1 U5235 ( .A1(n4666), .A2(n4665), .ZN(n4667) );
  NOR4_X1 U5236 ( .A1(n4670), .A2(n4669), .A3(n4668), .A4(n4667), .ZN(n4684)
         );
  INV_X1 U5237 ( .A(IR_REG_8__SCAN_IN), .ZN(n4671) );
  XOR2_X1 U5238 ( .A(n4671), .B(keyinput126), .Z(n4676) );
  INV_X1 U5239 ( .A(IR_REG_22__SCAN_IN), .ZN(n4672) );
  XOR2_X1 U5240 ( .A(n4672), .B(keyinput16), .Z(n4675) );
  XNOR2_X1 U5241 ( .A(IR_REG_21__SCAN_IN), .B(keyinput55), .ZN(n4674) );
  XNOR2_X1 U5242 ( .A(IR_REG_16__SCAN_IN), .B(keyinput36), .ZN(n4673) );
  NAND4_X1 U5243 ( .A1(n4676), .A2(n4675), .A3(n4674), .A4(n4673), .ZN(n4682)
         );
  XNOR2_X1 U5244 ( .A(IR_REG_11__SCAN_IN), .B(keyinput109), .ZN(n4680) );
  XNOR2_X1 U5245 ( .A(IR_REG_6__SCAN_IN), .B(keyinput113), .ZN(n4679) );
  XNOR2_X1 U5246 ( .A(IR_REG_13__SCAN_IN), .B(keyinput60), .ZN(n4678) );
  XNOR2_X1 U5247 ( .A(IR_REG_12__SCAN_IN), .B(keyinput122), .ZN(n4677) );
  NAND4_X1 U5248 ( .A1(n4680), .A2(n4679), .A3(n4678), .A4(n4677), .ZN(n4681)
         );
  NOR2_X1 U5249 ( .A1(n4682), .A2(n4681), .ZN(n4683) );
  NAND4_X1 U5250 ( .A1(n4686), .A2(n4685), .A3(n4684), .A4(n4683), .ZN(n4858)
         );
  AOI22_X1 U5251 ( .A1(n4689), .A2(keyinput69), .B1(keyinput59), .B2(n4688), 
        .ZN(n4687) );
  OAI221_X1 U5252 ( .B1(n4689), .B2(keyinput69), .C1(n4688), .C2(keyinput59), 
        .A(n4687), .ZN(n4700) );
  AOI22_X1 U5253 ( .A1(n4692), .A2(keyinput119), .B1(keyinput40), .B2(n4691), 
        .ZN(n4690) );
  OAI221_X1 U5254 ( .B1(n4692), .B2(keyinput119), .C1(n4691), .C2(keyinput40), 
        .A(n4690), .ZN(n4699) );
  XOR2_X1 U5255 ( .A(n4693), .B(keyinput42), .Z(n4697) );
  XNOR2_X1 U5256 ( .A(IR_REG_23__SCAN_IN), .B(keyinput86), .ZN(n4696) );
  XNOR2_X1 U5257 ( .A(IR_REG_24__SCAN_IN), .B(keyinput12), .ZN(n4695) );
  XNOR2_X1 U5258 ( .A(IR_REG_25__SCAN_IN), .B(keyinput103), .ZN(n4694) );
  NAND4_X1 U5259 ( .A1(n4697), .A2(n4696), .A3(n4695), .A4(n4694), .ZN(n4698)
         );
  NOR3_X1 U5260 ( .A1(n4700), .A2(n4699), .A3(n4698), .ZN(n4750) );
  AOI22_X1 U5261 ( .A1(n4703), .A2(keyinput72), .B1(keyinput116), .B2(n4702), 
        .ZN(n4701) );
  OAI221_X1 U5262 ( .B1(n4703), .B2(keyinput72), .C1(n4702), .C2(keyinput116), 
        .A(n4701), .ZN(n4716) );
  AOI22_X1 U5263 ( .A1(n4706), .A2(keyinput118), .B1(keyinput44), .B2(n4705), 
        .ZN(n4704) );
  OAI221_X1 U5264 ( .B1(n4706), .B2(keyinput118), .C1(n4705), .C2(keyinput44), 
        .A(n4704), .ZN(n4715) );
  AOI22_X1 U5265 ( .A1(n4709), .A2(keyinput39), .B1(keyinput95), .B2(n4708), 
        .ZN(n4707) );
  OAI221_X1 U5266 ( .B1(n4709), .B2(keyinput39), .C1(n4708), .C2(keyinput95), 
        .A(n4707), .ZN(n4714) );
  AOI22_X1 U5267 ( .A1(n4712), .A2(keyinput15), .B1(keyinput107), .B2(n4711), 
        .ZN(n4710) );
  OAI221_X1 U5268 ( .B1(n4712), .B2(keyinput15), .C1(n4711), .C2(keyinput107), 
        .A(n4710), .ZN(n4713) );
  NOR4_X1 U5269 ( .A1(n4716), .A2(n4715), .A3(n4714), .A4(n4713), .ZN(n4749)
         );
  AOI22_X1 U5270 ( .A1(n4719), .A2(keyinput3), .B1(n4718), .B2(keyinput18), 
        .ZN(n4717) );
  OAI221_X1 U5271 ( .B1(n4719), .B2(keyinput3), .C1(n4718), .C2(keyinput18), 
        .A(n4717), .ZN(n4732) );
  AOI22_X1 U5272 ( .A1(n4722), .A2(keyinput76), .B1(keyinput31), .B2(n4721), 
        .ZN(n4720) );
  OAI221_X1 U5273 ( .B1(n4722), .B2(keyinput76), .C1(n4721), .C2(keyinput31), 
        .A(n4720), .ZN(n4731) );
  AOI22_X1 U5274 ( .A1(n4725), .A2(keyinput41), .B1(n4724), .B2(keyinput35), 
        .ZN(n4723) );
  OAI221_X1 U5275 ( .B1(n4725), .B2(keyinput41), .C1(n4724), .C2(keyinput35), 
        .A(n4723), .ZN(n4730) );
  AOI22_X1 U5276 ( .A1(n4728), .A2(keyinput47), .B1(n4727), .B2(keyinput77), 
        .ZN(n4726) );
  OAI221_X1 U5277 ( .B1(n4728), .B2(keyinput47), .C1(n4727), .C2(keyinput77), 
        .A(n4726), .ZN(n4729) );
  NOR4_X1 U5278 ( .A1(n4732), .A2(n4731), .A3(n4730), .A4(n4729), .ZN(n4748)
         );
  AOI22_X1 U5279 ( .A1(n4862), .A2(keyinput46), .B1(n4734), .B2(keyinput45), 
        .ZN(n4733) );
  OAI221_X1 U5280 ( .B1(n4862), .B2(keyinput46), .C1(n4734), .C2(keyinput45), 
        .A(n4733), .ZN(n4746) );
  AOI22_X1 U5281 ( .A1(n4737), .A2(keyinput22), .B1(n4736), .B2(keyinput67), 
        .ZN(n4735) );
  OAI221_X1 U5282 ( .B1(n4737), .B2(keyinput22), .C1(n4736), .C2(keyinput67), 
        .A(n4735), .ZN(n4745) );
  AOI22_X1 U5283 ( .A1(n4861), .A2(keyinput4), .B1(n4739), .B2(keyinput21), 
        .ZN(n4738) );
  OAI221_X1 U5284 ( .B1(n4861), .B2(keyinput4), .C1(n4739), .C2(keyinput21), 
        .A(n4738), .ZN(n4744) );
  INV_X1 U5285 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4742) );
  AOI22_X1 U5286 ( .A1(n4742), .A2(keyinput120), .B1(n4741), .B2(keyinput78), 
        .ZN(n4740) );
  OAI221_X1 U5287 ( .B1(n4742), .B2(keyinput120), .C1(n4741), .C2(keyinput78), 
        .A(n4740), .ZN(n4743) );
  NOR4_X1 U5288 ( .A1(n4746), .A2(n4745), .A3(n4744), .A4(n4743), .ZN(n4747)
         );
  NAND4_X1 U5289 ( .A1(n4750), .A2(n4749), .A3(n4748), .A4(n4747), .ZN(n4857)
         );
  INV_X1 U5290 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4753) );
  AOI22_X1 U5291 ( .A1(n4753), .A2(keyinput49), .B1(keyinput1), .B2(n4752), 
        .ZN(n4751) );
  OAI221_X1 U5292 ( .B1(n4753), .B2(keyinput49), .C1(n4752), .C2(keyinput1), 
        .A(n4751), .ZN(n4762) );
  AOI22_X1 U5293 ( .A1(n4755), .A2(keyinput124), .B1(keyinput100), .B2(n4869), 
        .ZN(n4754) );
  OAI221_X1 U5294 ( .B1(n4755), .B2(keyinput124), .C1(n4869), .C2(keyinput100), 
        .A(n4754), .ZN(n4761) );
  INV_X1 U5295 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4757) );
  AOI22_X1 U5296 ( .A1(n4867), .A2(keyinput8), .B1(n4757), .B2(keyinput83), 
        .ZN(n4756) );
  OAI221_X1 U5297 ( .B1(n4867), .B2(keyinput8), .C1(n4757), .C2(keyinput83), 
        .A(n4756), .ZN(n4760) );
  AOI22_X1 U5298 ( .A1(n4868), .A2(keyinput114), .B1(keyinput73), .B2(n4866), 
        .ZN(n4758) );
  OAI221_X1 U5299 ( .B1(n4868), .B2(keyinput114), .C1(n4866), .C2(keyinput73), 
        .A(n4758), .ZN(n4759) );
  NOR4_X1 U5300 ( .A1(n4762), .A2(n4761), .A3(n4760), .A4(n4759), .ZN(n4802)
         );
  AOI22_X1 U5301 ( .A1(n4878), .A2(keyinput56), .B1(n4887), .B2(keyinput75), 
        .ZN(n4763) );
  OAI221_X1 U5302 ( .B1(n4878), .B2(keyinput56), .C1(n4887), .C2(keyinput75), 
        .A(n4763), .ZN(n4771) );
  AOI22_X1 U5303 ( .A1(n3104), .A2(keyinput121), .B1(n3158), .B2(keyinput87), 
        .ZN(n4764) );
  OAI221_X1 U5304 ( .B1(n3104), .B2(keyinput121), .C1(n3158), .C2(keyinput87), 
        .A(n4764), .ZN(n4770) );
  XOR2_X1 U5305 ( .A(n2213), .B(keyinput82), .Z(n4768) );
  XNOR2_X1 U5306 ( .A(REG1_REG_0__SCAN_IN), .B(keyinput98), .ZN(n4767) );
  XNOR2_X1 U5307 ( .A(REG1_REG_1__SCAN_IN), .B(keyinput43), .ZN(n4766) );
  XNOR2_X1 U5308 ( .A(REG1_REG_2__SCAN_IN), .B(keyinput102), .ZN(n4765) );
  NAND4_X1 U5309 ( .A1(n4768), .A2(n4767), .A3(n4766), .A4(n4765), .ZN(n4769)
         );
  NOR3_X1 U5310 ( .A1(n4771), .A2(n4770), .A3(n4769), .ZN(n4801) );
  AOI22_X1 U5311 ( .A1(n4774), .A2(keyinput48), .B1(n4773), .B2(keyinput32), 
        .ZN(n4772) );
  OAI221_X1 U5312 ( .B1(n4774), .B2(keyinput48), .C1(n4773), .C2(keyinput32), 
        .A(n4772), .ZN(n4786) );
  INV_X1 U5313 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4777) );
  AOI22_X1 U5314 ( .A1(n4777), .A2(keyinput17), .B1(n4776), .B2(keyinput28), 
        .ZN(n4775) );
  OAI221_X1 U5315 ( .B1(n4777), .B2(keyinput17), .C1(n4776), .C2(keyinput28), 
        .A(n4775), .ZN(n4785) );
  AOI22_X1 U5316 ( .A1(n4870), .A2(keyinput23), .B1(keyinput38), .B2(n4779), 
        .ZN(n4778) );
  OAI221_X1 U5317 ( .B1(n4870), .B2(keyinput23), .C1(n4779), .C2(keyinput38), 
        .A(n4778), .ZN(n4784) );
  INV_X1 U5318 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4781) );
  AOI22_X1 U5319 ( .A1(n4782), .A2(keyinput127), .B1(n4781), .B2(keyinput93), 
        .ZN(n4780) );
  OAI221_X1 U5320 ( .B1(n4782), .B2(keyinput127), .C1(n4781), .C2(keyinput93), 
        .A(n4780), .ZN(n4783) );
  NOR4_X1 U5321 ( .A1(n4786), .A2(n4785), .A3(n4784), .A4(n4783), .ZN(n4800)
         );
  INV_X1 U5322 ( .A(REG1_REG_29__SCAN_IN), .ZN(n4788) );
  AOI22_X1 U5323 ( .A1(n4789), .A2(keyinput105), .B1(n4788), .B2(keyinput101), 
        .ZN(n4787) );
  OAI221_X1 U5324 ( .B1(n4789), .B2(keyinput105), .C1(n4788), .C2(keyinput101), 
        .A(n4787), .ZN(n4798) );
  INV_X1 U5325 ( .A(REG2_REG_3__SCAN_IN), .ZN(n4791) );
  AOI22_X1 U5326 ( .A1(n2247), .A2(keyinput94), .B1(n4791), .B2(keyinput66), 
        .ZN(n4790) );
  OAI221_X1 U5327 ( .B1(n2247), .B2(keyinput94), .C1(n4791), .C2(keyinput66), 
        .A(n4790), .ZN(n4797) );
  AOI22_X1 U5328 ( .A1(n3289), .A2(keyinput90), .B1(n3406), .B2(keyinput27), 
        .ZN(n4792) );
  OAI221_X1 U5329 ( .B1(n3289), .B2(keyinput90), .C1(n3406), .C2(keyinput27), 
        .A(n4792), .ZN(n4796) );
  AOI22_X1 U5330 ( .A1(n4794), .A2(keyinput63), .B1(keyinput6), .B2(n4864), 
        .ZN(n4793) );
  OAI221_X1 U5331 ( .B1(n4794), .B2(keyinput63), .C1(n4864), .C2(keyinput6), 
        .A(n4793), .ZN(n4795) );
  NOR4_X1 U5332 ( .A1(n4798), .A2(n4797), .A3(n4796), .A4(n4795), .ZN(n4799)
         );
  NAND4_X1 U5333 ( .A1(n4802), .A2(n4801), .A3(n4800), .A4(n4799), .ZN(n4856)
         );
  INV_X1 U5334 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4804) );
  AOI22_X1 U5335 ( .A1(n4804), .A2(keyinput104), .B1(n4135), .B2(keyinput84), 
        .ZN(n4803) );
  OAI221_X1 U5336 ( .B1(n4804), .B2(keyinput104), .C1(n4135), .C2(keyinput84), 
        .A(n4803), .ZN(n4814) );
  INV_X1 U5337 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4806) );
  AOI22_X1 U5338 ( .A1(n4021), .A2(keyinput30), .B1(keyinput88), .B2(n4806), 
        .ZN(n4805) );
  OAI221_X1 U5339 ( .B1(n4021), .B2(keyinput30), .C1(n4806), .C2(keyinput88), 
        .A(n4805), .ZN(n4813) );
  AOI22_X1 U5340 ( .A1(n4863), .A2(keyinput50), .B1(keyinput29), .B2(n4808), 
        .ZN(n4807) );
  OAI221_X1 U5341 ( .B1(n4863), .B2(keyinput50), .C1(n4808), .C2(keyinput29), 
        .A(n4807), .ZN(n4812) );
  INV_X1 U5342 ( .A(ADDR_REG_10__SCAN_IN), .ZN(n4810) );
  AOI22_X1 U5343 ( .A1(n4916), .A2(keyinput11), .B1(keyinput91), .B2(n4810), 
        .ZN(n4809) );
  OAI221_X1 U5344 ( .B1(n4916), .B2(keyinput11), .C1(n4810), .C2(keyinput91), 
        .A(n4809), .ZN(n4811) );
  NOR4_X1 U5345 ( .A1(n4814), .A2(n4813), .A3(n4812), .A4(n4811), .ZN(n4854)
         );
  OAI22_X1 U5346 ( .A1(keyinput26), .A2(n3126), .B1(n4816), .B2(keyinput10), 
        .ZN(n4815) );
  AOI221_X1 U5347 ( .B1(n3126), .B2(keyinput26), .C1(n4816), .C2(keyinput10), 
        .A(n4815), .ZN(n4824) );
  INV_X1 U5348 ( .A(ADDR_REG_2__SCAN_IN), .ZN(n4914) );
  OAI22_X1 U5349 ( .A1(n4915), .A2(keyinput80), .B1(n4914), .B2(keyinput25), 
        .ZN(n4817) );
  AOI221_X1 U5350 ( .B1(n4915), .B2(keyinput80), .C1(keyinput25), .C2(n4914), 
        .A(n4817), .ZN(n4823) );
  INV_X1 U5351 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n4913) );
  OAI22_X1 U5352 ( .A1(keyinput58), .A2(n3088), .B1(n4913), .B2(keyinput34), 
        .ZN(n4818) );
  AOI221_X1 U5353 ( .B1(n3088), .B2(keyinput58), .C1(n4913), .C2(keyinput34), 
        .A(n4818), .ZN(n4822) );
  OAI22_X1 U5354 ( .A1(n4820), .A2(keyinput68), .B1(n4912), .B2(keyinput51), 
        .ZN(n4819) );
  AOI221_X1 U5355 ( .B1(n4820), .B2(keyinput68), .C1(keyinput51), .C2(n4912), 
        .A(n4819), .ZN(n4821) );
  AND4_X1 U5356 ( .A1(n4824), .A2(n4823), .A3(n4822), .A4(n4821), .ZN(n4853)
         );
  AOI22_X1 U5357 ( .A1(n4826), .A2(keyinput54), .B1(keyinput57), .B2(n4911), 
        .ZN(n4825) );
  OAI221_X1 U5358 ( .B1(n4826), .B2(keyinput54), .C1(n4911), .C2(keyinput57), 
        .A(n4825), .ZN(n4837) );
  INV_X1 U5359 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n4829) );
  AOI22_X1 U5360 ( .A1(n4829), .A2(keyinput61), .B1(keyinput74), .B2(n4828), 
        .ZN(n4827) );
  OAI221_X1 U5361 ( .B1(n4829), .B2(keyinput61), .C1(n4828), .C2(keyinput74), 
        .A(n4827), .ZN(n4836) );
  AOI22_X1 U5362 ( .A1(n4831), .A2(keyinput70), .B1(keyinput53), .B2(n4919), 
        .ZN(n4830) );
  OAI221_X1 U5363 ( .B1(n4831), .B2(keyinput70), .C1(n4919), .C2(keyinput53), 
        .A(n4830), .ZN(n4835) );
  AOI22_X1 U5364 ( .A1(n4918), .A2(keyinput20), .B1(keyinput9), .B2(n4833), 
        .ZN(n4832) );
  OAI221_X1 U5365 ( .B1(n4918), .B2(keyinput20), .C1(n4833), .C2(keyinput9), 
        .A(n4832), .ZN(n4834) );
  NOR4_X1 U5366 ( .A1(n4837), .A2(n4836), .A3(n4835), .A4(n4834), .ZN(n4852)
         );
  AOI22_X1 U5367 ( .A1(n4839), .A2(keyinput19), .B1(keyinput13), .B2(n4917), 
        .ZN(n4838) );
  OAI221_X1 U5368 ( .B1(n4839), .B2(keyinput19), .C1(n4917), .C2(keyinput13), 
        .A(n4838), .ZN(n4850) );
  AOI22_X1 U5369 ( .A1(n4920), .A2(keyinput5), .B1(keyinput81), .B2(n2372), 
        .ZN(n4840) );
  OAI221_X1 U5370 ( .B1(n4920), .B2(keyinput5), .C1(n2372), .C2(keyinput81), 
        .A(n4840), .ZN(n4849) );
  INV_X1 U5371 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4843) );
  AOI22_X1 U5372 ( .A1(n4843), .A2(keyinput65), .B1(n4842), .B2(keyinput85), 
        .ZN(n4841) );
  OAI221_X1 U5373 ( .B1(n4843), .B2(keyinput65), .C1(n4842), .C2(keyinput85), 
        .A(n4841), .ZN(n4848) );
  INV_X1 U5374 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4891) );
  XOR2_X1 U5375 ( .A(n4891), .B(keyinput62), .Z(n4846) );
  XNOR2_X1 U5376 ( .A(IR_REG_2__SCAN_IN), .B(keyinput117), .ZN(n4845) );
  NAND2_X1 U5377 ( .A1(n4846), .A2(n4845), .ZN(n4847) );
  NOR4_X1 U5378 ( .A1(n4850), .A2(n4849), .A3(n4848), .A4(n4847), .ZN(n4851)
         );
  NAND4_X1 U5379 ( .A1(n4854), .A2(n4853), .A3(n4852), .A4(n4851), .ZN(n4855)
         );
  NOR4_X1 U5380 ( .A1(n4858), .A2(n4857), .A3(n4856), .A4(n4855), .ZN(n4859)
         );
  XNOR2_X1 U5381 ( .A(n4860), .B(n4859), .ZN(n4938) );
  NAND4_X1 U5382 ( .A1(REG0_REG_12__SCAN_IN), .A2(REG0_REG_13__SCAN_IN), .A3(
        REG0_REG_8__SCAN_IN), .A4(n4861), .ZN(n4936) );
  NAND4_X1 U5383 ( .A1(REG0_REG_2__SCAN_IN), .A2(REG0_REG_5__SCAN_IN), .A3(
        REG0_REG_1__SCAN_IN), .A4(n4862), .ZN(n4935) );
  NAND4_X1 U5384 ( .A1(REG2_REG_18__SCAN_IN), .A2(REG2_REG_24__SCAN_IN), .A3(
        n4864), .A4(n4863), .ZN(n4865) );
  NOR3_X1 U5385 ( .A1(REG2_REG_28__SCAN_IN), .A2(REG2_REG_21__SCAN_IN), .A3(
        n4865), .ZN(n4876) );
  NAND4_X1 U5386 ( .A1(REG0_REG_27__SCAN_IN), .A2(n4868), .A3(n4867), .A4(
        n4866), .ZN(n4874) );
  NAND4_X1 U5387 ( .A1(REG0_REG_15__SCAN_IN), .A2(REG0_REG_20__SCAN_IN), .A3(
        REG0_REG_14__SCAN_IN), .A4(n4869), .ZN(n4873) );
  NAND4_X1 U5388 ( .A1(REG1_REG_28__SCAN_IN), .A2(REG1_REG_27__SCAN_IN), .A3(
        REG1_REG_25__SCAN_IN), .A4(REG1_REG_24__SCAN_IN), .ZN(n4872) );
  NAND4_X1 U5389 ( .A1(REG1_REG_20__SCAN_IN), .A2(REG1_REG_16__SCAN_IN), .A3(
        REG1_REG_18__SCAN_IN), .A4(n4870), .ZN(n4871) );
  NOR4_X1 U5390 ( .A1(n4874), .A2(n4873), .A3(n4872), .A4(n4871), .ZN(n4875)
         );
  NAND4_X1 U5391 ( .A1(REG1_REG_29__SCAN_IN), .A2(REG2_REG_16__SCAN_IN), .A3(
        n4876), .A4(n4875), .ZN(n4934) );
  NAND4_X1 U5392 ( .A1(REG2_REG_6__SCAN_IN), .A2(REG2_REG_8__SCAN_IN), .A3(
        REG2_REG_3__SCAN_IN), .A4(n2247), .ZN(n4885) );
  NAND4_X1 U5393 ( .A1(n4877), .A2(REG1_REG_4__SCAN_IN), .A3(
        REG3_REG_12__SCAN_IN), .A4(REG1_REG_12__SCAN_IN), .ZN(n4884) );
  INV_X1 U5394 ( .A(IR_REG_21__SCAN_IN), .ZN(n4880) );
  NAND4_X1 U5395 ( .A1(n4880), .A2(n4879), .A3(IR_REG_13__SCAN_IN), .A4(n4878), 
        .ZN(n4883) );
  NAND4_X1 U5396 ( .A1(n4881), .A2(IR_REG_25__SCAN_IN), .A3(IR_REG_22__SCAN_IN), .A4(IR_REG_23__SCAN_IN), .ZN(n4882) );
  NOR4_X1 U5397 ( .A1(n4885), .A2(n4884), .A3(n4883), .A4(n4882), .ZN(n4932)
         );
  AND4_X1 U5398 ( .A1(REG1_REG_7__SCAN_IN), .A2(REG1_REG_2__SCAN_IN), .A3(
        REG1_REG_1__SCAN_IN), .A4(n3104), .ZN(n4889) );
  INV_X1 U5399 ( .A(n4886), .ZN(n4888) );
  AND4_X1 U5400 ( .A1(n4889), .A2(n4888), .A3(n4887), .A4(n2319), .ZN(n4892)
         );
  NAND3_X1 U5401 ( .A1(n4892), .A2(n4891), .A3(n4890), .ZN(n4893) );
  NOR2_X1 U5402 ( .A1(IR_REG_2__SCAN_IN), .A2(n4893), .ZN(n4895) );
  AND4_X1 U5403 ( .A1(n4895), .A2(IR_REG_1__SCAN_IN), .A3(n4894), .A4(
        IR_REG_8__SCAN_IN), .ZN(n4931) );
  NOR4_X1 U5404 ( .A1(DATAI_19_), .A2(DATAI_13_), .A3(DATAI_10_), .A4(DATAI_9_), .ZN(n4896) );
  NAND3_X1 U5405 ( .A1(DATAI_23_), .A2(DATAI_22_), .A3(n4896), .ZN(n4909) );
  NAND4_X1 U5406 ( .A1(D_REG_1__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n4902) );
  NAND4_X1 U5407 ( .A1(REG3_REG_8__SCAN_IN), .A2(n4898), .A3(n2514), .A4(n4897), .ZN(n4901) );
  NAND4_X1 U5408 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n4900) );
  NAND4_X1 U5409 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n4899) );
  NOR4_X1 U5410 ( .A1(n4902), .A2(n4901), .A3(n4900), .A4(n4899), .ZN(n4907)
         );
  NOR4_X1 U5411 ( .A1(DATAI_6_), .A2(DATAI_5_), .A3(DATAI_8_), .A4(n4903), 
        .ZN(n4906) );
  AND4_X1 U5412 ( .A1(n4904), .A2(REG3_REG_23__SCAN_IN), .A3(DATAI_4_), .A4(
        DATAI_3_), .ZN(n4905) );
  NAND3_X1 U5413 ( .A1(n4907), .A2(n4906), .A3(n4905), .ZN(n4908) );
  NOR4_X1 U5414 ( .A1(DATAI_27_), .A2(n4910), .A3(n4909), .A4(n4908), .ZN(
        n4930) );
  NAND4_X1 U5415 ( .A1(DATAO_REG_9__SCAN_IN), .A2(DATAO_REG_17__SCAN_IN), .A3(
        DATAO_REG_18__SCAN_IN), .A4(n4911), .ZN(n4927) );
  NAND4_X1 U5416 ( .A1(DATAO_REG_0__SCAN_IN), .A2(DATAO_REG_3__SCAN_IN), .A3(
        n4913), .A4(n4912), .ZN(n4926) );
  NOR4_X1 U5417 ( .A1(n4915), .A2(n4914), .A3(n3088), .A4(ADDR_REG_5__SCAN_IN), 
        .ZN(n4924) );
  NOR4_X1 U5418 ( .A1(ADDR_REG_14__SCAN_IN), .A2(ADDR_REG_10__SCAN_IN), .A3(
        ADDR_REG_7__SCAN_IN), .A4(n4916), .ZN(n4923) );
  NOR4_X1 U5419 ( .A1(REG3_REG_11__SCAN_IN), .A2(REG3_REG_6__SCAN_IN), .A3(
        DATAO_REG_23__SCAN_IN), .A4(DATAO_REG_24__SCAN_IN), .ZN(n4922) );
  NOR4_X1 U5420 ( .A1(n4920), .A2(n4919), .A3(n4918), .A4(n4917), .ZN(n4921)
         );
  NAND4_X1 U5421 ( .A1(n4924), .A2(n4923), .A3(n4922), .A4(n4921), .ZN(n4925)
         );
  NOR4_X1 U5422 ( .A1(n4928), .A2(n4927), .A3(n4926), .A4(n4925), .ZN(n4929)
         );
  NAND4_X1 U5423 ( .A1(n4932), .A2(n4931), .A3(n4930), .A4(n4929), .ZN(n4933)
         );
  NOR4_X1 U5424 ( .A1(n4936), .A2(n4935), .A3(n4934), .A4(n4933), .ZN(n4937)
         );
  XNOR2_X1 U5425 ( .A(n4938), .B(n4937), .ZN(U3252) );
endmodule

