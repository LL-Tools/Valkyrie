

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091;

  AOI211_X1 U11146 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17384), .A(
        n17383), .B(n17382), .ZN(n17385) );
  INV_X2 U11147 ( .A(n19889), .ZN(n13187) );
  INV_X1 U11148 ( .A(n17723), .ZN(n17715) );
  NAND2_X1 U11149 ( .A1(n15195), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15197) );
  AND2_X1 U11150 ( .A1(n17377), .A2(n12625), .ZN(n15533) );
  BUF_X1 U11151 ( .A(n15766), .Z(n9737) );
  NOR2_X1 U11152 ( .A1(n13429), .A2(n13529), .ZN(n13527) );
  OAI21_X1 U11153 ( .B1(n20735), .B2(n12126), .A(n11944), .ZN(n13430) );
  NAND2_X1 U11154 ( .A1(n13301), .A2(n13300), .ZN(n13333) );
  AND2_X2 U11155 ( .A1(n10215), .A2(n19546), .ZN(n10991) );
  OR2_X1 U11156 ( .A1(n13206), .A2(n13308), .ZN(n13209) );
  INV_X1 U11157 ( .A(n17638), .ZN(n17636) );
  AND2_X1 U11159 ( .A1(n10287), .A2(n10289), .ZN(n10434) );
  CLKBUF_X2 U11161 ( .A(n10596), .Z(n9757) );
  CLKBUF_X1 U11162 ( .A(n12512), .Z(n17026) );
  CLKBUF_X3 U11163 ( .A(n12544), .Z(n17051) );
  CLKBUF_X2 U11165 ( .A(n12512), .Z(n17043) );
  CLKBUF_X1 U11166 ( .A(n12403), .Z(n9711) );
  INV_X1 U11167 ( .A(n12402), .ZN(n17017) );
  CLKBUF_X1 U11168 ( .A(n12543), .Z(n9709) );
  CLKBUF_X3 U11169 ( .A(n12450), .Z(n9717) );
  AND3_X1 U11170 ( .A1(n18709), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n18527), .ZN(n10056) );
  CLKBUF_X2 U11171 ( .A(n11338), .Z(n12173) );
  CLKBUF_X2 U11172 ( .A(n12206), .Z(n12155) );
  CLKBUF_X2 U11173 ( .A(n14301), .Z(n9708) );
  AND2_X2 U11174 ( .A1(n9759), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10372) );
  CLKBUF_X2 U11176 ( .A(n11438), .Z(n11305) );
  CLKBUF_X2 U11177 ( .A(n11337), .Z(n12214) );
  CLKBUF_X2 U11178 ( .A(n11863), .Z(n12207) );
  NOR2_X2 U11179 ( .A1(n10558), .A2(n9763), .ZN(n13914) );
  NOR2_X1 U11180 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14277) );
  NAND2_X1 U11181 ( .A1(n11267), .A2(n13436), .ZN(n11760) );
  AND4_X1 U11182 ( .A1(n11181), .A2(n11180), .A3(n11179), .A4(n11178), .ZN(
        n11182) );
  CLKBUF_X2 U11183 ( .A(n10137), .Z(n9733) );
  AND2_X1 U11184 ( .A1(n10031), .A2(n11159), .ZN(n11863) );
  AND2_X1 U11185 ( .A1(n11157), .A2(n13550), .ZN(n12206) );
  AND2_X1 U11186 ( .A1(n11151), .A2(n13552), .ZN(n12208) );
  NAND3_X1 U11187 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13503) );
  CLKBUF_X1 U11188 ( .A(n18492), .Z(n9702) );
  NOR2_X1 U11189 ( .A1(n18556), .A2(n18395), .ZN(n18492) );
  CLKBUF_X1 U11190 ( .A(n18491), .Z(n9703) );
  AND2_X1 U11191 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10143) );
  AOI21_X1 U11192 ( .B1(n10110), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n10143), .ZN(n10147) );
  XNOR2_X1 U11193 ( .A(n11402), .B(n11400), .ZN(n11920) );
  INV_X1 U11194 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10091) );
  NOR2_X1 U11195 ( .A1(n10195), .A2(n10558), .ZN(n10557) );
  XNOR2_X1 U11196 ( .A(n11538), .B(n11526), .ZN(n11915) );
  BUF_X1 U11197 ( .A(n11274), .Z(n13071) );
  NOR2_X2 U11199 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11159) );
  NAND2_X1 U11200 ( .A1(n9797), .A2(n9779), .ZN(n9879) );
  NAND2_X1 U11201 ( .A1(n10287), .A2(n10280), .ZN(n19380) );
  NAND2_X1 U11202 ( .A1(n18709), .A2(n18686), .ZN(n12370) );
  AND2_X1 U11203 ( .A1(n11335), .A2(n11333), .ZN(n11302) );
  XNOR2_X1 U11204 ( .A(n10757), .B(n10756), .ZN(n10761) );
  AND4_X1 U11205 ( .A1(n10596), .A2(n10558), .A3(n10195), .A4(n10193), .ZN(
        n13009) );
  NAND2_X1 U11207 ( .A1(n13944), .A2(n10478), .ZN(n10479) );
  AND2_X1 U11208 ( .A1(n9971), .A2(n9952), .ZN(n9951) );
  NOR2_X1 U11209 ( .A1(n12370), .A2(n12372), .ZN(n12535) );
  XNOR2_X1 U11211 ( .A(n14373), .B(n10065), .ZN(n15091) );
  XNOR2_X1 U11212 ( .A(n15187), .B(n15188), .ZN(n15203) );
  NOR2_X1 U11213 ( .A1(n10025), .A2(n14190), .ZN(n10083) );
  AND2_X1 U11214 ( .A1(n16442), .A2(n9710), .ZN(n16429) );
  AOI21_X1 U11215 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16496), .A(
        n16688), .ZN(n16484) );
  NOR2_X1 U11216 ( .A1(n17948), .A2(n18547), .ZN(n17971) );
  NAND2_X1 U11217 ( .A1(n17971), .A2(n18090), .ZN(n18037) );
  AND3_X1 U11218 ( .A1(n12401), .A2(n12400), .A3(n12399), .ZN(n18104) );
  INV_X1 U11219 ( .A(n13643), .ZN(n19978) );
  OR3_X1 U11220 ( .A1(n12388), .A2(n12389), .A3(n9848), .ZN(n16678) );
  INV_X1 U11221 ( .A(n17583), .ZN(n17530) );
  INV_X2 U11222 ( .A(n17731), .ZN(n17630) );
  OR2_X1 U11223 ( .A1(n15954), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n9704) );
  INV_X1 U11224 ( .A(n9713), .ZN(n9716) );
  INV_X1 U11225 ( .A(n9713), .ZN(n9715) );
  XOR2_X1 U11226 ( .A(n12358), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .Z(n9705) );
  AND4_X1 U11227 ( .A1(n11169), .A2(n11168), .A3(n11167), .A4(n11166), .ZN(
        n9706) );
  NOR2_X4 U11228 ( .A1(n10650), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10655) );
  OR3_X2 U11229 ( .A1(n15115), .A2(n15114), .A3(n18951), .ZN(n15076) );
  AND2_X4 U11230 ( .A1(n10304), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10296) );
  AND2_X4 U11231 ( .A1(n10304), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9755) );
  NAND2_X1 U11232 ( .A1(n10193), .A2(n9764), .ZN(n10205) );
  AND2_X4 U11233 ( .A1(n11157), .A2(n11160), .ZN(n9752) );
  NAND2_X2 U11234 ( .A1(n11626), .A2(n19978), .ZN(n13065) );
  AND3_X4 U11235 ( .A1(n11264), .A2(n13438), .A3(n11263), .ZN(n11626) );
  NAND2_X2 U11236 ( .A1(n13697), .A2(n13336), .ZN(n13337) );
  NOR2_X1 U11237 ( .A1(n18538), .A2(n12371), .ZN(n12546) );
  AND2_X1 U11238 ( .A1(n11160), .A2(n13270), .ZN(n11337) );
  AND2_X1 U11240 ( .A1(n9754), .A2(n10188), .ZN(n14301) );
  NOR2_X2 U11241 ( .A1(n16223), .A2(n17909), .ZN(n17799) );
  NOR2_X1 U11242 ( .A1(n18539), .A2(n12373), .ZN(n12543) );
  INV_X4 U11243 ( .A(n10088), .ZN(n15766) );
  INV_X2 U11244 ( .A(n9705), .ZN(n9710) );
  OAI21_X2 U11245 ( .B1(n17699), .B2(n12606), .A(n10074), .ZN(n17674) );
  AND2_X2 U11246 ( .A1(n14604), .A2(n14605), .ZN(n14557) );
  NOR2_X1 U11247 ( .A1(n18539), .A2(n12370), .ZN(n12403) );
  AND2_X2 U11249 ( .A1(n13312), .A2(n13700), .ZN(n13334) );
  NAND2_X2 U11251 ( .A1(n15186), .A2(n15185), .ZN(n15187) );
  XNOR2_X2 U11252 ( .A(n14309), .B(n14310), .ZN(n15109) );
  XNOR2_X2 U11253 ( .A(n11360), .B(n19932), .ZN(n13249) );
  INV_X1 U11254 ( .A(n12545), .ZN(n9712) );
  INV_X1 U11255 ( .A(n12545), .ZN(n9713) );
  INV_X4 U11256 ( .A(n9712), .ZN(n9714) );
  NOR2_X1 U11257 ( .A1(n18535), .A2(n12370), .ZN(n12545) );
  AND2_X2 U11258 ( .A1(n15224), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15303) );
  NAND2_X1 U11259 ( .A1(n15094), .A2(n14357), .ZN(n14373) );
  INV_X1 U11260 ( .A(n17107), .ZN(n17103) );
  CLKBUF_X1 U11261 ( .A(n15766), .Z(n9736) );
  NAND2_X1 U11262 ( .A1(n10453), .A2(n10452), .ZN(n10485) );
  BUF_X1 U11263 ( .A(n17724), .Z(n9765) );
  OR2_X1 U11264 ( .A1(n11134), .A2(n15149), .ZN(n15150) );
  NOR2_X1 U11265 ( .A1(n17176), .A2(n17358), .ZN(n17172) );
  NOR2_X1 U11266 ( .A1(n18896), .A2(n12969), .ZN(n15968) );
  BUF_X2 U11268 ( .A(n12777), .Z(n18896) );
  NAND3_X1 U11270 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19697), .A3(n19545), 
        .ZN(n16077) );
  INV_X2 U11271 ( .A(n18534), .ZN(n18549) );
  NAND2_X1 U11272 ( .A1(n12700), .A2(n12696), .ZN(n18534) );
  NAND2_X1 U11273 ( .A1(n19727), .A2(n13687), .ZN(n19447) );
  CLKBUF_X1 U11274 ( .A(n10648), .Z(n10638) );
  AOI21_X1 U11275 ( .B1(n9836), .B2(n14107), .A(n18579), .ZN(n15608) );
  NAND2_X1 U11276 ( .A1(n10229), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9981) );
  NAND2_X1 U11277 ( .A1(n10887), .A2(n9980), .ZN(n9982) );
  INV_X2 U11278 ( .A(n18119), .ZN(n17097) );
  CLKBUF_X3 U11280 ( .A(n10312), .Z(n19737) );
  INV_X1 U11281 ( .A(n10215), .ZN(n10312) );
  INV_X1 U11282 ( .A(n10193), .ZN(n19115) );
  INV_X2 U11284 ( .A(n10558), .ZN(n10203) );
  CLKBUF_X3 U11285 ( .A(n11271), .Z(n19992) );
  NAND2_X4 U11287 ( .A1(n10175), .A2(n10174), .ZN(n10215) );
  OR2_X2 U11288 ( .A1(n11214), .A2(n11213), .ZN(n19996) );
  INV_X4 U11289 ( .A(n12585), .ZN(n9719) );
  CLKBUF_X2 U11290 ( .A(n10353), .Z(n14264) );
  BUF_X2 U11291 ( .A(n10056), .Z(n12571) );
  NOR2_X1 U11292 ( .A1(n18535), .A2(n12373), .ZN(n16686) );
  CLKBUF_X2 U11293 ( .A(n11875), .Z(n12192) );
  INV_X2 U11294 ( .A(n12535), .ZN(n12560) );
  CLKBUF_X1 U11295 ( .A(n10110), .Z(n9742) );
  CLKBUF_X2 U11296 ( .A(n11339), .Z(n12216) );
  CLKBUF_X2 U11297 ( .A(n11224), .Z(n12135) );
  NOR2_X1 U11298 ( .A1(n12372), .A2(n12371), .ZN(n12544) );
  AND2_X2 U11299 ( .A1(n10297), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10352) );
  AND2_X2 U11300 ( .A1(n14277), .A2(n13500), .ZN(n10374) );
  AND2_X1 U11301 ( .A1(n11930), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11151) );
  INV_X4 U11302 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18709) );
  INV_X4 U11303 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n19597) );
  INV_X2 U11304 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n15945) );
  NOR2_X4 U11305 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11158) );
  INV_X4 U11306 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11150) );
  NOR2_X1 U11307 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11152) );
  AND2_X1 U11308 ( .A1(n9799), .A2(n10058), .ZN(n9895) );
  AND3_X1 U11309 ( .A1(n10055), .A2(n14250), .A3(n14249), .ZN(n9802) );
  NAND2_X1 U11310 ( .A1(n10035), .A2(n10034), .ZN(n12936) );
  OAI211_X1 U11311 ( .C1(n14237), .C2(n14236), .A(n14235), .B(n14234), .ZN(
        n14242) );
  AOI21_X1 U11312 ( .B1(n15257), .B2(n16153), .A(n9931), .ZN(n9930) );
  NAND2_X1 U11313 ( .A1(n9968), .A2(n9967), .ZN(n12947) );
  OR2_X1 U11314 ( .A1(n15236), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9968) );
  AND2_X1 U11315 ( .A1(n15303), .A2(n14198), .ZN(n15213) );
  AND2_X1 U11316 ( .A1(n15303), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16005) );
  OR2_X1 U11317 ( .A1(n14474), .A2(n19975), .ZN(n10054) );
  NOR2_X1 U11318 ( .A1(n15330), .A2(n15344), .ZN(n15236) );
  AND2_X1 U11319 ( .A1(n15248), .A2(n12320), .ZN(n12720) );
  NAND2_X1 U11320 ( .A1(n15365), .A2(n9955), .ZN(n15330) );
  AND2_X1 U11321 ( .A1(n16033), .A2(n16032), .ZN(n16108) );
  CLKBUF_X1 U11322 ( .A(n14187), .Z(n14188) );
  AOI21_X1 U11323 ( .B1(n14207), .B2(n14206), .A(n14205), .ZN(n15222) );
  AND2_X1 U11324 ( .A1(n12723), .A2(n12722), .ZN(n14207) );
  NAND2_X1 U11325 ( .A1(n15232), .A2(n15231), .ZN(n15230) );
  OR2_X1 U11326 ( .A1(n14134), .A2(n12825), .ZN(n15180) );
  XNOR2_X1 U11327 ( .A(n14134), .B(n14133), .ZN(n15976) );
  OAI21_X1 U11328 ( .B1(n15374), .B2(n12326), .A(n15372), .ZN(n15356) );
  AND2_X1 U11329 ( .A1(n12823), .A2(n12824), .ZN(n14134) );
  AND2_X1 U11330 ( .A1(n14373), .A2(n10065), .ZN(n14374) );
  NAND2_X1 U11331 ( .A1(n14024), .A2(n14025), .ZN(n14026) );
  NOR2_X1 U11332 ( .A1(n15024), .A2(n15009), .ZN(n15008) );
  OR2_X1 U11333 ( .A1(n15028), .A2(n10934), .ZN(n15188) );
  OR2_X1 U11334 ( .A1(n12810), .A2(n15022), .ZN(n15024) );
  NOR2_X1 U11335 ( .A1(n9803), .A2(n10052), .ZN(n10051) );
  OAI21_X1 U11336 ( .B1(n14025), .B2(n9889), .A(n9885), .ZN(n9884) );
  AND2_X1 U11337 ( .A1(n10736), .A2(n9979), .ZN(n9978) );
  AND2_X1 U11338 ( .A1(n14850), .A2(n14852), .ZN(n14835) );
  INV_X1 U11339 ( .A(n11106), .ZN(n15042) );
  INV_X1 U11340 ( .A(n19290), .ZN(n19306) );
  AND2_X1 U11341 ( .A1(n10635), .A2(n14027), .ZN(n14025) );
  OR3_X1 U11342 ( .A1(n14165), .A2(n14161), .A3(n14164), .ZN(n14847) );
  INV_X1 U11343 ( .A(n10480), .ZN(n13943) );
  OAI21_X1 U11344 ( .B1(n19088), .B2(n19126), .A(n19545), .ZN(n19129) );
  AND2_X1 U11345 ( .A1(n12728), .A2(n10834), .ZN(n14096) );
  AND2_X1 U11346 ( .A1(n10742), .A2(n20973), .ZN(n15301) );
  OAI21_X1 U11347 ( .B1(n14464), .B2(n14139), .A(n14463), .ZN(n14465) );
  OAI21_X1 U11348 ( .B1(n15498), .B2(n15497), .A(n15496), .ZN(n19531) );
  AND2_X1 U11349 ( .A1(n10819), .A2(n10018), .ZN(n12728) );
  OAI21_X1 U11350 ( .B1(n19352), .B2(n19331), .A(n19545), .ZN(n19354) );
  OR2_X1 U11351 ( .A1(n10606), .A2(n13936), .ZN(n10480) );
  INV_X1 U11352 ( .A(n10506), .ZN(n10508) );
  OR3_X1 U11353 ( .A1(n15540), .A2(n10934), .A3(n20973), .ZN(n15299) );
  NOR2_X2 U11354 ( .A1(n16851), .A2(n20981), .ZN(n16854) );
  AND2_X1 U11355 ( .A1(n14146), .A2(n12796), .ZN(n14454) );
  OR2_X1 U11356 ( .A1(n10485), .A2(n10484), .ZN(n10506) );
  XNOR2_X1 U11357 ( .A(n10485), .B(n10481), .ZN(n10627) );
  NAND2_X1 U11358 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17126), .ZN(n17125) );
  NAND2_X1 U11359 ( .A1(n10711), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14209) );
  INV_X1 U11360 ( .A(n10481), .ZN(n10484) );
  INV_X1 U11361 ( .A(n19327), .ZN(n19318) );
  NOR2_X1 U11362 ( .A1(n19132), .A2(n19083), .ZN(n19153) );
  AND2_X1 U11363 ( .A1(n14993), .A2(n14994), .ZN(n14996) );
  INV_X1 U11364 ( .A(n17130), .ZN(n17126) );
  INV_X1 U11365 ( .A(n19243), .ZN(n19245) );
  OR3_X1 U11366 ( .A1(n18796), .A2(n10934), .A3(n15317), .ZN(n14206) );
  AND2_X1 U11367 ( .A1(n13337), .A2(n9956), .ZN(n13520) );
  NAND2_X1 U11368 ( .A1(n19681), .A2(n18937), .ZN(n19405) );
  NAND2_X1 U11369 ( .A1(n10396), .A2(n9881), .ZN(n9880) );
  NAND2_X1 U11370 ( .A1(n11490), .A2(n11489), .ZN(n11518) );
  OR2_X1 U11371 ( .A1(n14101), .A2(n10934), .ZN(n10722) );
  AND2_X1 U11372 ( .A1(n9846), .A2(n10450), .ZN(n10452) );
  OR2_X1 U11373 ( .A1(n18805), .A2(n10934), .ZN(n10719) );
  AND2_X1 U11374 ( .A1(n10476), .A2(n10475), .ZN(n10481) );
  NOR2_X2 U11375 ( .A1(n15150), .A2(n14192), .ZN(n14191) );
  NAND2_X1 U11376 ( .A1(n10715), .A2(n10714), .ZN(n18805) );
  OR2_X1 U11377 ( .A1(n10464), .A2(n10463), .ZN(n10476) );
  NAND2_X1 U11378 ( .A1(n10674), .A2(n15983), .ZN(n10709) );
  AND2_X1 U11379 ( .A1(n14214), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15309) );
  MUX2_X1 U11380 ( .A(n10713), .B(n10712), .S(n9757), .Z(n10715) );
  NOR2_X1 U11381 ( .A1(n14550), .A2(n14539), .ZN(n14538) );
  INV_X1 U11382 ( .A(n10707), .ZN(n10674) );
  NOR2_X1 U11383 ( .A1(n12730), .A2(n10874), .ZN(n14214) );
  OR2_X1 U11384 ( .A1(n10713), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10714) );
  NAND2_X1 U11385 ( .A1(n11447), .A2(n20126), .ZN(n11476) );
  NOR2_X2 U11386 ( .A1(n12733), .A2(n12734), .ZN(n14091) );
  OR2_X1 U11387 ( .A1(n10725), .A2(n15376), .ZN(n15372) );
  NAND2_X1 U11388 ( .A1(n17172), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17171) );
  OR2_X1 U11389 ( .A1(n18835), .A2(n10934), .ZN(n10727) );
  INV_X1 U11390 ( .A(n10341), .ZN(n19221) );
  NAND2_X1 U11391 ( .A1(n9954), .A2(n10289), .ZN(n13678) );
  NAND3_X1 U11392 ( .A1(n12322), .A2(n12321), .A3(n15398), .ZN(n12323) );
  OR2_X1 U11393 ( .A1(n12340), .A2(n12341), .ZN(n12733) );
  NAND2_X1 U11394 ( .A1(n13219), .A2(n13218), .ZN(n13299) );
  AND2_X1 U11395 ( .A1(n13233), .A2(n13214), .ZN(n13223) );
  INV_X2 U11396 ( .A(n13302), .ZN(n10278) );
  NAND2_X1 U11397 ( .A1(n11446), .A2(n11445), .ZN(n20126) );
  NAND2_X1 U11398 ( .A1(n19931), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19932) );
  AND2_X1 U11399 ( .A1(n19064), .A2(n13005), .ZN(n10280) );
  AND2_X1 U11400 ( .A1(n13209), .A2(n13208), .ZN(n13234) );
  OR2_X2 U11401 ( .A1(n14669), .A2(n12903), .ZN(n14672) );
  OR2_X1 U11402 ( .A1(n11402), .A2(n11401), .ZN(n11403) );
  NAND2_X1 U11403 ( .A1(n11359), .A2(n11358), .ZN(n19931) );
  NAND2_X1 U11404 ( .A1(n13204), .A2(n13203), .ZN(n13228) );
  NAND2_X1 U11405 ( .A1(n10936), .A2(n10935), .ZN(n13204) );
  AND2_X1 U11406 ( .A1(n10593), .A2(n19731), .ZN(n10891) );
  AND2_X1 U11407 ( .A1(n10655), .A2(n18964), .ZN(n10657) );
  NOR2_X2 U11408 ( .A1(n19125), .A2(n19737), .ZN(n13769) );
  NOR3_X2 U11409 ( .A1(n17063), .A2(n16632), .A3(n17064), .ZN(n9792) );
  NAND3_X1 U11410 ( .A1(n10236), .A2(n10235), .A3(n10234), .ZN(n10276) );
  AOI21_X1 U11411 ( .B1(n12471), .B2(n14106), .A(n12473), .ZN(n12700) );
  NOR2_X1 U11412 ( .A1(n13107), .A2(n13038), .ZN(n13060) );
  NOR2_X1 U11413 ( .A1(n13152), .A2(n10913), .ZN(n13586) );
  NAND2_X1 U11414 ( .A1(n14108), .A2(n15608), .ZN(n17085) );
  AND2_X1 U11415 ( .A1(n10061), .A2(n10264), .ZN(n10757) );
  NAND2_X1 U11416 ( .A1(n12470), .A2(n12660), .ZN(n17308) );
  AOI21_X1 U11417 ( .B1(n9926), .B2(n10931), .A(n13142), .ZN(n9924) );
  INV_X1 U11418 ( .A(n11333), .ZN(n11334) );
  OR2_X1 U11419 ( .A1(n15516), .A2(n15517), .ZN(n9836) );
  AOI21_X1 U11420 ( .B1(n13324), .B2(n13323), .A(n10904), .ZN(n10912) );
  XNOR2_X1 U11421 ( .A(n13145), .B(n9945), .ZN(n13324) );
  OR2_X1 U11422 ( .A1(n10239), .A2(n10888), .ZN(n15475) );
  NAND4_X1 U11423 ( .A1(n11285), .A2(n11284), .A3(n9992), .A4(n11286), .ZN(
        n11785) );
  AND2_X1 U11424 ( .A1(n18109), .A2(n12695), .ZN(n17305) );
  AND2_X1 U11425 ( .A1(n13148), .A2(n13147), .ZN(n13145) );
  NOR2_X2 U11426 ( .A1(n17401), .A2(n17402), .ZN(n17390) );
  NAND2_X1 U11427 ( .A1(n10853), .A2(n9983), .ZN(n10237) );
  NAND2_X1 U11428 ( .A1(n11644), .A2(n14978), .ZN(n11284) );
  CLKBUF_X1 U11429 ( .A(n10252), .Z(n14129) );
  AND2_X1 U11430 ( .A1(n15609), .A2(n18119), .ZN(n12471) );
  CLKBUF_X2 U11431 ( .A(n9910), .Z(n9732) );
  NAND2_X1 U11432 ( .A1(n17447), .A2(n10080), .ZN(n17401) );
  INV_X1 U11433 ( .A(n13009), .ZN(n10865) );
  NAND2_X1 U11434 ( .A1(n19115), .A2(n10596), .ZN(n10214) );
  NAND2_X1 U11435 ( .A1(n11626), .A2(n13244), .ZN(n13288) );
  AOI211_X1 U11436 ( .C1(n12658), .C2(n12657), .A(n12656), .B(n12655), .ZN(
        n18516) );
  NOR2_X1 U11437 ( .A1(n13263), .A2(n11283), .ZN(n9992) );
  NAND2_X1 U11438 ( .A1(n11281), .A2(n11280), .ZN(n14978) );
  CLKBUF_X1 U11439 ( .A(n10849), .Z(n13135) );
  INV_X1 U11440 ( .A(n17098), .ZN(n18115) );
  INV_X1 U11441 ( .A(n11654), .ZN(n13244) );
  INV_X1 U11442 ( .A(n18090), .ZN(n18728) );
  INV_X1 U11443 ( .A(n20763), .ZN(n15572) );
  CLKBUF_X1 U11444 ( .A(n11653), .Z(n14497) );
  NAND2_X1 U11445 ( .A1(n10528), .A2(n10312), .ZN(n10533) );
  INV_X1 U11446 ( .A(n10551), .ZN(n12783) );
  AND2_X1 U11447 ( .A1(n12311), .A2(n20013), .ZN(n11296) );
  NOR2_X2 U11448 ( .A1(n12457), .A2(n12456), .ZN(n18090) );
  NAND2_X1 U11449 ( .A1(n11272), .A2(n11271), .ZN(n14495) );
  INV_X1 U11450 ( .A(n16237), .ZN(n18190) );
  OR2_X1 U11451 ( .A1(n10394), .A2(n10393), .ZN(n10552) );
  NAND2_X1 U11452 ( .A1(n11777), .A2(n11272), .ZN(n13076) );
  NAND2_X1 U11453 ( .A1(n10216), .A2(n9758), .ZN(n10551) );
  OR2_X1 U11454 ( .A1(n10311), .A2(n10310), .ZN(n10518) );
  NAND2_X2 U11455 ( .A1(n9781), .A2(n9791), .ZN(n12678) );
  OR2_X2 U11456 ( .A1(n11272), .A2(n13643), .ZN(n11744) );
  INV_X1 U11457 ( .A(n10212), .ZN(n10857) );
  INV_X1 U11458 ( .A(n11271), .ZN(n13256) );
  OR2_X1 U11459 ( .A1(n11349), .A2(n11348), .ZN(n11539) );
  OR2_X1 U11460 ( .A1(n11328), .A2(n11327), .ZN(n11415) );
  NAND2_X1 U11462 ( .A1(n10114), .A2(n10113), .ZN(n10212) );
  NAND2_X2 U11463 ( .A1(n9706), .A2(n9790), .ZN(n20013) );
  INV_X1 U11464 ( .A(n9721), .ZN(n11277) );
  AND4_X1 U11465 ( .A1(n11223), .A2(n11222), .A3(n11221), .A4(n11220), .ZN(
        n11240) );
  AND4_X1 U11466 ( .A1(n11232), .A2(n11231), .A3(n11230), .A4(n11229), .ZN(
        n11238) );
  AND4_X1 U11467 ( .A1(n11177), .A2(n11176), .A3(n11175), .A4(n11174), .ZN(
        n11183) );
  OR2_X2 U11468 ( .A1(n11203), .A2(n11202), .ZN(n11272) );
  AND4_X1 U11469 ( .A1(n10106), .A2(n10105), .A3(n10104), .A4(n10103), .ZN(
        n10107) );
  AND2_X1 U11470 ( .A1(n9950), .A2(n9949), .ZN(n10115) );
  AND4_X1 U11471 ( .A1(n11187), .A2(n11186), .A3(n11185), .A4(n11184), .ZN(
        n11193) );
  AND3_X1 U11472 ( .A1(n10152), .A2(n10151), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10155) );
  AND4_X1 U11473 ( .A1(n10096), .A2(n10095), .A3(n10094), .A4(n10093), .ZN(
        n10102) );
  AND4_X1 U11474 ( .A1(n11236), .A2(n11235), .A3(n11234), .A4(n11233), .ZN(
        n11237) );
  AND4_X1 U11475 ( .A1(n11245), .A2(n11244), .A3(n11243), .A4(n11242), .ZN(
        n11261) );
  INV_X2 U11476 ( .A(n16870), .ZN(n12590) );
  AND4_X1 U11477 ( .A1(n11257), .A2(n11256), .A3(n11255), .A4(n11254), .ZN(
        n11258) );
  INV_X1 U11478 ( .A(n16870), .ZN(n17032) );
  AND4_X1 U11479 ( .A1(n11228), .A2(n11227), .A3(n11226), .A4(n11225), .ZN(
        n11239) );
  NAND2_X2 U11480 ( .A1(n18719), .A2(n18607), .ZN(n18658) );
  BUF_X4 U11481 ( .A(n16686), .Z(n9718) );
  INV_X2 U11482 ( .A(n12451), .ZN(n17027) );
  AOI21_X1 U11483 ( .B1(n18555), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12474), .ZN(n12480) );
  INV_X2 U11484 ( .A(n16345), .ZN(U215) );
  NAND2_X2 U11485 ( .A1(n19665), .A2(n19621), .ZN(n19672) );
  NAND2_X2 U11486 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19665), .ZN(n19669) );
  CLKBUF_X1 U11487 ( .A(n9752), .Z(n12168) );
  AND2_X2 U11488 ( .A1(n11161), .A2(n11158), .ZN(n11338) );
  AND2_X2 U11489 ( .A1(n13550), .A2(n14985), .ZN(n11438) );
  AND2_X2 U11490 ( .A1(n11160), .A2(n11159), .ZN(n11875) );
  AND2_X1 U11491 ( .A1(n12654), .A2(n12652), .ZN(n12474) );
  AND2_X1 U11492 ( .A1(n17671), .A2(n12348), .ZN(n17660) );
  OR2_X1 U11493 ( .A1(n12369), .A2(n18538), .ZN(n12402) );
  OR2_X1 U11494 ( .A1(n12372), .A2(n12373), .ZN(n12451) );
  AND2_X2 U11495 ( .A1(n10303), .A2(n10091), .ZN(n9770) );
  INV_X2 U11496 ( .A(n16347), .ZN(n16349) );
  AND2_X2 U11497 ( .A1(n13550), .A2(n13270), .ZN(n12215) );
  AND2_X1 U11498 ( .A1(n11930), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11161) );
  NAND2_X1 U11499 ( .A1(n18686), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12373) );
  CLKBUF_X2 U11500 ( .A(n11159), .Z(n14985) );
  NAND2_X1 U11501 ( .A1(n18703), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n18539) );
  AND2_X2 U11502 ( .A1(n13552), .A2(n11152), .ZN(n9746) );
  AND2_X2 U11503 ( .A1(n13500), .A2(n10091), .ZN(n10297) );
  AND2_X1 U11504 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17671) );
  AND2_X2 U11505 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13270) );
  AND2_X2 U11506 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13552) );
  INV_X2 U11507 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18703) );
  INV_X1 U11508 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10188) );
  INV_X1 U11509 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18686) );
  AND2_X1 U11510 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13500) );
  CLKBUF_X1 U11511 ( .A(n11336), .Z(n11376) );
  NAND2_X1 U11512 ( .A1(n15203), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15272) );
  OR2_X1 U11513 ( .A1(n13643), .A2(n19992), .ZN(n20763) );
  CLKBUF_X1 U11514 ( .A(n11927), .Z(n20438) );
  NOR2_X2 U11515 ( .A1(n9722), .A2(n9723), .ZN(n9721) );
  NAND4_X1 U11516 ( .A1(n11156), .A2(n11155), .A3(n11154), .A4(n11153), .ZN(
        n9722) );
  NAND4_X1 U11517 ( .A1(n11165), .A2(n11164), .A3(n11163), .A4(n11162), .ZN(
        n9723) );
  NOR2_X1 U11518 ( .A1(n17389), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9724) );
  OR2_X1 U11519 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17636), .ZN(
        n9725) );
  OR2_X1 U11520 ( .A1(n17763), .A2(n12622), .ZN(n9726) );
  NAND3_X1 U11521 ( .A1(n9725), .A2(n9726), .A3(n12621), .ZN(n17389) );
  NOR2_X2 U11522 ( .A1(n17520), .A2(n9794), .ZN(n17510) );
  NOR2_X1 U11523 ( .A1(n17389), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17388) );
  XNOR2_X1 U11524 ( .A(n11335), .B(n11334), .ZN(n11929) );
  OAI21_X1 U11525 ( .B1(n11551), .B2(n11550), .A(n11549), .ZN(n14834) );
  INV_X1 U11527 ( .A(n15450), .ZN(n9728) );
  NAND2_X1 U11528 ( .A1(n10238), .A2(n13491), .ZN(n9729) );
  NAND2_X1 U11529 ( .A1(n10510), .A2(n10509), .ZN(n15438) );
  NAND2_X1 U11530 ( .A1(n10238), .A2(n13491), .ZN(n10888) );
  NAND2_X2 U11531 ( .A1(n10228), .A2(n10227), .ZN(n13491) );
  OAI22_X1 U11532 ( .A1(n10243), .A2(n13236), .B1(n19597), .B2(n10242), .ZN(
        n10244) );
  NAND2_X1 U11533 ( .A1(n11364), .A2(n11287), .ZN(n9730) );
  INV_X1 U11534 ( .A(n19996), .ZN(n9731) );
  NAND2_X1 U11535 ( .A1(n11364), .A2(n11287), .ZN(n11369) );
  INV_X1 U11536 ( .A(n19996), .ZN(n11777) );
  NOR2_X2 U11537 ( .A1(n16883), .A2(n16907), .ZN(n16896) );
  NOR2_X4 U11538 ( .A1(n15197), .A2(n14459), .ZN(n14246) );
  INV_X2 U11539 ( .A(n10298), .ZN(n14439) );
  NAND2_X2 U11540 ( .A1(n10575), .A2(n10092), .ZN(n10298) );
  AND2_X2 U11541 ( .A1(n10090), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10304) );
  NOR2_X1 U11542 ( .A1(n12370), .A2(n18538), .ZN(n12450) );
  NOR2_X1 U11543 ( .A1(n13069), .A2(n11771), .ZN(n9910) );
  AND2_X4 U11544 ( .A1(n15473), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10110) );
  NOR2_X2 U11545 ( .A1(n11272), .A2(n19996), .ZN(n13268) );
  AND2_X1 U11546 ( .A1(n13550), .A2(n14985), .ZN(n9734) );
  AND2_X1 U11547 ( .A1(n13550), .A2(n14985), .ZN(n9735) );
  INV_X4 U11548 ( .A(n9786), .ZN(n17050) );
  NAND2_X2 U11549 ( .A1(n10277), .A2(n10276), .ZN(n10275) );
  AOI21_X1 U11550 ( .B1(n10265), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10256), .ZN(n10258) );
  XNOR2_X2 U11551 ( .A(n10247), .B(n10248), .ZN(n10274) );
  NOR2_X2 U11552 ( .A1(n14573), .A2(n14572), .ZN(n14574) );
  AND2_X1 U11553 ( .A1(n13550), .A2(n13270), .ZN(n9738) );
  AND2_X1 U11554 ( .A1(n13550), .A2(n13270), .ZN(n9739) );
  AND2_X1 U11555 ( .A1(n11160), .A2(n11161), .ZN(n11868) );
  AND2_X1 U11556 ( .A1(n11160), .A2(n11161), .ZN(n9768) );
  AND2_X2 U11557 ( .A1(n11160), .A2(n11161), .ZN(n9767) );
  INV_X2 U11558 ( .A(n9719), .ZN(n9740) );
  AND2_X1 U11559 ( .A1(n11161), .A2(n11158), .ZN(n9741) );
  AND2_X4 U11560 ( .A1(n10092), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10303) );
  INV_X1 U11561 ( .A(n12571), .ZN(n9743) );
  AND2_X1 U11562 ( .A1(n11151), .A2(n13552), .ZN(n9744) );
  AND2_X2 U11563 ( .A1(n11151), .A2(n13552), .ZN(n9745) );
  AND2_X2 U11564 ( .A1(n13552), .A2(n11152), .ZN(n9747) );
  AND2_X2 U11565 ( .A1(n13552), .A2(n11152), .ZN(n11381) );
  AND2_X2 U11566 ( .A1(n13500), .A2(n10091), .ZN(n9748) );
  AND2_X2 U11567 ( .A1(n13500), .A2(n10091), .ZN(n9749) );
  AND2_X1 U11568 ( .A1(n11157), .A2(n13550), .ZN(n9750) );
  AND2_X1 U11569 ( .A1(n13550), .A2(n13270), .ZN(n9751) );
  BUF_X4 U11570 ( .A(n14433), .Z(n9753) );
  BUF_X4 U11571 ( .A(n14433), .Z(n9754) );
  AND3_X2 U11572 ( .A1(n15462), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        n10092), .ZN(n14433) );
  NAND2_X1 U11573 ( .A1(n11352), .A2(n11351), .ZN(n11391) );
  OR2_X2 U11574 ( .A1(n14005), .A2(n11545), .ZN(n14861) );
  NOR2_X2 U11575 ( .A1(n13575), .A2(n13605), .ZN(n13604) );
  NOR2_X1 U11576 ( .A1(n14847), .A2(n14849), .ZN(n11551) );
  XNOR2_X2 U11577 ( .A(n11422), .B(n11665), .ZN(n13384) );
  INV_X1 U11578 ( .A(n10298), .ZN(n9756) );
  CLKBUF_X1 U11579 ( .A(n14439), .Z(n9771) );
  XOR2_X2 U11580 ( .A(n12678), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n17722) );
  OAI211_X2 U11581 ( .C1(n11957), .C2(n12126), .A(n11956), .B(n11955), .ZN(
        n13576) );
  OR2_X1 U11582 ( .A1(n15335), .A2(n15363), .ZN(n15366) );
  AOI21_X2 U11583 ( .B1(n14395), .B2(n14394), .A(n14398), .ZN(n15083) );
  NAND2_X4 U11584 ( .A1(n11368), .A2(n20023), .ZN(n20508) );
  NAND2_X2 U11585 ( .A1(n11304), .A2(n11303), .ZN(n20023) );
  XNOR2_X2 U11586 ( .A(n10285), .B(n10275), .ZN(n13206) );
  OAI21_X2 U11587 ( .B1(n10606), .B2(n14238), .A(n18909), .ZN(n10624) );
  XNOR2_X2 U11588 ( .A(n11454), .B(n19961), .ZN(n13482) );
  NAND2_X2 U11589 ( .A1(n11424), .A2(n11423), .ZN(n11454) );
  INV_X2 U11590 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10092) );
  AND4_X2 U11591 ( .A1(n10218), .A2(n10849), .A3(n10557), .A4(n10217), .ZN(
        n10887) );
  NAND2_X1 U11592 ( .A1(n10175), .A2(n10174), .ZN(n9758) );
  INV_X2 U11593 ( .A(n10208), .ZN(n19100) );
  MUX2_X2 U11594 ( .A(n10124), .B(n10123), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10208) );
  NAND2_X2 U11595 ( .A1(n11563), .A2(n14935), .ZN(n14757) );
  INV_X2 U11596 ( .A(n13503), .ZN(n9759) );
  INV_X2 U11597 ( .A(n13503), .ZN(n9760) );
  NOR2_X2 U11598 ( .A1(n13705), .A2(n13834), .ZN(n13827) );
  NAND2_X2 U11599 ( .A1(n10053), .A2(n10051), .ZN(n11555) );
  AND2_X2 U11600 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10575) );
  AND2_X2 U11601 ( .A1(n10287), .A2(n10286), .ZN(n10433) );
  BUF_X2 U11602 ( .A(n13216), .Z(n9761) );
  NAND2_X2 U11603 ( .A1(n10270), .A2(n10261), .ZN(n10760) );
  OAI211_X1 U11604 ( .C1(n12307), .C2(n9996), .A(n9994), .B(n9993), .ZN(n14500) );
  NAND2_X1 U11605 ( .A1(n12838), .A2(n12307), .ZN(n14474) );
  AOI21_X1 U11606 ( .B1(n12308), .B2(n12307), .A(n12894), .ZN(n14754) );
  BUF_X4 U11609 ( .A(n10204), .Z(n9764) );
  NAND2_X2 U11610 ( .A1(n10150), .A2(n10149), .ZN(n10204) );
  AND3_X2 U11611 ( .A1(n9843), .A2(n9841), .A3(n9842), .ZN(n9788) );
  AND2_X2 U11612 ( .A1(n14276), .A2(n14275), .ZN(n14309) );
  OAI21_X2 U11613 ( .B1(n16094), .B2(n14238), .A(n13623), .ZN(n16093) );
  NOR2_X2 U11614 ( .A1(n15109), .A2(n15108), .ZN(n15107) );
  XNOR2_X1 U11615 ( .A(n11922), .B(n11317), .ZN(n14970) );
  NOR2_X2 U11616 ( .A1(n15335), .A2(n12868), .ZN(n15195) );
  NOR2_X2 U11617 ( .A1(n13611), .A2(n9962), .ZN(n14276) );
  NAND2_X2 U11618 ( .A1(n13536), .A2(n13535), .ZN(n13611) );
  NAND2_X2 U11619 ( .A1(n15375), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15335) );
  NOR2_X2 U11620 ( .A1(n15408), .A2(n15379), .ZN(n15375) );
  AND2_X1 U11621 ( .A1(n13302), .A2(n9761), .ZN(n10288) );
  AND2_X1 U11622 ( .A1(n13226), .A2(n13302), .ZN(n9954) );
  OAI21_X1 U11623 ( .B1(n13302), .B2(n13308), .A(n13307), .ZN(n13335) );
  NOR2_X2 U11624 ( .A1(n15104), .A2(n15103), .ZN(n14354) );
  NOR2_X2 U11625 ( .A1(n15107), .A2(n14311), .ZN(n15104) );
  AND2_X2 U11626 ( .A1(n10303), .A2(n10091), .ZN(n9769) );
  AND2_X2 U11627 ( .A1(n10303), .A2(n10091), .ZN(n10295) );
  NAND3_X1 U11628 ( .A1(n9814), .A2(n9981), .A3(n9982), .ZN(n9773) );
  NAND3_X1 U11629 ( .A1(n9814), .A2(n9981), .A3(n9982), .ZN(n9774) );
  AND2_X1 U11630 ( .A1(n15473), .A2(n10092), .ZN(n9775) );
  AND2_X1 U11631 ( .A1(n15473), .A2(n10092), .ZN(n10137) );
  AND2_X2 U11632 ( .A1(n10303), .A2(n14277), .ZN(n10373) );
  AND2_X1 U11633 ( .A1(n12231), .A2(n14631), .ZN(n10006) );
  INV_X1 U11634 ( .A(n14620), .ZN(n12231) );
  INV_X1 U11635 ( .A(n12300), .ZN(n12892) );
  INV_X1 U11637 ( .A(n11491), .ZN(n11489) );
  INV_X1 U11638 ( .A(n12840), .ZN(n11373) );
  NAND2_X1 U11639 ( .A1(n11785), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11287) );
  NOR2_X2 U11640 ( .A1(n11587), .A2(n13073), .ZN(n11617) );
  NAND2_X1 U11641 ( .A1(n19100), .A2(n10212), .ZN(n9984) );
  INV_X1 U11642 ( .A(n14392), .ZN(n13221) );
  INV_X1 U11643 ( .A(n14643), .ZN(n12149) );
  AND2_X1 U11644 ( .A1(n20244), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12891) );
  AND2_X1 U11645 ( .A1(n10088), .A2(n9835), .ZN(n10052) );
  AND2_X1 U11646 ( .A1(n20006), .A2(n19992), .ZN(n11642) );
  AND2_X1 U11647 ( .A1(n11428), .A2(n20640), .ZN(n20285) );
  NAND2_X1 U11648 ( .A1(n10637), .A2(n10636), .ZN(n10648) );
  INV_X1 U11649 ( .A(n10255), .ZN(n9877) );
  NAND2_X1 U11650 ( .A1(n14354), .A2(n14356), .ZN(n14357) );
  NAND2_X1 U11651 ( .A1(n10780), .A2(n10017), .ZN(n10016) );
  INV_X1 U11652 ( .A(n13512), .ZN(n10017) );
  AND2_X1 U11653 ( .A1(n13210), .A2(n10215), .ZN(n14392) );
  INV_X1 U11654 ( .A(n13424), .ZN(n10780) );
  AND3_X1 U11655 ( .A1(n10851), .A2(n9776), .A3(n10215), .ZN(n10213) );
  NOR2_X1 U11656 ( .A1(n12624), .A2(n9918), .ZN(n9917) );
  OR2_X1 U11657 ( .A1(n20758), .A2(n13636), .ZN(n19773) );
  NAND2_X1 U11658 ( .A1(n14538), .A2(n9827), .ZN(n14494) );
  INV_X1 U11659 ( .A(n14476), .ZN(n9901) );
  AND2_X1 U11660 ( .A1(n12205), .A2(n12204), .ZN(n14631) );
  XNOR2_X1 U11661 ( .A(n12942), .B(n14504), .ZN(n13644) );
  NOR2_X1 U11662 ( .A1(n12941), .A2(n14752), .ZN(n12942) );
  AOI21_X1 U11663 ( .B1(n12306), .B2(n12305), .A(n12304), .ZN(n12837) );
  AND2_X1 U11664 ( .A1(n10009), .A2(n10008), .ZN(n10007) );
  INV_X1 U11665 ( .A(n14518), .ZN(n10008) );
  AND2_X1 U11666 ( .A1(n9766), .A2(n20438), .ZN(n20506) );
  AND2_X1 U11667 ( .A1(n12737), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12773) );
  AND2_X1 U11668 ( .A1(n10830), .A2(n10829), .ZN(n12729) );
  INV_X1 U11669 ( .A(n15395), .ZN(n10718) );
  NAND2_X1 U11670 ( .A1(n17217), .A2(n12583), .ZN(n16260) );
  OR2_X1 U11671 ( .A1(n11488), .A2(n11487), .ZN(n11497) );
  OR2_X1 U11672 ( .A1(n11387), .A2(n11386), .ZN(n11413) );
  OR2_X1 U11673 ( .A1(n13643), .A2(n15945), .ZN(n11587) );
  OR2_X1 U11674 ( .A1(n11315), .A2(n11314), .ZN(n11414) );
  INV_X1 U11675 ( .A(n11413), .ZN(n11412) );
  NAND2_X1 U11676 ( .A1(n13643), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11431) );
  AND2_X1 U11677 ( .A1(n20006), .A2(n11262), .ZN(n11215) );
  AOI22_X1 U11678 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9756), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U11679 ( .A1(n10865), .A2(n10850), .ZN(n10231) );
  AND2_X1 U11680 ( .A1(n13206), .A2(n13005), .ZN(n10279) );
  NOR2_X1 U11681 ( .A1(n17101), .A2(n18115), .ZN(n12645) );
  NOR2_X1 U11682 ( .A1(n12467), .A2(n12642), .ZN(n12695) );
  NAND2_X1 U11683 ( .A1(n11293), .A2(n11292), .ZN(n11335) );
  NOR2_X1 U11684 ( .A1(n14545), .A2(n10011), .ZN(n10010) );
  INV_X1 U11685 ( .A(n14558), .ZN(n10011) );
  INV_X1 U11686 ( .A(n12234), .ZN(n12297) );
  OR2_X1 U11687 ( .A1(n14978), .A2(n15945), .ZN(n12234) );
  AND2_X1 U11688 ( .A1(n14677), .A2(n14158), .ZN(n14156) );
  NAND2_X1 U11689 ( .A1(n12028), .A2(n14153), .ZN(n14157) );
  NAND2_X1 U11690 ( .A1(n13071), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12126) );
  INV_X1 U11691 ( .A(n12126), .ZN(n12057) );
  NAND2_X1 U11692 ( .A1(n14828), .A2(n9832), .ZN(n10050) );
  INV_X1 U11693 ( .A(n10050), .ZN(n10045) );
  NAND2_X1 U11694 ( .A1(n11554), .A2(n15766), .ZN(n10046) );
  NAND2_X1 U11695 ( .A1(n14861), .A2(n11546), .ZN(n14159) );
  NAND2_X1 U11696 ( .A1(n11332), .A2(n11331), .ZN(n11360) );
  INV_X1 U11697 ( .A(n11414), .ZN(n11396) );
  OAI21_X1 U11698 ( .B1(n20764), .B2(n15941), .A(n20726), .ZN(n19977) );
  AND2_X1 U11699 ( .A1(n12756), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12737) );
  MUX2_X1 U11700 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n10594), .S(n9764), .Z(n10614) );
  INV_X1 U11701 ( .A(n13949), .ZN(n10021) );
  INV_X1 U11702 ( .A(n13854), .ZN(n10818) );
  NAND2_X1 U11703 ( .A1(n9960), .A2(n9959), .ZN(n9958) );
  NAND2_X1 U11704 ( .A1(n14374), .A2(n9960), .ZN(n9957) );
  INV_X1 U11705 ( .A(n15090), .ZN(n9959) );
  NAND2_X1 U11706 ( .A1(n14091), .A2(n9828), .ZN(n11134) );
  NOR2_X1 U11707 ( .A1(n10533), .A2(n9984), .ZN(n10853) );
  NOR2_X1 U11708 ( .A1(n15204), .A2(n9865), .ZN(n9864) );
  NOR2_X1 U11709 ( .A1(n18778), .A2(n9862), .ZN(n9861) );
  NOR2_X1 U11710 ( .A1(n10029), .A2(n10028), .ZN(n10027) );
  INV_X1 U11711 ( .A(n13733), .ZN(n10028) );
  NOR2_X1 U11712 ( .A1(n10789), .A2(n9875), .ZN(n9874) );
  INV_X1 U11713 ( .A(n12765), .ZN(n9869) );
  NOR2_X1 U11714 ( .A1(n10763), .A2(n9871), .ZN(n9870) );
  AND4_X1 U11715 ( .A1(n10493), .A2(n10492), .A3(n10491), .A4(n10490), .ZN(
        n10500) );
  AND4_X1 U11716 ( .A1(n10497), .A2(n10496), .A3(n10495), .A4(n10494), .ZN(
        n10499) );
  NOR2_X1 U11717 ( .A1(n15025), .A2(n9944), .ZN(n9943) );
  INV_X1 U11718 ( .A(n11138), .ZN(n9944) );
  NAND2_X1 U11719 ( .A1(n10718), .A2(n9839), .ZN(n9842) );
  INV_X1 U11720 ( .A(n10845), .ZN(n10024) );
  AND2_X1 U11721 ( .A1(n9816), .A2(n12335), .ZN(n10020) );
  NAND2_X1 U11722 ( .A1(n12327), .A2(n15354), .ZN(n9892) );
  NOR2_X1 U11723 ( .A1(n15387), .A2(n9940), .ZN(n9939) );
  INV_X1 U11724 ( .A(n13544), .ZN(n9940) );
  AND2_X1 U11725 ( .A1(n9939), .A2(n13630), .ZN(n9938) );
  NAND2_X1 U11726 ( .A1(n10803), .A2(n10030), .ZN(n10029) );
  INV_X1 U11727 ( .A(n15383), .ZN(n10030) );
  AND2_X1 U11728 ( .A1(n10062), .A2(n10646), .ZN(n9985) );
  NAND2_X1 U11729 ( .A1(n12983), .A2(n12984), .ZN(n12985) );
  NAND2_X1 U11730 ( .A1(n14024), .A2(n9805), .ZN(n9986) );
  NAND2_X1 U11731 ( .A1(n9948), .A2(n13238), .ZN(n9947) );
  INV_X1 U11732 ( .A(n13229), .ZN(n9948) );
  NAND2_X1 U11733 ( .A1(n9927), .A2(n13933), .ZN(n9926) );
  INV_X1 U11734 ( .A(n13693), .ZN(n9927) );
  NAND2_X1 U11735 ( .A1(n10396), .A2(n10395), .ZN(n10398) );
  INV_X1 U11736 ( .A(n9880), .ZN(n9878) );
  NOR2_X1 U11737 ( .A1(n10366), .A2(n10365), .ZN(n10893) );
  AND2_X1 U11738 ( .A1(n10851), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9980) );
  INV_X1 U11739 ( .A(n9984), .ZN(n10851) );
  OR2_X1 U11740 ( .A1(n13221), .A2(n13220), .ZN(n13297) );
  NAND2_X1 U11741 ( .A1(n9954), .A2(n10279), .ZN(n10345) );
  NAND2_X1 U11742 ( .A1(n10129), .A2(n10188), .ZN(n10136) );
  BUF_X1 U11743 ( .A(n10430), .Z(n19536) );
  OR2_X1 U11744 ( .A1(n11080), .A2(n16214), .ZN(n13687) );
  OR3_X1 U11745 ( .A1(n10540), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n16204), .ZN(n10566) );
  NOR2_X1 U11746 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18709), .ZN(
        n12652) );
  NAND2_X1 U11747 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n9849) );
  NOR2_X1 U11748 ( .A1(n12369), .A2(n12372), .ZN(n12512) );
  NAND2_X1 U11749 ( .A1(n18709), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12371) );
  NOR2_X1 U11750 ( .A1(n17222), .A2(n12607), .ZN(n12583) );
  AND2_X1 U11751 ( .A1(n18529), .A2(n12645), .ZN(n14106) );
  NOR2_X1 U11752 ( .A1(n12599), .A2(n17708), .ZN(n12601) );
  AOI21_X1 U11753 ( .B1(n12480), .B2(n12479), .A(n12478), .ZN(n12656) );
  AOI211_X1 U11754 ( .C1(n18548), .C2(n18104), .A(n12462), .B(n12461), .ZN(
        n12463) );
  NOR2_X1 U11755 ( .A1(n18109), .A2(n12640), .ZN(n12661) );
  INV_X1 U11756 ( .A(n18519), .ZN(n15508) );
  NAND2_X1 U11757 ( .A1(n12695), .A2(n18530), .ZN(n15516) );
  NAND2_X1 U11758 ( .A1(n9732), .A2(n11655), .ZN(n11659) );
  INV_X1 U11759 ( .A(n11628), .ZN(n13436) );
  NAND2_X1 U11760 ( .A1(n12290), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12302) );
  AND2_X1 U11761 ( .A1(n10006), .A2(n10005), .ZN(n10004) );
  INV_X1 U11762 ( .A(n14614), .ZN(n10005) );
  NOR2_X1 U11763 ( .A1(n12165), .A2(n14822), .ZN(n12185) );
  AND2_X1 U11764 ( .A1(n14676), .A2(n14677), .ZN(n14678) );
  NOR2_X1 U11765 ( .A1(n11959), .A2(n19819), .ZN(n11958) );
  NOR2_X1 U11766 ( .A1(n20835), .A2(n11939), .ZN(n11948) );
  NAND2_X1 U11767 ( .A1(n15766), .A2(n14889), .ZN(n10034) );
  NAND2_X1 U11768 ( .A1(n14784), .A2(n10033), .ZN(n10035) );
  AND2_X1 U11769 ( .A1(n14772), .A2(n9819), .ZN(n10033) );
  OAI21_X1 U11770 ( .B1(n11555), .B2(n11558), .A(n10088), .ZN(n14935) );
  NAND2_X1 U11771 ( .A1(n15781), .A2(n15783), .ZN(n10032) );
  AND2_X1 U11772 ( .A1(n11798), .A2(n11797), .ZN(n15881) );
  NAND2_X1 U11773 ( .A1(n11430), .A2(n11429), .ZN(n20127) );
  NOR2_X1 U11774 ( .A1(n20511), .A2(n20135), .ZN(n20364) );
  NOR2_X1 U11775 ( .A1(n20136), .A2(n20135), .ZN(n20522) );
  NAND2_X1 U11776 ( .A1(n15945), .A2(n19977), .ZN(n20135) );
  AND2_X1 U11777 ( .A1(n11625), .A2(n11624), .ZN(n13280) );
  OR2_X1 U11778 ( .A1(n11588), .A2(n11577), .ZN(n11625) );
  NAND2_X1 U11779 ( .A1(n20957), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15579) );
  AND2_X1 U11780 ( .A1(n10542), .A2(n10541), .ZN(n10572) );
  OR2_X1 U11781 ( .A1(n10540), .A2(n10539), .ZN(n10542) );
  AND2_X1 U11782 ( .A1(n11105), .A2(n10689), .ZN(n11106) );
  AND2_X1 U11783 ( .A1(n11122), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12752) );
  NAND2_X1 U11784 ( .A1(n10675), .A2(n10835), .ZN(n10740) );
  INV_X1 U11785 ( .A(n10709), .ZN(n10675) );
  INV_X1 U11786 ( .A(n13778), .ZN(n10014) );
  AND2_X1 U11787 ( .A1(n16183), .A2(n19731), .ZN(n12997) );
  NAND2_X1 U11788 ( .A1(n10251), .A2(n10250), .ZN(n10272) );
  AND3_X1 U11789 ( .A1(n11007), .A2(n11006), .A3(n11005), .ZN(n13806) );
  NOR2_X1 U11790 ( .A1(n12747), .A2(n15175), .ZN(n12746) );
  OR2_X1 U11791 ( .A1(n12749), .A2(n12871), .ZN(n12747) );
  NAND2_X1 U11792 ( .A1(n12773), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12774) );
  NAND2_X1 U11793 ( .A1(n12760), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12770) );
  AND2_X1 U11794 ( .A1(n10796), .A2(n10795), .ZN(n13800) );
  NAND2_X1 U11795 ( .A1(n9777), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12767) );
  CLKBUF_X1 U11796 ( .A(n10632), .Z(n14238) );
  NAND2_X1 U11797 ( .A1(n9987), .A2(n9988), .ZN(n12920) );
  AOI21_X1 U11798 ( .B1(n12858), .B2(n9834), .A(n9991), .ZN(n9988) );
  INV_X1 U11799 ( .A(n15188), .ZN(n9838) );
  AND2_X1 U11800 ( .A1(n11111), .A2(n11110), .ZN(n15100) );
  NAND2_X1 U11801 ( .A1(n14084), .A2(n15305), .ZN(n10843) );
  NAND2_X1 U11802 ( .A1(n10718), .A2(n10717), .ZN(n9976) );
  AND2_X1 U11803 ( .A1(n11048), .A2(n11047), .ZN(n13852) );
  NAND2_X1 U11804 ( .A1(n9886), .A2(n9883), .ZN(n12325) );
  INV_X1 U11805 ( .A(n9884), .ZN(n9883) );
  AND3_X1 U11806 ( .A1(n10979), .A2(n10978), .A3(n10977), .ZN(n13785) );
  NAND2_X1 U11807 ( .A1(n10168), .A2(n10188), .ZN(n10175) );
  NAND2_X1 U11808 ( .A1(n10173), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10174) );
  NOR2_X1 U11809 ( .A1(n10215), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13007) );
  OAI21_X1 U11810 ( .B1(n13005), .B2(n13308), .A(n13004), .ZN(n13212) );
  XNOR2_X1 U11811 ( .A(n13299), .B(n13297), .ZN(n13222) );
  OR3_X1 U11812 ( .A1(n19281), .A2(n19303), .A3(n19732), .ZN(n19285) );
  NOR2_X1 U11813 ( .A1(n15488), .A2(n19698), .ZN(n13725) );
  NAND2_X1 U11814 ( .A1(n15488), .A2(n19698), .ZN(n19132) );
  NAND2_X1 U11815 ( .A1(n19692), .A2(n19698), .ZN(n19439) );
  NAND2_X1 U11816 ( .A1(n19681), .A2(n19710), .ZN(n19440) );
  NAND2_X1 U11817 ( .A1(n18745), .A2(n16678), .ZN(n12492) );
  INV_X2 U11818 ( .A(n12451), .ZN(n16755) );
  NAND2_X1 U11819 ( .A1(n9915), .A2(n9917), .ZN(n17378) );
  AND2_X1 U11820 ( .A1(n17638), .A2(n17858), .ZN(n12615) );
  AND2_X1 U11821 ( .A1(n17521), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12616) );
  INV_X1 U11822 ( .A(n17215), .ZN(n16252) );
  NAND2_X1 U11823 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18697), .ZN(
        n18538) );
  INV_X1 U11824 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20516) );
  AND2_X1 U11825 ( .A1(n19773), .A2(n13637), .ZN(n19821) );
  INV_X1 U11826 ( .A(n19816), .ZN(n15641) );
  NAND2_X1 U11827 ( .A1(n9903), .A2(n9902), .ZN(n14499) );
  INV_X1 U11828 ( .A(n14494), .ZN(n14475) );
  NAND2_X1 U11829 ( .A1(n12315), .A2(n13183), .ZN(n14669) );
  NAND2_X1 U11830 ( .A1(n13284), .A2(n12314), .ZN(n12315) );
  INV_X1 U11831 ( .A(n14669), .ZN(n14682) );
  NAND2_X1 U11832 ( .A1(n12308), .A2(n9995), .ZN(n9993) );
  NAND2_X1 U11833 ( .A1(n9997), .A2(n12893), .ZN(n9996) );
  NAND2_X1 U11834 ( .A1(n12307), .A2(n9995), .ZN(n9994) );
  OR2_X1 U11835 ( .A1(n19938), .A2(n12841), .ZN(n15795) );
  INV_X1 U11836 ( .A(n19964), .ZN(n15909) );
  INV_X1 U11837 ( .A(n11920), .ZN(n11922) );
  CLKBUF_X1 U11838 ( .A(n14973), .Z(n14974) );
  INV_X1 U11839 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20746) );
  NAND2_X1 U11840 ( .A1(n9856), .A2(n9853), .ZN(n12969) );
  NAND2_X1 U11841 ( .A1(n12777), .A2(n9857), .ZN(n9856) );
  NAND2_X1 U11842 ( .A1(n15538), .A2(n9854), .ZN(n9853) );
  INV_X1 U11843 ( .A(n12971), .ZN(n9857) );
  AND2_X2 U11844 ( .A1(n13010), .A2(n19731), .ZN(n18965) );
  OR2_X1 U11845 ( .A1(n13498), .A2(n13501), .ZN(n13010) );
  INV_X1 U11846 ( .A(n19710), .ZN(n18937) );
  AOI21_X1 U11847 ( .B1(n18799), .B2(n19063), .A(n12741), .ZN(n12742) );
  OR2_X1 U11848 ( .A1(n18757), .A2(n19737), .ZN(n16084) );
  NAND2_X1 U11849 ( .A1(n18757), .A2(n11081), .ZN(n16100) );
  INV_X1 U11850 ( .A(n16090), .ZN(n19061) );
  INV_X1 U11851 ( .A(n16077), .ZN(n19063) );
  OR2_X1 U11852 ( .A1(n14996), .A2(n14995), .ZN(n15253) );
  NAND2_X1 U11853 ( .A1(n15255), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9934) );
  NAND2_X1 U11854 ( .A1(n9933), .A2(n16143), .ZN(n9932) );
  OAI21_X1 U11855 ( .B1(n16005), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15214), .ZN(n11079) );
  NAND2_X1 U11856 ( .A1(n9978), .A2(n9973), .ZN(n9972) );
  NAND2_X1 U11857 ( .A1(n10718), .A2(n10717), .ZN(n9973) );
  XNOR2_X1 U11858 ( .A(n12725), .B(n9815), .ZN(n12743) );
  OAI21_X1 U11859 ( .B1(n12720), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15223), .ZN(n12736) );
  INV_X1 U11860 ( .A(n12720), .ZN(n9967) );
  AND2_X1 U11861 ( .A1(n10891), .A2(n19719), .ZN(n19069) );
  NAND2_X1 U11862 ( .A1(n10891), .A2(n19720), .ZN(n19074) );
  INV_X1 U11863 ( .A(n19069), .ZN(n16163) );
  INV_X1 U11864 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19708) );
  INV_X1 U11865 ( .A(n15488), .ZN(n19692) );
  INV_X1 U11866 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19689) );
  AND2_X1 U11867 ( .A1(n13303), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19585) );
  INV_X1 U11868 ( .A(n16731), .ZN(n16706) );
  INV_X1 U11869 ( .A(n16725), .ZN(n16693) );
  AOI211_X1 U11870 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18728), .A(n12488), .B(
        n12492), .ZN(n16732) );
  INV_X1 U11871 ( .A(n17040), .ZN(n17012) );
  NOR2_X1 U11872 ( .A1(n17135), .A2(n18119), .ZN(n17131) );
  NAND2_X1 U11873 ( .A1(n17131), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17130) );
  NAND2_X1 U11874 ( .A1(n12884), .A2(n17980), .ZN(n12715) );
  NOR2_X2 U11875 ( .A1(n12626), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17377) );
  NOR2_X1 U11876 ( .A1(n17388), .A2(n12624), .ZN(n12626) );
  INV_X1 U11877 ( .A(n17907), .ZN(n17980) );
  NOR2_X1 U11878 ( .A1(n18521), .A2(n18050), .ZN(n18048) );
  OR2_X1 U11879 ( .A1(n11598), .A2(n11597), .ZN(n11614) );
  AND2_X1 U11880 ( .A1(n10436), .A2(n10435), .ZN(n9847) );
  OAI22_X1 U11881 ( .A1(n10345), .A2(n13211), .B1(n10344), .B2(n10343), .ZN(
        n10346) );
  AOI22_X1 U11882 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10314), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10291) );
  OR2_X1 U11883 ( .A1(n12479), .A2(n12480), .ZN(n12475) );
  OR2_X1 U11884 ( .A1(n11466), .A2(n11465), .ZN(n11494) );
  AND2_X2 U11885 ( .A1(n11149), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11157) );
  INV_X1 U11886 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11149) );
  OR3_X1 U11887 ( .A1(n11613), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n19973), .ZN(n11615) );
  NAND2_X1 U11888 ( .A1(n11432), .A2(n11431), .ZN(n11598) );
  NOR2_X2 U11889 ( .A1(n10694), .A2(n10693), .ZN(n10692) );
  INV_X1 U11890 ( .A(n14394), .ZN(n9960) );
  AND4_X1 U11891 ( .A1(n10489), .A2(n10488), .A3(n10487), .A4(n10486), .ZN(
        n10501) );
  NAND2_X1 U11892 ( .A1(n9975), .A2(n15299), .ZN(n9974) );
  OR2_X1 U11893 ( .A1(n10448), .A2(n10447), .ZN(n10602) );
  AND2_X1 U11894 ( .A1(n10395), .A2(n10313), .ZN(n9881) );
  INV_X1 U11895 ( .A(n10552), .ZN(n10907) );
  AND2_X1 U11896 ( .A1(n19737), .A2(n10176), .ZN(n9882) );
  OR2_X1 U11897 ( .A1(n10380), .A2(n10379), .ZN(n10595) );
  AND2_X1 U11898 ( .A1(n10555), .A2(n10203), .ZN(n10207) );
  NAND2_X1 U11899 ( .A1(n10290), .A2(n10286), .ZN(n10316) );
  NAND2_X1 U11900 ( .A1(n10575), .A2(n9807), .ZN(n9949) );
  NOR2_X1 U11901 ( .A1(n17230), .A2(n12584), .ZN(n12602) );
  AND2_X1 U11902 ( .A1(n12678), .A2(n17730), .ZN(n12674) );
  NAND2_X1 U11903 ( .A1(n11301), .A2(n9789), .ZN(n11333) );
  NAND2_X1 U11904 ( .A1(n11744), .A2(n14495), .ZN(n11653) );
  NAND2_X1 U11905 ( .A1(n11262), .A2(n20013), .ZN(n11628) );
  AND2_X1 U11906 ( .A1(n11812), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12290) );
  AND2_X1 U11907 ( .A1(n10010), .A2(n12283), .ZN(n10009) );
  NOR2_X1 U11908 ( .A1(n12258), .A2(n14796), .ZN(n12268) );
  INV_X1 U11909 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12041) );
  NAND2_X1 U11910 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11939) );
  NOR2_X1 U11911 ( .A1(n9909), .A2(n9908), .ZN(n9907) );
  INV_X1 U11912 ( .A(n14629), .ZN(n9908) );
  INV_X1 U11913 ( .A(n14633), .ZN(n9909) );
  NOR2_X1 U11914 ( .A1(n14654), .A2(n9899), .ZN(n9898) );
  INV_X1 U11915 ( .A(n14073), .ZN(n9899) );
  OR2_X1 U11916 ( .A1(n11687), .A2(n9913), .ZN(n9912) );
  INV_X1 U11917 ( .A(n13837), .ZN(n9913) );
  AND2_X1 U11918 ( .A1(n11521), .A2(n11520), .ZN(n11522) );
  OR2_X1 U11919 ( .A1(n11273), .A2(n14495), .ZN(n11778) );
  AND2_X1 U11920 ( .A1(n13280), .A2(n11786), .ZN(n12310) );
  NAND2_X1 U11921 ( .A1(n11929), .A2(n15945), .ZN(n11352) );
  AND2_X1 U11922 ( .A1(n11399), .A2(n11398), .ZN(n11400) );
  OAI211_X1 U11923 ( .C1(n19987), .C2(n11373), .A(n11372), .B(n11371), .ZN(
        n11374) );
  NAND2_X1 U11924 ( .A1(n11370), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11372) );
  XNOR2_X1 U11925 ( .A(n10041), .B(n11389), .ZN(n11408) );
  NAND2_X1 U11926 ( .A1(n10039), .A2(n9817), .ZN(n10041) );
  NAND2_X1 U11927 ( .A1(n11274), .A2(n20006), .ZN(n11278) );
  NOR2_X1 U11928 ( .A1(n19992), .A2(n20006), .ZN(n11265) );
  AND2_X2 U11929 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13550) );
  INV_X1 U11930 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20284) );
  NAND2_X1 U11931 ( .A1(n11289), .A2(n11288), .ZN(n11290) );
  AOI22_X1 U11932 ( .A1(n11339), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_7__6__SCAN_IN), .B2(n12213), .ZN(n11178) );
  OR2_X1 U11933 ( .A1(n11613), .A2(n11574), .ZN(n11576) );
  NAND2_X1 U11934 ( .A1(n11617), .A2(n11642), .ZN(n11588) );
  NAND2_X1 U11935 ( .A1(n10533), .A2(n10551), .ZN(n10849) );
  INV_X1 U11936 ( .A(n12857), .ZN(n12861) );
  NAND2_X1 U11937 ( .A1(n10148), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10149) );
  NAND2_X1 U11938 ( .A1(n10142), .A2(n10188), .ZN(n10150) );
  NAND2_X1 U11939 ( .A1(n10657), .A2(n13541), .ZN(n10667) );
  OR2_X1 U11940 ( .A1(n10474), .A2(n10473), .ZN(n10628) );
  NAND2_X1 U11941 ( .A1(n9963), .A2(n13868), .ZN(n9962) );
  OR2_X1 U11942 ( .A1(n11094), .A2(n11093), .ZN(n9841) );
  AND2_X1 U11943 ( .A1(n13967), .A2(n9888), .ZN(n9887) );
  AOI21_X1 U11944 ( .B1(n9888), .B2(n16071), .A(n12323), .ZN(n9885) );
  NAND2_X1 U11945 ( .A1(n15438), .A2(n9833), .ZN(n15408) );
  NOR2_X1 U11946 ( .A1(n16114), .A2(n20889), .ZN(n9961) );
  AND3_X1 U11947 ( .A1(n10924), .A2(n10923), .A3(n10922), .ZN(n13693) );
  INV_X1 U11948 ( .A(n10595), .ZN(n10900) );
  XNOR2_X1 U11949 ( .A(n10912), .B(n10911), .ZN(n13154) );
  NAND2_X1 U11950 ( .A1(n13003), .A2(n19546), .ZN(n13306) );
  OR2_X1 U11951 ( .A1(n13221), .A2(n13211), .ZN(n13213) );
  AND2_X1 U11952 ( .A1(n13914), .A2(n10193), .ZN(n9983) );
  NAND2_X1 U11953 ( .A1(n10287), .A2(n10279), .ZN(n10340) );
  NAND2_X1 U11954 ( .A1(n10290), .A2(n10280), .ZN(n10326) );
  NOR2_X1 U11955 ( .A1(n17097), .A2(n12434), .ZN(n12468) );
  NAND2_X1 U11956 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12369) );
  NAND2_X1 U11957 ( .A1(n18746), .A2(n16358), .ZN(n15510) );
  NAND2_X1 U11958 ( .A1(n15510), .A2(n17308), .ZN(n12473) );
  AND2_X1 U11959 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12609), .ZN(
        n12610) );
  OAI21_X1 U11960 ( .B1(n12582), .B2(n16252), .A(n17636), .ZN(n12612) );
  XNOR2_X1 U11961 ( .A(n17235), .B(n12678), .ZN(n12598) );
  NOR2_X1 U11962 ( .A1(n15611), .A2(n12465), .ZN(n12647) );
  NAND3_X1 U11963 ( .A1(n12444), .A2(n12443), .A3(n12442), .ZN(n12640) );
  AOI211_X1 U11964 ( .C1(n9718), .C2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n12441), .B(n12440), .ZN(n12442) );
  INV_X1 U11965 ( .A(n15512), .ZN(n15610) );
  OAI21_X1 U11966 ( .B1(n15519), .B2(n15511), .A(n15513), .ZN(n15512) );
  INV_X1 U11967 ( .A(n17308), .ZN(n15511) );
  INV_X1 U11968 ( .A(n12239), .ZN(n11811) );
  NAND2_X1 U11969 ( .A1(n13647), .A2(n13649), .ZN(n19845) );
  INV_X1 U11970 ( .A(n19773), .ZN(n19803) );
  NAND2_X1 U11971 ( .A1(n19773), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13642) );
  OR2_X1 U11972 ( .A1(n14494), .A2(n9904), .ZN(n9903) );
  INV_X1 U11973 ( .A(n14496), .ZN(n9904) );
  NAND2_X1 U11974 ( .A1(n14634), .A2(n9907), .ZN(n14628) );
  AND2_X1 U11975 ( .A1(n14634), .A2(n14633), .ZN(n14636) );
  AND2_X1 U11976 ( .A1(n11699), .A2(n11698), .ZN(n13928) );
  NAND2_X1 U11977 ( .A1(n13398), .A2(n13244), .ZN(n9914) );
  NAND2_X1 U11978 ( .A1(n15728), .A2(n13436), .ZN(n13439) );
  INV_X1 U11979 ( .A(n19976), .ZN(n19974) );
  INV_X1 U11980 ( .A(n12308), .ZN(n9997) );
  INV_X1 U11981 ( .A(n12893), .ZN(n9995) );
  OR2_X1 U11982 ( .A1(n12294), .A2(n12293), .ZN(n14518) );
  OR2_X1 U11983 ( .A1(n12272), .A2(n12271), .ZN(n14545) );
  AOI21_X1 U11984 ( .B1(n12261), .B2(n12260), .A(n12259), .ZN(n14558) );
  AND2_X1 U11985 ( .A1(n14800), .A2(n12303), .ZN(n12259) );
  NOR2_X1 U11986 ( .A1(n12203), .A2(n12199), .ZN(n12228) );
  NAND2_X1 U11987 ( .A1(n12228), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12239) );
  AND2_X1 U11988 ( .A1(n12187), .A2(n12186), .ZN(n14637) );
  NAND2_X1 U11989 ( .A1(n12146), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12165) );
  AND2_X1 U11990 ( .A1(n12130), .A2(n14156), .ZN(n10012) );
  AND2_X1 U11991 ( .A1(n14072), .A2(n14069), .ZN(n12130) );
  NOR2_X1 U11992 ( .A1(n12097), .A2(n12096), .ZN(n12093) );
  NAND2_X1 U11993 ( .A1(n12093), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12092) );
  AND2_X1 U11994 ( .A1(n14157), .A2(n14156), .ZN(n14070) );
  NAND2_X1 U11995 ( .A1(n12112), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12097) );
  INV_X1 U11996 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12096) );
  OR2_X1 U11997 ( .A1(n14666), .A2(n14589), .ZN(n14651) );
  OR2_X1 U11998 ( .A1(n14664), .A2(n14663), .ZN(n14666) );
  OR2_X1 U11999 ( .A1(n12040), .A2(n12041), .ZN(n12058) );
  AND2_X1 U12000 ( .A1(n11995), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12025) );
  NAND2_X1 U12001 ( .A1(n12025), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12040) );
  NOR2_X1 U12002 ( .A1(n11981), .A2(n19779), .ZN(n11995) );
  NAND2_X1 U12003 ( .A1(n11966), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11981) );
  AND2_X1 U12004 ( .A1(n11980), .A2(n11979), .ZN(n13834) );
  NAND2_X1 U12005 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n11958), .ZN(
        n11912) );
  AOI21_X1 U12006 ( .B1(n11964), .B2(n12057), .A(n11963), .ZN(n13605) );
  INV_X1 U12007 ( .A(n11947), .ZN(n11954) );
  NAND2_X1 U12008 ( .A1(n11954), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11959) );
  AOI21_X1 U12009 ( .B1(n11953), .B2(n12057), .A(n11952), .ZN(n13529) );
  CLKBUF_X1 U12010 ( .A(n13527), .Z(n13528) );
  AOI21_X1 U12011 ( .B1(n11919), .B2(n12126), .A(n10002), .ZN(n10001) );
  INV_X1 U12012 ( .A(n11938), .ZN(n10002) );
  OR2_X1 U12013 ( .A1(n14565), .A2(n14548), .ZN(n14550) );
  AND2_X1 U12014 ( .A1(n14616), .A2(n14607), .ZN(n14609) );
  NAND2_X1 U12015 ( .A1(n14609), .A2(n14563), .ZN(n14565) );
  NAND2_X1 U12016 ( .A1(n14634), .A2(n9905), .ZN(n14624) );
  NOR2_X1 U12017 ( .A1(n14622), .A2(n9906), .ZN(n9905) );
  INV_X1 U12018 ( .A(n9907), .ZN(n9906) );
  NOR2_X1 U12019 ( .A1(n14624), .A2(n14617), .ZN(n14616) );
  NAND2_X1 U12020 ( .A1(n10044), .A2(n10048), .ZN(n14936) );
  INV_X1 U12021 ( .A(n10049), .ZN(n10048) );
  OAI21_X1 U12022 ( .B1(n10051), .B2(n10050), .A(n9737), .ZN(n10049) );
  NOR2_X1 U12023 ( .A1(n14647), .A2(n14576), .ZN(n14634) );
  NAND2_X1 U12024 ( .A1(n10047), .A2(n10046), .ZN(n10053) );
  NAND2_X1 U12025 ( .A1(n11715), .A2(n9896), .ZN(n14647) );
  NOR2_X1 U12026 ( .A1(n9897), .A2(n14644), .ZN(n9896) );
  INV_X1 U12027 ( .A(n9898), .ZN(n9897) );
  NAND2_X1 U12028 ( .A1(n11715), .A2(n9898), .ZN(n14645) );
  AND2_X1 U12029 ( .A1(n11715), .A2(n9900), .ZN(n14656) );
  AND2_X1 U12030 ( .A1(n14983), .A2(n15945), .ZN(n12840) );
  OR2_X1 U12031 ( .A1(n15766), .A2(n11548), .ZN(n14850) );
  AND2_X1 U12032 ( .A1(n11711), .A2(n11710), .ZN(n14667) );
  INV_X1 U12033 ( .A(n11715), .ZN(n14655) );
  AND2_X1 U12034 ( .A1(n15766), .A2(n14162), .ZN(n14164) );
  OR2_X1 U12035 ( .A1(n13927), .A2(n13928), .ZN(n14014) );
  NOR2_X1 U12036 ( .A1(n14014), .A2(n14015), .ZN(n14674) );
  OR2_X1 U12037 ( .A1(n13711), .A2(n9911), .ZN(n13927) );
  OR2_X1 U12038 ( .A1(n9912), .A2(n13830), .ZN(n9911) );
  OR2_X1 U12039 ( .A1(n13711), .A2(n9912), .ZN(n13836) );
  NOR2_X1 U12040 ( .A1(n13711), .A2(n11687), .ZN(n13838) );
  NAND2_X1 U12041 ( .A1(n11679), .A2(n11678), .ZN(n13711) );
  NOR2_X1 U12042 ( .A1(n13579), .A2(n13578), .ZN(n11678) );
  INV_X1 U12043 ( .A(n13580), .ZN(n11679) );
  NAND2_X1 U12044 ( .A1(n13387), .A2(n13433), .ZN(n13580) );
  NAND2_X1 U12045 ( .A1(n11421), .A2(n11420), .ZN(n13385) );
  NAND2_X1 U12046 ( .A1(n11795), .A2(n15548), .ZN(n15848) );
  BUF_X1 U12047 ( .A(n11425), .Z(n13314) );
  OR2_X1 U12048 ( .A1(n20092), .A2(n9766), .ZN(n20022) );
  INV_X1 U12049 ( .A(n20742), .ZN(n20409) );
  INV_X1 U12050 ( .A(n20438), .ZN(n20470) );
  NOR2_X1 U12051 ( .A1(n20588), .A2(n9766), .ZN(n20476) );
  INV_X1 U12052 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20579) );
  AND3_X1 U12053 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n15945), .A3(n19977), 
        .ZN(n20014) );
  NAND2_X1 U12054 ( .A1(n9766), .A2(n20470), .ZN(n20253) );
  OR2_X1 U12055 ( .A1(n14974), .A2(n19979), .ZN(n20588) );
  AOI21_X1 U12056 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20471), .A(n20135), 
        .ZN(n20589) );
  OAI21_X1 U12057 ( .B1(n10552), .B2(n10551), .A(n10550), .ZN(n10594) );
  NAND2_X1 U12058 ( .A1(n15953), .A2(n12848), .ZN(n12855) );
  NOR2_X1 U12059 ( .A1(n12971), .A2(n9855), .ZN(n9854) );
  INV_X1 U12060 ( .A(n16010), .ZN(n9855) );
  INV_X1 U12061 ( .A(n18870), .ZN(n12777) );
  NAND2_X1 U12062 ( .A1(n10737), .A2(n10738), .ZN(n10744) );
  NAND2_X1 U12063 ( .A1(n10680), .A2(n10673), .ZN(n10707) );
  AND2_X1 U12064 ( .A1(n10652), .A2(n10651), .ZN(n18865) );
  OAI21_X1 U12065 ( .B1(n9763), .B2(P2_EBX_REG_5__SCAN_IN), .A(n10925), .ZN(
        n10603) );
  CLKBUF_X1 U12066 ( .A(n10607), .Z(n10620) );
  NAND2_X1 U12067 ( .A1(n9876), .A2(n10257), .ZN(n10260) );
  NOR2_X1 U12068 ( .A1(n18896), .A2(n15049), .ZN(n15064) );
  NAND2_X1 U12069 ( .A1(n10819), .A2(n10020), .ZN(n12334) );
  AND2_X1 U12070 ( .A1(n10819), .A2(n9816), .ZN(n13951) );
  AND2_X1 U12071 ( .A1(n10817), .A2(n10816), .ZN(n13854) );
  NAND2_X1 U12072 ( .A1(n10819), .A2(n10818), .ZN(n13950) );
  AND2_X1 U12073 ( .A1(n13614), .A2(n9964), .ZN(n9963) );
  INV_X1 U12074 ( .A(n18952), .ZN(n9964) );
  NOR2_X1 U12075 ( .A1(n13613), .A2(n13612), .ZN(n13614) );
  INV_X1 U12076 ( .A(n13611), .ZN(n9965) );
  AND2_X1 U12077 ( .A1(n10785), .A2(n10784), .ZN(n13512) );
  NOR2_X1 U12078 ( .A1(n15089), .A2(n14374), .ZN(n14395) );
  AND2_X1 U12079 ( .A1(n14309), .A2(n14310), .ZN(n14311) );
  OR2_X1 U12080 ( .A1(n15980), .A2(n15979), .ZN(n15982) );
  OR2_X1 U12081 ( .A1(n15982), .A2(n14271), .ZN(n15164) );
  AND2_X1 U12082 ( .A1(n11054), .A2(n11053), .ZN(n12734) );
  OR2_X1 U12083 ( .A1(n18944), .A2(n18943), .ZN(n18946) );
  AND3_X1 U12084 ( .A1(n11033), .A2(n11032), .A3(n11031), .ZN(n15387) );
  AND3_X1 U12085 ( .A1(n10952), .A2(n10951), .A3(n10950), .ZN(n13229) );
  INV_X1 U12086 ( .A(n12965), .ZN(n13917) );
  NAND2_X1 U12087 ( .A1(n12752), .A2(n9785), .ZN(n12749) );
  NAND2_X1 U12088 ( .A1(n12752), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12750) );
  NAND2_X1 U12089 ( .A1(n12773), .A2(n9784), .ZN(n12776) );
  NOR2_X1 U12090 ( .A1(n12770), .A2(n10809), .ZN(n12758) );
  NAND2_X1 U12091 ( .A1(n9874), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9873) );
  INV_X1 U12092 ( .A(n12768), .ZN(n9872) );
  NOR2_X1 U12093 ( .A1(n12768), .A2(n10789), .ZN(n12769) );
  NAND2_X1 U12094 ( .A1(n12761), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12768) );
  AND2_X1 U12095 ( .A1(n10779), .A2(n10778), .ZN(n13424) );
  NAND2_X1 U12096 ( .A1(n10015), .A2(n10780), .ZN(n13513) );
  INV_X1 U12097 ( .A(n13406), .ZN(n10015) );
  NOR2_X1 U12098 ( .A1(n9868), .A2(n14032), .ZN(n9867) );
  INV_X1 U12099 ( .A(n9870), .ZN(n9868) );
  NOR2_X1 U12100 ( .A1(n12765), .A2(n10763), .ZN(n12766) );
  AND2_X1 U12101 ( .A1(n10766), .A2(n10765), .ZN(n13340) );
  NAND2_X1 U12102 ( .A1(n12763), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12765) );
  NAND2_X1 U12103 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12764) );
  INV_X1 U12104 ( .A(n10761), .ZN(n10269) );
  AND2_X1 U12105 ( .A1(n9943), .A2(n9942), .ZN(n9941) );
  INV_X1 U12106 ( .A(n15010), .ZN(n9942) );
  INV_X1 U12107 ( .A(n15256), .ZN(n9933) );
  NAND2_X1 U12108 ( .A1(n14191), .A2(n9943), .ZN(n15027) );
  NOR2_X1 U12109 ( .A1(n15042), .A2(n11107), .ZN(n14185) );
  AND2_X1 U12110 ( .A1(n9824), .A2(n10023), .ZN(n10022) );
  INV_X1 U12111 ( .A(n15100), .ZN(n10023) );
  NAND2_X1 U12112 ( .A1(n14084), .A2(n9824), .ZN(n15101) );
  INV_X1 U12113 ( .A(n15301), .ZN(n9979) );
  AND2_X1 U12114 ( .A1(n14091), .A2(n14090), .ZN(n14093) );
  AND2_X1 U12115 ( .A1(n10833), .A2(n10832), .ZN(n14094) );
  AND2_X1 U12116 ( .A1(n10020), .A2(n10019), .ZN(n10018) );
  INV_X1 U12117 ( .A(n12729), .ZN(n10019) );
  NOR2_X2 U12118 ( .A1(n15335), .A2(n10511), .ZN(n15224) );
  AOI21_X1 U12119 ( .B1(n15356), .B2(n9893), .A(n9891), .ZN(n15232) );
  NOR2_X1 U12120 ( .A1(n15242), .A2(n9894), .ZN(n9893) );
  INV_X1 U12121 ( .A(n15354), .ZN(n9894) );
  AND2_X1 U12122 ( .A1(n12331), .A2(n12330), .ZN(n15231) );
  AND2_X1 U12123 ( .A1(n9938), .A2(n9937), .ZN(n9936) );
  INV_X1 U12124 ( .A(n13852), .ZN(n9937) );
  AND2_X1 U12125 ( .A1(n10808), .A2(n10807), .ZN(n15383) );
  INV_X1 U12126 ( .A(n13800), .ZN(n10797) );
  NAND2_X1 U12127 ( .A1(n10026), .A2(n10803), .ZN(n15384) );
  NAND2_X1 U12128 ( .A1(n9986), .A2(n9985), .ZN(n12324) );
  OR2_X1 U12129 ( .A1(n9947), .A2(n13785), .ZN(n9946) );
  NAND2_X1 U12130 ( .A1(n13932), .A2(n10931), .ZN(n13143) );
  NAND2_X1 U12131 ( .A1(n13944), .A2(n10480), .ZN(n10477) );
  OR2_X1 U12132 ( .A1(n13587), .A2(n9926), .ZN(n13932) );
  AND2_X1 U12133 ( .A1(n10755), .A2(n10754), .ZN(n13746) );
  NAND2_X1 U12134 ( .A1(n9951), .A2(n9953), .ZN(n16096) );
  INV_X1 U12135 ( .A(n9825), .ZN(n9952) );
  NAND2_X1 U12136 ( .A1(n9953), .A2(n9971), .ZN(n16094) );
  AND2_X1 U12137 ( .A1(n10216), .A2(n19115), .ZN(n10013) );
  OAI21_X1 U12138 ( .B1(n10908), .B2(n18928), .A(n10898), .ZN(n13148) );
  OAI211_X1 U12139 ( .C1(n10899), .C2(n10893), .A(n10905), .B(n10895), .ZN(
        n13147) );
  AND2_X1 U12140 ( .A1(n10230), .A2(n10233), .ZN(n10234) );
  AND2_X1 U12141 ( .A1(n9982), .A2(n10219), .ZN(n10220) );
  XNOR2_X1 U12142 ( .A(n13212), .B(n13213), .ZN(n13235) );
  INV_X1 U12143 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15462) );
  INV_X1 U12144 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10090) );
  AND3_X1 U12145 ( .A1(n10864), .A2(n10863), .A3(n10862), .ZN(n15461) );
  NAND2_X1 U12146 ( .A1(n10587), .A2(n10547), .ZN(n16187) );
  NAND2_X1 U12147 ( .A1(n9776), .A2(n10572), .ZN(n10547) );
  INV_X1 U12148 ( .A(n10345), .ZN(n19090) );
  NAND2_X1 U12149 ( .A1(n10288), .A2(n10286), .ZN(n19254) );
  INV_X1 U12150 ( .A(n19120), .ZN(n19123) );
  INV_X1 U12151 ( .A(n19119), .ZN(n19121) );
  NOR2_X2 U12152 ( .A1(n13913), .A2(n16077), .ZN(n19120) );
  NOR2_X2 U12153 ( .A1(n13917), .A2(n16077), .ZN(n19119) );
  INV_X1 U12154 ( .A(n13725), .ZN(n19084) );
  AND2_X1 U12155 ( .A1(n19407), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13303) );
  NOR2_X1 U12156 ( .A1(n10572), .A2(n10571), .ZN(n16183) );
  AND2_X1 U12157 ( .A1(n10570), .A2(n10569), .ZN(n10571) );
  NOR2_X1 U12158 ( .A1(n15519), .A2(n12473), .ZN(n18518) );
  AOI21_X1 U12159 ( .B1(n12484), .B2(n12656), .A(n12655), .ZN(n18519) );
  NAND2_X1 U12160 ( .A1(n16862), .A2(P3_EBX_REG_25__SCAN_IN), .ZN(n16851) );
  NAND2_X1 U12161 ( .A1(n16945), .A2(P3_EBX_REG_18__SCAN_IN), .ZN(n16909) );
  NAND3_X1 U12162 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16985), .A3(n15503), 
        .ZN(n16944) );
  NAND3_X1 U12163 ( .A1(n12433), .A2(n12432), .A3(n12431), .ZN(n17098) );
  OAI211_X1 U12164 ( .C1(n12553), .C2(n12552), .A(n12551), .B(n9793), .ZN(
        n12554) );
  NOR2_X1 U12165 ( .A1(n15510), .A2(n15509), .ZN(n17247) );
  NAND2_X1 U12166 ( .A1(n17724), .A2(n17215), .ZN(n17600) );
  AND2_X1 U12167 ( .A1(n9916), .A2(n9917), .ZN(n15534) );
  NOR2_X1 U12168 ( .A1(n12651), .A2(n12649), .ZN(n16253) );
  INV_X1 U12169 ( .A(n16241), .ZN(n16256) );
  NAND2_X1 U12170 ( .A1(n17428), .A2(n12619), .ZN(n17417) );
  NAND2_X1 U12171 ( .A1(n12618), .A2(n10057), .ZN(n12619) );
  NAND2_X1 U12172 ( .A1(n12620), .A2(n17777), .ZN(n12618) );
  NOR3_X1 U12173 ( .A1(n17596), .A2(n9920), .A3(n9921), .ZN(n9919) );
  INV_X1 U12174 ( .A(n17878), .ZN(n9920) );
  INV_X1 U12175 ( .A(n18037), .ZN(n18515) );
  NAND2_X1 U12176 ( .A1(n17558), .A2(n9922), .ZN(n9921) );
  NOR2_X1 U12177 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n9922) );
  NAND2_X1 U12178 ( .A1(n12614), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17566) );
  NAND2_X1 U12179 ( .A1(n17651), .A2(n9787), .ZN(n12614) );
  NOR2_X1 U12180 ( .A1(n12640), .A2(n12466), .ZN(n18529) );
  AND3_X1 U12181 ( .A1(n17651), .A2(n9796), .A3(n9928), .ZN(n17608) );
  NOR2_X1 U12182 ( .A1(n17638), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9928) );
  INV_X1 U12183 ( .A(n17908), .ZN(n17935) );
  INV_X1 U12184 ( .A(n18545), .ZN(n17866) );
  INV_X1 U12185 ( .A(n17933), .ZN(n17909) );
  INV_X1 U12186 ( .A(n17566), .ZN(n17559) );
  OR2_X1 U12187 ( .A1(n17688), .A2(n12603), .ZN(n12606) );
  NOR2_X1 U12188 ( .A1(n18746), .A2(n15516), .ZN(n18545) );
  INV_X1 U12189 ( .A(n12640), .ZN(n18094) );
  NOR2_X1 U12190 ( .A1(n12423), .A2(n12422), .ZN(n18109) );
  INV_X1 U12191 ( .A(n18426), .ZN(n18189) );
  INV_X1 U12192 ( .A(n14495), .ZN(n13033) );
  AND2_X1 U12193 ( .A1(n19773), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19858) );
  AND2_X1 U12194 ( .A1(n19773), .A2(n13645), .ZN(n19865) );
  AND2_X1 U12195 ( .A1(n14494), .A2(n14477), .ZN(n14878) );
  NAND2_X1 U12196 ( .A1(n13245), .A2(n13244), .ZN(n13247) );
  XNOR2_X1 U12197 ( .A(n11663), .B(n13398), .ZN(n13245) );
  NAND2_X1 U12198 ( .A1(n12902), .A2(n13183), .ZN(n15717) );
  OR2_X1 U12199 ( .A1(n13287), .A2(n12901), .ZN(n12902) );
  INV_X1 U12200 ( .A(n15726), .ZN(n14747) );
  INV_X1 U12201 ( .A(n15725), .ZN(n14744) );
  AND2_X1 U12202 ( .A1(n13186), .A2(n13185), .ZN(n19897) );
  INV_X2 U12203 ( .A(n19888), .ZN(n19896) );
  OR2_X1 U12204 ( .A1(n12836), .A2(n12837), .ZN(n12838) );
  AND2_X1 U12205 ( .A1(n14613), .A2(n14621), .ZN(n15730) );
  INV_X1 U12206 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14841) );
  NOR2_X1 U12207 ( .A1(n14653), .A2(n14652), .ZN(n15745) );
  AND2_X1 U12208 ( .A1(n14651), .A2(n14650), .ZN(n14652) );
  INV_X1 U12209 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14177) );
  AOI21_X1 U12210 ( .B1(n14680), .B2(n14679), .A(n14678), .ZN(n15761) );
  INV_X1 U12211 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20835) );
  AND2_X1 U12212 ( .A1(n15795), .A2(n19935), .ZN(n15791) );
  INV_X1 U12213 ( .A(n15795), .ZN(n19936) );
  INV_X1 U12214 ( .A(n12940), .ZN(n19975) );
  AND2_X1 U12215 ( .A1(n13290), .A2(n12835), .ZN(n19938) );
  NAND2_X1 U12216 ( .A1(n10037), .A2(n10036), .ZN(n12939) );
  NAND2_X1 U12217 ( .A1(n12936), .A2(n10038), .ZN(n10037) );
  AND2_X1 U12218 ( .A1(n11803), .A2(n15882), .ZN(n15591) );
  INV_X1 U12219 ( .A(n19939), .ZN(n15908) );
  NAND2_X1 U12220 ( .A1(n10032), .A2(n15782), .ZN(n15775) );
  NAND2_X1 U12221 ( .A1(n11795), .A2(n13273), .ZN(n15865) );
  AND2_X1 U12222 ( .A1(n11795), .A2(n11761), .ZN(n19964) );
  AND2_X1 U12223 ( .A1(n11795), .A2(n11652), .ZN(n19965) );
  INV_X1 U12224 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19973) );
  OAI21_X1 U12225 ( .B1(n13567), .B2(n15947), .A(n20135), .ZN(n20747) );
  CLKBUF_X1 U12226 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n20732) );
  INV_X1 U12227 ( .A(n15582), .ZN(n20726) );
  CLKBUF_X1 U12228 ( .A(n12895), .Z(n12896) );
  NOR2_X1 U12229 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14983) );
  OAI211_X1 U12230 ( .C1(n10066), .C2(n20446), .A(n20364), .B(n19984), .ZN(
        n20019) );
  OR2_X1 U12231 ( .A1(n20092), .A2(n20049), .ZN(n20120) );
  OAI21_X1 U12232 ( .B1(n20138), .B2(n20137), .A(n20522), .ZN(n20163) );
  OAI22_X1 U12233 ( .A1(n20214), .A2(n20213), .B1(n20212), .B2(n20447), .ZN(
        n20238) );
  OAI211_X1 U12234 ( .C1(n20293), .C2(n20446), .A(n20364), .B(n20292), .ZN(
        n20318) );
  INV_X1 U12235 ( .A(n20469), .ZN(n20440) );
  OAI211_X1 U12236 ( .C1(n10081), .C2(n20446), .A(n20522), .B(n20445), .ZN(
        n20466) );
  NOR2_X1 U12237 ( .A1(n19985), .A2(n20135), .ZN(n20514) );
  NOR2_X1 U12238 ( .A1(n19997), .A2(n20135), .ZN(n20535) );
  NOR2_X1 U12239 ( .A1(n20000), .A2(n20135), .ZN(n20541) );
  NOR2_X1 U12240 ( .A1(n20007), .A2(n20135), .ZN(n20553) );
  NOR2_X1 U12241 ( .A1(n20010), .A2(n20135), .ZN(n20559) );
  INV_X1 U12242 ( .A(n20524), .ZN(n20570) );
  NOR2_X1 U12243 ( .A1(n20017), .A2(n20135), .ZN(n20566) );
  INV_X1 U12244 ( .A(n20514), .ZN(n20584) );
  INV_X1 U12245 ( .A(n20529), .ZN(n20596) );
  INV_X1 U12246 ( .A(n20535), .ZN(n20603) );
  INV_X1 U12247 ( .A(n20547), .ZN(n20617) );
  INV_X1 U12248 ( .A(n20553), .ZN(n20624) );
  INV_X1 U12249 ( .A(n20559), .ZN(n20631) );
  INV_X1 U12250 ( .A(n20566), .ZN(n20638) );
  NOR2_X1 U12251 ( .A1(n20446), .A2(n13280), .ZN(n15582) );
  INV_X1 U12252 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20957) );
  INV_X1 U12253 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20446) );
  AND2_X1 U12254 ( .A1(n9729), .A2(n12997), .ZN(n18753) );
  NOR2_X1 U12255 ( .A1(n15000), .A2(n18896), .ZN(n12778) );
  OAI21_X1 U12256 ( .B1(n15006), .B2(n9859), .A(n9858), .ZN(n15000) );
  NAND2_X1 U12257 ( .A1(n9860), .A2(n15194), .ZN(n9859) );
  NAND2_X1 U12258 ( .A1(n18896), .A2(n9860), .ZN(n9858) );
  INV_X1 U12259 ( .A(n15001), .ZN(n9860) );
  NOR2_X1 U12260 ( .A1(n15006), .A2(n15007), .ZN(n15005) );
  NOR2_X1 U12261 ( .A1(n18896), .A2(n15043), .ZN(n15950) );
  NOR2_X1 U12262 ( .A1(n15546), .A2(n12777), .ZN(n12970) );
  NAND2_X1 U12263 ( .A1(n18870), .A2(n9798), .ZN(n15538) );
  AND2_X1 U12264 ( .A1(n15538), .A2(n16010), .ZN(n15546) );
  INV_X1 U12265 ( .A(n18923), .ZN(n18921) );
  INV_X1 U12266 ( .A(n18929), .ZN(n18912) );
  OR4_X1 U12267 ( .A1(n19044), .A2(n18917), .A3(n18753), .A4(n16210), .ZN(
        n18929) );
  AND2_X1 U12268 ( .A1(n18753), .A2(n16206), .ZN(n18923) );
  INV_X1 U12269 ( .A(n18900), .ZN(n18933) );
  INV_X1 U12270 ( .A(n18956), .ZN(n13613) );
  OR2_X1 U12271 ( .A1(n10949), .A2(n10948), .ZN(n13518) );
  AND2_X1 U12272 ( .A1(n9782), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n9956)
         );
  INV_X1 U12273 ( .A(n18951), .ZN(n18966) );
  CLKBUF_X1 U12274 ( .A(n13302), .Z(n16148) );
  INV_X1 U12275 ( .A(n19702), .ZN(n19698) );
  NAND2_X1 U12276 ( .A1(n18965), .A2(n10203), .ZN(n18951) );
  OR2_X1 U12277 ( .A1(n18995), .A2(n13915), .ZN(n15169) );
  OR2_X1 U12278 ( .A1(n18995), .A2(n10203), .ZN(n15994) );
  INV_X1 U12279 ( .A(n15169), .ZN(n18974) );
  AND2_X1 U12280 ( .A1(n18998), .A2(n15994), .ZN(n19004) );
  INV_X1 U12281 ( .A(n13632), .ZN(n18997) );
  INV_X1 U12282 ( .A(n15994), .ZN(n18980) );
  INV_X2 U12283 ( .A(n19016), .ZN(n19040) );
  OR2_X1 U12284 ( .A1(n13037), .A2(n13012), .ZN(n13133) );
  NOR2_X1 U12285 ( .A1(n15337), .A2(n15363), .ZN(n9955) );
  INV_X1 U12286 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16101) );
  INV_X1 U12287 ( .A(n16084), .ZN(n19056) );
  OAI21_X1 U12288 ( .B1(n14467), .B2(n16161), .A(n14466), .ZN(n14468) );
  NOR2_X1 U12289 ( .A1(n14460), .A2(n14465), .ZN(n14466) );
  NAND2_X1 U12290 ( .A1(n15272), .A2(n9837), .ZN(n15191) );
  NAND2_X1 U12291 ( .A1(n15187), .A2(n9838), .ZN(n9837) );
  NOR2_X1 U12292 ( .A1(n15213), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14229) );
  NAND2_X1 U12293 ( .A1(n9890), .A2(n15354), .ZN(n15243) );
  OR2_X1 U12294 ( .A1(n15356), .A2(n12327), .ZN(n9890) );
  AND2_X1 U12295 ( .A1(n16102), .A2(n10884), .ZN(n15364) );
  AND2_X1 U12296 ( .A1(n10868), .A2(n19070), .ZN(n13171) );
  NAND2_X1 U12297 ( .A1(n15454), .A2(n13008), .ZN(n19710) );
  INV_X1 U12298 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19696) );
  AOI221_X1 U12299 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16219), .C1(n19718), .C2(
        n16219), .A(n19545), .ZN(n19713) );
  INV_X1 U12300 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16204) );
  NAND2_X1 U12301 ( .A1(n13224), .A2(n13301), .ZN(n15488) );
  AND2_X1 U12302 ( .A1(n16187), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16214) );
  INV_X1 U12303 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16201) );
  INV_X1 U12304 ( .A(n19211), .ZN(n19201) );
  AND2_X1 U12305 ( .A1(n19219), .A2(n19218), .ZN(n19236) );
  INV_X1 U12306 ( .A(n19236), .ZN(n19247) );
  OAI21_X1 U12307 ( .B1(n19224), .B2(n19223), .A(n19222), .ZN(n19246) );
  AND2_X1 U12308 ( .A1(n19282), .A2(n19285), .ZN(n19290) );
  AOI21_X1 U12309 ( .B1(n19732), .B2(n19287), .A(n19286), .ZN(n19304) );
  INV_X1 U12310 ( .A(n19357), .ZN(n19347) );
  OR2_X1 U12311 ( .A1(n19440), .A2(n19132), .ZN(n19369) );
  INV_X1 U12312 ( .A(n19369), .ZN(n19370) );
  OAI21_X1 U12313 ( .B1(n19383), .B2(n19398), .A(n19545), .ZN(n19401) );
  INV_X1 U12314 ( .A(n19375), .ZN(n19400) );
  NOR2_X1 U12315 ( .A1(n19440), .A2(n19404), .ZN(n19427) );
  INV_X1 U12316 ( .A(n19561), .ZN(n19455) );
  OAI21_X1 U12317 ( .B1(n19468), .B2(n19546), .A(n19450), .ZN(n19471) );
  OAI22_X1 U12318 ( .A1(n19124), .A2(n19123), .B1(n19122), .B2(n19121), .ZN(
        n19502) );
  INV_X1 U12319 ( .A(n19555), .ZN(n19512) );
  OAI22_X1 U12320 ( .A1(n19114), .A2(n19123), .B1(n21048), .B2(n19121), .ZN(
        n19524) );
  OR2_X1 U12321 ( .A1(n19405), .A2(n19439), .ZN(n19535) );
  INV_X1 U12322 ( .A(n19488), .ZN(n19552) );
  OR2_X1 U12323 ( .A1(n19405), .A2(n19084), .ZN(n19577) );
  INV_X1 U12324 ( .A(n19593), .ZN(n19574) );
  INV_X1 U12325 ( .A(n19467), .ZN(n19580) );
  INV_X1 U12326 ( .A(n19524), .ZN(n19583) );
  INV_X1 U12327 ( .A(n19577), .ZN(n19589) );
  NOR2_X1 U12328 ( .A1(n9823), .A2(n19538), .ZN(n19587) );
  INV_X1 U12329 ( .A(n19502), .ZN(n19594) );
  AND2_X1 U12330 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10592), .ZN(n19731) );
  NOR2_X1 U12331 ( .A1(n15609), .A2(n14108), .ZN(n18746) );
  INV_X1 U12332 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18732) );
  NAND2_X1 U12333 ( .A1(n9850), .A2(n18726), .ZN(n16359) );
  INV_X1 U12334 ( .A(n18524), .ZN(n9850) );
  INV_X1 U12335 ( .A(n16733), .ZN(n16720) );
  INV_X1 U12336 ( .A(n16692), .ZN(n16721) );
  NOR2_X2 U12337 ( .A1(n18573), .A2(n12492), .ZN(n16723) );
  NAND4_X1 U12338 ( .A1(n17892), .A2(n16677), .A3(n18588), .A4(n18577), .ZN(
        n16733) );
  AND2_X1 U12339 ( .A1(n16868), .A2(P3_EBX_REG_24__SCAN_IN), .ZN(n16862) );
  NOR2_X1 U12340 ( .A1(n16837), .A2(n16882), .ZN(n16863) );
  AND2_X1 U12341 ( .A1(n16863), .A2(P3_EBX_REG_23__SCAN_IN), .ZN(n16868) );
  NAND2_X1 U12342 ( .A1(n16921), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n16907) );
  NOR2_X1 U12343 ( .A1(n16909), .A2(n20935), .ZN(n16921) );
  NOR2_X1 U12344 ( .A1(n16944), .A2(n16527), .ZN(n16945) );
  INV_X1 U12345 ( .A(n16997), .ZN(n16985) );
  NAND2_X1 U12346 ( .A1(n16998), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n16997) );
  NAND2_X1 U12347 ( .A1(n9792), .A2(P3_EBX_REG_9__SCAN_IN), .ZN(n17040) );
  NAND2_X1 U12348 ( .A1(n17070), .A2(n9829), .ZN(n17063) );
  NOR2_X1 U12349 ( .A1(n17085), .A2(n17074), .ZN(n17070) );
  NOR2_X2 U12350 ( .A1(n17258), .A2(n17125), .ZN(n17120) );
  NOR2_X1 U12351 ( .A1(n17269), .A2(n17159), .ZN(n17154) );
  NOR2_X2 U12352 ( .A1(n17101), .A2(n17234), .ZN(n17170) );
  INV_X1 U12353 ( .A(n17145), .ZN(n17169) );
  AOI211_X1 U12354 ( .C1(n12590), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n12379), .B(n12378), .ZN(n12380) );
  NOR2_X1 U12355 ( .A1(n12518), .A2(n12517), .ZN(n17222) );
  AND2_X1 U12356 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17233), .ZN(n17228) );
  INV_X1 U12357 ( .A(n17243), .ZN(n17234) );
  NOR2_X1 U12358 ( .A1(n17304), .A2(n17182), .ZN(n17240) );
  NOR2_X1 U12359 ( .A1(n17097), .A2(n17096), .ZN(n17243) );
  INV_X1 U12360 ( .A(n17239), .ZN(n17241) );
  NOR2_X1 U12361 ( .A1(n17354), .A2(n18090), .ZN(n17355) );
  NOR2_X1 U12362 ( .A1(n17881), .A2(n16225), .ZN(n16257) );
  NAND2_X1 U12363 ( .A1(n17397), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17386) );
  AND2_X1 U12364 ( .A1(n17516), .A2(n9844), .ZN(n17397) );
  NOR2_X1 U12365 ( .A1(n17759), .A2(n17364), .ZN(n9844) );
  NOR2_X1 U12366 ( .A1(n17598), .A2(n16223), .ZN(n17516) );
  INV_X1 U12367 ( .A(n17516), .ZN(n17536) );
  INV_X1 U12368 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17553) );
  INV_X1 U12369 ( .A(n17600), .ZN(n17640) );
  BUF_X1 U12370 ( .A(n16237), .Z(n18460) );
  NOR2_X1 U12371 ( .A1(n16359), .A2(n18090), .ZN(n17724) );
  NAND2_X1 U12372 ( .A1(n17508), .A2(n17583), .ZN(n17723) );
  OAI21_X1 U12373 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18725), .A(n16359), 
        .ZN(n17731) );
  XNOR2_X1 U12374 ( .A(n17380), .B(n17638), .ZN(n17750) );
  AND2_X1 U12375 ( .A1(n9852), .A2(n9851), .ZN(n17941) );
  NAND2_X1 U12376 ( .A1(n12700), .A2(n18529), .ZN(n9851) );
  INV_X1 U12377 ( .A(n18528), .ZN(n9852) );
  NAND2_X1 U12378 ( .A1(n17866), .A2(n18549), .ZN(n17948) );
  NOR2_X1 U12379 ( .A1(n17559), .A2(n12710), .ZN(n17981) );
  AND2_X1 U12380 ( .A1(n17651), .A2(n9796), .ZN(n12710) );
  INV_X1 U12381 ( .A(n17964), .ZN(n17979) );
  CLKBUF_X1 U12382 ( .A(n18044), .Z(n17892) );
  INV_X1 U12383 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18560) );
  INV_X1 U12384 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18087) );
  INV_X1 U12385 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20853) );
  OR2_X1 U12386 ( .A1(n16350), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18740) );
  AND2_X1 U12387 ( .A1(n12913), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n19976)
         );
  NAND2_X1 U12389 ( .A1(n14500), .A2(n19821), .ZN(n9999) );
  OAI22_X1 U12390 ( .A1(n14516), .A2(n14684), .B1(n12316), .B2(n14682), .ZN(
        n12317) );
  OAI21_X1 U12391 ( .B1(n11087), .B2(n16084), .A(n11086), .ZN(n11088) );
  AOI21_X1 U12392 ( .B1(n15111), .B2(n19063), .A(n11085), .ZN(n11086) );
  OAI21_X1 U12393 ( .B1(n12743), .B2(n16084), .A(n12742), .ZN(n12744) );
  OAI21_X1 U12394 ( .B1(n12947), .B2(n16083), .A(n9966), .ZN(P2_U2996) );
  INV_X1 U12395 ( .A(n12953), .ZN(n9966) );
  AOI21_X1 U12396 ( .B1(n15182), .B2(n16153), .A(n12933), .ZN(n12934) );
  OAI211_X1 U12397 ( .C1(n15258), .C2(n16163), .A(n9935), .B(n9930), .ZN(
        P2_U3017) );
  INV_X1 U12398 ( .A(n15254), .ZN(n9935) );
  OAI21_X1 U12399 ( .B1(n12743), .B2(n16163), .A(n9895), .ZN(P2_U3027) );
  OAI21_X1 U12400 ( .B1(n12952), .B2(n16163), .A(n12345), .ZN(n12346) );
  NOR2_X1 U12401 ( .A1(n12344), .A2(n10072), .ZN(n12345) );
  AOI211_X1 U12402 ( .C1(n16381), .C2(n16713), .A(n16380), .B(n16379), .ZN(
        n16384) );
  INV_X1 U12403 ( .A(n16998), .ZN(n17010) );
  OAI211_X1 U12404 ( .C1(n12885), .C2(n18055), .A(n12716), .B(n12715), .ZN(
        n12717) );
  NAND2_X2 U12405 ( .A1(n10136), .A2(n10135), .ZN(n10193) );
  AND2_X1 U12406 ( .A1(n10216), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9776) );
  AND2_X1 U12407 ( .A1(n9869), .A2(n9867), .ZN(n9777) );
  AND2_X1 U12408 ( .A1(n9965), .A2(n9963), .ZN(n9778) );
  NAND2_X1 U12409 ( .A1(n13542), .A2(n13544), .ZN(n13543) );
  AND4_X1 U12410 ( .A1(n10294), .A2(n10293), .A3(n10292), .A4(n10291), .ZN(
        n9779) );
  AND4_X1 U12411 ( .A1(n9812), .A2(n10162), .A3(n10150), .A4(n10161), .ZN(
        n9780) );
  AND2_X2 U12412 ( .A1(n9733), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10367) );
  AND2_X2 U12413 ( .A1(n14277), .A2(n10305), .ZN(n10360) );
  NOR2_X1 U12414 ( .A1(n12369), .A2(n18539), .ZN(n12530) );
  AND4_X1 U12415 ( .A1(n12534), .A2(n12533), .A3(n12532), .A4(n12531), .ZN(
        n9781) );
  AND2_X1 U12416 ( .A1(n14557), .A2(n10007), .ZN(n12836) );
  NAND2_X1 U12417 ( .A1(n14630), .A2(n10006), .ZN(n14613) );
  NAND2_X1 U12418 ( .A1(n9869), .A2(n9870), .ZN(n12762) );
  NAND2_X1 U12419 ( .A1(n9965), .A2(n13614), .ZN(n13731) );
  AND2_X1 U12420 ( .A1(n13542), .A2(n9939), .ZN(n13628) );
  AND2_X1 U12421 ( .A1(n14091), .A2(n9826), .ZN(n11065) );
  XNOR2_X1 U12422 ( .A(n14499), .B(n14498), .ZN(n14867) );
  AND2_X1 U12423 ( .A1(n13698), .A2(n9831), .ZN(n9782) );
  AND2_X1 U12424 ( .A1(n9841), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9783) );
  NAND2_X1 U12425 ( .A1(n9872), .A2(n9874), .ZN(n12759) );
  OR2_X1 U12426 ( .A1(n13228), .A2(n9947), .ZN(n13239) );
  INV_X1 U12427 ( .A(n9925), .ZN(n13694) );
  AND2_X1 U12428 ( .A1(n9861), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9784) );
  CLKBUF_X1 U12429 ( .A(n9733), .Z(n14313) );
  AND2_X1 U12430 ( .A1(n9864), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9785) );
  INV_X1 U12431 ( .A(n10254), .ZN(n14132) );
  NAND3_X4 U12432 ( .A1(n9814), .A2(n9981), .A3(n9982), .ZN(n10254) );
  OR2_X1 U12433 ( .A1(n18539), .A2(n12371), .ZN(n9786) );
  NAND2_X1 U12434 ( .A1(n13007), .A2(n9763), .ZN(n10899) );
  OR2_X1 U12435 ( .A1(n12613), .A2(n12612), .ZN(n9787) );
  OR2_X1 U12436 ( .A1(n13256), .A2(n13643), .ZN(n11654) );
  NAND2_X1 U12437 ( .A1(n9986), .A2(n10646), .ZN(n15415) );
  AND2_X1 U12438 ( .A1(n9769), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10382) );
  AND2_X1 U12440 ( .A1(n9727), .A2(n9961), .ZN(n15423) );
  AND2_X1 U12441 ( .A1(n14630), .A2(n10004), .ZN(n14604) );
  NAND2_X1 U12442 ( .A1(n14557), .A2(n10009), .ZN(n14517) );
  AND2_X1 U12443 ( .A1(n14557), .A2(n10010), .ZN(n14532) );
  NAND2_X1 U12444 ( .A1(n14630), .A2(n14631), .ZN(n14619) );
  NOR2_X1 U12445 ( .A1(n12764), .A2(n16101), .ZN(n12763) );
  AND4_X1 U12446 ( .A1(n11300), .A2(n9992), .A3(n11299), .A4(n11780), .ZN(
        n9789) );
  AND4_X1 U12447 ( .A1(n11173), .A2(n11172), .A3(n11171), .A4(n11170), .ZN(
        n9790) );
  AND4_X1 U12448 ( .A1(n12539), .A2(n12538), .A3(n12537), .A4(n12536), .ZN(
        n9791) );
  AND4_X1 U12449 ( .A1(n12550), .A2(n12549), .A3(n12548), .A4(n12547), .ZN(
        n9793) );
  OR2_X1 U12450 ( .A1(n12616), .A2(n12615), .ZN(n9794) );
  AND3_X1 U12451 ( .A1(n19115), .A2(n9780), .A3(n10216), .ZN(n9795) );
  NAND2_X1 U12452 ( .A1(n10272), .A2(n10271), .ZN(n10270) );
  NAND2_X1 U12453 ( .A1(n13966), .A2(n13967), .ZN(n14024) );
  AND2_X1 U12454 ( .A1(n9787), .A2(n9929), .ZN(n9796) );
  NAND2_X1 U12455 ( .A1(n9972), .A2(n15299), .ZN(n11095) );
  INV_X1 U12456 ( .A(n10177), .ZN(n16207) );
  NAND2_X1 U12457 ( .A1(n11555), .A2(n14828), .ZN(n14817) );
  AND4_X1 U12458 ( .A1(n10284), .A2(n10283), .A3(n10282), .A4(n10281), .ZN(
        n9797) );
  OR2_X1 U12459 ( .A1(n18785), .A2(n18784), .ZN(n9798) );
  OR2_X1 U12460 ( .A1(n12736), .A2(n19074), .ZN(n9799) );
  AND2_X1 U12461 ( .A1(n9773), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n9800) );
  INV_X1 U12462 ( .A(n11093), .ZN(n9975) );
  OR2_X1 U12463 ( .A1(n15180), .A2(n18900), .ZN(n9801) );
  OR2_X1 U12464 ( .A1(n11550), .A2(n14833), .ZN(n9803) );
  AND2_X1 U12465 ( .A1(n9795), .A2(n10176), .ZN(n9804) );
  AND2_X1 U12466 ( .A1(n14025), .A2(n10642), .ZN(n9805) );
  AND4_X1 U12467 ( .A1(n10426), .A2(n10429), .A3(n10428), .A4(n10437), .ZN(
        n9806) );
  NAND2_X1 U12468 ( .A1(n9727), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15437) );
  AND2_X1 U12469 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n9807) );
  AND2_X1 U12470 ( .A1(n10288), .A2(n10289), .ZN(n10314) );
  OR2_X1 U12471 ( .A1(n10016), .A2(n10014), .ZN(n9808) );
  AND2_X1 U12472 ( .A1(n14191), .A2(n9941), .ZN(n14993) );
  OAI21_X1 U12473 ( .B1(n15242), .B2(n9892), .A(n12329), .ZN(n9891) );
  AND2_X1 U12474 ( .A1(n15008), .A2(n12869), .ZN(n12823) );
  OR2_X1 U12475 ( .A1(n15251), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9809) );
  NOR2_X1 U12476 ( .A1(n15091), .A2(n15090), .ZN(n15089) );
  NOR2_X1 U12477 ( .A1(n15005), .A2(n18896), .ZN(n9811) );
  INV_X1 U12478 ( .A(n9889), .ZN(n9888) );
  NAND2_X1 U12479 ( .A1(n9985), .A2(n15396), .ZN(n9889) );
  AND2_X1 U12480 ( .A1(n10149), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9812) );
  OR2_X1 U12481 ( .A1(n12858), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9813) );
  INV_X1 U12482 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18540) );
  INV_X1 U12483 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18697) );
  NAND2_X1 U12484 ( .A1(n9795), .A2(n9882), .ZN(n9814) );
  AND2_X2 U12485 ( .A1(n11157), .A2(n10031), .ZN(n11336) );
  INV_X1 U12486 ( .A(n10908), .ZN(n14144) );
  NAND2_X1 U12487 ( .A1(n10040), .A2(n11425), .ZN(n13262) );
  AND2_X1 U12488 ( .A1(n13649), .A2(n13646), .ZN(n19863) );
  NOR2_X1 U12489 ( .A1(n12768), .A2(n9873), .ZN(n12760) );
  NOR2_X1 U12490 ( .A1(n12767), .A2(n10781), .ZN(n12761) );
  NAND2_X1 U12491 ( .A1(n14084), .A2(n10022), .ZN(n10025) );
  INV_X1 U12492 ( .A(n10689), .ZN(n11100) );
  NOR2_X1 U12493 ( .A1(n13802), .A2(n10029), .ZN(n13732) );
  AND2_X1 U12494 ( .A1(n11241), .A2(n11269), .ZN(n13079) );
  NOR2_X1 U12495 ( .A1(n12755), .A2(n15233), .ZN(n12756) );
  OAI21_X1 U12496 ( .B1(n13846), .B2(n11544), .A(n11543), .ZN(n14005) );
  AND2_X1 U12497 ( .A1(n14674), .A2(n14673), .ZN(n14172) );
  AND2_X1 U12498 ( .A1(n12721), .A2(n14206), .ZN(n9815) );
  NAND2_X1 U12499 ( .A1(n10270), .A2(n10273), .ZN(n13216) );
  INV_X1 U12500 ( .A(n9761), .ZN(n13226) );
  NOR2_X1 U12501 ( .A1(n12776), .A2(n12973), .ZN(n11121) );
  AND2_X1 U12502 ( .A1(n10818), .A2(n10021), .ZN(n9816) );
  OR2_X1 U12503 ( .A1(n11412), .A2(n11432), .ZN(n9817) );
  INV_X1 U12504 ( .A(n14654), .ZN(n9900) );
  AND2_X1 U12505 ( .A1(n11718), .A2(n11717), .ZN(n14654) );
  NAND2_X1 U12506 ( .A1(n10798), .A2(n10797), .ZN(n13802) );
  NAND2_X1 U12507 ( .A1(n14191), .A2(n11138), .ZN(n12788) );
  OR3_X1 U12508 ( .A1(n17596), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n9818) );
  INV_X1 U12509 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19727) );
  AND2_X1 U12510 ( .A1(n14096), .A2(n14085), .ZN(n14084) );
  OR2_X1 U12511 ( .A1(n15766), .A2(n14888), .ZN(n9819) );
  AND2_X1 U12512 ( .A1(n12773), .A2(n9861), .ZN(n9820) );
  AND2_X1 U12513 ( .A1(n11565), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9821) );
  NOR2_X1 U12514 ( .A1(n20736), .A2(n19982), .ZN(n9822) );
  INV_X1 U12515 ( .A(n19072), .ZN(n16143) );
  NAND2_X1 U12516 ( .A1(n13337), .A2(n13698), .ZN(n13345) );
  INV_X1 U12517 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9871) );
  NOR3_X1 U12518 ( .A1(n19536), .A2(n19585), .A3(n19732), .ZN(n9823) );
  OAI22_X2 U12519 ( .A1(n19727), .A2(n14139), .B1(n14244), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n18870) );
  NAND2_X1 U12520 ( .A1(n13337), .A2(n9782), .ZN(n13423) );
  NOR2_X1 U12521 ( .A1(n12985), .A2(n13806), .ZN(n13542) );
  AND2_X1 U12522 ( .A1(n13542), .A2(n9936), .ZN(n13851) );
  NOR2_X1 U12523 ( .A1(n13406), .A2(n10016), .ZN(n13514) );
  NOR2_X1 U12524 ( .A1(n13406), .A2(n9808), .ZN(n12988) );
  NOR2_X1 U12525 ( .A1(n13228), .A2(n13229), .ZN(n13230) );
  NAND2_X1 U12526 ( .A1(n13542), .A2(n9938), .ZN(n13629) );
  NOR2_X1 U12527 ( .A1(n13228), .A2(n9946), .ZN(n12983) );
  AND2_X1 U12528 ( .A1(n10024), .A2(n15305), .ZN(n9824) );
  NOR2_X1 U12529 ( .A1(n13338), .A2(n13347), .ZN(n13348) );
  XOR2_X1 U12530 ( .A(n10404), .B(n10262), .Z(n9825) );
  AND2_X1 U12531 ( .A1(n14038), .A2(n14090), .ZN(n9826) );
  AND2_X1 U12532 ( .A1(n13520), .A2(n13519), .ZN(n13536) );
  NAND2_X1 U12533 ( .A1(n14172), .A2(n14173), .ZN(n14171) );
  OR2_X1 U12534 ( .A1(n13587), .A2(n13693), .ZN(n9925) );
  AND2_X1 U12535 ( .A1(n9901), .A2(n14519), .ZN(n9827) );
  AND2_X1 U12536 ( .A1(n9826), .A2(n11064), .ZN(n9828) );
  AND2_X1 U12537 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .ZN(n9829) );
  OR2_X1 U12538 ( .A1(n11043), .A2(n11042), .ZN(n13868) );
  AND2_X1 U12539 ( .A1(n12752), .A2(n9864), .ZN(n9830) );
  INV_X1 U12540 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9862) );
  INV_X1 U12541 ( .A(n18579), .ZN(n18726) );
  AND2_X1 U12542 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9831) );
  NOR2_X1 U12543 ( .A1(n13388), .A2(n13389), .ZN(n13387) );
  INV_X1 U12544 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n9875) );
  INV_X1 U12545 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n9863) );
  INV_X1 U12546 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9865) );
  AND2_X1 U12547 ( .A1(n15586), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9832) );
  AND2_X1 U12548 ( .A1(n9961), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9833) );
  NAND2_X1 U12549 ( .A1(n15264), .A2(n12852), .ZN(n9834) );
  INV_X1 U12550 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9866) );
  OR2_X1 U12551 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9835) );
  INV_X1 U12552 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9918) );
  INV_X1 U12553 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n9929) );
  INV_X1 U12554 ( .A(n19447), .ZN(n19545) );
  AOI22_X2 U12555 ( .A1(DATAI_18_), .A2(n20016), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20015), .ZN(n20540) );
  AOI22_X2 U12556 ( .A1(DATAI_17_), .A2(n20016), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20015), .ZN(n20534) );
  AOI22_X2 U12557 ( .A1(DATAI_22_), .A2(n20016), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20015), .ZN(n20564) );
  AND2_X1 U12558 ( .A1(n19479), .A2(n19710), .ZN(n19212) );
  NAND2_X1 U12559 ( .A1(n19479), .A2(n18937), .ZN(n19250) );
  INV_X1 U12560 ( .A(n19479), .ZN(n19681) );
  AOI22_X2 U12561 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20015), .B1(DATAI_29_), 
        .B2(n20016), .ZN(n20630) );
  NOR2_X2 U12562 ( .A1(n18305), .A2(n18325), .ZN(n18390) );
  NOR2_X4 U12563 ( .A1(n20959), .A2(n20770), .ZN(n20713) );
  NOR2_X2 U12564 ( .A1(n19125), .A2(n19100), .ZN(n19562) );
  NAND2_X1 U12565 ( .A1(n16220), .A2(n13687), .ZN(n19125) );
  NOR2_X2 U12566 ( .A1(n18540), .A2(n18703), .ZN(n18527) );
  NOR2_X1 U12567 ( .A1(n12445), .A2(n12661), .ZN(n12467) );
  AND2_X2 U12568 ( .A1(n17025), .A2(P3_EBX_REG_11__SCAN_IN), .ZN(n16998) );
  NOR2_X1 U12569 ( .A1(n9977), .A2(n9974), .ZN(n9839) );
  OR2_X2 U12570 ( .A1(n9978), .A2(n9974), .ZN(n9843) );
  NAND2_X1 U12571 ( .A1(n9840), .A2(n15210), .ZN(n11102) );
  NAND3_X1 U12572 ( .A1(n9843), .A2(n9842), .A3(n9783), .ZN(n9840) );
  NAND2_X1 U12573 ( .A1(n18540), .A2(n18703), .ZN(n12372) );
  NAND2_X1 U12574 ( .A1(n9879), .A2(n10523), .ZN(n9845) );
  NOR2_X2 U12575 ( .A1(n9880), .A2(n9845), .ZN(n10453) );
  NAND4_X1 U12576 ( .A1(n9847), .A2(n10438), .A3(n9806), .A4(n10427), .ZN(
        n9846) );
  NOR2_X2 U12577 ( .A1(n18728), .A2(n16678), .ZN(n15609) );
  NAND3_X1 U12578 ( .A1(n12391), .A2(n12390), .A3(n9849), .ZN(n9848) );
  INV_X2 U12579 ( .A(n17941), .ZN(n18547) );
  INV_X1 U12580 ( .A(n10259), .ZN(n9876) );
  NOR2_X1 U12581 ( .A1(n9800), .A2(n9877), .ZN(n10259) );
  NAND2_X1 U12582 ( .A1(n9879), .A2(n10313), .ZN(n10397) );
  NAND2_X2 U12583 ( .A1(n9878), .A2(n9879), .ZN(n9971) );
  NAND2_X1 U12584 ( .A1(n13966), .A2(n9887), .ZN(n9886) );
  NAND2_X1 U12585 ( .A1(n14538), .A2(n14519), .ZN(n14521) );
  NAND2_X1 U12586 ( .A1(n14494), .A2(n14495), .ZN(n9902) );
  NAND2_X1 U12587 ( .A1(n9732), .A2(n11664), .ZN(n11668) );
  NAND2_X1 U12588 ( .A1(n9732), .A2(n20872), .ZN(n11723) );
  NAND2_X1 U12589 ( .A1(n9732), .A2(n14625), .ZN(n11736) );
  NAND2_X1 U12590 ( .A1(n9732), .A2(n14602), .ZN(n11747) );
  NAND2_X1 U12591 ( .A1(n9732), .A2(n15707), .ZN(n11699) );
  NAND2_X1 U12592 ( .A1(n9732), .A2(n11708), .ZN(n11711) );
  NAND2_X1 U12593 ( .A1(n9732), .A2(n14658), .ZN(n11718) );
  NAND2_X1 U12594 ( .A1(n9732), .A2(n14610), .ZN(n11741) );
  MUX2_X1 U12595 ( .A(n9732), .B(n11752), .S(P1_EBX_REG_4__SCAN_IN), .Z(n11673) );
  MUX2_X1 U12596 ( .A(n9732), .B(n11752), .S(P1_EBX_REG_6__SCAN_IN), .Z(n11680) );
  MUX2_X1 U12597 ( .A(n9732), .B(n11752), .S(P1_EBX_REG_8__SCAN_IN), .Z(n11688) );
  MUX2_X1 U12598 ( .A(n9732), .B(n11752), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n11702) );
  MUX2_X1 U12599 ( .A(n9732), .B(n11752), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n11727) );
  MUX2_X1 U12600 ( .A(n9732), .B(n11752), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n11753) );
  NAND2_X1 U12601 ( .A1(n11663), .A2(n9914), .ZN(n13388) );
  INV_X1 U12602 ( .A(n9724), .ZN(n9915) );
  NOR2_X1 U12603 ( .A1(n9724), .A2(n10075), .ZN(n9916) );
  NOR2_X1 U12604 ( .A1(n17596), .A2(n9921), .ZN(n17560) );
  NOR2_X1 U12605 ( .A1(n9919), .A2(n17638), .ZN(n17520) );
  NOR2_X1 U12606 ( .A1(n17596), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17565) );
  NAND2_X1 U12607 ( .A1(n13587), .A2(n10931), .ZN(n9923) );
  NAND2_X1 U12608 ( .A1(n9923), .A2(n9924), .ZN(n10936) );
  OR2_X2 U12609 ( .A1(n12596), .A2(n12595), .ZN(n17730) );
  NAND3_X1 U12610 ( .A1(n17651), .A2(n9796), .A3(n17636), .ZN(n17616) );
  NAND3_X1 U12611 ( .A1(n9809), .A2(n9934), .A3(n9932), .ZN(n9931) );
  INV_X1 U12612 ( .A(n10903), .ZN(n9945) );
  OAI21_X1 U12613 ( .B1(n10908), .B2(n19622), .A(n10892), .ZN(n10903) );
  NAND2_X1 U12614 ( .A1(n9756), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n9950) );
  NAND2_X1 U12615 ( .A1(n10397), .A2(n10398), .ZN(n9953) );
  NAND2_X1 U12616 ( .A1(n9954), .A2(n10286), .ZN(n10320) );
  NAND2_X1 U12617 ( .A1(n9954), .A2(n10280), .ZN(n19167) );
  INV_X1 U12618 ( .A(n15335), .ZN(n15365) );
  OAI21_X1 U12619 ( .B1(n15091), .B2(n9958), .A(n9957), .ZN(n14398) );
  NAND2_X1 U12620 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10061) );
  NAND2_X1 U12621 ( .A1(n9969), .A2(n10483), .ZN(n14021) );
  OAI21_X1 U12622 ( .B1(n10479), .B2(n9810), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U12623 ( .A1(n9970), .A2(n10482), .ZN(n13965) );
  NAND2_X1 U12624 ( .A1(n10483), .A2(n10479), .ZN(n9970) );
  INV_X1 U12625 ( .A(n10482), .ZN(n9810) );
  NAND2_X1 U12626 ( .A1(n9971), .A2(n10921), .ZN(n10418) );
  INV_X1 U12627 ( .A(n10717), .ZN(n9977) );
  NAND2_X1 U12628 ( .A1(n9976), .A2(n10736), .ZN(n15298) );
  NOR2_X4 U12629 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15473) );
  NAND2_X1 U12630 ( .A1(n10887), .A2(n10851), .ZN(n10846) );
  NAND3_X1 U12631 ( .A1(n12847), .A2(n9813), .A3(n9989), .ZN(n9987) );
  NAND2_X1 U12632 ( .A1(n12847), .A2(n12846), .ZN(n15186) );
  NOR2_X1 U12633 ( .A1(n12851), .A2(n9990), .ZN(n9989) );
  INV_X1 U12634 ( .A(n12846), .ZN(n9990) );
  INV_X1 U12635 ( .A(n15185), .ZN(n9991) );
  NAND2_X1 U12636 ( .A1(n11368), .A2(n11367), .ZN(n11375) );
  NAND2_X2 U12637 ( .A1(n20090), .A2(n11302), .ZN(n11368) );
  NAND3_X1 U12638 ( .A1(n11368), .A2(n11367), .A3(n10042), .ZN(n10040) );
  NAND2_X1 U12639 ( .A1(n14874), .A2(n19863), .ZN(n9998) );
  NOR2_X1 U12640 ( .A1(n12307), .A2(n12308), .ZN(n12894) );
  NAND3_X1 U12641 ( .A1(n9999), .A2(n14506), .A3(n9998), .ZN(P1_U2809) );
  NAND2_X1 U12642 ( .A1(n14973), .A2(n11919), .ZN(n10000) );
  NAND2_X1 U12643 ( .A1(n10000), .A2(n10001), .ZN(n13415) );
  NAND2_X1 U12644 ( .A1(n10003), .A2(n11937), .ZN(n13412) );
  INV_X1 U12645 ( .A(n13415), .ZN(n10003) );
  NAND2_X1 U12646 ( .A1(n14557), .A2(n14558), .ZN(n14543) );
  NAND2_X1 U12647 ( .A1(n14157), .A2(n10012), .ZN(n14071) );
  INV_X1 U12648 ( .A(n14071), .ZN(n12150) );
  NAND3_X1 U12649 ( .A1(n10176), .A2(n13914), .A3(n10013), .ZN(n10238) );
  NAND3_X1 U12650 ( .A1(n10176), .A2(n13914), .A3(n19115), .ZN(n10177) );
  INV_X1 U12651 ( .A(n13802), .ZN(n10026) );
  NAND2_X1 U12652 ( .A1(n10026), .A2(n10027), .ZN(n13734) );
  NAND2_X1 U12653 ( .A1(n13745), .A2(n10762), .ZN(n13749) );
  NAND2_X1 U12654 ( .A1(n10760), .A2(n10761), .ZN(n13745) );
  AND2_X2 U12655 ( .A1(n10031), .A2(n13270), .ZN(n12213) );
  AND2_X2 U12656 ( .A1(n11150), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10031) );
  NAND3_X1 U12657 ( .A1(n11269), .A2(n11241), .A3(n13256), .ZN(n12895) );
  NAND3_X1 U12658 ( .A1(n10032), .A2(n15782), .A3(n11533), .ZN(n15777) );
  NAND2_X1 U12659 ( .A1(n14784), .A2(n14772), .ZN(n12832) );
  NAND2_X1 U12660 ( .A1(n12832), .A2(n11565), .ZN(n12937) );
  NAND2_X1 U12661 ( .A1(n12832), .A2(n9821), .ZN(n10036) );
  AND2_X1 U12662 ( .A1(n12935), .A2(n12938), .ZN(n10038) );
  NAND3_X1 U12663 ( .A1(n10040), .A2(n11425), .A3(n15945), .ZN(n10039) );
  INV_X1 U12664 ( .A(n11374), .ZN(n10042) );
  AND2_X1 U12665 ( .A1(n14935), .A2(n11559), .ZN(n10043) );
  NAND2_X1 U12666 ( .A1(n10043), .A2(n11563), .ZN(n14793) );
  INV_X1 U12667 ( .A(n14793), .ZN(n11561) );
  INV_X1 U12668 ( .A(n14159), .ZN(n10047) );
  NAND3_X1 U12669 ( .A1(n10047), .A2(n10046), .A3(n10045), .ZN(n10044) );
  AND2_X2 U12670 ( .A1(n10278), .A2(n13226), .ZN(n10287) );
  AND2_X1 U12671 ( .A1(n10606), .A2(n13936), .ZN(n13941) );
  NAND2_X1 U12672 ( .A1(n11478), .A2(n11477), .ZN(n11492) );
  AOI211_X1 U12673 ( .C1(n19063), .C2(n15097), .A(n14231), .B(n14230), .ZN(
        n14232) );
  INV_X4 U12674 ( .A(n14128), .ZN(n12819) );
  INV_X2 U12675 ( .A(n10243), .ZN(n14128) );
  AOI21_X1 U12676 ( .B1(n14471), .B2(n16153), .A(n14470), .ZN(n14472) );
  INV_X1 U12677 ( .A(n13734), .ZN(n10819) );
  XNOR2_X1 U12678 ( .A(n13333), .B(n13334), .ZN(n19479) );
  INV_X1 U12679 ( .A(n12989), .ZN(n10798) );
  NOR2_X2 U12680 ( .A1(n18019), .A2(n17700), .ZN(n17699) );
  NAND2_X1 U12681 ( .A1(n13216), .A2(n13215), .ZN(n13219) );
  OR2_X1 U12682 ( .A1(n12347), .A2(n12346), .ZN(P2_U3028) );
  XNOR2_X1 U12683 ( .A(n12920), .B(n10063), .ZN(n15258) );
  NOR2_X1 U12684 ( .A1(n12622), .A2(n17636), .ZN(n17408) );
  OAI21_X1 U12685 ( .B1(n13235), .B2(n13234), .A(n13233), .ZN(n19702) );
  NAND2_X1 U12686 ( .A1(n11296), .A2(n11276), .ZN(n11640) );
  NAND2_X2 U12687 ( .A1(n11183), .A2(n11182), .ZN(n11262) );
  INV_X1 U12688 ( .A(n10316), .ZN(n19475) );
  NAND2_X1 U12689 ( .A1(n13223), .A2(n13222), .ZN(n13301) );
  OR2_X1 U12690 ( .A1(n13223), .A2(n13222), .ZN(n13224) );
  INV_X1 U12691 ( .A(n20006), .ZN(n13072) );
  OR2_X2 U12692 ( .A1(n11651), .A2(n11268), .ZN(n10089) );
  NAND2_X1 U12693 ( .A1(n10865), .A2(n19100), .ZN(n10209) );
  CLKBUF_X1 U12694 ( .A(n13270), .Z(n14984) );
  INV_X1 U12695 ( .A(n10216), .ZN(n10528) );
  INV_X1 U12696 ( .A(n11640), .ZN(n11772) );
  XNOR2_X1 U12697 ( .A(n14354), .B(n14355), .ZN(n15096) );
  CLKBUF_X1 U12698 ( .A(n14159), .Z(n15765) );
  NAND2_X1 U12699 ( .A1(n10183), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10191) );
  NAND2_X1 U12700 ( .A1(n15096), .A2(n15095), .ZN(n15094) );
  NAND2_X1 U12701 ( .A1(n12836), .A2(n12837), .ZN(n12307) );
  OR2_X1 U12702 ( .A1(n14669), .A2(n20013), .ZN(n14684) );
  OR2_X1 U12703 ( .A1(n20013), .A2(n20244), .ZN(n12300) );
  AND3_X1 U12704 ( .A1(n11765), .A2(n13640), .A3(n11767), .ZN(n11285) );
  NAND2_X1 U12705 ( .A1(n15902), .A2(n13252), .ZN(n15900) );
  OR2_X1 U12706 ( .A1(n15976), .A2(n16077), .ZN(n10055) );
  INV_X1 U12707 ( .A(n12546), .ZN(n12519) );
  INV_X1 U12708 ( .A(n9719), .ZN(n12570) );
  OR3_X1 U12709 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17441), .ZN(n10057) );
  INV_X2 U12710 ( .A(n17272), .ZN(n17300) );
  NOR2_X1 U12711 ( .A1(n12735), .A2(n10073), .ZN(n10058) );
  OR2_X1 U12712 ( .A1(n11128), .A2(n19074), .ZN(n10059) );
  OR2_X1 U12713 ( .A1(n15180), .A2(n19072), .ZN(n10060) );
  NOR2_X1 U12714 ( .A1(n15416), .A2(n10660), .ZN(n10062) );
  AND2_X1 U12715 ( .A1(n14234), .A2(n12919), .ZN(n10063) );
  OR2_X1 U12716 ( .A1(n9764), .A2(n18947), .ZN(n10064) );
  AND2_X1 U12717 ( .A1(n14372), .A2(n14392), .ZN(n10065) );
  CLKBUF_X3 U12718 ( .A(n12542), .Z(n17049) );
  INV_X1 U12719 ( .A(n17231), .ZN(n17218) );
  NOR2_X1 U12720 ( .A1(n20439), .A2(n20050), .ZN(n10066) );
  OR2_X1 U12721 ( .A1(n16693), .A2(n12880), .ZN(n10067) );
  AND2_X1 U12722 ( .A1(n15728), .A2(n12903), .ZN(n10068) );
  NOR2_X1 U12723 ( .A1(n18592), .A2(n17630), .ZN(n17476) );
  INV_X1 U12724 ( .A(n17476), .ZN(n17508) );
  AND3_X1 U12725 ( .A1(n14206), .A2(n10706), .A3(n12330), .ZN(n10069) );
  OR2_X1 U12726 ( .A1(n14497), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10070) );
  OR2_X1 U12727 ( .A1(n14492), .A2(n13255), .ZN(n19928) );
  AND2_X1 U12728 ( .A1(n11147), .A2(n11146), .ZN(n10071) );
  AND2_X1 U12729 ( .A1(n13997), .A2(n19067), .ZN(n10072) );
  AND2_X1 U12730 ( .A1(n18800), .A2(n19067), .ZN(n10073) );
  NAND2_X1 U12731 ( .A1(n12605), .A2(n17690), .ZN(n10074) );
  OR2_X1 U12732 ( .A1(n17636), .A2(n17366), .ZN(n10075) );
  OR2_X1 U12733 ( .A1(n19803), .A2(n14546), .ZN(n10076) );
  INV_X1 U12734 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13318) );
  NAND2_X1 U12735 ( .A1(n17390), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12349) );
  OR2_X1 U12736 ( .A1(n14497), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10077) );
  OR3_X1 U12737 ( .A1(n12497), .A2(n12496), .A3(n12495), .ZN(P3_U2640) );
  INV_X1 U12738 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13274) );
  INV_X1 U12739 ( .A(n13678), .ZN(n10432) );
  AND2_X1 U12740 ( .A1(n12453), .A2(n12452), .ZN(n10079) );
  INV_X1 U12741 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19819) );
  INV_X1 U12742 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17718) );
  INV_X1 U12743 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17704) );
  NAND2_X1 U12744 ( .A1(n12720), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15223) );
  AND3_X1 U12745 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10080) );
  INV_X1 U12746 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19779) );
  NOR2_X1 U12747 ( .A1(n20439), .A2(n20578), .ZN(n10081) );
  AND3_X1 U12748 ( .A1(n10109), .A2(n10108), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10082) );
  INV_X1 U12749 ( .A(n14532), .ZN(n14544) );
  INV_X2 U12750 ( .A(n17089), .ZN(n17079) );
  AND3_X1 U12751 ( .A1(n12889), .A2(n12888), .A3(n12887), .ZN(n10084) );
  INV_X1 U12752 ( .A(n17537), .ZN(n17735) );
  NOR2_X1 U12753 ( .A1(n18728), .A2(n16359), .ZN(n17537) );
  AND2_X1 U12754 ( .A1(n11127), .A2(n11126), .ZN(n10085) );
  OR2_X1 U12755 ( .A1(n12736), .A2(n16083), .ZN(n10086) );
  OR2_X1 U12756 ( .A1(n11128), .A2(n16083), .ZN(n10087) );
  INV_X1 U12757 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11930) );
  AND2_X4 U12758 ( .A1(n11538), .A2(n11537), .ZN(n10088) );
  AND2_X1 U12759 ( .A1(n11598), .A2(n11582), .ZN(n11604) );
  AOI21_X1 U12760 ( .B1(n10252), .B2(P2_REIP_REG_1__SCAN_IN), .A(n10244), .ZN(
        n10245) );
  NAND2_X1 U12761 ( .A1(n10430), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10324) );
  AOI22_X1 U12762 ( .A1(n15475), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n10266), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U12763 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10432), .B1(
        n10433), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10292) );
  AND2_X1 U12764 ( .A1(n20471), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11592) );
  OR2_X1 U12765 ( .A1(n11514), .A2(n11513), .ZN(n11528) );
  NAND2_X1 U12766 ( .A1(n11778), .A2(n11282), .ZN(n13263) );
  NAND2_X1 U12767 ( .A1(n13073), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11432) );
  AND2_X1 U12768 ( .A1(n13144), .A2(n10312), .ZN(n10850) );
  INV_X1 U12769 ( .A(n16071), .ZN(n10642) );
  OR2_X1 U12770 ( .A1(n10417), .A2(n10416), .ZN(n10523) );
  OAI21_X1 U12771 ( .B1(n10214), .B2(n10216), .A(n19100), .ZN(n10218) );
  OR2_X1 U12772 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19973), .ZN(
        n11575) );
  AND2_X2 U12773 ( .A1(n11157), .A2(n11158), .ZN(n11437) );
  INV_X1 U12774 ( .A(n14534), .ZN(n12283) );
  INV_X1 U12775 ( .A(n13924), .ZN(n12012) );
  NOR2_X1 U12776 ( .A1(n11353), .A2(n15945), .ZN(n11536) );
  INV_X1 U12777 ( .A(n11262), .ZN(n11274) );
  OR2_X1 U12778 ( .A1(n11444), .A2(n11443), .ZN(n11451) );
  INV_X1 U12779 ( .A(n14355), .ZN(n14356) );
  INV_X1 U12780 ( .A(n13340), .ZN(n10767) );
  INV_X1 U12781 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12852) );
  NOR2_X1 U12782 ( .A1(n16028), .A2(n10735), .ZN(n10717) );
  NAND2_X1 U12783 ( .A1(n10505), .A2(n10504), .ZN(n16066) );
  NAND2_X1 U12784 ( .A1(n10419), .A2(n10451), .ZN(n10454) );
  INV_X1 U12785 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n20819) );
  AND2_X1 U12786 ( .A1(n11576), .A2(n11575), .ZN(n11636) );
  NAND2_X1 U12787 ( .A1(n11369), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11293) );
  INV_X1 U12788 ( .A(n11744), .ZN(n11752) );
  AND2_X1 U12789 ( .A1(n14479), .A2(n12303), .ZN(n12304) );
  NAND2_X1 U12790 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11244) );
  INV_X1 U12791 ( .A(n14835), .ZN(n11550) );
  INV_X1 U12792 ( .A(n13414), .ZN(n11937) );
  INV_X1 U12793 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11559) );
  NAND2_X1 U12794 ( .A1(n20736), .A2(n15945), .ZN(n11446) );
  INV_X1 U12795 ( .A(n11350), .ZN(n11351) );
  NAND2_X1 U12797 ( .A1(n10268), .A2(n10267), .ZN(n10756) );
  AND2_X1 U12798 ( .A1(n15166), .A2(n11066), .ZN(n11064) );
  AND2_X1 U12799 ( .A1(n10772), .A2(n10771), .ZN(n13347) );
  OR3_X1 U12800 ( .A1(n15358), .A2(n20857), .A3(n12338), .ZN(n12730) );
  OR2_X1 U12801 ( .A1(n18819), .A2(n10934), .ZN(n10723) );
  AND2_X1 U12802 ( .A1(n18932), .A2(n10274), .ZN(n10289) );
  AND2_X1 U12803 ( .A1(n18932), .A2(n10285), .ZN(n10286) );
  INV_X1 U12804 ( .A(n17413), .ZN(n12365) );
  INV_X1 U12805 ( .A(n16686), .ZN(n12553) );
  AOI21_X1 U12806 ( .B1(n17636), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n12632), .ZN(n12633) );
  AND2_X1 U12807 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12604), .ZN(
        n12603) );
  OR2_X1 U12808 ( .A1(n12302), .A2(n12843), .ZN(n12941) );
  OR2_X1 U12809 ( .A1(n15576), .A2(n13635), .ZN(n13636) );
  NOR2_X1 U12810 ( .A1(n13069), .A2(n13033), .ZN(n11748) );
  NOR2_X1 U12811 ( .A1(n12092), .A2(n14841), .ZN(n12146) );
  INV_X1 U12812 ( .A(n12224), .ZN(n12303) );
  INV_X1 U12813 ( .A(n11912), .ZN(n11966) );
  NAND3_X1 U12814 ( .A1(n11564), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14792), .ZN(n14772) );
  INV_X1 U12815 ( .A(n15774), .ZN(n11533) );
  NAND2_X1 U12816 ( .A1(n11356), .A2(n11355), .ZN(n11390) );
  OR2_X1 U12817 ( .A1(n10870), .A2(n10869), .ZN(n16186) );
  INV_X1 U12818 ( .A(n10683), .ZN(n10690) );
  INV_X1 U12819 ( .A(n13610), .ZN(n10803) );
  INV_X1 U12820 ( .A(n16083), .ZN(n14248) );
  AND2_X1 U12821 ( .A1(n10260), .A2(n10261), .ZN(n10271) );
  AND2_X1 U12822 ( .A1(n15309), .A2(n14198), .ZN(n14194) );
  OR2_X1 U12823 ( .A1(n12974), .A2(n10934), .ZN(n10746) );
  INV_X1 U12824 ( .A(n12867), .ZN(n10511) );
  OR2_X1 U12825 ( .A1(n18847), .A2(n10934), .ZN(n10725) );
  INV_X1 U12826 ( .A(n15375), .ZN(n15410) );
  NOR2_X1 U12827 ( .A1(n16115), .A2(n10880), .ZN(n15402) );
  OR2_X1 U12828 ( .A1(n13781), .A2(n10934), .ZN(n10663) );
  AND2_X1 U12829 ( .A1(n10641), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16071) );
  INV_X1 U12830 ( .A(n16186), .ZN(n13134) );
  INV_X1 U12831 ( .A(n19254), .ZN(n19257) );
  OR3_X1 U12832 ( .A1(n19475), .A2(n19500), .A3(n19732), .ZN(n19481) );
  INV_X1 U12833 ( .A(n12633), .ZN(n12634) );
  OR2_X1 U12834 ( .A1(n17408), .A2(n12623), .ZN(n12624) );
  NAND2_X1 U12835 ( .A1(n12268), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12280) );
  AND2_X1 U12836 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n11811), .ZN(
        n12248) );
  AND2_X1 U12837 ( .A1(n11723), .A2(n11722), .ZN(n14644) );
  AND2_X1 U12838 ( .A1(n13644), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13637) );
  NOR2_X1 U12839 ( .A1(n13643), .A2(n13642), .ZN(n13649) );
  INV_X1 U12840 ( .A(n19751), .ZN(n13183) );
  NOR2_X1 U12841 ( .A1(n12058), .A2(n14177), .ZN(n12112) );
  AND2_X1 U12842 ( .A1(n12057), .A2(n12023), .ZN(n14152) );
  OR2_X1 U12843 ( .A1(n14848), .A2(n14847), .ZN(n15750) );
  NAND2_X1 U12844 ( .A1(n15777), .A2(n11535), .ZN(n13846) );
  AND2_X1 U12845 ( .A1(n11648), .A2(n13183), .ZN(n11795) );
  AND3_X1 U12846 ( .A1(n13294), .A2(n13293), .A3(n13292), .ZN(n13562) );
  AND2_X1 U12847 ( .A1(n20131), .A2(n20130), .ZN(n20160) );
  AND2_X1 U12848 ( .A1(n20170), .A2(n20169), .ZN(n20199) );
  AND2_X1 U12849 ( .A1(n20287), .A2(n20286), .ZN(n20314) );
  OR2_X1 U12850 ( .A1(n20735), .A2(n11410), .ZN(n20742) );
  AND2_X1 U12851 ( .A1(n20474), .A2(n20473), .ZN(n20499) );
  INV_X1 U12852 ( .A(n20541), .ZN(n20610) );
  OR2_X1 U12853 ( .A1(n10638), .A2(n9757), .ZN(n10689) );
  INV_X1 U12854 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14032) );
  AND2_X1 U12855 ( .A1(n10750), .A2(n10749), .ZN(n10845) );
  AND2_X1 U12856 ( .A1(n10823), .A2(n10822), .ZN(n13949) );
  OR2_X1 U12857 ( .A1(n11004), .A2(n11003), .ZN(n18956) );
  AND2_X1 U12858 ( .A1(n10933), .A2(n10932), .ZN(n13142) );
  NAND2_X2 U12859 ( .A1(n10191), .A2(n10190), .ZN(n10216) );
  AOI21_X1 U12860 ( .B1(n16143), .B2(n15088), .A(n11145), .ZN(n11146) );
  AND2_X1 U12861 ( .A1(n10802), .A2(n10801), .ZN(n13610) );
  AND2_X1 U12862 ( .A1(n16113), .A2(n10881), .ZN(n16102) );
  XNOR2_X1 U12863 ( .A(n10506), .B(n10934), .ZN(n14022) );
  NAND2_X1 U12864 ( .A1(n10891), .A2(n10848), .ZN(n19072) );
  AND2_X1 U12865 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19407) );
  INV_X1 U12866 ( .A(n10344), .ZN(n19281) );
  OR3_X1 U12867 ( .A1(n10314), .A2(n19333), .A3(n19732), .ZN(n13723) );
  OR2_X1 U12868 ( .A1(n10434), .A2(n19408), .ZN(n19414) );
  NOR2_X1 U12869 ( .A1(n12696), .A2(n12472), .ZN(n15519) );
  NOR2_X1 U12870 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16620), .ZN(n16609) );
  NOR2_X1 U12871 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16642), .ZN(n16628) );
  AOI211_X1 U12872 ( .C1(n9717), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n12430), .B(n12429), .ZN(n12431) );
  INV_X1 U12873 ( .A(n18109), .ZN(n17101) );
  AOI21_X1 U12874 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17476), .A(
        n18460), .ZN(n17572) );
  NAND2_X1 U12875 ( .A1(n12693), .A2(n17628), .ZN(n17933) );
  NAND2_X1 U12876 ( .A1(n17559), .A2(n17842), .ZN(n17521) );
  NAND2_X1 U12877 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n12711), .ZN(
        n17908) );
  INV_X1 U12878 ( .A(n17651), .ZN(n17652) );
  XNOR2_X1 U12879 ( .A(n12598), .B(n18043), .ZN(n17709) );
  INV_X1 U12880 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18555) );
  INV_X1 U12881 ( .A(n16678), .ZN(n18084) );
  NOR2_X1 U12882 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18082), .ZN(n18426) );
  INV_X1 U12883 ( .A(n15519), .ZN(n15520) );
  INV_X1 U12884 ( .A(n13280), .ZN(n13290) );
  OR2_X1 U12885 ( .A1(n15579), .A2(n15945), .ZN(n19751) );
  NAND2_X1 U12886 ( .A1(n12248), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12258) );
  INV_X1 U12887 ( .A(n19845), .ZN(n19853) );
  NOR2_X1 U12888 ( .A1(n19754), .A2(n19803), .ZN(n19836) );
  NAND2_X1 U12889 ( .A1(n11948), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11947) );
  INV_X1 U12891 ( .A(n14684), .ZN(n14670) );
  INV_X1 U12892 ( .A(n15723), .ZN(n14731) );
  INV_X1 U12893 ( .A(n14740), .ZN(n15726) );
  INV_X1 U12894 ( .A(n13360), .ZN(n13470) );
  NAND2_X1 U12895 ( .A1(n12185), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12203) );
  AND2_X1 U12896 ( .A1(n14666), .A2(n14665), .ZN(n15755) );
  NAND2_X1 U12897 ( .A1(n14774), .A2(n14773), .ZN(n14776) );
  OR2_X1 U12898 ( .A1(n15591), .A2(n11805), .ZN(n15796) );
  OR2_X1 U12899 ( .A1(n14164), .A2(n14163), .ZN(n15759) );
  INV_X1 U12900 ( .A(n15908), .ZN(n19953) );
  OR2_X1 U12901 ( .A1(n19967), .A2(n19969), .ZN(n15907) );
  AND2_X1 U12902 ( .A1(n12840), .A2(n20244), .ZN(n19939) );
  OAI22_X1 U12903 ( .A1(n19989), .A2(n19988), .B1(n20366), .B2(n20129), .ZN(
        n20018) );
  INV_X1 U12904 ( .A(n20086), .ZN(n20053) );
  OAI22_X1 U12905 ( .A1(n20059), .A2(n20058), .B1(n20366), .B2(n20212), .ZN(
        n20082) );
  INV_X1 U12906 ( .A(n20166), .ZN(n20157) );
  INV_X1 U12907 ( .A(n20236), .ZN(n20195) );
  NOR2_X1 U12908 ( .A1(n20249), .A2(n9766), .ZN(n20176) );
  INV_X1 U12909 ( .A(n20276), .ZN(n20317) );
  INV_X1 U12910 ( .A(n20395), .ZN(n20355) );
  OAI22_X1 U12911 ( .A1(n20368), .A2(n20367), .B1(n20366), .B2(n20509), .ZN(
        n20391) );
  NOR2_X1 U12912 ( .A1(n20742), .A2(n9766), .ZN(n20331) );
  OAI22_X1 U12913 ( .A1(n20450), .A2(n20449), .B1(n20448), .B2(n20447), .ZN(
        n20465) );
  INV_X1 U12914 ( .A(n20253), .ZN(n20408) );
  AND2_X1 U12915 ( .A1(n20476), .A2(n20438), .ZN(n20502) );
  NOR2_X1 U12916 ( .A1(n19993), .A2(n20135), .ZN(n20529) );
  NOR2_X1 U12917 ( .A1(n20003), .A2(n20135), .ZN(n20547) );
  OAI211_X1 U12918 ( .C1(n20567), .C2(n20523), .A(n20522), .B(n20521), .ZN(
        n20571) );
  NOR2_X2 U12919 ( .A1(n20588), .A2(n20253), .ZN(n20644) );
  NOR2_X1 U12920 ( .A1(n18896), .A2(n15032), .ZN(n15006) );
  INV_X1 U12921 ( .A(n18885), .ZN(n18927) );
  AND2_X1 U12922 ( .A1(n12826), .A2(n12784), .ZN(n18885) );
  AND2_X1 U12923 ( .A1(n18753), .A2(n12801), .ZN(n18922) );
  INV_X1 U12924 ( .A(n19602), .ZN(n18917) );
  INV_X1 U12925 ( .A(n18908), .ZN(n18939) );
  INV_X1 U12926 ( .A(n11065), .ZN(n14039) );
  INV_X1 U12927 ( .A(n15168), .ZN(n18995) );
  AND2_X1 U12928 ( .A1(n13015), .A2(n13014), .ZN(n19029) );
  INV_X1 U12929 ( .A(n13133), .ZN(n13107) );
  INV_X1 U12930 ( .A(n13112), .ZN(n13130) );
  AOI21_X1 U12931 ( .B1(n18809), .B2(n19063), .A(n12950), .ZN(n12951) );
  AND2_X1 U12932 ( .A1(n16100), .A2(n14257), .ZN(n16090) );
  INV_X1 U12933 ( .A(n16100), .ZN(n19055) );
  INV_X1 U12934 ( .A(n11071), .ZN(n11072) );
  AND2_X1 U12935 ( .A1(n14209), .A2(n14208), .ZN(n15221) );
  INV_X1 U12936 ( .A(n11123), .ZN(n19044) );
  INV_X1 U12937 ( .A(n19074), .ZN(n16153) );
  INV_X1 U12938 ( .A(n16161), .ZN(n19067) );
  NAND2_X1 U12939 ( .A1(n19092), .A2(n19091), .ZN(n19128) );
  INV_X1 U12940 ( .A(n19404), .ZN(n13682) );
  NAND2_X1 U12941 ( .A1(n15488), .A2(n19702), .ZN(n19404) );
  AND2_X1 U12942 ( .A1(n19212), .A2(n19252), .ZN(n21079) );
  NOR2_X1 U12943 ( .A1(n19250), .A2(n19439), .ZN(n19305) );
  AND2_X1 U12944 ( .A1(n13723), .A2(n13722), .ZN(n19323) );
  NAND2_X1 U12945 ( .A1(n19336), .A2(n19335), .ZN(n19353) );
  AND2_X1 U12946 ( .A1(n19414), .A2(n19410), .ZN(n19434) );
  NOR2_X1 U12947 ( .A1(n19440), .A2(n19439), .ZN(n19503) );
  INV_X1 U12948 ( .A(n19535), .ZN(n19525) );
  INV_X1 U12949 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19732) );
  NOR2_X1 U12950 ( .A1(n18090), .A2(n18084), .ZN(n14108) );
  AOI22_X1 U12951 ( .A1(n18516), .A2(n18515), .B1(n18520), .B2(n16253), .ZN(
        n18524) );
  NOR2_X1 U12952 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16501), .ZN(n16488) );
  NOR2_X1 U12953 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16526), .ZN(n16509) );
  NOR2_X1 U12954 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16549), .ZN(n16530) );
  NOR2_X1 U12955 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16593), .ZN(n16580) );
  NOR2_X1 U12956 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16665), .ZN(n16650) );
  INV_X1 U12957 ( .A(n16723), .ZN(n16704) );
  NOR2_X2 U12958 ( .A1(n18678), .A2(n16720), .ZN(n16725) );
  NAND2_X1 U12959 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17120), .ZN(n17116) );
  NOR3_X1 U12960 ( .A1(n18119), .A2(n17171), .A3(n17273), .ZN(n17163) );
  NOR2_X1 U12961 ( .A1(n17199), .A2(n17203), .ZN(n17198) );
  NOR2_X1 U12962 ( .A1(n18109), .A2(n17098), .ZN(n18548) );
  AOI22_X1 U12963 ( .A1(n18726), .A2(n15610), .B1(n15609), .B2(n15608), .ZN(
        n17096) );
  NAND2_X1 U12964 ( .A1(n18726), .A2(n18519), .ZN(n17307) );
  INV_X1 U12965 ( .A(n17357), .ZN(n17348) );
  NAND2_X1 U12966 ( .A1(n17935), .A2(n17842), .ZN(n17881) );
  INV_X1 U12967 ( .A(n17799), .ZN(n17883) );
  INV_X1 U12968 ( .A(n17627), .ZN(n17639) );
  INV_X1 U12969 ( .A(n18057), .ZN(n18050) );
  OR2_X1 U12970 ( .A1(n18742), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18044) );
  AOI21_X2 U12971 ( .B1(n15515), .B2(n12665), .A(n18579), .ZN(n18057) );
  INV_X1 U12972 ( .A(n18225), .ZN(n18231) );
  INV_X1 U12973 ( .A(n18252), .ZN(n18254) );
  INV_X1 U12974 ( .A(n18415), .ZN(n18416) );
  INV_X1 U12975 ( .A(U212), .ZN(n16304) );
  NAND2_X1 U12976 ( .A1(n13290), .A2(n13031), .ZN(n14492) );
  NAND2_X1 U12977 ( .A1(n14491), .A2(n14492), .ZN(n20758) );
  XOR2_X1 U12978 ( .A(n14496), .B(n11759), .Z(n14516) );
  INV_X1 U12979 ( .A(n19858), .ZN(n19840) );
  INV_X1 U12980 ( .A(n19863), .ZN(n19791) );
  INV_X1 U12981 ( .A(n19821), .ZN(n15629) );
  INV_X1 U12982 ( .A(n19865), .ZN(n19851) );
  OR2_X1 U12983 ( .A1(n13439), .A2(n19974), .ZN(n15723) );
  INV_X1 U12984 ( .A(n15755), .ZN(n14743) );
  NAND2_X1 U12985 ( .A1(n15728), .A2(n13437), .ZN(n14740) );
  INV_X2 U12986 ( .A(n15717), .ZN(n15728) );
  OR2_X1 U12987 ( .A1(n19897), .A2(n13187), .ZN(n19888) );
  INV_X1 U12988 ( .A(n19897), .ZN(n19895) );
  INV_X1 U12989 ( .A(n19928), .ZN(n13360) );
  INV_X1 U12990 ( .A(n12944), .ZN(n12945) );
  OAI21_X1 U12991 ( .B1(n14575), .B2(n14642), .A(n14638), .ZN(n14827) );
  INV_X1 U12992 ( .A(n15791), .ZN(n15787) );
  INV_X1 U12993 ( .A(n19938), .ZN(n19757) );
  INV_X1 U12994 ( .A(n19965), .ZN(n15872) );
  INV_X1 U12995 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20471) );
  OR2_X1 U12996 ( .A1(n20022), .A2(n20470), .ZN(n20048) );
  OR2_X1 U12997 ( .A1(n20022), .A2(n20438), .ZN(n20086) );
  OR2_X1 U12998 ( .A1(n20092), .A2(n20253), .ZN(n20166) );
  NAND2_X1 U12999 ( .A1(n20176), .A2(n20438), .ZN(n20198) );
  NAND2_X1 U13000 ( .A1(n20176), .A2(n20470), .ZN(n20236) );
  NAND2_X1 U13001 ( .A1(n20254), .A2(n20506), .ZN(n20283) );
  NAND2_X1 U13002 ( .A1(n20331), .A2(n20438), .ZN(n20359) );
  NAND2_X1 U13003 ( .A1(n20331), .A2(n20470), .ZN(n20395) );
  NAND2_X1 U13004 ( .A1(n20409), .A2(n20506), .ZN(n20427) );
  NAND2_X1 U13005 ( .A1(n20409), .A2(n20408), .ZN(n20469) );
  NAND2_X1 U13006 ( .A1(n20476), .A2(n20470), .ZN(n20524) );
  NAND2_X1 U13007 ( .A1(n20507), .A2(n20506), .ZN(n20648) );
  INV_X1 U13008 ( .A(n20724), .ZN(n20720) );
  AND2_X1 U13009 ( .A1(n12829), .A2(n9801), .ZN(n12830) );
  OR2_X1 U13010 ( .A1(n12828), .A2(n12827), .ZN(n18900) );
  OR2_X1 U13011 ( .A1(n13996), .A2(n13995), .ZN(n15988) );
  AND2_X1 U13012 ( .A1(n13140), .A2(n19731), .ZN(n15168) );
  OR2_X1 U13013 ( .A1(n18995), .A2(n13144), .ZN(n18998) );
  OR2_X1 U13014 ( .A1(n19029), .A2(n19041), .ZN(n19016) );
  INV_X1 U13015 ( .A(n19029), .ZN(n19043) );
  INV_X1 U13016 ( .A(n13060), .ZN(n13112) );
  OAI21_X1 U13017 ( .B1(n12952), .B2(n16084), .A(n12951), .ZN(n12953) );
  INV_X1 U13018 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18853) );
  OR2_X1 U13019 ( .A1(n18757), .A2(n10215), .ZN(n16083) );
  INV_X1 U13020 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19715) );
  INV_X1 U13021 ( .A(n19153), .ZN(n19162) );
  NAND2_X1 U13022 ( .A1(n19212), .A2(n13682), .ZN(n19211) );
  OR2_X1 U13023 ( .A1(n19250), .A2(n19404), .ZN(n19243) );
  INV_X1 U13024 ( .A(n21079), .ZN(n19273) );
  INV_X1 U13025 ( .A(n19305), .ZN(n21086) );
  OR2_X1 U13026 ( .A1(n19250), .A2(n19084), .ZN(n19357) );
  INV_X1 U13027 ( .A(n19372), .ZN(n19364) );
  OR2_X1 U13028 ( .A1(n19405), .A2(n19132), .ZN(n19375) );
  INV_X1 U13029 ( .A(n19564), .ZN(n19424) );
  INV_X1 U13030 ( .A(n19427), .ZN(n19438) );
  INV_X1 U13031 ( .A(n19503), .ZN(n19499) );
  INV_X1 U13032 ( .A(n19532), .ZN(n19529) );
  OR2_X1 U13033 ( .A1(n19440), .A2(n19084), .ZN(n19593) );
  NOR2_X1 U13034 ( .A1(n18518), .A2(n17307), .ZN(n18745) );
  INV_X1 U13035 ( .A(n16732), .ZN(n16692) );
  NOR2_X1 U13036 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16576), .ZN(n16566) );
  NOR2_X1 U13037 ( .A1(n12581), .A2(n12580), .ZN(n17215) );
  NOR2_X1 U13038 ( .A1(n12529), .A2(n12528), .ZN(n17230) );
  NAND2_X1 U13039 ( .A1(n17287), .A2(n17303), .ZN(n17272) );
  NAND2_X1 U13040 ( .A1(n17248), .A2(n17247), .ZN(n17303) );
  AOI221_X1 U13041 ( .B1(n18730), .B2(n18572), .C1(n17308), .C2(n18572), .A(
        n17307), .ZN(n17311) );
  INV_X1 U13042 ( .A(n17355), .ZN(n17350) );
  NAND2_X1 U13043 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17728), .ZN(n17583) );
  NAND2_X1 U13044 ( .A1(n16252), .A2(n9765), .ZN(n17627) );
  INV_X1 U13045 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17695) );
  NOR2_X1 U13046 ( .A1(n17630), .A2(n17705), .ZN(n17728) );
  NAND2_X1 U13047 ( .A1(n16252), .A2(n18048), .ZN(n17964) );
  INV_X1 U13048 ( .A(n18060), .ZN(n18055) );
  INV_X1 U13049 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18564) );
  INV_X1 U13050 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18525) );
  INV_X1 U13051 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18107) );
  INV_X1 U13052 ( .A(n18129), .ZN(n18470) );
  INV_X1 U13053 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18678) );
  INV_X1 U13054 ( .A(n18675), .ZN(n18672) );
  INV_X1 U13055 ( .A(n18740), .ZN(n18719) );
  INV_X1 U13056 ( .A(n16310), .ZN(n16313) );
  OAI21_X1 U13057 ( .B1(n14690), .B2(n14672), .A(n12318), .ZN(P1_U2842) );
  OAI211_X1 U13058 ( .C1(n14887), .C2(n19757), .A(n10054), .B(n12845), .ZN(
        P1_U2970) );
  NAND2_X1 U13059 ( .A1(n10087), .A2(n10085), .ZN(P2_U2988) );
  NAND2_X1 U13060 ( .A1(n10086), .A2(n12745), .ZN(P2_U2995) );
  NAND2_X1 U13061 ( .A1(n10059), .A2(n10071), .ZN(P2_U3020) );
  AOI22_X1 U13062 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n9755), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10096) );
  AOI22_X1 U13063 ( .A1(n10110), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U13064 ( .A1(n9775), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(n9749), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10094) );
  AOI22_X1 U13065 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(n9756), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10093) );
  AOI22_X1 U13066 ( .A1(n10110), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10100) );
  AOI22_X1 U13067 ( .A1(n9733), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10297), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10099) );
  AOI22_X1 U13068 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10098) );
  AOI22_X1 U13069 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14439), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10097) );
  AND4_X1 U13070 ( .A1(n10100), .A2(n10099), .A3(n10098), .A4(n10097), .ZN(
        n10101) );
  MUX2_X2 U13071 ( .A(n10102), .B(n10101), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10195) );
  AOI22_X1 U13072 ( .A1(n10295), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9775), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10106) );
  AOI22_X1 U13073 ( .A1(n10110), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10105) );
  AOI22_X1 U13074 ( .A1(n9755), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10297), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10104) );
  AOI22_X1 U13075 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(n9756), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10103) );
  NAND2_X1 U13076 ( .A1(n10107), .A2(n10188), .ZN(n10114) );
  AOI22_X1 U13077 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9756), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10109) );
  AOI22_X1 U13078 ( .A1(n9748), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10108) );
  AOI22_X1 U13079 ( .A1(n9755), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9775), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U13080 ( .A1(n10295), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10110), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10111) );
  NAND3_X1 U13081 ( .A1(n10082), .A2(n10112), .A3(n10111), .ZN(n10113) );
  AOI22_X1 U13082 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n9755), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10118) );
  AOI22_X1 U13083 ( .A1(n10110), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10117) );
  AOI22_X1 U13084 ( .A1(n9775), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10297), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10116) );
  NAND4_X1 U13085 ( .A1(n10118), .A2(n10117), .A3(n10116), .A4(n10115), .ZN(
        n10124) );
  AOI22_X1 U13086 ( .A1(n10295), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9755), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10122) );
  AOI22_X1 U13087 ( .A1(n10110), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10121) );
  AOI22_X1 U13088 ( .A1(n9733), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10297), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10120) );
  AOI22_X1 U13089 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14439), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10119) );
  NAND4_X1 U13090 ( .A1(n10122), .A2(n10121), .A3(n10120), .A4(n10119), .ZN(
        n10123) );
  AOI22_X1 U13092 ( .A1(n9775), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9749), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10128) );
  AOI22_X1 U13093 ( .A1(n10110), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10127) );
  AOI22_X1 U13094 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9755), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10126) );
  AOI22_X1 U13095 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14439), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10125) );
  NAND4_X1 U13096 ( .A1(n10128), .A2(n10127), .A3(n10126), .A4(n10125), .ZN(
        n10129) );
  AOI22_X1 U13097 ( .A1(n10110), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U13098 ( .A1(n9733), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10297), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10132) );
  AOI22_X1 U13099 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10131) );
  AOI22_X1 U13100 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14439), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10130) );
  NAND4_X1 U13101 ( .A1(n10133), .A2(n10132), .A3(n10131), .A4(n10130), .ZN(
        n10134) );
  NAND2_X1 U13102 ( .A1(n10134), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10135) );
  AOI22_X1 U13103 ( .A1(n10295), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10141) );
  AOI22_X1 U13104 ( .A1(n10110), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10140) );
  AOI22_X1 U13105 ( .A1(n9733), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9749), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10139) );
  AOI22_X1 U13106 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14439), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10138) );
  NAND4_X1 U13107 ( .A1(n10141), .A2(n10140), .A3(n10139), .A4(n10138), .ZN(
        n10142) );
  AOI22_X1 U13108 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9755), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U13109 ( .A1(n9775), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9748), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10145) );
  NAND4_X1 U13110 ( .A1(n10147), .A2(n10146), .A3(n10145), .A4(n10144), .ZN(
        n10148) );
  AOI22_X1 U13111 ( .A1(n10110), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10152) );
  AOI22_X1 U13112 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9756), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U13113 ( .A1(n9733), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9748), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10154) );
  AOI22_X1 U13114 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10153) );
  NAND3_X1 U13115 ( .A1(n10155), .A2(n10154), .A3(n10153), .ZN(n10162) );
  AOI22_X1 U13116 ( .A1(n10110), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U13117 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14439), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10156) );
  AND3_X1 U13118 ( .A1(n10157), .A2(n10156), .A3(n10188), .ZN(n10160) );
  AOI22_X1 U13119 ( .A1(n9755), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10297), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U13120 ( .A1(n10295), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9733), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10158) );
  NAND3_X1 U13121 ( .A1(n10160), .A2(n10159), .A3(n10158), .ZN(n10161) );
  NOR2_X1 U13122 ( .A1(n10205), .A2(n10558), .ZN(n10163) );
  AND2_X2 U13123 ( .A1(n10176), .A2(n10163), .ZN(n16189) );
  AOI22_X1 U13124 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U13125 ( .A1(n10110), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10166) );
  AOI22_X1 U13126 ( .A1(n9775), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(n9748), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U13127 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(n9756), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10164) );
  NAND4_X1 U13128 ( .A1(n10167), .A2(n10166), .A3(n10165), .A4(n10164), .ZN(
        n10168) );
  AOI22_X1 U13129 ( .A1(n10296), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10110), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U13130 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14439), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10171) );
  AOI22_X1 U13131 ( .A1(n9733), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(n9754), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U13132 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10297), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10169) );
  NAND4_X1 U13133 ( .A1(n10172), .A2(n10171), .A3(n10170), .A4(n10169), .ZN(
        n10173) );
  NAND2_X1 U13134 ( .A1(n13724), .A2(n10215), .ZN(n10178) );
  OAI21_X1 U13135 ( .B1(n16189), .B2(n10178), .A(n10177), .ZN(n10886) );
  INV_X1 U13136 ( .A(n10886), .ZN(n10192) );
  AOI22_X1 U13137 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10110), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U13138 ( .A1(n10296), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9733), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10181) );
  AOI22_X1 U13139 ( .A1(n9749), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U13140 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14439), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10179) );
  NAND4_X1 U13141 ( .A1(n10182), .A2(n10181), .A3(n10180), .A4(n10179), .ZN(
        n10183) );
  AOI22_X1 U13142 ( .A1(n10295), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9775), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U13143 ( .A1(n9755), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n9749), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10186) );
  AOI22_X1 U13144 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14439), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U13145 ( .A1(n10110), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10184) );
  NAND4_X1 U13146 ( .A1(n10187), .A2(n10186), .A3(n10185), .A4(n10184), .ZN(
        n10189) );
  NAND2_X1 U13147 ( .A1(n10189), .A2(n10188), .ZN(n10190) );
  NAND2_X1 U13148 ( .A1(n10192), .A2(n9776), .ZN(n10201) );
  NAND2_X2 U13149 ( .A1(n19115), .A2(n9763), .ZN(n13144) );
  NAND4_X1 U13150 ( .A1(n10203), .A2(n10857), .A3(n10195), .A4(n9764), .ZN(
        n10226) );
  NAND2_X1 U13151 ( .A1(n10205), .A2(n13724), .ZN(n10194) );
  NAND2_X1 U13152 ( .A1(n10226), .A2(n10194), .ZN(n10199) );
  INV_X1 U13153 ( .A(n10557), .ZN(n10197) );
  INV_X1 U13154 ( .A(n10195), .ZN(n10202) );
  NAND2_X1 U13155 ( .A1(n10195), .A2(n10193), .ZN(n10196) );
  NAND2_X1 U13156 ( .A1(n10197), .A2(n10196), .ZN(n10198) );
  NAND2_X1 U13157 ( .A1(n13144), .A2(n10208), .ZN(n10217) );
  NAND3_X1 U13158 ( .A1(n10199), .A2(n10198), .A3(n10217), .ZN(n10856) );
  NOR2_X1 U13159 ( .A1(n10216), .A2(n19727), .ZN(n19735) );
  OAI21_X1 U13160 ( .B1(n10231), .B2(n10856), .A(n19735), .ZN(n10200) );
  AND2_X2 U13161 ( .A1(n10201), .A2(n10200), .ZN(n10230) );
  NAND2_X1 U13162 ( .A1(n13144), .A2(n10202), .ZN(n10555) );
  NAND2_X1 U13163 ( .A1(n10214), .A2(n10205), .ZN(n10561) );
  INV_X1 U13164 ( .A(n10561), .ZN(n10206) );
  NAND2_X1 U13165 ( .A1(n10206), .A2(n10195), .ZN(n10563) );
  NAND2_X1 U13166 ( .A1(n10207), .A2(n10563), .ZN(n10859) );
  NAND2_X1 U13167 ( .A1(n10859), .A2(n10208), .ZN(n10210) );
  NAND2_X1 U13168 ( .A1(n10210), .A2(n10209), .ZN(n10232) );
  NAND2_X1 U13169 ( .A1(n10232), .A2(n9776), .ZN(n10211) );
  NAND2_X2 U13170 ( .A1(n10230), .A2(n10211), .ZN(n10265) );
  NAND2_X2 U13171 ( .A1(n10213), .A2(n13009), .ZN(n10243) );
  OAI22_X1 U13172 ( .A1(n10265), .A2(n10213), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14128), .ZN(n10221) );
  NOR2_X1 U13173 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10266) );
  NAND2_X1 U13174 ( .A1(n10266), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10219) );
  NAND2_X1 U13175 ( .A1(n10221), .A2(n10220), .ZN(n10277) );
  AND2_X2 U13176 ( .A1(n9804), .A2(n10215), .ZN(n10252) );
  INV_X1 U13177 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n10224) );
  INV_X1 U13178 ( .A(n10266), .ZN(n10223) );
  NAND2_X1 U13179 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10222) );
  OAI211_X1 U13180 ( .C1(n10243), .C2(n10224), .A(n10223), .B(n10222), .ZN(
        n10225) );
  AOI21_X1 U13181 ( .B1(n10252), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10225), .ZN(
        n10236) );
  INV_X1 U13182 ( .A(n10226), .ZN(n10228) );
  AND3_X1 U13183 ( .A1(n19100), .A2(n10528), .A3(n10193), .ZN(n10227) );
  NAND2_X1 U13184 ( .A1(n10237), .A2(n13491), .ZN(n10229) );
  NAND2_X1 U13185 ( .A1(n9774), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10235) );
  NAND3_X1 U13186 ( .A1(n10232), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10231), 
        .ZN(n10233) );
  NAND2_X1 U13187 ( .A1(n10265), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10241) );
  INV_X1 U13188 ( .A(n10237), .ZN(n10239) );
  INV_X1 U13189 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13236) );
  INV_X1 U13190 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10242) );
  INV_X1 U13191 ( .A(n10245), .ZN(n10246) );
  AOI21_X2 U13192 ( .B1(n9774), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10246), .ZN(n10248) );
  NAND2_X1 U13193 ( .A1(n10275), .A2(n10274), .ZN(n10251) );
  INV_X1 U13194 ( .A(n10247), .ZN(n10249) );
  NAND2_X1 U13195 ( .A1(n10249), .A2(n10248), .ZN(n10250) );
  INV_X1 U13196 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13225) );
  INV_X1 U13197 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15057) );
  OAI22_X1 U13198 ( .A1(n10243), .A2(n13225), .B1(n19597), .B2(n15057), .ZN(
        n10253) );
  AOI21_X1 U13199 ( .B1(n10252), .B2(P2_REIP_REG_2__SCAN_IN), .A(n10253), .ZN(
        n10255) );
  OAI21_X1 U13200 ( .B1(n19696), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n19597), 
        .ZN(n10256) );
  INV_X1 U13201 ( .A(n10258), .ZN(n10257) );
  NAND2_X1 U13202 ( .A1(n10259), .A2(n10258), .ZN(n10261) );
  INV_X1 U13203 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10262) );
  INV_X1 U13204 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10598) );
  OAI22_X1 U13205 ( .A1(n12819), .A2(n10598), .B1(n19597), .B2(n16101), .ZN(
        n10263) );
  AOI21_X1 U13206 ( .B1(n10252), .B2(P2_REIP_REG_3__SCAN_IN), .A(n10263), .ZN(
        n10264) );
  NAND2_X1 U13207 ( .A1(n10265), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10268) );
  NAND2_X1 U13208 ( .A1(n10266), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10267) );
  XNOR2_X2 U13209 ( .A(n10760), .B(n10269), .ZN(n13302) );
  OR2_X2 U13210 ( .A1(n10272), .A2(n10271), .ZN(n10273) );
  AND2_X2 U13211 ( .A1(n10278), .A2(n9761), .ZN(n10290) );
  INV_X1 U13212 ( .A(n10274), .ZN(n10285) );
  XNOR2_X2 U13213 ( .A(n10277), .B(n10276), .ZN(n13005) );
  NAND2_X1 U13214 ( .A1(n10290), .A2(n10279), .ZN(n10328) );
  INV_X1 U13215 ( .A(n10328), .ZN(n19443) );
  INV_X1 U13216 ( .A(n13206), .ZN(n19064) );
  INV_X1 U13217 ( .A(n10326), .ZN(n15495) );
  AOI22_X1 U13218 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19443), .B1(
        n15495), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10284) );
  INV_X1 U13219 ( .A(n10340), .ZN(n19334) );
  NAND2_X1 U13220 ( .A1(n10288), .A2(n10280), .ZN(n10344) );
  AOI22_X1 U13221 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19334), .B1(
        n19281), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10283) );
  INV_X1 U13222 ( .A(n19167), .ZN(n10425) );
  AOI22_X1 U13223 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19090), .B1(
        n10425), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10282) );
  NAND2_X1 U13224 ( .A1(n10288), .A2(n10279), .ZN(n10341) );
  INV_X1 U13225 ( .A(n19380), .ZN(n10424) );
  AOI22_X1 U13226 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19221), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10281) );
  INV_X1 U13227 ( .A(n13005), .ZN(n18932) );
  INV_X1 U13228 ( .A(n10320), .ZN(n10431) );
  AOI22_X1 U13229 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19475), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10294) );
  AOI22_X1 U13230 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19257), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10293) );
  AND2_X2 U13231 ( .A1(n10290), .A2(n10289), .ZN(n10430) );
  AND2_X2 U13232 ( .A1(n10296), .A2(n10188), .ZN(n10354) );
  AOI22_X1 U13233 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10302) );
  AND2_X2 U13234 ( .A1(n10110), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10355) );
  AOI22_X1 U13235 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10301) );
  AND2_X2 U13236 ( .A1(n9755), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10406) );
  AOI22_X1 U13237 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10300) );
  AND2_X2 U13238 ( .A1(n14439), .A2(n10188), .ZN(n10383) );
  AND2_X2 U13239 ( .A1(n14439), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10407) );
  AOI22_X1 U13240 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10407), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10299) );
  NAND4_X1 U13241 ( .A1(n10302), .A2(n10301), .A3(n10300), .A4(n10299), .ZN(
        n10311) );
  AND2_X2 U13242 ( .A1(n9760), .A2(n10188), .ZN(n14294) );
  AOI22_X1 U13243 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10309) );
  AND2_X1 U13244 ( .A1(n9754), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10353) );
  AOI22_X1 U13245 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10308) );
  AND2_X2 U13246 ( .A1(n10304), .A2(n14277), .ZN(n10388) );
  AOI22_X1 U13247 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10307) );
  NOR2_X1 U13248 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U13249 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10306) );
  NAND4_X1 U13250 ( .A1(n10309), .A2(n10308), .A3(n10307), .A4(n10306), .ZN(
        n10310) );
  INV_X1 U13251 ( .A(n10518), .ZN(n10919) );
  NAND2_X1 U13252 ( .A1(n10919), .A2(n19737), .ZN(n10313) );
  INV_X1 U13253 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10318) );
  INV_X1 U13254 ( .A(n10314), .ZN(n10317) );
  INV_X1 U13255 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10315) );
  OAI22_X1 U13256 ( .A1(n10318), .A2(n10317), .B1(n10316), .B2(n10315), .ZN(
        n10323) );
  INV_X1 U13257 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10321) );
  INV_X1 U13258 ( .A(n10433), .ZN(n10319) );
  INV_X1 U13259 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13772) );
  OAI22_X1 U13260 ( .A1(n10321), .A2(n10320), .B1(n10319), .B2(n13772), .ZN(
        n10322) );
  NOR2_X1 U13261 ( .A1(n10323), .A2(n10322), .ZN(n10351) );
  INV_X1 U13262 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10325) );
  OAI211_X1 U13263 ( .C1(n10326), .C2(n10325), .A(n10324), .B(n10215), .ZN(
        n10331) );
  INV_X1 U13264 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10329) );
  INV_X1 U13265 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10327) );
  OAI22_X1 U13266 ( .A1(n10329), .A2(n19167), .B1(n10328), .B2(n10327), .ZN(
        n10330) );
  NOR2_X1 U13267 ( .A1(n10331), .A2(n10330), .ZN(n10350) );
  INV_X1 U13268 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10334) );
  INV_X1 U13269 ( .A(n10434), .ZN(n10333) );
  INV_X1 U13270 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10332) );
  OAI22_X1 U13271 ( .A1(n10334), .A2(n10333), .B1(n19380), .B2(n10332), .ZN(
        n10338) );
  INV_X1 U13272 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10336) );
  INV_X1 U13273 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10335) );
  OAI22_X1 U13274 ( .A1(n10336), .A2(n13678), .B1(n19254), .B2(n10335), .ZN(
        n10337) );
  NOR2_X1 U13275 ( .A1(n10338), .A2(n10337), .ZN(n10349) );
  INV_X1 U13276 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10342) );
  INV_X1 U13277 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10339) );
  OAI22_X1 U13278 ( .A1(n10342), .A2(n10341), .B1(n10340), .B2(n10339), .ZN(
        n10347) );
  INV_X1 U13279 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13211) );
  INV_X1 U13280 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10343) );
  NOR2_X1 U13281 ( .A1(n10347), .A2(n10346), .ZN(n10348) );
  NAND4_X1 U13282 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        n10396) );
  AOI22_X1 U13283 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10359) );
  AOI22_X1 U13284 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U13285 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U13286 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14294), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10356) );
  NAND4_X1 U13287 ( .A1(n10359), .A2(n10358), .A3(n10357), .A4(n10356), .ZN(
        n10366) );
  AOI22_X1 U13288 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U13289 ( .A1(n10388), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U13290 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U13291 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9707), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10361) );
  NAND4_X1 U13292 ( .A1(n10364), .A2(n10363), .A3(n10362), .A4(n10361), .ZN(
        n10365) );
  AOI22_X1 U13293 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10382), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10371) );
  AOI22_X1 U13294 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10406), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U13295 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10369) );
  AOI22_X1 U13296 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n14294), .B1(
        n10407), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10368) );
  NAND4_X1 U13297 ( .A1(n10371), .A2(n10370), .A3(n10369), .A4(n10368), .ZN(
        n10380) );
  AOI22_X1 U13298 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10372), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U13299 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n14301), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U13300 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10373), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U13301 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10360), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10375) );
  NAND4_X1 U13302 ( .A1(n10378), .A2(n10377), .A3(n10376), .A4(n10375), .ZN(
        n10379) );
  NAND2_X1 U13303 ( .A1(n19737), .A2(n10595), .ZN(n10381) );
  OR2_X1 U13304 ( .A1(n10893), .A2(n10381), .ZN(n10399) );
  AOI22_X1 U13305 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U13306 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10355), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13307 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10385) );
  AOI22_X1 U13308 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10384) );
  NAND4_X1 U13309 ( .A1(n10387), .A2(n10386), .A3(n10385), .A4(n10384), .ZN(
        n10394) );
  AOI22_X1 U13310 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10392) );
  AOI22_X1 U13311 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U13312 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U13313 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10389) );
  NAND4_X1 U13314 ( .A1(n10392), .A2(n10391), .A3(n10390), .A4(n10389), .ZN(
        n10393) );
  NAND2_X1 U13315 ( .A1(n10399), .A2(n10907), .ZN(n10395) );
  XOR2_X1 U13316 ( .A(n10907), .B(n10399), .Z(n13163) );
  OR2_X1 U13317 ( .A1(n10893), .A2(n10215), .ZN(n14254) );
  NAND2_X1 U13318 ( .A1(n14254), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14253) );
  XOR2_X1 U13319 ( .A(n10893), .B(n10595), .Z(n10400) );
  NOR2_X1 U13320 ( .A1(n14253), .A2(n10400), .ZN(n10401) );
  INV_X1 U13321 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19059) );
  XNOR2_X1 U13322 ( .A(n14253), .B(n10400), .ZN(n19058) );
  NOR2_X1 U13323 ( .A1(n19059), .A2(n19058), .ZN(n19057) );
  NOR2_X1 U13324 ( .A1(n10401), .A2(n19057), .ZN(n10402) );
  XOR2_X1 U13325 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10402), .Z(
        n13162) );
  NOR2_X1 U13326 ( .A1(n13163), .A2(n13162), .ZN(n13161) );
  INV_X1 U13327 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13172) );
  NOR2_X1 U13328 ( .A1(n10402), .A2(n13172), .ZN(n10403) );
  OR2_X1 U13329 ( .A1(n13161), .A2(n10403), .ZN(n10404) );
  NAND2_X1 U13330 ( .A1(n10404), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10405) );
  NAND2_X1 U13331 ( .A1(n16096), .A2(n10405), .ZN(n10421) );
  NAND2_X1 U13332 ( .A1(n10421), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10420) );
  AOI22_X1 U13333 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10382), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10411) );
  AOI22_X1 U13334 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n10406), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10410) );
  AOI22_X1 U13335 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U13336 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10407), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10408) );
  NAND4_X1 U13337 ( .A1(n10411), .A2(n10410), .A3(n10409), .A4(n10408), .ZN(
        n10417) );
  AOI22_X1 U13338 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n14294), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10415) );
  AOI22_X1 U13339 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n9708), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U13340 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10373), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U13341 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10360), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10412) );
  NAND4_X1 U13342 ( .A1(n10415), .A2(n10414), .A3(n10413), .A4(n10412), .ZN(
        n10416) );
  INV_X1 U13343 ( .A(n10523), .ZN(n10921) );
  INV_X1 U13344 ( .A(n10453), .ZN(n10419) );
  NAND2_X1 U13345 ( .A1(n10419), .A2(n10418), .ZN(n13741) );
  NAND2_X1 U13346 ( .A1(n10420), .A2(n13741), .ZN(n10423) );
  INV_X1 U13347 ( .A(n10421), .ZN(n13743) );
  INV_X1 U13348 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13935) );
  NAND2_X1 U13349 ( .A1(n13743), .A2(n13935), .ZN(n10422) );
  NAND2_X1 U13350 ( .A1(n10423), .A2(n10422), .ZN(n13940) );
  AOI22_X1 U13351 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19221), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U13352 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19281), .B1(
        n19334), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10428) );
  AOI22_X1 U13353 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19090), .B1(
        n10425), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U13354 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19443), .B1(
        n15495), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10426) );
  AOI22_X1 U13355 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n10314), .B1(
        n19536), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10438) );
  AOI22_X1 U13356 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n10431), .B1(
        n19475), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10437) );
  AOI22_X1 U13357 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n10432), .B1(
        n10433), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U13358 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19257), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10435) );
  AOI22_X1 U13359 ( .A1(n14293), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10406), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10442) );
  AOI22_X1 U13360 ( .A1(n10354), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10441) );
  AOI22_X1 U13361 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10355), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U13362 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10439) );
  NAND4_X1 U13363 ( .A1(n10442), .A2(n10441), .A3(n10440), .A4(n10439), .ZN(
        n10448) );
  AOI22_X1 U13364 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U13365 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10445) );
  AOI22_X1 U13366 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10444) );
  AOI22_X1 U13367 ( .A1(n10388), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10443) );
  NAND4_X1 U13368 ( .A1(n10446), .A2(n10445), .A3(n10444), .A4(n10443), .ZN(
        n10447) );
  INV_X1 U13369 ( .A(n10602), .ZN(n10449) );
  NAND2_X1 U13370 ( .A1(n10449), .A2(n19737), .ZN(n10450) );
  INV_X1 U13371 ( .A(n10452), .ZN(n10451) );
  NAND2_X1 U13372 ( .A1(n10454), .A2(n10485), .ZN(n10606) );
  INV_X1 U13373 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13936) );
  OR2_X2 U13374 ( .A1(n13940), .A2(n13941), .ZN(n13944) );
  AOI22_X1 U13375 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10314), .B1(
        n19536), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U13376 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10431), .B1(
        n19475), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U13377 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10432), .B1(
        n10433), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U13378 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19257), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10455) );
  NAND4_X1 U13379 ( .A1(n10458), .A2(n10457), .A3(n10456), .A4(n10455), .ZN(
        n10464) );
  AOI22_X1 U13380 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19221), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10462) );
  AOI22_X1 U13381 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19281), .B1(
        n19334), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10461) );
  AOI22_X1 U13382 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19090), .B1(
        n10425), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10460) );
  AOI22_X1 U13383 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19443), .B1(
        n15495), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10459) );
  NAND4_X1 U13384 ( .A1(n10462), .A2(n10461), .A3(n10460), .A4(n10459), .ZN(
        n10463) );
  AOI22_X1 U13385 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10468) );
  AOI22_X1 U13386 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10355), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10467) );
  AOI22_X1 U13387 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U13388 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10407), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10465) );
  NAND4_X1 U13389 ( .A1(n10468), .A2(n10467), .A3(n10466), .A4(n10465), .ZN(
        n10474) );
  AOI22_X1 U13390 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13391 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10471) );
  AOI22_X1 U13392 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10470) );
  AOI22_X1 U13393 ( .A1(n10388), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10469) );
  NAND4_X1 U13394 ( .A1(n10472), .A2(n10471), .A3(n10470), .A4(n10469), .ZN(
        n10473) );
  INV_X1 U13395 ( .A(n10628), .ZN(n10930) );
  NAND2_X1 U13396 ( .A1(n10930), .A2(n19737), .ZN(n10475) );
  INV_X1 U13397 ( .A(n10627), .ZN(n10478) );
  NAND2_X1 U13398 ( .A1(n10477), .A2(n10627), .ZN(n10483) );
  NAND2_X1 U13399 ( .A1(n13943), .A2(n10484), .ZN(n10482) );
  NAND2_X1 U13400 ( .A1(n14293), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10489) );
  NAND2_X1 U13401 ( .A1(n10354), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10488) );
  NAND2_X1 U13402 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10487) );
  NAND2_X1 U13403 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10486) );
  AOI22_X1 U13404 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10493) );
  AOI22_X1 U13405 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10492) );
  NAND2_X1 U13406 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10491) );
  NAND2_X1 U13407 ( .A1(n14264), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10490) );
  NAND2_X1 U13408 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10497) );
  NAND2_X1 U13409 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10496) );
  NAND2_X1 U13410 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10495) );
  NAND2_X1 U13411 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10494) );
  AOI22_X1 U13412 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10498) );
  NAND4_X1 U13413 ( .A1(n10501), .A2(n10500), .A3(n10499), .A4(n10498), .ZN(
        n10632) );
  INV_X1 U13414 ( .A(n10632), .ZN(n10934) );
  INV_X1 U13415 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10871) );
  NAND2_X1 U13416 ( .A1(n14022), .A2(n10871), .ZN(n10502) );
  NAND2_X1 U13417 ( .A1(n14021), .A2(n10502), .ZN(n10505) );
  INV_X1 U13418 ( .A(n14022), .ZN(n10503) );
  NAND2_X1 U13419 ( .A1(n10503), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10504) );
  NAND2_X1 U13420 ( .A1(n10508), .A2(n14238), .ZN(n10507) );
  XNOR2_X1 U13421 ( .A(n10507), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16067) );
  NAND2_X1 U13422 ( .A1(n16066), .A2(n16067), .ZN(n10510) );
  NAND3_X1 U13423 ( .A1(n10508), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n14238), .ZN(n10509) );
  INV_X1 U13424 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16114) );
  NAND2_X1 U13425 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15379) );
  INV_X1 U13426 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15376) );
  INV_X1 U13427 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15344) );
  INV_X1 U13428 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15337) );
  INV_X1 U13429 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15363) );
  NOR3_X1 U13430 ( .A1(n15344), .A2(n15337), .A3(n15363), .ZN(n12337) );
  AND4_X1 U13431 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(n12337), .ZN(n12867) );
  NAND2_X1 U13432 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11090) );
  INV_X1 U13433 ( .A(n11090), .ZN(n15287) );
  NAND2_X1 U13434 ( .A1(n15303), .A2(n15287), .ZN(n15214) );
  NOR2_X1 U13435 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19616) );
  AOI211_X1 U13436 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n19616), .ZN(n13014) );
  INV_X1 U13437 ( .A(n13014), .ZN(n19739) );
  NAND2_X1 U13438 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19726) );
  INV_X1 U13439 ( .A(n19726), .ZN(n19733) );
  NOR2_X1 U13440 ( .A1(n19739), .A2(n19733), .ZN(n13492) );
  NAND2_X1 U13441 ( .A1(n10857), .A2(n13492), .ZN(n10591) );
  XNOR2_X1 U13442 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10548) );
  NAND2_X1 U13443 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19715), .ZN(
        n10529) );
  INV_X1 U13444 ( .A(n10529), .ZN(n10512) );
  NAND2_X1 U13445 ( .A1(n10548), .A2(n10512), .ZN(n10514) );
  NAND2_X1 U13446 ( .A1(n19708), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10513) );
  NAND2_X1 U13447 ( .A1(n10514), .A2(n10513), .ZN(n10526) );
  XNOR2_X1 U13448 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10524) );
  NAND2_X1 U13449 ( .A1(n10526), .A2(n10524), .ZN(n10516) );
  NAND2_X1 U13450 ( .A1(n19696), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10515) );
  NAND2_X1 U13451 ( .A1(n10516), .A2(n10515), .ZN(n10520) );
  XNOR2_X1 U13452 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10519) );
  INV_X1 U13453 ( .A(n10519), .ZN(n10517) );
  XNOR2_X1 U13454 ( .A(n10520), .B(n10517), .ZN(n10568) );
  MUX2_X1 U13455 ( .A(n10518), .B(n10568), .S(n10551), .Z(n10599) );
  NAND2_X1 U13456 ( .A1(n10520), .A2(n10519), .ZN(n10522) );
  NAND2_X1 U13457 ( .A1(n19689), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10521) );
  NAND2_X1 U13458 ( .A1(n10522), .A2(n10521), .ZN(n10540) );
  MUX2_X1 U13459 ( .A(n10523), .B(n10566), .S(n10551), .Z(n10600) );
  AND2_X1 U13460 ( .A1(n10599), .A2(n10600), .ZN(n10553) );
  INV_X1 U13461 ( .A(n10524), .ZN(n10525) );
  XNOR2_X1 U13462 ( .A(n10526), .B(n10525), .ZN(n10567) );
  INV_X1 U13463 ( .A(n10567), .ZN(n10549) );
  INV_X1 U13464 ( .A(n10548), .ZN(n10527) );
  OAI21_X1 U13465 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19715), .A(
        n10529), .ZN(n10580) );
  OAI21_X1 U13466 ( .B1(n10527), .B2(n10580), .A(n12783), .ZN(n10532) );
  INV_X1 U13467 ( .A(n10580), .ZN(n10530) );
  XNOR2_X1 U13468 ( .A(n10548), .B(n10529), .ZN(n10570) );
  OAI211_X1 U13469 ( .C1(n10215), .C2(n10530), .A(n10528), .B(n10570), .ZN(
        n10531) );
  OAI211_X1 U13470 ( .C1(n10533), .C2(n10549), .A(n10532), .B(n10531), .ZN(
        n10534) );
  INV_X1 U13471 ( .A(n10534), .ZN(n10537) );
  NOR2_X1 U13472 ( .A1(n9776), .A2(n19737), .ZN(n10535) );
  MUX2_X1 U13473 ( .A(n10535), .B(n12783), .S(n10567), .Z(n10536) );
  OAI21_X1 U13474 ( .B1(n10537), .B2(n10536), .A(n10568), .ZN(n10538) );
  OAI21_X1 U13475 ( .B1(n10553), .B2(n12783), .A(n10538), .ZN(n10545) );
  INV_X1 U13476 ( .A(n10566), .ZN(n10543) );
  AND2_X1 U13477 ( .A1(n16204), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10539) );
  NAND2_X1 U13478 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16201), .ZN(
        n10541) );
  AOI21_X1 U13479 ( .B1(n12783), .B2(n10543), .A(n10572), .ZN(n10544) );
  NAND2_X1 U13480 ( .A1(n10545), .A2(n10544), .ZN(n10546) );
  MUX2_X1 U13481 ( .A(n10546), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19727), .Z(n10587) );
  NAND2_X1 U13482 ( .A1(n16187), .A2(n10215), .ZN(n13495) );
  MUX2_X1 U13483 ( .A(n10893), .B(n10580), .S(n10551), .Z(n10610) );
  NAND2_X1 U13484 ( .A1(n10551), .A2(n10549), .ZN(n10550) );
  OAI21_X1 U13485 ( .B1(n10610), .B2(n10527), .A(n10594), .ZN(n10554) );
  AOI21_X1 U13486 ( .B1(n10554), .B2(n10553), .A(n10572), .ZN(n19717) );
  AND2_X1 U13487 ( .A1(n19737), .A2(n10216), .ZN(n12798) );
  AND2_X1 U13488 ( .A1(n16189), .A2(n12798), .ZN(n19720) );
  NAND2_X1 U13489 ( .A1(n19717), .A2(n19720), .ZN(n11077) );
  NAND2_X1 U13490 ( .A1(n10555), .A2(n13724), .ZN(n10556) );
  NAND2_X1 U13491 ( .A1(n13491), .A2(n10556), .ZN(n10565) );
  NAND2_X1 U13492 ( .A1(n10557), .A2(n19737), .ZN(n10869) );
  OAI21_X1 U13493 ( .B1(n10528), .B2(n10558), .A(n13724), .ZN(n10559) );
  INV_X1 U13494 ( .A(n10559), .ZN(n10560) );
  AOI21_X1 U13495 ( .B1(n10869), .B2(n10560), .A(n10851), .ZN(n10564) );
  NAND2_X1 U13496 ( .A1(n10561), .A2(n10203), .ZN(n10562) );
  NAND2_X1 U13497 ( .A1(n10562), .A2(n12798), .ZN(n10860) );
  NAND4_X1 U13498 ( .A1(n10565), .A2(n10564), .A3(n10563), .A4(n10860), .ZN(
        n10870) );
  NAND3_X1 U13499 ( .A1(n10568), .A2(n10567), .A3(n10566), .ZN(n10579) );
  INV_X1 U13500 ( .A(n10579), .ZN(n10569) );
  AND3_X1 U13501 ( .A1(n16207), .A2(n16183), .A3(n13492), .ZN(n10573) );
  NOR2_X1 U13502 ( .A1(n10870), .A2(n10573), .ZN(n13493) );
  MUX2_X1 U13503 ( .A(n16207), .B(n10857), .S(n19737), .Z(n10574) );
  NAND3_X1 U13504 ( .A1(n10574), .A2(n16183), .A3(n19726), .ZN(n10585) );
  NAND2_X1 U13505 ( .A1(n10575), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10576) );
  NAND2_X1 U13506 ( .A1(n10576), .A2(n16201), .ZN(n16193) );
  INV_X1 U13507 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n10577) );
  OAI21_X1 U13508 ( .B1(n10406), .B2(n16193), .A(n10577), .ZN(n10578) );
  NAND2_X1 U13509 ( .A1(n10578), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19709) );
  OAI21_X1 U13510 ( .B1(n10580), .B2(n10579), .A(n16183), .ZN(n10581) );
  INV_X1 U13511 ( .A(n10581), .ZN(n10582) );
  NAND2_X1 U13512 ( .A1(n19597), .A2(n10582), .ZN(n10583) );
  NAND2_X1 U13513 ( .A1(n19709), .A2(n10583), .ZN(n16211) );
  NAND3_X1 U13514 ( .A1(n16189), .A2(n10215), .A3(n16211), .ZN(n10584) );
  AND3_X1 U13515 ( .A1(n13493), .A2(n10585), .A3(n10584), .ZN(n10586) );
  AND2_X1 U13516 ( .A1(n11077), .A2(n10586), .ZN(n10590) );
  AOI21_X1 U13517 ( .B1(n10587), .B2(n10528), .A(n10195), .ZN(n10588) );
  NAND2_X1 U13518 ( .A1(n13495), .A2(n10588), .ZN(n10589) );
  OAI211_X1 U13519 ( .C1(n10591), .C2(n13495), .A(n10590), .B(n10589), .ZN(
        n10593) );
  NAND2_X1 U13520 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19597), .ZN(n12786) );
  INV_X1 U13521 ( .A(n12786), .ZN(n10592) );
  NOR2_X1 U13522 ( .A1(n11079), .A2(n19074), .ZN(n11075) );
  NAND2_X1 U13523 ( .A1(n13236), .A2(n10224), .ZN(n10597) );
  MUX2_X1 U13524 ( .A(n10900), .B(n10597), .S(n10596), .Z(n10613) );
  NOR2_X2 U13525 ( .A1(n10614), .A2(n10613), .ZN(n10609) );
  MUX2_X1 U13526 ( .A(n10599), .B(n10598), .S(n9757), .Z(n10608) );
  NAND2_X1 U13527 ( .A1(n10609), .A2(n10608), .ZN(n10607) );
  INV_X1 U13528 ( .A(n10600), .ZN(n10601) );
  MUX2_X1 U13529 ( .A(n10601), .B(P2_EBX_REG_4__SCAN_IN), .S(n9757), .Z(n10619) );
  NOR2_X2 U13530 ( .A1(n10607), .A2(n10619), .ZN(n10604) );
  NAND2_X1 U13531 ( .A1(n10602), .A2(n9764), .ZN(n10925) );
  AND2_X2 U13532 ( .A1(n10604), .A2(n10603), .ZN(n10631) );
  NOR2_X1 U13533 ( .A1(n10604), .A2(n10603), .ZN(n10605) );
  OR2_X1 U13534 ( .A1(n10631), .A2(n10605), .ZN(n18909) );
  XNOR2_X1 U13535 ( .A(n10624), .B(n13936), .ZN(n13930) );
  OAI21_X1 U13536 ( .B1(n10609), .B2(n10608), .A(n10620), .ZN(n13623) );
  MUX2_X1 U13537 ( .A(n10610), .B(n10224), .S(n9757), .Z(n18926) );
  INV_X1 U13538 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14251) );
  OR2_X1 U13539 ( .A1(n18926), .A2(n14251), .ZN(n19052) );
  NAND3_X1 U13540 ( .A1(n9757), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10611) );
  NAND2_X1 U13541 ( .A1(n10613), .A2(n10611), .ZN(n19053) );
  NOR2_X1 U13542 ( .A1(n19052), .A2(n19053), .ZN(n10612) );
  NAND2_X1 U13543 ( .A1(n19052), .A2(n19053), .ZN(n19051) );
  OAI21_X1 U13544 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10612), .A(
        n19051), .ZN(n13165) );
  XNOR2_X1 U13545 ( .A(n10614), .B(n10613), .ZN(n10615) );
  XNOR2_X1 U13546 ( .A(n10615), .B(n13172), .ZN(n13164) );
  OR2_X1 U13547 ( .A1(n13165), .A2(n13164), .ZN(n13178) );
  INV_X1 U13548 ( .A(n10615), .ZN(n15054) );
  NAND2_X1 U13549 ( .A1(n15054), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10616) );
  NAND2_X1 U13550 ( .A1(n13178), .A2(n10616), .ZN(n16091) );
  OAI21_X1 U13551 ( .B1(n16093), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n16091), .ZN(n10618) );
  NAND2_X1 U13552 ( .A1(n16093), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10617) );
  NAND2_X1 U13553 ( .A1(n10618), .A2(n10617), .ZN(n13739) );
  XNOR2_X1 U13554 ( .A(n10620), .B(n10619), .ZN(n10621) );
  XNOR2_X1 U13555 ( .A(n10621), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13740) );
  NAND2_X1 U13556 ( .A1(n13739), .A2(n13740), .ZN(n10623) );
  INV_X1 U13557 ( .A(n10621), .ZN(n13821) );
  NAND2_X1 U13558 ( .A1(n13821), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10622) );
  NAND2_X1 U13559 ( .A1(n10623), .A2(n10622), .ZN(n13931) );
  NAND2_X1 U13560 ( .A1(n13930), .A2(n13931), .ZN(n10626) );
  NAND2_X1 U13561 ( .A1(n10624), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10625) );
  NAND2_X1 U13562 ( .A1(n10626), .A2(n10625), .ZN(n13966) );
  NAND2_X1 U13563 ( .A1(n10627), .A2(n10934), .ZN(n10629) );
  INV_X1 U13564 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n10769) );
  MUX2_X1 U13565 ( .A(n10769), .B(n10628), .S(n9764), .Z(n10630) );
  XNOR2_X1 U13566 ( .A(n10631), .B(n10630), .ZN(n18893) );
  NAND2_X1 U13567 ( .A1(n10629), .A2(n18893), .ZN(n10634) );
  INV_X1 U13568 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13978) );
  XNOR2_X1 U13569 ( .A(n10634), .B(n13978), .ZN(n13967) );
  AND2_X2 U13570 ( .A1(n10631), .A2(n10630), .ZN(n10637) );
  INV_X1 U13571 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13409) );
  MUX2_X1 U13572 ( .A(n13409), .B(n10632), .S(n9763), .Z(n10636) );
  INV_X1 U13573 ( .A(n10636), .ZN(n10633) );
  XNOR2_X1 U13574 ( .A(n10637), .B(n10633), .ZN(n18886) );
  AND2_X1 U13575 ( .A1(n18886), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14029) );
  INV_X1 U13576 ( .A(n14029), .ZN(n10635) );
  NAND2_X1 U13577 ( .A1(n10634), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14027) );
  NAND3_X1 U13578 ( .A1(n10638), .A2(n9757), .A3(P2_EBX_REG_8__SCAN_IN), .ZN(
        n10640) );
  OR2_X1 U13579 ( .A1(n10638), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10639) );
  AND3_X1 U13580 ( .A1(n10689), .A2(n10640), .A3(n10639), .ZN(n13797) );
  NAND2_X1 U13581 ( .A1(n13797), .A2(n14238), .ZN(n10644) );
  INV_X1 U13582 ( .A(n10644), .ZN(n10641) );
  INV_X1 U13583 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10643) );
  NAND2_X1 U13584 ( .A1(n10644), .A2(n10643), .ZN(n16070) );
  INV_X1 U13585 ( .A(n18886), .ZN(n10645) );
  NAND2_X1 U13586 ( .A1(n10645), .A2(n10871), .ZN(n16069) );
  AND2_X1 U13587 ( .A1(n16070), .A2(n16069), .ZN(n10646) );
  NAND2_X1 U13588 ( .A1(n9757), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10649) );
  INV_X1 U13589 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n13426) );
  NOR2_X1 U13590 ( .A1(n9764), .A2(n13426), .ZN(n10647) );
  OR2_X2 U13591 ( .A1(n10648), .A2(n10647), .ZN(n10650) );
  MUX2_X1 U13592 ( .A(n9757), .B(n10649), .S(n10650), .Z(n10652) );
  INV_X1 U13593 ( .A(n10655), .ZN(n10651) );
  AOI21_X1 U13594 ( .B1(n18865), .B2(n14238), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16047) );
  NAND2_X1 U13595 ( .A1(n9757), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10653) );
  MUX2_X1 U13596 ( .A(n10653), .B(P2_EBX_REG_10__SCAN_IN), .S(n10655), .Z(
        n10654) );
  NAND2_X1 U13597 ( .A1(n10654), .A2(n10689), .ZN(n13781) );
  AND2_X1 U13598 ( .A1(n10663), .A2(n16114), .ZN(n16052) );
  OR2_X1 U13599 ( .A1(n16047), .A2(n16052), .ZN(n15416) );
  INV_X1 U13600 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n18964) );
  NAND2_X1 U13601 ( .A1(n9757), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10656) );
  OR2_X1 U13602 ( .A1(n10657), .A2(n10656), .ZN(n10659) );
  INV_X1 U13603 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13541) );
  NAND2_X2 U13604 ( .A1(n10667), .A2(n10689), .ZN(n10665) );
  INV_X1 U13605 ( .A(n10665), .ZN(n10658) );
  NAND2_X1 U13606 ( .A1(n10659), .A2(n10658), .ZN(n12987) );
  INV_X1 U13607 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15427) );
  OAI21_X1 U13608 ( .B1(n12987), .B2(n10934), .A(n15427), .ZN(n15420) );
  INV_X1 U13609 ( .A(n15420), .ZN(n10660) );
  INV_X1 U13610 ( .A(n12987), .ZN(n10662) );
  AND2_X1 U13611 ( .A1(n14238), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10661) );
  NAND2_X1 U13612 ( .A1(n10662), .A2(n10661), .ZN(n15419) );
  NAND3_X1 U13613 ( .A1(n18865), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n14238), .ZN(n16048) );
  OR2_X1 U13614 ( .A1(n16114), .A2(n10663), .ZN(n16050) );
  NAND2_X1 U13615 ( .A1(n16048), .A2(n16050), .ZN(n15417) );
  INV_X1 U13616 ( .A(n15417), .ZN(n10664) );
  AND2_X1 U13617 ( .A1(n15419), .A2(n10664), .ZN(n12322) );
  NAND2_X1 U13618 ( .A1(n12324), .A2(n12322), .ZN(n15395) );
  NAND2_X1 U13619 ( .A1(n9757), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10666) );
  NAND2_X2 U13620 ( .A1(n10665), .A2(n10666), .ZN(n10694) );
  INV_X1 U13621 ( .A(n10666), .ZN(n10668) );
  NAND2_X1 U13622 ( .A1(n10668), .A2(n10667), .ZN(n10669) );
  NAND2_X1 U13623 ( .A1(n10694), .A2(n10669), .ZN(n13809) );
  NAND2_X1 U13624 ( .A1(n14238), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10670) );
  NOR2_X1 U13625 ( .A1(n13809), .A2(n10670), .ZN(n16028) );
  INV_X1 U13626 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10799) );
  NOR2_X1 U13627 ( .A1(n9763), .A2(n10799), .ZN(n10693) );
  NAND2_X1 U13628 ( .A1(n9757), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10697) );
  NAND2_X1 U13629 ( .A1(n10692), .A2(n10697), .ZN(n10684) );
  INV_X1 U13630 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10810) );
  NOR2_X1 U13631 ( .A1(n9764), .A2(n10810), .ZN(n10685) );
  NOR2_X2 U13632 ( .A1(n10684), .A2(n10685), .ZN(n10683) );
  INV_X1 U13633 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n18947) );
  NAND2_X1 U13634 ( .A1(n10683), .A2(n10064), .ZN(n10703) );
  INV_X1 U13635 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10820) );
  NOR2_X1 U13636 ( .A1(n9763), .A2(n10820), .ZN(n10702) );
  NOR2_X2 U13637 ( .A1(n10703), .A2(n10702), .ZN(n10680) );
  INV_X1 U13638 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n15987) );
  INV_X1 U13639 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10671) );
  NAND2_X1 U13640 ( .A1(n15987), .A2(n10671), .ZN(n10672) );
  NAND2_X1 U13641 ( .A1(n9757), .A2(n10672), .ZN(n10673) );
  INV_X1 U13642 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n15983) );
  INV_X1 U13643 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10835) );
  NOR2_X1 U13644 ( .A1(n9763), .A2(n10835), .ZN(n10676) );
  AOI21_X1 U13645 ( .B1(n10709), .B2(n10676), .A(n11100), .ZN(n10677) );
  NAND2_X1 U13646 ( .A1(n10740), .A2(n10677), .ZN(n18781) );
  INV_X1 U13647 ( .A(n18781), .ZN(n10678) );
  NAND2_X1 U13648 ( .A1(n10678), .A2(n14238), .ZN(n10721) );
  INV_X1 U13649 ( .A(n10721), .ZN(n10679) );
  NAND2_X1 U13650 ( .A1(n10679), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14203) );
  INV_X1 U13651 ( .A(n10680), .ZN(n10713) );
  NOR2_X1 U13652 ( .A1(n9764), .A2(n10671), .ZN(n10681) );
  NAND2_X1 U13653 ( .A1(n10714), .A2(n10681), .ZN(n10682) );
  NAND2_X1 U13654 ( .A1(n10682), .A2(n10707), .ZN(n18796) );
  INV_X1 U13655 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15317) );
  NAND2_X1 U13656 ( .A1(n10701), .A2(n10685), .ZN(n10686) );
  NAND2_X1 U13657 ( .A1(n10690), .A2(n10686), .ZN(n18835) );
  INV_X1 U13658 ( .A(n10727), .ZN(n10687) );
  NAND2_X1 U13659 ( .A1(n10687), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15355) );
  NAND3_X1 U13660 ( .A1(n10690), .A2(n9757), .A3(P2_EBX_REG_16__SCAN_IN), .ZN(
        n10688) );
  OAI211_X1 U13661 ( .C1(n10690), .C2(P2_EBX_REG_16__SCAN_IN), .A(n10689), .B(
        n10688), .ZN(n13856) );
  NAND2_X1 U13662 ( .A1(n14238), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10691) );
  OR2_X1 U13663 ( .A1(n13856), .A2(n10691), .ZN(n12329) );
  INV_X1 U13664 ( .A(n10692), .ZN(n10699) );
  NAND2_X1 U13665 ( .A1(n10694), .A2(n10693), .ZN(n10695) );
  NAND2_X1 U13666 ( .A1(n10699), .A2(n10695), .ZN(n18854) );
  NAND2_X1 U13667 ( .A1(n14238), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10696) );
  OR2_X1 U13668 ( .A1(n18854), .A2(n10696), .ZN(n15398) );
  INV_X1 U13669 ( .A(n10697), .ZN(n10698) );
  NAND2_X1 U13670 ( .A1(n10699), .A2(n10698), .ZN(n10700) );
  NAND2_X1 U13671 ( .A1(n10701), .A2(n10700), .ZN(n18847) );
  AND4_X1 U13672 ( .A1(n15355), .A2(n12329), .A3(n15398), .A4(n15372), .ZN(
        n10706) );
  NAND2_X1 U13673 ( .A1(n10703), .A2(n10702), .ZN(n10704) );
  NAND2_X1 U13674 ( .A1(n10713), .A2(n10704), .ZN(n18819) );
  NAND2_X1 U13675 ( .A1(n14238), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10705) );
  OR2_X1 U13676 ( .A1(n18819), .A2(n10705), .ZN(n12330) );
  NAND2_X1 U13677 ( .A1(n9757), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10708) );
  MUX2_X1 U13678 ( .A(n9757), .B(n10708), .S(n10707), .Z(n10710) );
  NAND2_X1 U13679 ( .A1(n10710), .A2(n10709), .ZN(n14101) );
  INV_X1 U13680 ( .A(n10722), .ZN(n10711) );
  NAND2_X1 U13681 ( .A1(n10713), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10712) );
  INV_X1 U13682 ( .A(n10719), .ZN(n10716) );
  NAND2_X1 U13683 ( .A1(n10716), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12722) );
  NAND4_X1 U13684 ( .A1(n14203), .A2(n10069), .A3(n14209), .A4(n12722), .ZN(
        n10735) );
  INV_X1 U13685 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n20857) );
  NAND2_X1 U13686 ( .A1(n10719), .A2(n20857), .ZN(n12332) );
  OR2_X1 U13687 ( .A1(n18796), .A2(n10934), .ZN(n10720) );
  NAND2_X1 U13688 ( .A1(n10720), .A2(n15317), .ZN(n12721) );
  AND2_X1 U13689 ( .A1(n12332), .A2(n12721), .ZN(n14204) );
  INV_X1 U13690 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10875) );
  NAND2_X1 U13691 ( .A1(n10721), .A2(n10875), .ZN(n14202) );
  INV_X1 U13692 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15318) );
  NAND2_X1 U13693 ( .A1(n10722), .A2(n15318), .ZN(n14208) );
  NAND2_X1 U13694 ( .A1(n10723), .A2(n15344), .ZN(n12331) );
  OR2_X1 U13695 ( .A1(n13856), .A2(n10934), .ZN(n10724) );
  XNOR2_X1 U13696 ( .A(n10724), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12328) );
  NAND2_X1 U13697 ( .A1(n10725), .A2(n15376), .ZN(n15371) );
  OR2_X1 U13698 ( .A1(n18854), .A2(n10934), .ZN(n10726) );
  INV_X1 U13699 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15409) );
  NAND2_X1 U13700 ( .A1(n10726), .A2(n15409), .ZN(n15399) );
  AND2_X1 U13701 ( .A1(n15371), .A2(n15399), .ZN(n10728) );
  NAND2_X1 U13702 ( .A1(n10727), .A2(n15363), .ZN(n15354) );
  AND4_X1 U13703 ( .A1(n12331), .A2(n12328), .A3(n10728), .A4(n15354), .ZN(
        n10729) );
  AND2_X1 U13704 ( .A1(n14208), .A2(n10729), .ZN(n10730) );
  AND3_X1 U13705 ( .A1(n14204), .A2(n14202), .A3(n10730), .ZN(n10733) );
  OR2_X1 U13706 ( .A1(n13809), .A2(n10934), .ZN(n10732) );
  INV_X1 U13707 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10731) );
  NAND2_X1 U13708 ( .A1(n10732), .A2(n10731), .ZN(n15396) );
  AND2_X1 U13709 ( .A1(n10733), .A2(n15396), .ZN(n10734) );
  OR2_X2 U13710 ( .A1(n10735), .A2(n10734), .ZN(n10736) );
  NAND2_X1 U13711 ( .A1(n10740), .A2(n10689), .ZN(n10737) );
  NAND2_X1 U13712 ( .A1(n9757), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10738) );
  INV_X1 U13713 ( .A(n10738), .ZN(n10739) );
  NAND2_X1 U13714 ( .A1(n10740), .A2(n10739), .ZN(n10741) );
  NAND2_X1 U13715 ( .A1(n10744), .A2(n10741), .ZN(n15540) );
  OR2_X1 U13716 ( .A1(n15540), .A2(n10934), .ZN(n10742) );
  INV_X1 U13717 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n20973) );
  INV_X1 U13718 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10747) );
  NOR2_X1 U13719 ( .A1(n9764), .A2(n10747), .ZN(n10743) );
  OR2_X2 U13720 ( .A1(n10744), .A2(n10743), .ZN(n11096) );
  NAND2_X1 U13721 ( .A1(n10744), .A2(n10743), .ZN(n10745) );
  NAND2_X1 U13722 ( .A1(n11096), .A2(n10745), .ZN(n12974) );
  XNOR2_X1 U13723 ( .A(n10746), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11094) );
  XNOR2_X1 U13724 ( .A(n11095), .B(n11094), .ZN(n11087) );
  AND2_X1 U13725 ( .A1(n16189), .A2(n12783), .ZN(n19719) );
  NAND2_X1 U13726 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10750) );
  INV_X1 U13727 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12973) );
  OAI22_X1 U13728 ( .A1(n12819), .A2(n10747), .B1(n19597), .B2(n12973), .ZN(
        n10748) );
  AOI21_X1 U13729 ( .B1(n14129), .B2(P2_REIP_REG_23__SCAN_IN), .A(n10748), 
        .ZN(n10749) );
  NAND2_X1 U13730 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10755) );
  INV_X1 U13731 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n10752) );
  INV_X1 U13732 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10751) );
  OAI22_X1 U13733 ( .A1(n12819), .A2(n10752), .B1(n19597), .B2(n10751), .ZN(
        n10753) );
  AOI21_X1 U13734 ( .B1(n10252), .B2(P2_REIP_REG_4__SCAN_IN), .A(n10753), .ZN(
        n10754) );
  INV_X1 U13735 ( .A(n10756), .ZN(n10758) );
  NAND2_X1 U13736 ( .A1(n10758), .A2(n10757), .ZN(n13744) );
  INV_X1 U13737 ( .A(n13744), .ZN(n10759) );
  NOR2_X1 U13738 ( .A1(n13746), .A2(n10759), .ZN(n10762) );
  INV_X1 U13739 ( .A(n13749), .ZN(n10768) );
  NAND2_X1 U13740 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10766) );
  INV_X1 U13741 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n18907) );
  INV_X1 U13742 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10763) );
  OAI22_X1 U13743 ( .A1(n12819), .A2(n18907), .B1(n19597), .B2(n10763), .ZN(
        n10764) );
  AOI21_X1 U13744 ( .B1(n14129), .B2(P2_REIP_REG_5__SCAN_IN), .A(n10764), .ZN(
        n10765) );
  NAND2_X1 U13745 ( .A1(n10768), .A2(n10767), .ZN(n13338) );
  NAND2_X1 U13746 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10772) );
  OAI22_X1 U13747 ( .A1(n12819), .A2(n10769), .B1(n19597), .B2(n9871), .ZN(
        n10770) );
  AOI21_X1 U13748 ( .B1(n14129), .B2(P2_REIP_REG_6__SCAN_IN), .A(n10770), .ZN(
        n10771) );
  NAND2_X1 U13749 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10775) );
  OAI22_X1 U13750 ( .A1(n12819), .A2(n13409), .B1(n19597), .B2(n14032), .ZN(
        n10773) );
  AOI21_X1 U13751 ( .B1(n14129), .B2(P2_REIP_REG_7__SCAN_IN), .A(n10773), .ZN(
        n10774) );
  NAND2_X1 U13752 ( .A1(n10775), .A2(n10774), .ZN(n13407) );
  NAND2_X1 U13753 ( .A1(n13348), .A2(n13407), .ZN(n13406) );
  NAND2_X1 U13754 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10779) );
  INV_X1 U13755 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10776) );
  OAI22_X1 U13756 ( .A1(n12819), .A2(n13426), .B1(n19597), .B2(n10776), .ZN(
        n10777) );
  AOI21_X1 U13757 ( .B1(n10252), .B2(P2_REIP_REG_8__SCAN_IN), .A(n10777), .ZN(
        n10778) );
  NAND2_X1 U13758 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10785) );
  INV_X1 U13759 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10782) );
  INV_X1 U13760 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10781) );
  OAI22_X1 U13761 ( .A1(n12819), .A2(n10782), .B1(n19597), .B2(n10781), .ZN(
        n10783) );
  AOI21_X1 U13762 ( .B1(n10252), .B2(P2_REIP_REG_9__SCAN_IN), .A(n10783), .ZN(
        n10784) );
  NAND2_X1 U13763 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10788) );
  INV_X1 U13764 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13780) );
  OAI22_X1 U13765 ( .A1(n12819), .A2(n18964), .B1(n19597), .B2(n13780), .ZN(
        n10786) );
  AOI21_X1 U13766 ( .B1(n10252), .B2(P2_REIP_REG_10__SCAN_IN), .A(n10786), 
        .ZN(n10787) );
  NAND2_X1 U13767 ( .A1(n10788), .A2(n10787), .ZN(n13778) );
  NAND2_X1 U13768 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10792) );
  INV_X1 U13769 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10789) );
  OAI22_X1 U13770 ( .A1(n12819), .A2(n13541), .B1(n19597), .B2(n10789), .ZN(
        n10790) );
  AOI21_X1 U13771 ( .B1(n10252), .B2(P2_REIP_REG_11__SCAN_IN), .A(n10790), 
        .ZN(n10791) );
  NAND2_X1 U13772 ( .A1(n10792), .A2(n10791), .ZN(n12990) );
  NAND2_X1 U13773 ( .A1(n12988), .A2(n12990), .ZN(n12989) );
  NAND2_X1 U13774 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10796) );
  INV_X1 U13775 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n10793) );
  OAI22_X1 U13776 ( .A1(n12819), .A2(n10793), .B1(n19597), .B2(n9875), .ZN(
        n10794) );
  AOI21_X1 U13777 ( .B1(n10252), .B2(P2_REIP_REG_12__SCAN_IN), .A(n10794), 
        .ZN(n10795) );
  NAND2_X1 U13778 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10802) );
  OAI22_X1 U13779 ( .A1(n12819), .A2(n10799), .B1(n19597), .B2(n18853), .ZN(
        n10800) );
  AOI21_X1 U13780 ( .B1(n10252), .B2(P2_REIP_REG_13__SCAN_IN), .A(n10800), 
        .ZN(n10801) );
  NAND2_X1 U13781 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10808) );
  INV_X1 U13782 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n10805) );
  INV_X1 U13783 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10804) );
  OAI22_X1 U13784 ( .A1(n12819), .A2(n10805), .B1(n19597), .B2(n10804), .ZN(
        n10806) );
  AOI21_X1 U13785 ( .B1(n10252), .B2(P2_REIP_REG_14__SCAN_IN), .A(n10806), 
        .ZN(n10807) );
  NAND2_X1 U13786 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10813) );
  INV_X1 U13787 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10809) );
  OAI22_X1 U13788 ( .A1(n12819), .A2(n10810), .B1(n19597), .B2(n10809), .ZN(
        n10811) );
  AOI21_X1 U13789 ( .B1(n10252), .B2(P2_REIP_REG_15__SCAN_IN), .A(n10811), 
        .ZN(n10812) );
  NAND2_X1 U13790 ( .A1(n10813), .A2(n10812), .ZN(n13733) );
  NAND2_X1 U13791 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10817) );
  INV_X1 U13792 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10814) );
  OAI22_X1 U13793 ( .A1(n12819), .A2(n18947), .B1(n19597), .B2(n10814), .ZN(
        n10815) );
  AOI21_X1 U13794 ( .B1(n10252), .B2(P2_REIP_REG_16__SCAN_IN), .A(n10815), 
        .ZN(n10816) );
  NAND2_X1 U13795 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10823) );
  INV_X1 U13796 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15233) );
  OAI22_X1 U13797 ( .A1(n12819), .A2(n10820), .B1(n19597), .B2(n15233), .ZN(
        n10821) );
  AOI21_X1 U13798 ( .B1(n10252), .B2(P2_REIP_REG_17__SCAN_IN), .A(n10821), 
        .ZN(n10822) );
  NAND2_X1 U13799 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10827) );
  INV_X1 U13800 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10824) );
  OAI22_X1 U13801 ( .A1(n12819), .A2(n15987), .B1(n19597), .B2(n10824), .ZN(
        n10825) );
  AOI21_X1 U13802 ( .B1(n10252), .B2(P2_REIP_REG_18__SCAN_IN), .A(n10825), 
        .ZN(n10826) );
  NAND2_X1 U13803 ( .A1(n10827), .A2(n10826), .ZN(n12335) );
  NAND2_X1 U13804 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10830) );
  INV_X1 U13805 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18795) );
  OAI22_X1 U13806 ( .A1(n12819), .A2(n10671), .B1(n19597), .B2(n18795), .ZN(
        n10828) );
  AOI21_X1 U13807 ( .B1(n10252), .B2(P2_REIP_REG_19__SCAN_IN), .A(n10828), 
        .ZN(n10829) );
  NAND2_X1 U13808 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10833) );
  OAI22_X1 U13809 ( .A1(n12819), .A2(n15983), .B1(n19597), .B2(n9862), .ZN(
        n10831) );
  AOI21_X1 U13810 ( .B1(n14129), .B2(P2_REIP_REG_20__SCAN_IN), .A(n10831), 
        .ZN(n10832) );
  INV_X1 U13811 ( .A(n14094), .ZN(n10834) );
  NAND2_X1 U13812 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10838) );
  INV_X1 U13813 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18778) );
  OAI22_X1 U13814 ( .A1(n12819), .A2(n10835), .B1(n19597), .B2(n18778), .ZN(
        n10836) );
  AOI21_X1 U13815 ( .B1(n14129), .B2(P2_REIP_REG_21__SCAN_IN), .A(n10836), 
        .ZN(n10837) );
  NAND2_X1 U13816 ( .A1(n10838), .A2(n10837), .ZN(n14085) );
  NAND2_X1 U13817 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10842) );
  INV_X1 U13818 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n10839) );
  OAI22_X1 U13819 ( .A1(n12819), .A2(n10839), .B1(n19597), .B2(n9863), .ZN(
        n10840) );
  AOI21_X1 U13820 ( .B1(n14129), .B2(P2_REIP_REG_22__SCAN_IN), .A(n10840), 
        .ZN(n10841) );
  NAND2_X1 U13821 ( .A1(n10842), .A2(n10841), .ZN(n15305) );
  INV_X1 U13822 ( .A(n15101), .ZN(n10844) );
  AOI21_X1 U13823 ( .B1(n10845), .B2(n10843), .A(n10844), .ZN(n15111) );
  NAND2_X1 U13824 ( .A1(n9728), .A2(n19737), .ZN(n10847) );
  NAND2_X1 U13825 ( .A1(n10847), .A2(n10846), .ZN(n10848) );
  NAND2_X1 U13826 ( .A1(n15111), .A2(n16143), .ZN(n11073) );
  OAI21_X1 U13827 ( .B1(n13009), .B2(n10850), .A(n13135), .ZN(n10852) );
  NAND2_X1 U13828 ( .A1(n10852), .A2(n10851), .ZN(n10854) );
  NAND2_X1 U13829 ( .A1(n10853), .A2(n13009), .ZN(n13138) );
  OAI211_X1 U13830 ( .C1(n10195), .C2(n13135), .A(n10854), .B(n13138), .ZN(
        n10855) );
  INV_X1 U13831 ( .A(n10855), .ZN(n10864) );
  MUX2_X1 U13832 ( .A(n10857), .B(n10856), .S(n10528), .Z(n10858) );
  INV_X1 U13833 ( .A(n10858), .ZN(n10863) );
  NAND2_X1 U13834 ( .A1(n10859), .A2(n10215), .ZN(n15448) );
  NAND2_X1 U13835 ( .A1(n15448), .A2(n10860), .ZN(n10861) );
  NAND2_X1 U13836 ( .A1(n10861), .A2(n10208), .ZN(n10862) );
  NAND2_X1 U13837 ( .A1(n15461), .A2(n10865), .ZN(n10866) );
  NAND2_X1 U13838 ( .A1(n10891), .A2(n10866), .ZN(n15333) );
  NAND2_X1 U13839 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19079) );
  INV_X1 U13840 ( .A(n19079), .ZN(n10867) );
  OR2_X1 U13841 ( .A1(n15333), .A2(n10867), .ZN(n10868) );
  NOR2_X2 U13842 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19697) );
  NAND2_X1 U13843 ( .A1(n19697), .A2(n19597), .ZN(n18751) );
  OR2_X1 U13844 ( .A1(n18751), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11123) );
  INV_X1 U13845 ( .A(n11123), .ZN(n16060) );
  OR2_X1 U13846 ( .A1(n10891), .A2(n16060), .ZN(n19070) );
  NAND2_X1 U13847 ( .A1(n10891), .A2(n13134), .ZN(n13156) );
  NAND2_X1 U13848 ( .A1(n13156), .A2(n15333), .ZN(n19078) );
  INV_X1 U13849 ( .A(n19078), .ZN(n15285) );
  NAND2_X1 U13850 ( .A1(n13171), .A2(n15285), .ZN(n16130) );
  INV_X1 U13851 ( .A(n16130), .ZN(n13976) );
  NOR3_X1 U13852 ( .A1(n10262), .A2(n13936), .A3(n13935), .ZN(n13979) );
  NAND2_X1 U13853 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13979), .ZN(
        n16133) );
  NOR2_X1 U13854 ( .A1(n10871), .A2(n16133), .ZN(n16134) );
  NAND2_X1 U13855 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n16134), .ZN(
        n10878) );
  INV_X1 U13856 ( .A(n13156), .ZN(n15331) );
  NOR2_X1 U13857 ( .A1(n13172), .A2(n19079), .ZN(n10872) );
  NAND2_X1 U13858 ( .A1(n13172), .A2(n19079), .ZN(n10876) );
  OAI211_X1 U13859 ( .C1(n15331), .C2(n10872), .A(n10876), .B(n19078), .ZN(
        n16132) );
  NOR2_X1 U13860 ( .A1(n10878), .A2(n16132), .ZN(n15440) );
  NAND2_X1 U13861 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15440), .ZN(
        n16115) );
  AND2_X1 U13862 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15426) );
  INV_X1 U13863 ( .A(n15426), .ZN(n10880) );
  INV_X1 U13864 ( .A(n15379), .ZN(n10873) );
  AND2_X1 U13865 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n10873), .ZN(
        n10882) );
  NAND2_X1 U13866 ( .A1(n15402), .A2(n10882), .ZN(n15358) );
  INV_X1 U13867 ( .A(n12337), .ZN(n12338) );
  NAND2_X1 U13868 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10874) );
  NAND2_X1 U13869 ( .A1(n14214), .A2(n10875), .ZN(n10885) );
  INV_X1 U13870 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n20889) );
  OR2_X1 U13871 ( .A1(n13156), .A2(n10876), .ZN(n13160) );
  INV_X1 U13872 ( .A(n15333), .ZN(n10877) );
  NAND2_X1 U13873 ( .A1(n10877), .A2(n13172), .ZN(n13155) );
  NAND3_X1 U13874 ( .A1(n13171), .A2(n13160), .A3(n13155), .ZN(n16156) );
  NOR3_X1 U13875 ( .A1(n10878), .A2(n20889), .A3(n16156), .ZN(n10879) );
  OR2_X1 U13876 ( .A1(n10879), .A2(n13976), .ZN(n16113) );
  NAND2_X1 U13877 ( .A1(n16130), .A2(n10880), .ZN(n10881) );
  INV_X1 U13878 ( .A(n10882), .ZN(n10883) );
  NAND2_X1 U13879 ( .A1(n16130), .A2(n10883), .ZN(n10884) );
  OAI211_X1 U13880 ( .C1(n12867), .C2(n13976), .A(n10885), .B(n15364), .ZN(
        n14213) );
  INV_X1 U13881 ( .A(n14213), .ZN(n15311) );
  INV_X1 U13882 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11092) );
  NAND2_X1 U13883 ( .A1(n10886), .A2(n10887), .ZN(n16181) );
  NAND2_X1 U13884 ( .A1(n9729), .A2(n10215), .ZN(n10889) );
  NAND2_X1 U13885 ( .A1(n16181), .A2(n10889), .ZN(n10890) );
  NAND2_X1 U13886 ( .A1(n10891), .A2(n10890), .ZN(n16161) );
  NAND2_X1 U13887 ( .A1(n13914), .A2(n13007), .ZN(n10908) );
  INV_X1 U13888 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19622) );
  AND2_X2 U13889 ( .A1(n10558), .A2(n19546), .ZN(n11131) );
  AOI22_X1 U13890 ( .A1(n11131), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n10991), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10892) );
  MUX2_X1 U13891 ( .A(n10203), .B(n19715), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10895) );
  INV_X1 U13892 ( .A(n13144), .ZN(n10894) );
  NAND2_X1 U13893 ( .A1(n10894), .A2(n10991), .ZN(n10905) );
  INV_X1 U13894 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18928) );
  NAND2_X1 U13895 ( .A1(n10558), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10897) );
  AOI21_X1 U13896 ( .B1(n10215), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10896) );
  AND2_X1 U13897 ( .A1(n10897), .A2(n10896), .ZN(n10898) );
  AND2_X1 U13898 ( .A1(n13144), .A2(n10203), .ZN(n13141) );
  MUX2_X1 U13899 ( .A(n13141), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_3__SCAN_IN), .Z(n10902) );
  NOR2_X1 U13900 ( .A1(n10899), .A2(n10900), .ZN(n10901) );
  NOR2_X1 U13901 ( .A1(n10902), .A2(n10901), .ZN(n13323) );
  NOR2_X1 U13902 ( .A1(n13145), .A2(n10903), .ZN(n10904) );
  NAND2_X1 U13903 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10906) );
  OAI211_X1 U13904 ( .C1(n10899), .C2(n10907), .A(n10906), .B(n10905), .ZN(
        n10911) );
  INV_X1 U13905 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19624) );
  OR2_X1 U13906 ( .A1(n10908), .A2(n19624), .ZN(n10910) );
  AOI22_X1 U13907 ( .A1(n11131), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n10991), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10909) );
  NAND2_X1 U13908 ( .A1(n10910), .A2(n10909), .ZN(n13153) );
  NOR2_X1 U13909 ( .A1(n13154), .A2(n13153), .ZN(n13152) );
  NOR2_X1 U13910 ( .A1(n10912), .A2(n10911), .ZN(n10913) );
  INV_X1 U13911 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n10914) );
  OR2_X1 U13912 ( .A1(n10908), .A2(n10914), .ZN(n10918) );
  AOI22_X1 U13913 ( .A1(n10991), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n10916) );
  NAND2_X1 U13914 ( .A1(n11131), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10915) );
  AND2_X1 U13915 ( .A1(n10916), .A2(n10915), .ZN(n10917) );
  OAI211_X1 U13916 ( .C1(n10919), .C2(n10899), .A(n10918), .B(n10917), .ZN(
        n13585) );
  NAND2_X1 U13917 ( .A1(n13586), .A2(n13585), .ZN(n13587) );
  INV_X1 U13918 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10920) );
  OR2_X1 U13919 ( .A1(n10908), .A2(n10920), .ZN(n10924) );
  AOI22_X1 U13920 ( .A1(n11131), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n10991), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10923) );
  OR2_X1 U13921 ( .A1(n10899), .A2(n10921), .ZN(n10922) );
  INV_X1 U13922 ( .A(n13007), .ZN(n10926) );
  OAI22_X1 U13923 ( .A1(n10908), .A2(n19628), .B1(n10926), .B2(n10925), .ZN(
        n10927) );
  INV_X1 U13924 ( .A(n10927), .ZN(n10929) );
  AOI22_X1 U13925 ( .A1(n11131), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n10991), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10928) );
  NAND2_X1 U13926 ( .A1(n10929), .A2(n10928), .ZN(n13933) );
  OR2_X1 U13927 ( .A1(n10899), .A2(n10930), .ZN(n10931) );
  INV_X1 U13928 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19630) );
  OR2_X1 U13929 ( .A1(n10908), .A2(n19630), .ZN(n10933) );
  AOI22_X1 U13930 ( .A1(n11131), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n10991), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10932) );
  OR2_X1 U13931 ( .A1(n10899), .A2(n10934), .ZN(n10935) );
  INV_X1 U13932 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19632) );
  OR2_X1 U13933 ( .A1(n10908), .A2(n19632), .ZN(n10938) );
  AOI22_X1 U13934 ( .A1(n11131), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n10991), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10937) );
  NAND2_X1 U13935 ( .A1(n10938), .A2(n10937), .ZN(n13203) );
  INV_X1 U13936 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n10939) );
  OR2_X1 U13937 ( .A1(n10908), .A2(n10939), .ZN(n10952) );
  AOI22_X1 U13938 ( .A1(n11131), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n10991), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10951) );
  AOI22_X1 U13939 ( .A1(n14293), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U13940 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U13941 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U13942 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10407), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10940) );
  NAND4_X1 U13943 ( .A1(n10943), .A2(n10942), .A3(n10941), .A4(n10940), .ZN(
        n10949) );
  AOI22_X1 U13944 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10947) );
  AOI22_X1 U13945 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10946) );
  AOI22_X1 U13946 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10945) );
  AOI22_X1 U13947 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10944) );
  NAND4_X1 U13948 ( .A1(n10947), .A2(n10946), .A3(n10945), .A4(n10944), .ZN(
        n10948) );
  INV_X1 U13949 ( .A(n13518), .ZN(n13522) );
  OR2_X1 U13950 ( .A1(n10899), .A2(n13522), .ZN(n10950) );
  AOI22_X1 U13951 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n14293), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10956) );
  AOI22_X1 U13952 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10406), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10955) );
  AOI22_X1 U13953 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10954) );
  AOI22_X1 U13954 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10372), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10953) );
  NAND4_X1 U13955 ( .A1(n10956), .A2(n10955), .A3(n10954), .A4(n10953), .ZN(
        n10962) );
  AOI22_X1 U13956 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10407), .B1(
        n14294), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U13957 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9708), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U13958 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10373), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U13959 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10374), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10957) );
  NAND4_X1 U13960 ( .A1(n10960), .A2(n10959), .A3(n10958), .A4(n10957), .ZN(
        n10961) );
  OR2_X1 U13961 ( .A1(n10962), .A2(n10961), .ZN(n13517) );
  INV_X1 U13962 ( .A(n13517), .ZN(n13521) );
  INV_X1 U13963 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n10963) );
  OR2_X1 U13964 ( .A1(n10908), .A2(n10963), .ZN(n10965) );
  AOI22_X1 U13965 ( .A1(n11131), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n10991), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10964) );
  OAI211_X1 U13966 ( .C1(n13521), .C2(n10899), .A(n10965), .B(n10964), .ZN(
        n13238) );
  INV_X1 U13967 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n10966) );
  OR2_X1 U13968 ( .A1(n10908), .A2(n10966), .ZN(n10979) );
  AOI22_X1 U13969 ( .A1(n11131), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10978) );
  AOI22_X1 U13970 ( .A1(n14293), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10406), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U13971 ( .A1(n10354), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10355), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10969) );
  AOI22_X1 U13972 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10968) );
  AOI22_X1 U13973 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10967) );
  NAND4_X1 U13974 ( .A1(n10970), .A2(n10969), .A3(n10968), .A4(n10967), .ZN(
        n10976) );
  AOI22_X1 U13975 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U13976 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10973) );
  AOI22_X1 U13977 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10972) );
  AOI22_X1 U13978 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10971) );
  NAND4_X1 U13979 ( .A1(n10974), .A2(n10973), .A3(n10972), .A4(n10971), .ZN(
        n10975) );
  OR2_X1 U13980 ( .A1(n10976), .A2(n10975), .ZN(n13534) );
  INV_X1 U13981 ( .A(n13534), .ZN(n18960) );
  OR2_X1 U13982 ( .A1(n10899), .A2(n18960), .ZN(n10977) );
  AOI22_X1 U13983 ( .A1(n14293), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10983) );
  AOI22_X1 U13984 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10982) );
  AOI22_X1 U13985 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10981) );
  AOI22_X1 U13986 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10407), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10980) );
  NAND4_X1 U13987 ( .A1(n10983), .A2(n10982), .A3(n10981), .A4(n10980), .ZN(
        n10989) );
  AOI22_X1 U13988 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10987) );
  AOI22_X1 U13989 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U13990 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10985) );
  AOI22_X1 U13991 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10984) );
  NAND4_X1 U13992 ( .A1(n10987), .A2(n10986), .A3(n10985), .A4(n10984), .ZN(
        n10988) );
  OR2_X1 U13993 ( .A1(n10989), .A2(n10988), .ZN(n13533) );
  INV_X1 U13994 ( .A(n13533), .ZN(n13531) );
  INV_X1 U13995 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n10990) );
  OR2_X1 U13996 ( .A1(n10908), .A2(n10990), .ZN(n10993) );
  AOI22_X1 U13997 ( .A1(n11131), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10992) );
  OAI211_X1 U13998 ( .C1(n13531), .C2(n10899), .A(n10993), .B(n10992), .ZN(
        n12984) );
  INV_X1 U13999 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n10994) );
  OR2_X1 U14000 ( .A1(n10908), .A2(n10994), .ZN(n11007) );
  AOI22_X1 U14001 ( .A1(n11131), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U14002 ( .A1(n14293), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U14003 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10997) );
  AOI22_X1 U14004 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10355), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10996) );
  AOI22_X1 U14005 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10995) );
  NAND4_X1 U14006 ( .A1(n10998), .A2(n10997), .A3(n10996), .A4(n10995), .ZN(
        n11004) );
  AOI22_X1 U14007 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10383), .B1(
        n10407), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U14008 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U14009 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U14010 ( .A1(n10388), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10999) );
  NAND4_X1 U14011 ( .A1(n11002), .A2(n11001), .A3(n11000), .A4(n10999), .ZN(
        n11003) );
  OR2_X1 U14012 ( .A1(n10899), .A2(n13613), .ZN(n11005) );
  AOI22_X1 U14013 ( .A1(n14293), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11011) );
  AOI22_X1 U14014 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11010) );
  AOI22_X1 U14015 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11009) );
  AOI22_X1 U14016 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10407), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11008) );
  NAND4_X1 U14017 ( .A1(n11011), .A2(n11010), .A3(n11009), .A4(n11008), .ZN(
        n11017) );
  AOI22_X1 U14018 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11015) );
  AOI22_X1 U14019 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11014) );
  AOI22_X1 U14020 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11013) );
  AOI22_X1 U14021 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11012) );
  NAND4_X1 U14022 ( .A1(n11015), .A2(n11014), .A3(n11013), .A4(n11012), .ZN(
        n11016) );
  NOR2_X1 U14023 ( .A1(n11017), .A2(n11016), .ZN(n13612) );
  NAND2_X1 U14024 ( .A1(n14144), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U14025 ( .A1(n11131), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11018) );
  OAI211_X1 U14026 ( .C1(n13612), .C2(n10899), .A(n11019), .B(n11018), .ZN(
        n13544) );
  INV_X1 U14027 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11020) );
  OR2_X1 U14028 ( .A1(n10908), .A2(n11020), .ZN(n11033) );
  AOI22_X1 U14029 ( .A1(n11131), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11032) );
  AOI22_X1 U14030 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11024) );
  AOI22_X1 U14031 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11023) );
  AOI22_X1 U14032 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U14033 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11021) );
  NAND4_X1 U14034 ( .A1(n11024), .A2(n11023), .A3(n11022), .A4(n11021), .ZN(
        n11030) );
  AOI22_X1 U14035 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11028) );
  AOI22_X1 U14036 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U14037 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11026) );
  AOI22_X1 U14038 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11025) );
  NAND4_X1 U14039 ( .A1(n11028), .A2(n11027), .A3(n11026), .A4(n11025), .ZN(
        n11029) );
  NOR2_X1 U14040 ( .A1(n11030), .A2(n11029), .ZN(n18952) );
  OR2_X1 U14041 ( .A1(n10899), .A2(n18952), .ZN(n11031) );
  INV_X1 U14042 ( .A(n10899), .ZN(n11044) );
  AOI22_X1 U14043 ( .A1(n14293), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11037) );
  AOI22_X1 U14044 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11036) );
  AOI22_X1 U14045 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11035) );
  AOI22_X1 U14046 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10407), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11034) );
  NAND4_X1 U14047 ( .A1(n11037), .A2(n11036), .A3(n11035), .A4(n11034), .ZN(
        n11043) );
  AOI22_X1 U14048 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11041) );
  AOI22_X1 U14049 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U14050 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11039) );
  AOI22_X1 U14051 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11038) );
  NAND4_X1 U14052 ( .A1(n11041), .A2(n11040), .A3(n11039), .A4(n11038), .ZN(
        n11042) );
  AOI22_X1 U14053 ( .A1(n14144), .A2(P2_REIP_REG_15__SCAN_IN), .B1(n11044), 
        .B2(n13868), .ZN(n11046) );
  AOI22_X1 U14054 ( .A1(n11131), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11045) );
  NAND2_X1 U14055 ( .A1(n11046), .A2(n11045), .ZN(n13630) );
  INV_X1 U14056 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15346) );
  OR2_X1 U14057 ( .A1(n10908), .A2(n15346), .ZN(n11048) );
  AOI22_X1 U14058 ( .A1(n11131), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11047) );
  INV_X1 U14059 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19644) );
  OR2_X1 U14060 ( .A1(n10908), .A2(n19644), .ZN(n11050) );
  AOI22_X1 U14061 ( .A1(n11131), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11049) );
  NAND2_X1 U14062 ( .A1(n11050), .A2(n11049), .ZN(n13956) );
  NAND2_X1 U14063 ( .A1(n13851), .A2(n13956), .ZN(n12340) );
  INV_X1 U14064 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19646) );
  OR2_X1 U14065 ( .A1(n10908), .A2(n19646), .ZN(n11052) );
  AOI22_X1 U14066 ( .A1(n11131), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11051) );
  AND2_X1 U14067 ( .A1(n11052), .A2(n11051), .ZN(n12341) );
  INV_X1 U14068 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19648) );
  OR2_X1 U14069 ( .A1(n10908), .A2(n19648), .ZN(n11054) );
  AOI22_X1 U14070 ( .A1(n11131), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11053) );
  OR2_X1 U14071 ( .A1(n10908), .A2(n19650), .ZN(n11056) );
  AOI22_X1 U14072 ( .A1(n11131), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11055) );
  NAND2_X1 U14073 ( .A1(n11056), .A2(n11055), .ZN(n14090) );
  INV_X1 U14074 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19652) );
  OR2_X1 U14075 ( .A1(n10908), .A2(n19652), .ZN(n11058) );
  AOI22_X1 U14076 ( .A1(n11131), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11057) );
  NAND2_X1 U14077 ( .A1(n11058), .A2(n11057), .ZN(n14038) );
  INV_X1 U14078 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n11059) );
  OR2_X1 U14079 ( .A1(n10908), .A2(n11059), .ZN(n11061) );
  AOI22_X1 U14080 ( .A1(n11131), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11060) );
  NAND2_X1 U14081 ( .A1(n11061), .A2(n11060), .ZN(n15166) );
  INV_X1 U14082 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19655) );
  OR2_X1 U14083 ( .A1(n10908), .A2(n19655), .ZN(n11063) );
  AOI22_X1 U14084 ( .A1(n11131), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11062) );
  NAND2_X1 U14085 ( .A1(n11063), .A2(n11062), .ZN(n11066) );
  INV_X1 U14086 ( .A(n11134), .ZN(n15152) );
  AOI21_X1 U14087 ( .B1(n15166), .B2(n11065), .A(n11066), .ZN(n11067) );
  NOR2_X1 U14088 ( .A1(n15152), .A2(n11067), .ZN(n15160) );
  NAND2_X1 U14089 ( .A1(n16060), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11083) );
  INV_X1 U14090 ( .A(n11083), .ZN(n11068) );
  AOI21_X1 U14091 ( .B1(n19067), .B2(n15160), .A(n11068), .ZN(n11070) );
  OAI211_X1 U14092 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15309), .B(n11090), .ZN(
        n11069) );
  OAI211_X1 U14093 ( .C1(n15311), .C2(n11092), .A(n11070), .B(n11069), .ZN(
        n11071) );
  OAI211_X1 U14094 ( .C1(n11087), .C2(n16163), .A(n11073), .B(n11072), .ZN(
        n11074) );
  OR2_X1 U14095 ( .A1(n11075), .A2(n11074), .ZN(P2_U3023) );
  NAND2_X1 U14096 ( .A1(n19719), .A2(n16211), .ZN(n11076) );
  NAND2_X1 U14097 ( .A1(n11077), .A2(n11076), .ZN(n11078) );
  NAND2_X1 U14098 ( .A1(n11078), .A2(n19731), .ZN(n18757) );
  NOR2_X1 U14099 ( .A1(n11079), .A2(n16083), .ZN(n11089) );
  NAND2_X1 U14100 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n13490) );
  AOI21_X1 U14101 ( .B1(n19732), .B2(n19597), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19742) );
  AND2_X1 U14102 ( .A1(n13490), .A2(n19742), .ZN(n11080) );
  NOR2_X1 U14103 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19596) );
  OR2_X1 U14104 ( .A1(n19697), .A2(n19596), .ZN(n19701) );
  NAND2_X1 U14105 ( .A1(n19701), .A2(n19727), .ZN(n11081) );
  NAND2_X1 U14106 ( .A1(n19727), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13308) );
  INV_X1 U14107 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19738) );
  NAND2_X1 U14108 ( .A1(n19738), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11082) );
  NAND2_X1 U14109 ( .A1(n13308), .A2(n11082), .ZN(n14257) );
  NAND2_X1 U14110 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n12758), .ZN(
        n12755) );
  AOI21_X1 U14111 ( .B1(n12973), .B2(n12776), .A(n11121), .ZN(n12971) );
  NAND2_X1 U14112 ( .A1(n16090), .A2(n12971), .ZN(n11084) );
  OAI211_X1 U14113 ( .C1(n12973), .C2(n16100), .A(n11084), .B(n11083), .ZN(
        n11085) );
  OR2_X1 U14114 ( .A1(n11089), .A2(n11088), .ZN(P2_U2991) );
  INV_X1 U14115 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14196) );
  INV_X1 U14116 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15286) );
  NOR2_X1 U14117 ( .A1(n11090), .A2(n15286), .ZN(n14198) );
  INV_X1 U14118 ( .A(n14198), .ZN(n11130) );
  NOR2_X1 U14119 ( .A1(n14196), .A2(n11130), .ZN(n11091) );
  AND2_X2 U14120 ( .A1(n11091), .A2(n15303), .ZN(n14228) );
  NAND2_X1 U14121 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11141) );
  INV_X1 U14122 ( .A(n11141), .ZN(n12928) );
  AND2_X1 U14123 ( .A1(n12928), .A2(n14198), .ZN(n12863) );
  NAND2_X1 U14124 ( .A1(n15303), .A2(n12863), .ZN(n15201) );
  OAI21_X1 U14125 ( .B1(n14228), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15201), .ZN(n11128) );
  NOR2_X2 U14126 ( .A1(n11096), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11103) );
  INV_X1 U14127 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n11112) );
  NAND2_X1 U14128 ( .A1(n11103), .A2(n11112), .ZN(n15954) );
  NAND2_X2 U14129 ( .A1(n10689), .A2(n9704), .ZN(n15953) );
  NOR2_X1 U14130 ( .A1(n15953), .A2(n10934), .ZN(n12859) );
  XOR2_X1 U14131 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n12859), .Z(
        n12846) );
  NOR3_X1 U14132 ( .A1(n12974), .A2(n10934), .A3(n11092), .ZN(n11093) );
  INV_X1 U14133 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n11098) );
  NOR2_X1 U14134 ( .A1(n9763), .A2(n11098), .ZN(n11099) );
  INV_X1 U14135 ( .A(n11096), .ZN(n11097) );
  MUX2_X1 U14136 ( .A(n11099), .B(n11098), .S(n11097), .Z(n11101) );
  NOR2_X1 U14137 ( .A1(n11101), .A2(n11100), .ZN(n15963) );
  NAND2_X1 U14138 ( .A1(n15963), .A2(n14238), .ZN(n15210) );
  OAI21_X1 U14139 ( .B1(n9788), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11102), .ZN(n14187) );
  NAND2_X1 U14140 ( .A1(n9757), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11104) );
  MUX2_X1 U14141 ( .A(n11104), .B(P2_EBX_REG_25__SCAN_IN), .S(n11103), .Z(
        n11105) );
  AOI21_X1 U14142 ( .B1(n11106), .B2(n14238), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14186) );
  NOR2_X2 U14143 ( .A1(n14187), .A2(n14186), .ZN(n12847) );
  NAND2_X1 U14144 ( .A1(n14238), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11107) );
  NOR2_X1 U14145 ( .A1(n12847), .A2(n14185), .ZN(n11108) );
  XOR2_X1 U14146 ( .A(n12846), .B(n11108), .Z(n11129) );
  OR2_X1 U14147 ( .A1(n11129), .A2(n16084), .ZN(n11127) );
  NAND2_X1 U14148 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11111) );
  INV_X1 U14149 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15215) );
  OAI22_X1 U14150 ( .A1(n12819), .A2(n11098), .B1(n19597), .B2(n15215), .ZN(
        n11109) );
  AOI21_X1 U14151 ( .B1(n14129), .B2(P2_REIP_REG_24__SCAN_IN), .A(n11109), 
        .ZN(n11110) );
  NAND2_X1 U14152 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11115) );
  INV_X1 U14153 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15038) );
  OAI22_X1 U14154 ( .A1(n12819), .A2(n11112), .B1(n19597), .B2(n15038), .ZN(
        n11113) );
  AOI21_X1 U14155 ( .B1(n14129), .B2(P2_REIP_REG_25__SCAN_IN), .A(n11113), 
        .ZN(n11114) );
  AND2_X1 U14156 ( .A1(n11115), .A2(n11114), .ZN(n14190) );
  NAND2_X1 U14157 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11118) );
  INV_X1 U14158 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n15952) );
  OAI22_X1 U14159 ( .A1(n12819), .A2(n15952), .B1(n19597), .B2(n9865), .ZN(
        n11116) );
  AOI21_X1 U14160 ( .B1(n14129), .B2(P2_REIP_REG_26__SCAN_IN), .A(n11116), 
        .ZN(n11117) );
  NAND2_X1 U14161 ( .A1(n11118), .A2(n11117), .ZN(n11119) );
  OR2_X1 U14162 ( .A1(n10083), .A2(n11119), .ZN(n11120) );
  NAND2_X1 U14163 ( .A1(n10083), .A2(n11119), .ZN(n12810) );
  AND2_X1 U14164 ( .A1(n11120), .A2(n12810), .ZN(n15088) );
  NAND2_X1 U14165 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n11121), .ZN(
        n12753) );
  INV_X1 U14166 ( .A(n12753), .ZN(n11122) );
  OAI21_X1 U14167 ( .B1(n12752), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n12750), .ZN(n12751) );
  INV_X1 U14168 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19661) );
  NOR2_X1 U14169 ( .A1(n11123), .A2(n19661), .ZN(n11140) );
  AOI21_X1 U14170 ( .B1(n19055), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n11140), .ZN(n11124) );
  OAI21_X1 U14171 ( .B1(n19061), .B2(n12751), .A(n11124), .ZN(n11125) );
  AOI21_X1 U14172 ( .B1(n15088), .B2(n19063), .A(n11125), .ZN(n11126) );
  OR2_X1 U14173 ( .A1(n11129), .A2(n16163), .ZN(n11147) );
  AOI21_X1 U14174 ( .B1(n11130), .B2(n19078), .A(n14213), .ZN(n14197) );
  INV_X1 U14175 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11144) );
  INV_X1 U14176 ( .A(n11131), .ZN(n14142) );
  INV_X1 U14177 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n11132) );
  INV_X1 U14178 ( .A(n10991), .ZN(n14140) );
  OAI22_X1 U14179 ( .A1(n14142), .A2(n11132), .B1(n14140), .B2(n15286), .ZN(
        n11133) );
  AOI21_X1 U14180 ( .B1(n14144), .B2(P2_REIP_REG_24__SCAN_IN), .A(n11133), 
        .ZN(n15149) );
  INV_X1 U14181 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15139) );
  OAI22_X1 U14182 ( .A1(n14142), .A2(n15139), .B1(n14140), .B2(n14196), .ZN(
        n11135) );
  AOI21_X1 U14183 ( .B1(n14144), .B2(P2_REIP_REG_25__SCAN_IN), .A(n11135), 
        .ZN(n14192) );
  OR2_X1 U14184 ( .A1(n10908), .A2(n19661), .ZN(n11137) );
  AOI22_X1 U14185 ( .A1(n11131), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U14186 ( .A1(n11137), .A2(n11136), .ZN(n11138) );
  OR2_X1 U14187 ( .A1(n14191), .A2(n11138), .ZN(n11139) );
  AND2_X1 U14188 ( .A1(n12788), .A2(n11139), .ZN(n15961) );
  AOI21_X1 U14189 ( .B1(n19067), .B2(n15961), .A(n11140), .ZN(n11143) );
  OAI211_X1 U14190 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n14194), .B(n11141), .ZN(
        n11142) );
  OAI211_X1 U14191 ( .C1(n14197), .C2(n11144), .A(n11143), .B(n11142), .ZN(
        n11145) );
  INV_X1 U14192 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11148) );
  AND2_X2 U14193 ( .A1(n11148), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11160) );
  AND2_X2 U14194 ( .A1(n11158), .A2(n13270), .ZN(n11339) );
  AOI22_X1 U14195 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11156) );
  AOI22_X1 U14196 ( .A1(n11437), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11438), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11155) );
  AOI22_X1 U14197 ( .A1(n11337), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11154) );
  AOI22_X1 U14198 ( .A1(n12208), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9747), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11153) );
  AOI22_X1 U14199 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9751), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11165) );
  AND2_X2 U14200 ( .A1(n11158), .A2(n11159), .ZN(n11224) );
  AOI22_X1 U14201 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11164) );
  AOI22_X1 U14202 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11163) );
  AOI22_X1 U14203 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11338), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11162) );
  AOI22_X1 U14204 ( .A1(n9768), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12213), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11169) );
  AOI22_X1 U14205 ( .A1(n11336), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11168) );
  AOI22_X1 U14206 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11167) );
  AOI22_X1 U14207 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11166) );
  AOI22_X1 U14208 ( .A1(n11437), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11173) );
  AOI22_X1 U14209 ( .A1(n11337), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11863), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11172) );
  AOI22_X1 U14210 ( .A1(n12208), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11381), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11171) );
  AOI22_X1 U14211 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11438), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11170) );
  NAND2_X1 U14212 ( .A1(n11277), .A2(n20013), .ZN(n11279) );
  AOI22_X1 U14213 ( .A1(n11437), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11177) );
  AOI22_X1 U14214 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11438), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11176) );
  AOI22_X1 U14215 ( .A1(n12208), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9747), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11175) );
  AOI22_X1 U14216 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11174) );
  AOI22_X1 U14217 ( .A1(n11337), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11338), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11181) );
  AOI22_X1 U14218 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11180) );
  AOI22_X1 U14219 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11179) );
  NAND2_X1 U14220 ( .A1(n11279), .A2(n11628), .ZN(n11204) );
  AOI22_X1 U14221 ( .A1(n11437), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11187) );
  AOI22_X1 U14222 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11438), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11186) );
  AOI22_X1 U14223 ( .A1(n9744), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11381), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11185) );
  AOI22_X1 U14224 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9739), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11184) );
  AOI22_X1 U14225 ( .A1(n12213), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11191) );
  AOI22_X1 U14226 ( .A1(n11337), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11338), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11190) );
  AOI22_X1 U14227 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11189) );
  AOI22_X1 U14228 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11188) );
  AND4_X2 U14229 ( .A1(n11191), .A2(n11190), .A3(n11189), .A4(n11188), .ZN(
        n11192) );
  NAND2_X4 U14230 ( .A1(n11193), .A2(n11192), .ZN(n20006) );
  AOI22_X1 U14231 ( .A1(n12213), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11197) );
  AOI22_X1 U14232 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11196) );
  AOI22_X1 U14233 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11195) );
  AOI22_X1 U14234 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11194) );
  NAND4_X1 U14235 ( .A1(n11197), .A2(n11196), .A3(n11195), .A4(n11194), .ZN(
        n11203) );
  AOI22_X1 U14236 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11338), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11201) );
  AOI22_X1 U14237 ( .A1(n11337), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11200) );
  AOI22_X1 U14238 ( .A1(n11437), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9735), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11199) );
  AOI22_X1 U14239 ( .A1(n12208), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9747), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11198) );
  NAND4_X1 U14240 ( .A1(n11201), .A2(n11200), .A3(n11199), .A4(n11198), .ZN(
        n11202) );
  NAND2_X1 U14241 ( .A1(n11278), .A2(n11272), .ZN(n11294) );
  NAND2_X1 U14242 ( .A1(n11204), .A2(n11294), .ZN(n11219) );
  AOI22_X1 U14243 ( .A1(n9768), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11208) );
  AOI22_X1 U14244 ( .A1(n11337), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11207) );
  AOI22_X1 U14245 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11206) );
  AOI22_X1 U14246 ( .A1(n12213), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11205) );
  NAND4_X1 U14247 ( .A1(n11208), .A2(n11207), .A3(n11206), .A4(n11205), .ZN(
        n11214) );
  AOI22_X1 U14248 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9734), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14249 ( .A1(n11437), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9750), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U14250 ( .A1(n12208), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11210) );
  AOI22_X1 U14251 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9738), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11209) );
  NAND4_X1 U14252 ( .A1(n11212), .A2(n11211), .A3(n11210), .A4(n11209), .ZN(
        n11213) );
  NAND2_X1 U14253 ( .A1(n11215), .A2(n9731), .ZN(n11217) );
  NAND2_X2 U14254 ( .A1(n20006), .A2(n9721), .ZN(n11273) );
  NAND2_X1 U14255 ( .A1(n11273), .A2(n19996), .ZN(n11216) );
  NAND2_X1 U14256 ( .A1(n11217), .A2(n11216), .ZN(n11218) );
  NOR2_X2 U14257 ( .A1(n11219), .A2(n11218), .ZN(n11269) );
  NAND2_X1 U14258 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11223) );
  NAND2_X1 U14259 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11222) );
  NAND2_X1 U14260 ( .A1(n11437), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11221) );
  NAND2_X1 U14261 ( .A1(n9751), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11220) );
  NAND2_X1 U14262 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11228) );
  NAND2_X1 U14263 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11227) );
  NAND2_X1 U14264 ( .A1(n11336), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11226) );
  NAND2_X1 U14265 ( .A1(n11224), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11225) );
  NAND2_X1 U14266 ( .A1(n11337), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11232) );
  NAND2_X1 U14267 ( .A1(n12213), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11231) );
  NAND2_X1 U14268 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11230) );
  NAND2_X1 U14269 ( .A1(n11339), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11229) );
  NAND2_X1 U14270 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11236) );
  NAND2_X1 U14271 ( .A1(n12208), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11235) );
  NAND2_X1 U14272 ( .A1(n11438), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11234) );
  NAND2_X1 U14273 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11233) );
  AND4_X4 U14274 ( .A1(n11240), .A2(n11239), .A3(n11238), .A4(n11237), .ZN(
        n13643) );
  NOR2_X1 U14275 ( .A1(n11273), .A2(n19978), .ZN(n11241) );
  NAND2_X1 U14276 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11245) );
  NAND2_X1 U14277 ( .A1(n12213), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11243) );
  NAND2_X1 U14278 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11242) );
  NAND2_X1 U14279 ( .A1(n11337), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11249) );
  NAND2_X1 U14280 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11248) );
  NAND2_X1 U14281 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11247) );
  NAND2_X1 U14282 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11246) );
  AND4_X1 U14283 ( .A1(n11249), .A2(n11248), .A3(n11247), .A4(n11246), .ZN(
        n11260) );
  NAND2_X1 U14284 ( .A1(n11437), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11253) );
  NAND2_X1 U14285 ( .A1(n9735), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11252) );
  NAND2_X1 U14286 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11251) );
  NAND2_X1 U14287 ( .A1(n12208), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11250) );
  AND4_X1 U14288 ( .A1(n11253), .A2(n11252), .A3(n11251), .A4(n11250), .ZN(
        n11259) );
  NAND2_X1 U14289 ( .A1(n11336), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11257) );
  NAND2_X1 U14290 ( .A1(n11224), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11256) );
  NAND2_X1 U14291 ( .A1(n11339), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11255) );
  NAND2_X1 U14292 ( .A1(n12215), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11254) );
  INV_X1 U14293 ( .A(n13076), .ZN(n11264) );
  AND2_X2 U14294 ( .A1(n13072), .A2(n20013), .ZN(n13438) );
  NOR2_X1 U14295 ( .A1(n11277), .A2(n11262), .ZN(n11263) );
  NAND2_X1 U14296 ( .A1(n12895), .A2(n13288), .ZN(n11651) );
  NAND2_X1 U14297 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20660) );
  OAI21_X1 U14298 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n20660), .ZN(n11627) );
  NAND2_X1 U14299 ( .A1(n13268), .A2(n13643), .ZN(n11767) );
  INV_X1 U14300 ( .A(n11767), .ZN(n11266) );
  NAND2_X1 U14301 ( .A1(n11266), .A2(n11265), .ZN(n13265) );
  INV_X1 U14302 ( .A(n13265), .ZN(n11267) );
  OAI21_X1 U14303 ( .B1(n13065), .B2(n11627), .A(n11760), .ZN(n11268) );
  NAND2_X2 U14304 ( .A1(n10089), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11364) );
  INV_X1 U14305 ( .A(n11269), .ZN(n11270) );
  NAND2_X1 U14306 ( .A1(n11270), .A2(n13643), .ZN(n11286) );
  NAND2_X1 U14307 ( .A1(n11653), .A2(n13076), .ZN(n11765) );
  NAND2_X1 U14308 ( .A1(n13643), .A2(n19992), .ZN(n13640) );
  NAND2_X1 U14309 ( .A1(n13072), .A2(n11262), .ZN(n12311) );
  INV_X1 U14310 ( .A(n11273), .ZN(n11275) );
  NAND2_X1 U14311 ( .A1(n11275), .A2(n13071), .ZN(n11276) );
  OR2_X2 U14312 ( .A1(n11640), .A2(n11277), .ZN(n11644) );
  INV_X1 U14313 ( .A(n11278), .ZN(n11281) );
  INV_X1 U14314 ( .A(n11279), .ZN(n11280) );
  NAND2_X1 U14315 ( .A1(n19978), .A2(n19996), .ZN(n11282) );
  NOR2_X1 U14316 ( .A1(n20763), .A2(n13073), .ZN(n11283) );
  NAND2_X1 U14317 ( .A1(n9730), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11289) );
  NAND2_X1 U14318 ( .A1(n20579), .A2(n20471), .ZN(n20439) );
  NAND2_X1 U14319 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n15552) );
  NAND2_X1 U14320 ( .A1(n20439), .A2(n15552), .ZN(n20362) );
  INV_X1 U14321 ( .A(n20362), .ZN(n20057) );
  AND2_X1 U14322 ( .A1(n15579), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11366) );
  AOI21_X1 U14323 ( .B1(n20057), .B2(n12840), .A(n11366), .ZN(n11288) );
  XNOR2_X2 U14324 ( .A(n11290), .B(n11364), .ZN(n20090) );
  INV_X1 U14325 ( .A(n15579), .ZN(n11291) );
  MUX2_X1 U14326 ( .A(n11291), .B(n11373), .S(n20471), .Z(n11292) );
  NAND2_X1 U14327 ( .A1(n11294), .A2(n11771), .ZN(n11295) );
  NAND2_X1 U14328 ( .A1(n13643), .A2(n13256), .ZN(n13638) );
  MUX2_X1 U14329 ( .A(n11269), .B(n11295), .S(n13638), .Z(n11301) );
  NAND3_X1 U14330 ( .A1(n11644), .A2(n14978), .A3(n19992), .ZN(n11300) );
  INV_X1 U14331 ( .A(n11296), .ZN(n11298) );
  NAND3_X1 U14332 ( .A1(n13640), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n14983), 
        .ZN(n11297) );
  AOI21_X1 U14333 ( .B1(n15572), .B2(n11298), .A(n11297), .ZN(n11299) );
  OR2_X1 U14334 ( .A1(n11767), .A2(n11262), .ZN(n11780) );
  INV_X1 U14335 ( .A(n20090), .ZN(n11304) );
  INV_X1 U14336 ( .A(n11302), .ZN(n11303) );
  AOI22_X1 U14337 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14338 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11318), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11308) );
  AOI22_X1 U14339 ( .A1(n13548), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11307) );
  AOI22_X1 U14340 ( .A1(n11339), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11306) );
  NAND4_X1 U14341 ( .A1(n11309), .A2(n11308), .A3(n11307), .A4(n11306), .ZN(
        n11315) );
  AOI22_X1 U14342 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11313) );
  AOI22_X1 U14343 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11312) );
  AOI22_X1 U14344 ( .A1(n11376), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11311) );
  AOI22_X1 U14345 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11310) );
  NAND4_X1 U14346 ( .A1(n11313), .A2(n11312), .A3(n11311), .A4(n11310), .ZN(
        n11314) );
  OR2_X1 U14347 ( .A1(n11432), .A2(n11396), .ZN(n11316) );
  OAI21_X2 U14348 ( .B1(n20508), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11316), 
        .ZN(n11317) );
  INV_X1 U14349 ( .A(n11317), .ZN(n11921) );
  NAND2_X1 U14350 ( .A1(n11921), .A2(n19992), .ZN(n11332) );
  AOI22_X1 U14351 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11322) );
  BUF_X1 U14352 ( .A(n11437), .Z(n11318) );
  AOI22_X1 U14353 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11318), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14354 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11381), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11320) );
  AOI22_X1 U14355 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11319) );
  NAND4_X1 U14356 ( .A1(n11322), .A2(n11321), .A3(n11320), .A4(n11319), .ZN(
        n11328) );
  AOI22_X1 U14357 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14358 ( .A1(n11376), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14359 ( .A1(n12213), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U14360 ( .A1(n11338), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11323) );
  NAND4_X1 U14361 ( .A1(n11326), .A2(n11325), .A3(n11324), .A4(n11323), .ZN(
        n11327) );
  XNOR2_X1 U14362 ( .A(n11396), .B(n11415), .ZN(n11330) );
  NAND2_X1 U14363 ( .A1(n9731), .A2(n20006), .ZN(n11329) );
  AOI21_X1 U14364 ( .B1(n15572), .B2(n11330), .A(n11329), .ZN(n11331) );
  AOI22_X1 U14365 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14366 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11338), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14367 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11341) );
  INV_X1 U14368 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n20953) );
  AOI22_X1 U14369 ( .A1(n12213), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11340) );
  NAND4_X1 U14370 ( .A1(n11343), .A2(n11342), .A3(n11341), .A4(n11340), .ZN(
        n11349) );
  AOI22_X1 U14371 ( .A1(n11318), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U14372 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14373 ( .A1(n12208), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9747), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U14374 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11344) );
  NAND4_X1 U14375 ( .A1(n11347), .A2(n11346), .A3(n11345), .A4(n11344), .ZN(
        n11348) );
  NAND2_X1 U14376 ( .A1(n13073), .A2(n11539), .ZN(n11353) );
  NOR2_X1 U14377 ( .A1(n11432), .A2(n11539), .ZN(n11394) );
  MUX2_X1 U14378 ( .A(n11536), .B(n11394), .S(n11415), .Z(n11350) );
  NAND2_X1 U14379 ( .A1(n11617), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11356) );
  OAI21_X1 U14380 ( .B1(n15945), .B2(n11415), .A(n11587), .ZN(n11354) );
  AND2_X1 U14381 ( .A1(n11354), .A2(n11353), .ZN(n11355) );
  XNOR2_X1 U14382 ( .A(n11391), .B(n11390), .ZN(n11927) );
  INV_X1 U14383 ( .A(n11642), .ZN(n11500) );
  OR2_X1 U14384 ( .A1(n11927), .A2(n11500), .ZN(n11359) );
  NAND2_X1 U14385 ( .A1(n13643), .A2(n11272), .ZN(n11417) );
  OAI21_X1 U14386 ( .B1(n20763), .B2(n11415), .A(n11417), .ZN(n11357) );
  INV_X1 U14387 ( .A(n11357), .ZN(n11358) );
  NAND2_X1 U14388 ( .A1(n13249), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11363) );
  INV_X1 U14389 ( .A(n19932), .ZN(n11361) );
  NAND2_X1 U14390 ( .A1(n11361), .A2(n11360), .ZN(n11362) );
  NAND2_X2 U14391 ( .A1(n11363), .A2(n11362), .ZN(n11422) );
  INV_X1 U14392 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11665) );
  INV_X1 U14393 ( .A(n11364), .ZN(n11365) );
  OAI21_X1 U14394 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11366), .A(
        n11365), .ZN(n11367) );
  XNOR2_X1 U14395 ( .A(n15552), .B(n20284), .ZN(n19987) );
  BUF_X1 U14396 ( .A(n11369), .Z(n11370) );
  NAND2_X1 U14397 ( .A1(n15579), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11371) );
  NAND2_X1 U14398 ( .A1(n11375), .A2(n11374), .ZN(n11425) );
  AOI22_X1 U14399 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11380) );
  AOI22_X1 U14400 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U14401 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14402 ( .A1(n12213), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11377) );
  NAND4_X1 U14403 ( .A1(n11380), .A2(n11379), .A3(n11378), .A4(n11377), .ZN(
        n11387) );
  AOI22_X1 U14404 ( .A1(n11318), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11385) );
  AOI22_X1 U14405 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U14406 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9747), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14407 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11382) );
  NAND4_X1 U14408 ( .A1(n11385), .A2(n11384), .A3(n11383), .A4(n11382), .ZN(
        n11386) );
  INV_X1 U14409 ( .A(n11617), .ZN(n11609) );
  INV_X1 U14410 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11388) );
  OAI22_X1 U14411 ( .A1(n11609), .A2(n11388), .B1(n11412), .B2(n11431), .ZN(
        n11389) );
  INV_X1 U14412 ( .A(n11408), .ZN(n11406) );
  NAND2_X1 U14413 ( .A1(n11391), .A2(n11390), .ZN(n11393) );
  INV_X1 U14414 ( .A(n11536), .ZN(n11392) );
  NAND2_X1 U14415 ( .A1(n11617), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11399) );
  INV_X1 U14416 ( .A(n11394), .ZN(n11395) );
  OAI21_X1 U14417 ( .B1(n11396), .B2(n11431), .A(n11395), .ZN(n11397) );
  INV_X1 U14418 ( .A(n11397), .ZN(n11398) );
  NAND2_X1 U14419 ( .A1(n11921), .A2(n11920), .ZN(n11404) );
  INV_X1 U14420 ( .A(n11400), .ZN(n11401) );
  NAND2_X1 U14421 ( .A1(n11404), .A2(n11403), .ZN(n11407) );
  INV_X1 U14422 ( .A(n11407), .ZN(n11405) );
  NAND2_X1 U14423 ( .A1(n11406), .A2(n11405), .ZN(n11448) );
  NAND2_X1 U14424 ( .A1(n11408), .A2(n11407), .ZN(n11409) );
  NAND2_X1 U14425 ( .A1(n11448), .A2(n11409), .ZN(n14973) );
  INV_X1 U14426 ( .A(n14973), .ZN(n11410) );
  NAND2_X1 U14427 ( .A1(n11410), .A2(n11642), .ZN(n11421) );
  NAND2_X1 U14428 ( .A1(n11414), .A2(n11415), .ZN(n11411) );
  NAND2_X1 U14429 ( .A1(n11412), .A2(n11411), .ZN(n11450) );
  NAND3_X1 U14430 ( .A1(n11415), .A2(n11414), .A3(n11413), .ZN(n11416) );
  NAND2_X1 U14431 ( .A1(n11450), .A2(n11416), .ZN(n11419) );
  INV_X1 U14432 ( .A(n11417), .ZN(n11418) );
  AOI21_X1 U14433 ( .B1(n15572), .B2(n11419), .A(n11418), .ZN(n11420) );
  NAND2_X1 U14434 ( .A1(n13384), .A2(n13385), .ZN(n11424) );
  NAND2_X1 U14435 ( .A1(n11422), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11423) );
  INV_X1 U14436 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19961) );
  INV_X1 U14437 ( .A(n11448), .ZN(n11447) );
  NAND2_X1 U14438 ( .A1(n11370), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11430) );
  INV_X1 U14439 ( .A(n15552), .ZN(n20398) );
  NAND2_X1 U14440 ( .A1(n20746), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20206) );
  INV_X1 U14441 ( .A(n20206), .ZN(n11426) );
  NAND2_X1 U14442 ( .A1(n20398), .A2(n11426), .ZN(n20278) );
  NAND2_X1 U14443 ( .A1(n20278), .A2(n20746), .ZN(n11428) );
  NAND2_X1 U14444 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20578) );
  INV_X1 U14445 ( .A(n20578), .ZN(n11427) );
  NAND2_X1 U14446 ( .A1(n20398), .A2(n11427), .ZN(n20640) );
  AOI22_X1 U14447 ( .A1(n20285), .A2(n12840), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15579), .ZN(n11429) );
  XNOR2_X2 U14448 ( .A(n13314), .B(n20127), .ZN(n20736) );
  AOI22_X1 U14449 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U14450 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14451 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14452 ( .A1(n13548), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11433) );
  NAND4_X1 U14453 ( .A1(n11436), .A2(n11435), .A3(n11434), .A4(n11433), .ZN(
        n11444) );
  AOI22_X1 U14454 ( .A1(n11318), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11442) );
  AOI22_X1 U14455 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U14456 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11440) );
  AOI22_X1 U14457 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9739), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11439) );
  NAND4_X1 U14458 ( .A1(n11442), .A2(n11441), .A3(n11440), .A4(n11439), .ZN(
        n11443) );
  AOI22_X1 U14459 ( .A1(n11617), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11598), .B2(n11451), .ZN(n11445) );
  INV_X1 U14460 ( .A(n20126), .ZN(n19979) );
  NAND2_X1 U14461 ( .A1(n11448), .A2(n19979), .ZN(n11449) );
  NAND2_X1 U14462 ( .A1(n11476), .A2(n11449), .ZN(n20735) );
  OR2_X1 U14463 ( .A1(n20735), .A2(n11500), .ZN(n11453) );
  NAND2_X1 U14464 ( .A1(n11450), .A2(n11451), .ZN(n11496) );
  OAI211_X1 U14465 ( .C1(n11451), .C2(n11450), .A(n11496), .B(n15572), .ZN(
        n11452) );
  NAND2_X1 U14466 ( .A1(n11453), .A2(n11452), .ZN(n13483) );
  NAND2_X1 U14467 ( .A1(n13482), .A2(n13483), .ZN(n11456) );
  NAND2_X1 U14468 ( .A1(n11454), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11455) );
  NAND2_X1 U14469 ( .A1(n11456), .A2(n11455), .ZN(n13598) );
  NAND2_X1 U14470 ( .A1(n11617), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11468) );
  AOI22_X1 U14471 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n9767), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14472 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12214), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11459) );
  AOI22_X1 U14473 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11458) );
  AOI22_X1 U14474 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13548), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11457) );
  NAND4_X1 U14475 ( .A1(n11460), .A2(n11459), .A3(n11458), .A4(n11457), .ZN(
        n11466) );
  AOI22_X1 U14476 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12155), .B1(
        n11318), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U14477 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U14478 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U14479 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11461) );
  NAND4_X1 U14480 ( .A1(n11464), .A2(n11463), .A3(n11462), .A4(n11461), .ZN(
        n11465) );
  NAND2_X1 U14481 ( .A1(n11598), .A2(n11494), .ZN(n11467) );
  NAND2_X1 U14482 ( .A1(n11468), .A2(n11467), .ZN(n11477) );
  XNOR2_X1 U14483 ( .A(n11476), .B(n11477), .ZN(n11953) );
  NAND2_X1 U14484 ( .A1(n11953), .A2(n11642), .ZN(n11471) );
  XNOR2_X1 U14485 ( .A(n11496), .B(n11494), .ZN(n11469) );
  NAND2_X1 U14486 ( .A1(n11469), .A2(n15572), .ZN(n11470) );
  NAND2_X1 U14487 ( .A1(n11471), .A2(n11470), .ZN(n11473) );
  INV_X1 U14488 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11472) );
  XNOR2_X1 U14489 ( .A(n11473), .B(n11472), .ZN(n13599) );
  NAND2_X1 U14490 ( .A1(n13598), .A2(n13599), .ZN(n11475) );
  NAND2_X1 U14491 ( .A1(n11473), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11474) );
  NAND2_X1 U14492 ( .A1(n11475), .A2(n11474), .ZN(n15788) );
  INV_X1 U14493 ( .A(n11476), .ZN(n11478) );
  INV_X1 U14494 ( .A(n11492), .ZN(n11490) );
  AOI22_X1 U14495 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U14496 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14497 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14498 ( .A1(n12213), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11479) );
  NAND4_X1 U14499 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(
        n11488) );
  AOI22_X1 U14500 ( .A1(n11318), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U14501 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14502 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11381), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14503 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11483) );
  NAND4_X1 U14504 ( .A1(n11486), .A2(n11485), .A3(n11484), .A4(n11483), .ZN(
        n11487) );
  AOI22_X1 U14505 ( .A1(n11617), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11598), .B2(n11497), .ZN(n11491) );
  NAND2_X1 U14506 ( .A1(n11492), .A2(n11491), .ZN(n11493) );
  NAND2_X1 U14507 ( .A1(n11518), .A2(n11493), .ZN(n11957) );
  INV_X1 U14508 ( .A(n11494), .ZN(n11495) );
  NOR2_X1 U14509 ( .A1(n11496), .A2(n11495), .ZN(n11498) );
  NAND2_X1 U14510 ( .A1(n11498), .A2(n11497), .ZN(n11527) );
  OAI211_X1 U14511 ( .C1(n11498), .C2(n11497), .A(n11527), .B(n15572), .ZN(
        n11499) );
  OAI21_X1 U14512 ( .B1(n11957), .B2(n11500), .A(n11499), .ZN(n11502) );
  INV_X1 U14513 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11501) );
  XNOR2_X1 U14514 ( .A(n11502), .B(n11501), .ZN(n15789) );
  NAND2_X1 U14515 ( .A1(n15788), .A2(n15789), .ZN(n11504) );
  NAND2_X1 U14516 ( .A1(n11502), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11503) );
  NAND2_X1 U14517 ( .A1(n11504), .A2(n11503), .ZN(n15781) );
  INV_X1 U14518 ( .A(n11518), .ZN(n11516) );
  AOI22_X1 U14519 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U14520 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11507) );
  INV_X1 U14521 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n21012) );
  AOI22_X1 U14522 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U14523 ( .A1(n13548), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11505) );
  NAND4_X1 U14524 ( .A1(n11508), .A2(n11507), .A3(n11506), .A4(n11505), .ZN(
        n11514) );
  AOI22_X1 U14525 ( .A1(n11318), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14526 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14527 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9747), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14528 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11509) );
  NAND4_X1 U14529 ( .A1(n11512), .A2(n11511), .A3(n11510), .A4(n11509), .ZN(
        n11513) );
  AOI22_X1 U14530 ( .A1(n11617), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11598), .B2(n11528), .ZN(n11517) );
  INV_X1 U14531 ( .A(n11517), .ZN(n11515) );
  NAND2_X2 U14532 ( .A1(n11516), .A2(n11515), .ZN(n11538) );
  NAND2_X1 U14533 ( .A1(n11518), .A2(n11517), .ZN(n11964) );
  NAND3_X1 U14534 ( .A1(n11538), .A2(n11642), .A3(n11964), .ZN(n11521) );
  XNOR2_X1 U14535 ( .A(n11527), .B(n11528), .ZN(n11519) );
  NAND2_X1 U14536 ( .A1(n11519), .A2(n15572), .ZN(n11520) );
  INV_X1 U14537 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15912) );
  NAND2_X1 U14538 ( .A1(n11522), .A2(n15912), .ZN(n15783) );
  INV_X1 U14539 ( .A(n11522), .ZN(n11523) );
  NAND2_X1 U14540 ( .A1(n11523), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15782) );
  INV_X1 U14541 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11525) );
  NAND2_X1 U14542 ( .A1(n11598), .A2(n11539), .ZN(n11524) );
  OAI21_X1 U14543 ( .B1(n11609), .B2(n11525), .A(n11524), .ZN(n11526) );
  NAND2_X1 U14544 ( .A1(n11915), .A2(n11642), .ZN(n11532) );
  INV_X1 U14545 ( .A(n11527), .ZN(n11529) );
  NAND2_X1 U14546 ( .A1(n11529), .A2(n11528), .ZN(n11541) );
  XNOR2_X1 U14547 ( .A(n11541), .B(n11539), .ZN(n11530) );
  NAND2_X1 U14548 ( .A1(n11530), .A2(n15572), .ZN(n11531) );
  NAND2_X1 U14549 ( .A1(n11532), .A2(n11531), .ZN(n11534) );
  XNOR2_X1 U14550 ( .A(n11534), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15774) );
  OR2_X1 U14551 ( .A1(n11534), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11535) );
  AND2_X1 U14552 ( .A1(n11536), .A2(n11642), .ZN(n11537) );
  NAND2_X1 U14553 ( .A1(n15572), .A2(n11539), .ZN(n11540) );
  OR2_X1 U14554 ( .A1(n11541), .A2(n11540), .ZN(n11542) );
  NAND2_X1 U14555 ( .A1(n15766), .A2(n11542), .ZN(n13844) );
  NOR2_X1 U14556 ( .A1(n13844), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11544) );
  NAND2_X1 U14557 ( .A1(n13844), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11543) );
  INV_X1 U14558 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14006) );
  NOR2_X1 U14559 ( .A1(n9736), .A2(n14006), .ZN(n11545) );
  NAND2_X1 U14560 ( .A1(n9736), .A2(n14006), .ZN(n11546) );
  INV_X1 U14561 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15751) );
  XNOR2_X1 U14562 ( .A(n15766), .B(n15751), .ZN(n14165) );
  NAND2_X1 U14563 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11547) );
  AND2_X1 U14564 ( .A1(n15766), .A2(n11547), .ZN(n14161) );
  INV_X1 U14565 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14162) );
  INV_X1 U14566 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21043) );
  AND2_X1 U14567 ( .A1(n9736), .A2(n21043), .ZN(n14849) );
  NOR2_X1 U14568 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11548) );
  INV_X1 U14569 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15831) );
  OR2_X1 U14570 ( .A1(n15766), .A2(n15831), .ZN(n14852) );
  XNOR2_X1 U14571 ( .A(n9737), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14959) );
  NAND2_X1 U14572 ( .A1(n9736), .A2(n15831), .ZN(n14957) );
  AND2_X1 U14573 ( .A1(n14959), .A2(n14957), .ZN(n11549) );
  INV_X1 U14574 ( .A(n14834), .ZN(n11552) );
  NAND2_X1 U14575 ( .A1(n11552), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11554) );
  NOR2_X1 U14576 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14160) );
  AND2_X1 U14577 ( .A1(n14160), .A2(n14162), .ZN(n11553) );
  NOR2_X1 U14578 ( .A1(n9736), .A2(n11553), .ZN(n14833) );
  XNOR2_X1 U14579 ( .A(n9737), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14828) );
  AND2_X1 U14580 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15586) );
  NAND2_X1 U14581 ( .A1(n14936), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11563) );
  INV_X1 U14582 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11557) );
  INV_X1 U14583 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14947) );
  INV_X1 U14584 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11556) );
  INV_X1 U14585 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15816) );
  NAND4_X1 U14586 ( .A1(n11557), .A2(n14947), .A3(n11556), .A4(n15816), .ZN(
        n11558) );
  INV_X1 U14587 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14929) );
  INV_X1 U14588 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14917) );
  NAND2_X1 U14589 ( .A1(n14929), .A2(n14917), .ZN(n14760) );
  INV_X1 U14590 ( .A(n14760), .ZN(n11560) );
  NAND2_X1 U14591 ( .A1(n11561), .A2(n11560), .ZN(n11562) );
  NAND2_X1 U14592 ( .A1(n11562), .A2(n10088), .ZN(n14784) );
  NAND3_X1 U14593 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14907) );
  NAND2_X1 U14594 ( .A1(n14757), .A2(n14907), .ZN(n11564) );
  NAND2_X1 U14595 ( .A1(n11563), .A2(n9737), .ZN(n14792) );
  NOR2_X1 U14596 ( .A1(n15766), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12935) );
  NOR2_X1 U14597 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14888) );
  NAND2_X1 U14598 ( .A1(n12935), .A2(n14888), .ZN(n11566) );
  AND2_X1 U14599 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14880) );
  INV_X1 U14600 ( .A(n14880), .ZN(n14889) );
  INV_X1 U14601 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14879) );
  NOR2_X1 U14602 ( .A1(n14889), .A2(n14879), .ZN(n11791) );
  AND2_X1 U14603 ( .A1(n15766), .A2(n11791), .ZN(n11565) );
  OAI21_X1 U14604 ( .B1(n12832), .B2(n11566), .A(n12937), .ZN(n11567) );
  XNOR2_X1 U14605 ( .A(n11567), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14756) );
  XNOR2_X1 U14606 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11593) );
  NAND2_X1 U14607 ( .A1(n11592), .A2(n11593), .ZN(n11569) );
  NAND2_X1 U14608 ( .A1(n20579), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11568) );
  NAND2_X1 U14609 ( .A1(n11569), .A2(n11568), .ZN(n11581) );
  XNOR2_X1 U14610 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11580) );
  NAND2_X1 U14611 ( .A1(n11581), .A2(n11580), .ZN(n11571) );
  NAND2_X1 U14612 ( .A1(n20284), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11570) );
  NAND2_X1 U14613 ( .A1(n11571), .A2(n11570), .ZN(n11579) );
  XNOR2_X1 U14614 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11578) );
  NAND2_X1 U14615 ( .A1(n11579), .A2(n11578), .ZN(n11573) );
  NAND2_X1 U14616 ( .A1(n20746), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11572) );
  NAND2_X1 U14617 ( .A1(n11573), .A2(n11572), .ZN(n11613) );
  NOR2_X1 U14618 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13318), .ZN(
        n11574) );
  INV_X1 U14619 ( .A(n11636), .ZN(n11577) );
  NAND2_X1 U14620 ( .A1(n11636), .A2(n11598), .ZN(n11623) );
  INV_X1 U14621 ( .A(n11588), .ZN(n11612) );
  XNOR2_X1 U14622 ( .A(n11579), .B(n11578), .ZN(n11633) );
  XNOR2_X1 U14623 ( .A(n11581), .B(n11580), .ZN(n11632) );
  INV_X1 U14624 ( .A(n11632), .ZN(n11582) );
  OR2_X1 U14625 ( .A1(n20006), .A2(n13643), .ZN(n11583) );
  NAND2_X1 U14626 ( .A1(n11583), .A2(n13256), .ZN(n11605) );
  INV_X1 U14627 ( .A(n11605), .ZN(n11584) );
  AOI211_X1 U14628 ( .C1(n11617), .C2(n11632), .A(n11604), .B(n11584), .ZN(
        n11608) );
  INV_X1 U14629 ( .A(n11592), .ZN(n11585) );
  OAI21_X1 U14630 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20471), .A(
        n11585), .ZN(n11589) );
  INV_X1 U14631 ( .A(n11589), .ZN(n11586) );
  OAI211_X1 U14632 ( .C1(n11273), .C2(n11587), .A(n11586), .B(n11605), .ZN(
        n11591) );
  INV_X1 U14633 ( .A(n11598), .ZN(n11594) );
  OAI21_X1 U14634 ( .B1(n11594), .B2(n11589), .A(n11588), .ZN(n11590) );
  NAND2_X1 U14635 ( .A1(n11591), .A2(n11590), .ZN(n11599) );
  INV_X1 U14636 ( .A(n11599), .ZN(n11603) );
  XNOR2_X1 U14637 ( .A(n11593), .B(n11592), .ZN(n11631) );
  NAND2_X1 U14638 ( .A1(n13072), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11596) );
  OAI21_X1 U14639 ( .B1(n11594), .B2(n13256), .A(n11596), .ZN(n11595) );
  AOI21_X1 U14640 ( .B1(n11617), .B2(n11631), .A(n11595), .ZN(n11600) );
  INV_X1 U14641 ( .A(n11600), .ZN(n11602) );
  NAND2_X1 U14642 ( .A1(n11596), .A2(n19992), .ZN(n11597) );
  AOI22_X1 U14643 ( .A1(n11631), .A2(n11614), .B1(n11600), .B2(n11599), .ZN(
        n11601) );
  AOI21_X1 U14644 ( .B1(n11603), .B2(n11602), .A(n11601), .ZN(n11607) );
  INV_X1 U14645 ( .A(n11604), .ZN(n11606) );
  OAI22_X1 U14646 ( .A1(n11608), .A2(n11607), .B1(n11606), .B2(n11605), .ZN(
        n11611) );
  NAND2_X1 U14647 ( .A1(n11609), .A2(n11633), .ZN(n11610) );
  AOI22_X1 U14648 ( .A1(n11612), .A2(n11633), .B1(n11611), .B2(n11610), .ZN(
        n11620) );
  NOR2_X1 U14649 ( .A1(n11617), .A2(n11615), .ZN(n11619) );
  INV_X1 U14650 ( .A(n11614), .ZN(n11616) );
  INV_X1 U14651 ( .A(n11615), .ZN(n11634) );
  NAND3_X1 U14652 ( .A1(n11617), .A2(n11616), .A3(n11634), .ZN(n11618) );
  OAI21_X1 U14653 ( .B1(n11620), .B2(n11619), .A(n11618), .ZN(n11621) );
  AOI21_X1 U14654 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n15945), .A(
        n11621), .ZN(n11622) );
  NAND2_X1 U14655 ( .A1(n11623), .A2(n11622), .ZN(n11624) );
  NAND2_X1 U14656 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20760) );
  OR2_X1 U14657 ( .A1(n11627), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n15604) );
  NAND2_X1 U14658 ( .A1(n13256), .A2(n15604), .ZN(n13641) );
  NAND3_X1 U14659 ( .A1(n11626), .A2(n20760), .A3(n13641), .ZN(n11629) );
  NAND3_X1 U14660 ( .A1(n11629), .A2(n19978), .A3(n11628), .ZN(n11630) );
  NAND2_X1 U14661 ( .A1(n13290), .A2(n11630), .ZN(n11639) );
  NOR4_X1 U14662 ( .A1(n11634), .A2(n11633), .A3(n11632), .A4(n11631), .ZN(
        n11635) );
  NOR2_X1 U14663 ( .A1(n11636), .A2(n11635), .ZN(n13077) );
  INV_X1 U14664 ( .A(n20760), .ZN(n20662) );
  AOI21_X1 U14665 ( .B1(n19992), .B2(n15604), .A(n20662), .ZN(n11637) );
  NAND2_X1 U14666 ( .A1(n13077), .A2(n11637), .ZN(n11638) );
  MUX2_X1 U14667 ( .A(n11639), .B(n11638), .S(n19996), .Z(n11647) );
  AOI21_X1 U14668 ( .B1(n14978), .B2(n13643), .A(n13076), .ZN(n11641) );
  NAND2_X1 U14669 ( .A1(n11641), .A2(n11772), .ZN(n12897) );
  INV_X1 U14670 ( .A(n12897), .ZN(n11645) );
  AND2_X1 U14671 ( .A1(n11642), .A2(n13071), .ZN(n11786) );
  NOR2_X1 U14672 ( .A1(n11786), .A2(n13643), .ZN(n11643) );
  NAND2_X1 U14673 ( .A1(n11644), .A2(n11643), .ZN(n11774) );
  OAI21_X1 U14674 ( .B1(n13079), .B2(n11645), .A(n11774), .ZN(n13283) );
  NOR2_X1 U14675 ( .A1(n13283), .A2(n12310), .ZN(n11646) );
  NAND2_X1 U14676 ( .A1(n11647), .A2(n11646), .ZN(n11648) );
  AND2_X1 U14677 ( .A1(n11273), .A2(n13638), .ZN(n11649) );
  OR2_X1 U14678 ( .A1(n12897), .A2(n11649), .ZN(n13074) );
  OAI21_X1 U14679 ( .B1(n13073), .B2(n11760), .A(n13074), .ZN(n11650) );
  OR2_X1 U14680 ( .A1(n11651), .A2(n11650), .ZN(n11652) );
  AOI22_X1 U14681 ( .A1(n14497), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n13069), .ZN(n14496) );
  INV_X1 U14682 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n11655) );
  INV_X1 U14683 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11656) );
  NAND2_X1 U14684 ( .A1(n11744), .A2(n11656), .ZN(n11657) );
  OAI211_X1 U14685 ( .C1(n13069), .C2(P1_EBX_REG_1__SCAN_IN), .A(n11657), .B(
        n11771), .ZN(n11658) );
  NAND2_X1 U14686 ( .A1(n11659), .A2(n11658), .ZN(n11663) );
  NAND2_X1 U14687 ( .A1(n11744), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11662) );
  INV_X1 U14688 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n11660) );
  NAND2_X1 U14689 ( .A1(n11771), .A2(n11660), .ZN(n11661) );
  NAND2_X1 U14690 ( .A1(n11662), .A2(n11661), .ZN(n13398) );
  INV_X1 U14691 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n11664) );
  NAND2_X1 U14692 ( .A1(n11744), .A2(n11665), .ZN(n11666) );
  OAI211_X1 U14693 ( .C1(n13069), .C2(P1_EBX_REG_2__SCAN_IN), .A(n11666), .B(
        n14495), .ZN(n11667) );
  AND2_X1 U14694 ( .A1(n11668), .A2(n11667), .ZN(n13389) );
  MUX2_X1 U14695 ( .A(n11748), .B(n13033), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n11670) );
  NOR2_X1 U14696 ( .A1(n14497), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11669) );
  NOR2_X1 U14697 ( .A1(n11670), .A2(n11669), .ZN(n13433) );
  NAND2_X1 U14698 ( .A1(n11752), .A2(n13069), .ZN(n11729) );
  NAND2_X1 U14699 ( .A1(n13069), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11671) );
  NAND2_X1 U14700 ( .A1(n11729), .A2(n11671), .ZN(n11672) );
  NOR2_X1 U14701 ( .A1(n11673), .A2(n11672), .ZN(n13579) );
  INV_X1 U14702 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n11674) );
  NAND2_X1 U14703 ( .A1(n11748), .A2(n11674), .ZN(n11677) );
  NAND2_X1 U14704 ( .A1(n11771), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11675) );
  OAI211_X1 U14705 ( .C1(n13069), .C2(P1_EBX_REG_5__SCAN_IN), .A(n11744), .B(
        n11675), .ZN(n11676) );
  NAND2_X1 U14706 ( .A1(n11677), .A2(n11676), .ZN(n13578) );
  INV_X1 U14707 ( .A(n11680), .ZN(n11683) );
  NAND2_X1 U14708 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13069), .ZN(
        n11681) );
  AND2_X1 U14709 ( .A1(n11729), .A2(n11681), .ZN(n11682) );
  NAND2_X1 U14710 ( .A1(n11683), .A2(n11682), .ZN(n13713) );
  INV_X1 U14711 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13716) );
  NAND2_X1 U14712 ( .A1(n11748), .A2(n13716), .ZN(n11686) );
  NAND2_X1 U14713 ( .A1(n14495), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11684) );
  OAI211_X1 U14714 ( .C1(n13069), .C2(P1_EBX_REG_7__SCAN_IN), .A(n11744), .B(
        n11684), .ZN(n11685) );
  AND2_X1 U14715 ( .A1(n11686), .A2(n11685), .ZN(n13712) );
  NAND2_X1 U14716 ( .A1(n13713), .A2(n13712), .ZN(n11687) );
  INV_X1 U14717 ( .A(n11688), .ZN(n11691) );
  NAND2_X1 U14718 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n13069), .ZN(
        n11689) );
  AND2_X1 U14719 ( .A1(n11729), .A2(n11689), .ZN(n11690) );
  NAND2_X1 U14720 ( .A1(n11691), .A2(n11690), .ZN(n13837) );
  INV_X1 U14721 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n11692) );
  NAND2_X1 U14722 ( .A1(n11748), .A2(n11692), .ZN(n11695) );
  NAND2_X1 U14723 ( .A1(n11771), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11693) );
  OAI211_X1 U14724 ( .C1(n13069), .C2(P1_EBX_REG_9__SCAN_IN), .A(n11744), .B(
        n11693), .ZN(n11694) );
  NAND2_X1 U14725 ( .A1(n11695), .A2(n11694), .ZN(n13830) );
  INV_X1 U14726 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15707) );
  INV_X1 U14727 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11696) );
  NAND2_X1 U14728 ( .A1(n11744), .A2(n11696), .ZN(n11697) );
  OAI211_X1 U14729 ( .C1(n13069), .C2(P1_EBX_REG_10__SCAN_IN), .A(n11697), .B(
        n11771), .ZN(n11698) );
  MUX2_X1 U14730 ( .A(n11748), .B(n13033), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n11700) );
  INV_X1 U14731 ( .A(n11700), .ZN(n11701) );
  NAND2_X1 U14732 ( .A1(n11701), .A2(n10070), .ZN(n14015) );
  INV_X1 U14733 ( .A(n11702), .ZN(n11705) );
  NAND2_X1 U14734 ( .A1(n13069), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11703) );
  AND2_X1 U14735 ( .A1(n11729), .A2(n11703), .ZN(n11704) );
  NAND2_X1 U14736 ( .A1(n11705), .A2(n11704), .ZN(n14673) );
  MUX2_X1 U14737 ( .A(n11748), .B(n13033), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n11707) );
  NOR2_X1 U14738 ( .A1(n14497), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11706) );
  NOR2_X1 U14739 ( .A1(n11707), .A2(n11706), .ZN(n14173) );
  INV_X1 U14740 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n11708) );
  NAND2_X1 U14741 ( .A1(n11744), .A2(n21043), .ZN(n11709) );
  OAI211_X1 U14742 ( .C1(n13069), .C2(P1_EBX_REG_14__SCAN_IN), .A(n11709), .B(
        n11771), .ZN(n11710) );
  MUX2_X1 U14743 ( .A(n11748), .B(n13033), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11712) );
  INV_X1 U14744 ( .A(n11712), .ZN(n11714) );
  INV_X1 U14745 ( .A(n14497), .ZN(n13400) );
  NAND2_X1 U14746 ( .A1(n13400), .A2(n15831), .ZN(n11713) );
  NAND2_X1 U14747 ( .A1(n11714), .A2(n11713), .ZN(n14594) );
  NOR3_X2 U14748 ( .A1(n14171), .A2(n14667), .A3(n14594), .ZN(n11715) );
  INV_X1 U14749 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14658) );
  INV_X1 U14750 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14832) );
  NAND2_X1 U14751 ( .A1(n11744), .A2(n14832), .ZN(n11716) );
  OAI211_X1 U14752 ( .C1(n13069), .C2(P1_EBX_REG_16__SCAN_IN), .A(n11716), .B(
        n11771), .ZN(n11717) );
  MUX2_X1 U14753 ( .A(n11748), .B(n13033), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n11720) );
  NOR2_X1 U14754 ( .A1(n14497), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11719) );
  NOR2_X1 U14755 ( .A1(n11720), .A2(n11719), .ZN(n14073) );
  INV_X1 U14756 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n20872) );
  NAND2_X1 U14757 ( .A1(n11744), .A2(n15816), .ZN(n11721) );
  OAI211_X1 U14758 ( .C1(n13069), .C2(P1_EBX_REG_18__SCAN_IN), .A(n11721), .B(
        n11771), .ZN(n11722) );
  INV_X1 U14759 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14583) );
  NAND2_X1 U14760 ( .A1(n11748), .A2(n14583), .ZN(n11726) );
  NAND2_X1 U14761 ( .A1(n11771), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11724) );
  OAI211_X1 U14762 ( .C1(n13069), .C2(P1_EBX_REG_19__SCAN_IN), .A(n11744), .B(
        n11724), .ZN(n11725) );
  NAND2_X1 U14763 ( .A1(n11726), .A2(n11725), .ZN(n14576) );
  INV_X1 U14764 ( .A(n11727), .ZN(n11731) );
  NAND2_X1 U14765 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n13069), .ZN(
        n11728) );
  AND2_X1 U14766 ( .A1(n11729), .A2(n11728), .ZN(n11730) );
  NAND2_X1 U14767 ( .A1(n11731), .A2(n11730), .ZN(n14633) );
  MUX2_X1 U14768 ( .A(n11748), .B(n13033), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n11733) );
  NOR2_X1 U14769 ( .A1(n14497), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11732) );
  NOR2_X1 U14770 ( .A1(n11733), .A2(n11732), .ZN(n14629) );
  INV_X1 U14771 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14625) );
  INV_X1 U14772 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14944) );
  NAND2_X1 U14773 ( .A1(n11744), .A2(n14944), .ZN(n11734) );
  OAI211_X1 U14774 ( .C1(n13069), .C2(P1_EBX_REG_22__SCAN_IN), .A(n11734), .B(
        n11771), .ZN(n11735) );
  AND2_X1 U14775 ( .A1(n11736), .A2(n11735), .ZN(n14622) );
  MUX2_X1 U14776 ( .A(n11748), .B(n13033), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n11737) );
  INV_X1 U14777 ( .A(n11737), .ZN(n11738) );
  NAND2_X1 U14778 ( .A1(n11738), .A2(n10077), .ZN(n14617) );
  INV_X1 U14779 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14610) );
  NAND2_X1 U14780 ( .A1(n11744), .A2(n14929), .ZN(n11739) );
  OAI211_X1 U14781 ( .C1(n13069), .C2(P1_EBX_REG_24__SCAN_IN), .A(n11739), .B(
        n11771), .ZN(n11740) );
  NAND2_X1 U14782 ( .A1(n11741), .A2(n11740), .ZN(n14607) );
  MUX2_X1 U14783 ( .A(n11748), .B(n13033), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n11743) );
  NOR2_X1 U14784 ( .A1(n14497), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11742) );
  NOR2_X1 U14785 ( .A1(n11743), .A2(n11742), .ZN(n14563) );
  INV_X1 U14786 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14602) );
  INV_X1 U14787 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14906) );
  NAND2_X1 U14788 ( .A1(n11744), .A2(n14906), .ZN(n11745) );
  OAI211_X1 U14789 ( .C1(n13069), .C2(P1_EBX_REG_26__SCAN_IN), .A(n11745), .B(
        n11771), .ZN(n11746) );
  AND2_X1 U14790 ( .A1(n11747), .A2(n11746), .ZN(n14548) );
  MUX2_X1 U14791 ( .A(n11748), .B(n13033), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n11749) );
  INV_X1 U14792 ( .A(n11749), .ZN(n11751) );
  INV_X1 U14793 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14775) );
  NAND2_X1 U14794 ( .A1(n13400), .A2(n14775), .ZN(n11750) );
  NAND2_X1 U14795 ( .A1(n11751), .A2(n11750), .ZN(n14539) );
  INV_X1 U14796 ( .A(n11753), .ZN(n11755) );
  NAND2_X1 U14797 ( .A1(n13069), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11754) );
  NAND2_X1 U14798 ( .A1(n11755), .A2(n11754), .ZN(n14519) );
  INV_X1 U14799 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n11756) );
  NAND2_X1 U14800 ( .A1(n13244), .A2(n11756), .ZN(n11757) );
  OAI21_X1 U14801 ( .B1(n14497), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11757), .ZN(n11758) );
  MUX2_X1 U14802 ( .A(n11757), .B(n11758), .S(n11771), .Z(n14476) );
  OAI22_X1 U14803 ( .A1(n14475), .A2(n11771), .B1(n14521), .B2(n11758), .ZN(
        n11759) );
  OR2_X1 U14804 ( .A1(n13065), .A2(n19992), .ZN(n13181) );
  OAI21_X1 U14805 ( .B1(n11760), .B2(n11277), .A(n13181), .ZN(n11761) );
  NAND2_X1 U14806 ( .A1(n19939), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14750) );
  OAI21_X1 U14807 ( .B1(n14516), .B2(n15909), .A(n14750), .ZN(n11762) );
  INV_X1 U14808 ( .A(n11762), .ZN(n11810) );
  NAND3_X1 U14809 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15810) );
  NOR3_X1 U14810 ( .A1(n15816), .A2(n21043), .A3(n15810), .ZN(n11793) );
  AND2_X1 U14811 ( .A1(n13079), .A2(n19992), .ZN(n15548) );
  INV_X1 U14812 ( .A(n13640), .ZN(n11763) );
  NAND2_X1 U14813 ( .A1(n11763), .A2(n11273), .ZN(n11764) );
  AND2_X1 U14814 ( .A1(n11765), .A2(n11764), .ZN(n11770) );
  INV_X1 U14815 ( .A(n20013), .ZN(n12903) );
  AOI21_X1 U14816 ( .B1(n13071), .B2(n19996), .A(n12903), .ZN(n11766) );
  NAND2_X1 U14817 ( .A1(n11767), .A2(n11766), .ZN(n11768) );
  NAND2_X1 U14818 ( .A1(n11768), .A2(n19992), .ZN(n11769) );
  OAI211_X1 U14819 ( .C1(n11772), .C2(n11771), .A(n11770), .B(n11769), .ZN(
        n11773) );
  INV_X1 U14820 ( .A(n11773), .ZN(n11775) );
  OAI211_X1 U14821 ( .C1(n11269), .C2(n13638), .A(n11775), .B(n11774), .ZN(
        n11776) );
  INV_X1 U14822 ( .A(n11776), .ZN(n13267) );
  MUX2_X1 U14823 ( .A(n11778), .B(n9731), .S(n19978), .Z(n11779) );
  NAND3_X1 U14824 ( .A1(n13267), .A2(n11780), .A3(n11779), .ZN(n11781) );
  NAND2_X1 U14825 ( .A1(n11795), .A2(n11781), .ZN(n15840) );
  NAND2_X1 U14826 ( .A1(n15848), .A2(n15840), .ZN(n15902) );
  INV_X1 U14827 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19933) );
  NAND2_X1 U14828 ( .A1(n19933), .A2(n15848), .ZN(n13252) );
  INV_X1 U14829 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11782) );
  INV_X1 U14830 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15915) );
  INV_X1 U14831 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15921) );
  NOR3_X1 U14832 ( .A1(n15915), .A2(n15921), .A3(n15912), .ZN(n15885) );
  NAND3_X1 U14833 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n15885), .ZN(n15863) );
  NOR2_X1 U14834 ( .A1(n11782), .A2(n15863), .ZN(n15868) );
  NAND2_X1 U14835 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15868), .ZN(
        n11784) );
  NAND2_X1 U14836 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19942) );
  INV_X1 U14837 ( .A(n19942), .ZN(n15901) );
  NAND4_X1 U14838 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A4(n15901), .ZN(n15862) );
  NOR2_X1 U14839 ( .A1(n11784), .A2(n15862), .ZN(n15853) );
  NAND2_X1 U14840 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15853), .ZN(
        n14961) );
  AOI21_X1 U14841 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19944) );
  NAND2_X1 U14842 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15901), .ZN(
        n11783) );
  NOR2_X1 U14843 ( .A1(n19944), .A2(n11783), .ZN(n15884) );
  INV_X1 U14844 ( .A(n11784), .ZN(n11792) );
  NAND2_X1 U14845 ( .A1(n15884), .A2(n11792), .ZN(n15843) );
  INV_X1 U14846 ( .A(n11786), .ZN(n11787) );
  NOR2_X1 U14847 ( .A1(n11785), .A2(n11787), .ZN(n13273) );
  INV_X1 U14848 ( .A(n15840), .ZN(n11794) );
  NAND3_X1 U14849 ( .A1(n11794), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n15853), .ZN(n11788) );
  OAI21_X1 U14850 ( .B1(n15843), .B2(n15865), .A(n11788), .ZN(n15839) );
  NAND2_X1 U14851 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15839), .ZN(
        n14949) );
  OAI21_X1 U14852 ( .B1(n15900), .B2(n14961), .A(n14949), .ZN(n14956) );
  NAND2_X1 U14853 ( .A1(n11793), .A2(n14956), .ZN(n15808) );
  INV_X1 U14854 ( .A(n15586), .ZN(n11789) );
  NOR2_X1 U14855 ( .A1(n15808), .A2(n11789), .ZN(n15593) );
  NAND3_X1 U14856 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n15593), .ZN(n15802) );
  INV_X1 U14857 ( .A(n15802), .ZN(n14916) );
  NAND2_X1 U14858 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n14916), .ZN(
        n11790) );
  NOR2_X1 U14859 ( .A1(n14907), .A2(n11790), .ZN(n14898) );
  NAND2_X1 U14860 ( .A1(n14898), .A2(n11791), .ZN(n14872) );
  INV_X1 U14861 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12938) );
  NAND2_X1 U14862 ( .A1(n14872), .A2(n12938), .ZN(n11808) );
  NAND2_X1 U14863 ( .A1(n15865), .A2(n15840), .ZN(n19967) );
  INV_X1 U14864 ( .A(n15848), .ZN(n19969) );
  INV_X1 U14865 ( .A(n15907), .ZN(n11807) );
  INV_X1 U14866 ( .A(n15884), .ZN(n14962) );
  NAND2_X1 U14867 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n11792), .ZN(
        n15833) );
  INV_X1 U14868 ( .A(n11793), .ZN(n11799) );
  NOR3_X1 U14869 ( .A1(n14962), .A2(n15833), .A3(n11799), .ZN(n11801) );
  NAND2_X1 U14870 ( .A1(n11794), .A2(n19933), .ZN(n11798) );
  INV_X1 U14871 ( .A(n11795), .ZN(n11796) );
  NAND2_X1 U14872 ( .A1(n11796), .A2(n15908), .ZN(n11797) );
  OAI21_X1 U14873 ( .B1(n11799), .B2(n14961), .A(n15902), .ZN(n11800) );
  OAI211_X1 U14874 ( .C1(n11801), .C2(n15865), .A(n15881), .B(n11800), .ZN(
        n15803) );
  INV_X1 U14875 ( .A(n15803), .ZN(n11802) );
  NAND2_X1 U14876 ( .A1(n11802), .A2(n15586), .ZN(n11803) );
  NAND2_X1 U14877 ( .A1(n11807), .A2(n15881), .ZN(n15882) );
  NOR2_X1 U14878 ( .A1(n11557), .A2(n14944), .ZN(n14938) );
  INV_X1 U14879 ( .A(n14938), .ZN(n11804) );
  AND2_X1 U14880 ( .A1(n15907), .A2(n11804), .ZN(n11805) );
  AND2_X1 U14881 ( .A1(n15907), .A2(n14907), .ZN(n11806) );
  NOR2_X1 U14882 ( .A1(n15796), .A2(n11806), .ZN(n14915) );
  NAND2_X1 U14883 ( .A1(n14915), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14912) );
  OAI21_X1 U14884 ( .B1(n14912), .B2(n14889), .A(n15882), .ZN(n14877) );
  OAI211_X1 U14885 ( .C1(n11807), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14877), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14868) );
  NAND2_X1 U14886 ( .A1(n11808), .A2(n14868), .ZN(n11809) );
  OAI211_X1 U14887 ( .C1(n14756), .C2(n15872), .A(n11810), .B(n11809), .ZN(
        P1_U3001) );
  NAND2_X1 U14888 ( .A1(n20244), .A2(n20516), .ZN(n12224) );
  INV_X1 U14889 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14822) );
  INV_X1 U14890 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12199) );
  INV_X1 U14891 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14796) );
  INV_X1 U14892 ( .A(n12280), .ZN(n11812) );
  INV_X1 U14893 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12843) );
  INV_X1 U14894 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14752) );
  XNOR2_X1 U14895 ( .A(n12941), .B(n14752), .ZN(n14748) );
  AOI22_X1 U14896 ( .A1(n12168), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U14897 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U14898 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U14899 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11813) );
  NAND4_X1 U14900 ( .A1(n11816), .A2(n11815), .A3(n11814), .A4(n11813), .ZN(
        n11822) );
  AOI22_X1 U14901 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11820) );
  AOI22_X1 U14902 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11819) );
  AOI22_X1 U14903 ( .A1(n11437), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11381), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11818) );
  AOI22_X1 U14904 ( .A1(n11305), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11817) );
  NAND4_X1 U14905 ( .A1(n11820), .A2(n11819), .A3(n11818), .A4(n11817), .ZN(
        n11821) );
  NOR2_X1 U14906 ( .A1(n11822), .A2(n11821), .ZN(n11907) );
  AOI22_X1 U14907 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U14908 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U14909 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U14910 ( .A1(n11437), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9739), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11823) );
  NAND4_X1 U14911 ( .A1(n11826), .A2(n11825), .A3(n11824), .A4(n11823), .ZN(
        n11832) );
  AOI22_X1 U14912 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U14913 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U14914 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U14915 ( .A1(n12168), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11827) );
  NAND4_X1 U14916 ( .A1(n11830), .A2(n11829), .A3(n11828), .A4(n11827), .ZN(
        n11831) );
  NOR2_X1 U14917 ( .A1(n11832), .A2(n11831), .ZN(n12295) );
  AOI22_X1 U14918 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12192), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U14919 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12168), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U14920 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n9746), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11834) );
  AOI22_X1 U14921 ( .A1(n12213), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11833) );
  NAND4_X1 U14922 ( .A1(n11836), .A2(n11835), .A3(n11834), .A4(n11833), .ZN(
        n11842) );
  AOI22_X1 U14923 ( .A1(n11437), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U14924 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12155), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U14925 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n9767), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U14926 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11837) );
  NAND4_X1 U14927 ( .A1(n11840), .A2(n11839), .A3(n11838), .A4(n11837), .ZN(
        n11841) );
  NOR2_X1 U14928 ( .A1(n11842), .A2(n11841), .ZN(n12273) );
  AOI22_X1 U14929 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U14930 ( .A1(n12168), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U14931 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U14932 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11843) );
  NAND4_X1 U14933 ( .A1(n11846), .A2(n11845), .A3(n11844), .A4(n11843), .ZN(
        n11852) );
  AOI22_X1 U14934 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U14935 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U14936 ( .A1(n11305), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U14937 ( .A1(n11318), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9747), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11847) );
  NAND4_X1 U14938 ( .A1(n11850), .A2(n11849), .A3(n11848), .A4(n11847), .ZN(
        n11851) );
  NOR2_X1 U14939 ( .A1(n11852), .A2(n11851), .ZN(n12254) );
  AOI22_X1 U14940 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U14941 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11855) );
  AOI22_X1 U14942 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n9746), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U14943 ( .A1(n11305), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11853) );
  NAND4_X1 U14944 ( .A1(n11856), .A2(n11855), .A3(n11854), .A4(n11853), .ZN(
        n11862) );
  AOI22_X1 U14945 ( .A1(n12168), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11318), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U14946 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11859) );
  AOI22_X1 U14947 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11858) );
  AOI22_X1 U14948 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11857) );
  NAND4_X1 U14949 ( .A1(n11860), .A2(n11859), .A3(n11858), .A4(n11857), .ZN(
        n11861) );
  NOR2_X1 U14950 ( .A1(n11862), .A2(n11861), .ZN(n12232) );
  AOI22_X1 U14951 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U14952 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U14953 ( .A1(n12168), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U14954 ( .A1(n11318), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11864) );
  NAND4_X1 U14955 ( .A1(n11867), .A2(n11866), .A3(n11865), .A4(n11864), .ZN(
        n11874) );
  AOI22_X1 U14956 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U14957 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U14958 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U14959 ( .A1(n12216), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9747), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11869) );
  NAND4_X1 U14960 ( .A1(n11872), .A2(n11871), .A3(n11870), .A4(n11869), .ZN(
        n11873) );
  NOR2_X1 U14961 ( .A1(n11874), .A2(n11873), .ZN(n12233) );
  NOR2_X1 U14962 ( .A1(n12232), .A2(n12233), .ZN(n12244) );
  AOI22_X1 U14963 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U14964 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U14965 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U14966 ( .A1(n12213), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11876) );
  NAND4_X1 U14967 ( .A1(n11879), .A2(n11878), .A3(n11877), .A4(n11876), .ZN(
        n11885) );
  AOI22_X1 U14968 ( .A1(n11318), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U14969 ( .A1(n12168), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U14970 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n9746), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U14971 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11880) );
  NAND4_X1 U14972 ( .A1(n11883), .A2(n11882), .A3(n11881), .A4(n11880), .ZN(
        n11884) );
  OR2_X1 U14973 ( .A1(n11885), .A2(n11884), .ZN(n12242) );
  NAND2_X1 U14974 ( .A1(n12244), .A2(n12242), .ZN(n12255) );
  NOR2_X1 U14975 ( .A1(n12254), .A2(n12255), .ZN(n12264) );
  AOI22_X1 U14976 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11889) );
  INV_X1 U14977 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n20867) );
  AOI22_X1 U14978 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11888) );
  AOI22_X1 U14979 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11887) );
  AOI22_X1 U14980 ( .A1(n12213), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11886) );
  NAND4_X1 U14981 ( .A1(n11889), .A2(n11888), .A3(n11887), .A4(n11886), .ZN(
        n11895) );
  AOI22_X1 U14982 ( .A1(n11437), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U14983 ( .A1(n12168), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U14984 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11381), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14985 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11890) );
  NAND4_X1 U14986 ( .A1(n11893), .A2(n11892), .A3(n11891), .A4(n11890), .ZN(
        n11894) );
  OR2_X1 U14987 ( .A1(n11895), .A2(n11894), .ZN(n12262) );
  NAND2_X1 U14988 ( .A1(n12264), .A2(n12262), .ZN(n12274) );
  NOR2_X1 U14989 ( .A1(n12273), .A2(n12274), .ZN(n12286) );
  AOI22_X1 U14990 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U14991 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11898) );
  AOI22_X1 U14992 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U14993 ( .A1(n12213), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11896) );
  NAND4_X1 U14994 ( .A1(n11899), .A2(n11898), .A3(n11897), .A4(n11896), .ZN(
        n11905) );
  AOI22_X1 U14995 ( .A1(n11318), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11903) );
  AOI22_X1 U14996 ( .A1(n12168), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11902) );
  AOI22_X1 U14997 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11381), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11901) );
  AOI22_X1 U14998 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11900) );
  NAND4_X1 U14999 ( .A1(n11903), .A2(n11902), .A3(n11901), .A4(n11900), .ZN(
        n11904) );
  OR2_X1 U15000 ( .A1(n11905), .A2(n11904), .ZN(n12284) );
  NAND2_X1 U15001 ( .A1(n12286), .A2(n12284), .ZN(n12296) );
  NOR2_X1 U15002 ( .A1(n12295), .A2(n12296), .ZN(n11906) );
  XOR2_X1 U15003 ( .A(n11907), .B(n11906), .Z(n11910) );
  AOI21_X1 U15004 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20244), .A(
        n12303), .ZN(n11909) );
  INV_X1 U15005 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20244) );
  NAND2_X1 U15006 ( .A1(n12892), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n11908) );
  OAI211_X1 U15007 ( .C1(n11910), .C2(n12234), .A(n11909), .B(n11908), .ZN(
        n11911) );
  OAI21_X1 U15008 ( .B1(n13633), .B2(n14748), .A(n11911), .ZN(n12308) );
  INV_X1 U15009 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13709) );
  OAI21_X1 U15010 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11958), .A(
        n11912), .ZN(n19812) );
  AOI22_X1 U15011 ( .A1(n12303), .A2(n19812), .B1(n12891), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11913) );
  OAI21_X1 U15012 ( .B1(n12300), .B2(n13709), .A(n11913), .ZN(n11914) );
  AOI21_X1 U15013 ( .B1(n11915), .B2(n12057), .A(n11914), .ZN(n13706) );
  INV_X1 U15014 ( .A(n13706), .ZN(n11965) );
  AND2_X1 U15015 ( .A1(n13436), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11945) );
  INV_X1 U15016 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n11917) );
  XNOR2_X1 U15017 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13667) );
  AOI21_X1 U15018 ( .B1(n12303), .B2(n13667), .A(n12891), .ZN(n11916) );
  OAI21_X1 U15019 ( .B1(n12300), .B2(n11917), .A(n11916), .ZN(n11918) );
  AOI21_X1 U15020 ( .B1(n11945), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11918), .ZN(n11919) );
  NAND2_X1 U15021 ( .A1(n12891), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11938) );
  NAND2_X1 U15022 ( .A1(n14970), .A2(n12057), .ZN(n11926) );
  INV_X1 U15023 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n11923) );
  INV_X1 U15024 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13660) );
  OAI22_X1 U15025 ( .A1(n12300), .A2(n11923), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13660), .ZN(n11924) );
  AOI21_X1 U15026 ( .B1(n11945), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11924), .ZN(n11925) );
  NAND2_X1 U15027 ( .A1(n11926), .A2(n11925), .ZN(n13243) );
  NAND2_X1 U15028 ( .A1(n20438), .A2(n13071), .ZN(n11928) );
  NAND2_X1 U15029 ( .A1(n11928), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13401) );
  INV_X1 U15030 ( .A(n11945), .ZN(n11933) );
  NAND2_X1 U15031 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11932) );
  NAND2_X1 U15032 ( .A1(n12892), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11931) );
  OAI211_X1 U15033 ( .C1(n11933), .C2(n11930), .A(n11932), .B(n11931), .ZN(
        n11934) );
  AOI21_X1 U15034 ( .B1(n20089), .B2(n12057), .A(n11934), .ZN(n11935) );
  OR2_X1 U15035 ( .A1(n13401), .A2(n11935), .ZN(n13402) );
  INV_X1 U15036 ( .A(n11935), .ZN(n13403) );
  OR2_X1 U15037 ( .A1(n13403), .A2(n12224), .ZN(n11936) );
  NAND2_X1 U15038 ( .A1(n13402), .A2(n11936), .ZN(n13242) );
  NAND2_X1 U15039 ( .A1(n13243), .A2(n13242), .ZN(n13414) );
  NAND2_X1 U15040 ( .A1(n13412), .A2(n11938), .ZN(n13431) );
  INV_X1 U15041 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n13440) );
  INV_X1 U15042 ( .A(n11939), .ZN(n11941) );
  INV_X1 U15043 ( .A(n11948), .ZN(n11940) );
  OAI21_X1 U15044 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11941), .A(
        n11940), .ZN(n13485) );
  AOI22_X1 U15045 ( .A1(n12303), .A2(n13485), .B1(n12891), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11942) );
  OAI21_X1 U15046 ( .B1(n12300), .B2(n13440), .A(n11942), .ZN(n11943) );
  AOI21_X1 U15047 ( .B1(n11945), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11943), .ZN(n11944) );
  NAND2_X1 U15048 ( .A1(n13431), .A2(n13430), .ZN(n13429) );
  NAND2_X1 U15049 ( .A1(n11945), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11951) );
  INV_X1 U15050 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19839) );
  AOI21_X1 U15051 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n19839), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11946) );
  AOI21_X1 U15052 ( .B1(n12892), .B2(P1_EAX_REG_4__SCAN_IN), .A(n11946), .ZN(
        n11950) );
  OAI21_X1 U15053 ( .B1(n11948), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11947), .ZN(n19852) );
  NOR2_X1 U15054 ( .A1(n13633), .A2(n19852), .ZN(n11949) );
  AOI21_X1 U15055 ( .B1(n11951), .B2(n11950), .A(n11949), .ZN(n11952) );
  OAI21_X1 U15056 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11954), .A(
        n11959), .ZN(n19835) );
  AOI22_X1 U15057 ( .A1(n12303), .A2(n19835), .B1(n12891), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11956) );
  NAND2_X1 U15058 ( .A1(n12892), .A2(P1_EAX_REG_5__SCAN_IN), .ZN(n11955) );
  NAND2_X1 U15059 ( .A1(n13527), .A2(n13576), .ZN(n13575) );
  INV_X1 U15060 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11962) );
  AOI21_X1 U15061 ( .B1(n11959), .B2(n19819), .A(n11958), .ZN(n15780) );
  INV_X1 U15062 ( .A(n12891), .ZN(n12073) );
  OAI22_X1 U15063 ( .A1(n15780), .A2(n13633), .B1(n12073), .B2(n19819), .ZN(
        n11960) );
  INV_X1 U15064 ( .A(n11960), .ZN(n11961) );
  OAI21_X1 U15065 ( .B1(n12300), .B2(n11962), .A(n11961), .ZN(n11963) );
  NAND2_X1 U15066 ( .A1(n11965), .A2(n13604), .ZN(n13705) );
  INV_X1 U15067 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13842) );
  XNOR2_X1 U15068 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11966), .ZN(
        n19793) );
  AOI22_X1 U15069 ( .A1(n12303), .A2(n19793), .B1(n12891), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11967) );
  OAI21_X1 U15070 ( .B1(n12300), .B2(n13842), .A(n11967), .ZN(n11968) );
  INV_X1 U15071 ( .A(n11968), .ZN(n11980) );
  AOI22_X1 U15072 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11318), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U15073 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U15074 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n9747), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11970) );
  AOI22_X1 U15075 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11969) );
  NAND4_X1 U15076 ( .A1(n11972), .A2(n11971), .A3(n11970), .A4(n11969), .ZN(
        n11978) );
  AOI22_X1 U15077 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15078 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U15079 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U15080 ( .A1(n11305), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9739), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11973) );
  NAND4_X1 U15081 ( .A1(n11976), .A2(n11975), .A3(n11974), .A4(n11973), .ZN(
        n11977) );
  OAI21_X1 U15082 ( .B1(n11978), .B2(n11977), .A(n12057), .ZN(n11979) );
  XOR2_X1 U15083 ( .A(n19779), .B(n11981), .Z(n19783) );
  AOI22_X1 U15084 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U15085 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U15086 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U15087 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11381), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11982) );
  NAND4_X1 U15088 ( .A1(n11985), .A2(n11984), .A3(n11983), .A4(n11982), .ZN(
        n11991) );
  AOI22_X1 U15089 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U15090 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U15091 ( .A1(n11318), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U15092 ( .A1(n13548), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11986) );
  NAND4_X1 U15093 ( .A1(n11989), .A2(n11988), .A3(n11987), .A4(n11986), .ZN(
        n11990) );
  OR2_X1 U15094 ( .A1(n11991), .A2(n11990), .ZN(n11992) );
  AOI22_X1 U15095 ( .A1(n12057), .A2(n11992), .B1(n12891), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11994) );
  NAND2_X1 U15096 ( .A1(n12892), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11993) );
  OAI211_X1 U15097 ( .C1(n19783), .C2(n13633), .A(n11994), .B(n11993), .ZN(
        n13828) );
  NAND2_X1 U15098 ( .A1(n13827), .A2(n13828), .ZN(n12024) );
  XNOR2_X1 U15099 ( .A(n11995), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15709) );
  NAND2_X1 U15100 ( .A1(n15709), .A2(n12303), .ZN(n12011) );
  AOI22_X1 U15101 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U15102 ( .A1(n12168), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U15103 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(n9747), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U15104 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11996) );
  NAND4_X1 U15105 ( .A1(n11999), .A2(n11998), .A3(n11997), .A4(n11996), .ZN(
        n12005) );
  AOI22_X1 U15106 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U15107 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11318), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U15108 ( .A1(n11376), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U15109 ( .A1(n11305), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12000) );
  NAND4_X1 U15110 ( .A1(n12003), .A2(n12002), .A3(n12001), .A4(n12000), .ZN(
        n12004) );
  NOR2_X1 U15111 ( .A1(n12005), .A2(n12004), .ZN(n12008) );
  NAND2_X1 U15112 ( .A1(n12892), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12007) );
  NAND2_X1 U15113 ( .A1(n12891), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12006) );
  OAI211_X1 U15114 ( .C1(n12126), .C2(n12008), .A(n12007), .B(n12006), .ZN(
        n12009) );
  INV_X1 U15115 ( .A(n12009), .ZN(n12010) );
  NAND2_X1 U15116 ( .A1(n12011), .A2(n12010), .ZN(n13924) );
  NOR2_X2 U15117 ( .A1(n12024), .A2(n12012), .ZN(n13925) );
  AOI22_X1 U15118 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U15119 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U15120 ( .A1(n12168), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U15121 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11381), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12013) );
  NAND4_X1 U15122 ( .A1(n12016), .A2(n12015), .A3(n12014), .A4(n12013), .ZN(
        n12022) );
  AOI22_X1 U15123 ( .A1(n11318), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U15124 ( .A1(n13548), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U15125 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U15126 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12017) );
  NAND4_X1 U15127 ( .A1(n12020), .A2(n12019), .A3(n12018), .A4(n12017), .ZN(
        n12021) );
  OR2_X1 U15128 ( .A1(n12022), .A2(n12021), .ZN(n12023) );
  NAND2_X1 U15129 ( .A1(n13925), .A2(n14152), .ZN(n12028) );
  INV_X1 U15130 ( .A(n12024), .ZN(n13826) );
  INV_X1 U15131 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14019) );
  OAI21_X1 U15132 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12025), .A(
        n12040), .ZN(n15773) );
  AOI22_X1 U15133 ( .A1(n12303), .A2(n15773), .B1(n12891), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12026) );
  OAI21_X1 U15134 ( .B1(n12300), .B2(n14019), .A(n12026), .ZN(n14012) );
  AND2_X1 U15135 ( .A1(n13924), .A2(n14012), .ZN(n12027) );
  NAND2_X1 U15136 ( .A1(n13826), .A2(n12027), .ZN(n14153) );
  INV_X1 U15137 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U15138 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12168), .B1(
        n11318), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U15139 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U15140 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12207), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U15141 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(n9747), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12029) );
  NAND4_X1 U15142 ( .A1(n12032), .A2(n12031), .A3(n12030), .A4(n12029), .ZN(
        n12038) );
  AOI22_X1 U15143 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n9767), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U15144 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n13548), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U15145 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12173), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U15146 ( .A1(n12135), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12033) );
  NAND4_X1 U15147 ( .A1(n12036), .A2(n12035), .A3(n12034), .A4(n12033), .ZN(
        n12037) );
  OR2_X1 U15148 ( .A1(n12038), .A2(n12037), .ZN(n12039) );
  NAND2_X1 U15149 ( .A1(n12057), .A2(n12039), .ZN(n12044) );
  XNOR2_X1 U15150 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12040), .ZN(
        n15762) );
  OAI22_X1 U15151 ( .A1(n15762), .A2(n13633), .B1(n12073), .B2(n12041), .ZN(
        n12042) );
  INV_X1 U15152 ( .A(n12042), .ZN(n12043) );
  OAI211_X1 U15153 ( .C1(n12045), .C2(n12300), .A(n12044), .B(n12043), .ZN(
        n14677) );
  INV_X1 U15154 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15155 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15156 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12048) );
  AOI22_X1 U15157 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9739), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12047) );
  AOI22_X1 U15158 ( .A1(n12135), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12046) );
  NAND4_X1 U15159 ( .A1(n12049), .A2(n12048), .A3(n12047), .A4(n12046), .ZN(
        n12055) );
  AOI22_X1 U15160 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U15161 ( .A1(n11318), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U15162 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11381), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U15163 ( .A1(n12168), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12050) );
  NAND4_X1 U15164 ( .A1(n12053), .A2(n12052), .A3(n12051), .A4(n12050), .ZN(
        n12054) );
  OR2_X1 U15165 ( .A1(n12055), .A2(n12054), .ZN(n12056) );
  NAND2_X1 U15166 ( .A1(n12057), .A2(n12056), .ZN(n12061) );
  XNOR2_X1 U15167 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12058), .ZN(
        n14183) );
  OAI22_X1 U15168 ( .A1(n13633), .A2(n14183), .B1(n12073), .B2(n14177), .ZN(
        n12059) );
  INV_X1 U15169 ( .A(n12059), .ZN(n12060) );
  OAI211_X1 U15170 ( .C1(n12300), .C2(n12062), .A(n12061), .B(n12060), .ZN(
        n14158) );
  AOI22_X1 U15171 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9767), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U15172 ( .A1(n12168), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15173 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U15174 ( .A1(n12216), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9739), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12063) );
  NAND4_X1 U15175 ( .A1(n12066), .A2(n12065), .A3(n12064), .A4(n12063), .ZN(
        n12072) );
  AOI22_X1 U15176 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U15177 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15178 ( .A1(n11318), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15179 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n9746), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12067) );
  NAND4_X1 U15180 ( .A1(n12070), .A2(n12069), .A3(n12068), .A4(n12067), .ZN(
        n12071) );
  NOR2_X1 U15181 ( .A1(n12072), .A2(n12071), .ZN(n12076) );
  XNOR2_X1 U15182 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12092), .ZN(
        n14845) );
  OAI22_X1 U15183 ( .A1(n13633), .A2(n14845), .B1(n12073), .B2(n14841), .ZN(
        n12074) );
  AOI21_X1 U15184 ( .B1(n12892), .B2(P1_EAX_REG_17__SCAN_IN), .A(n12074), .ZN(
        n12075) );
  OAI21_X1 U15185 ( .B1(n12234), .B2(n12076), .A(n12075), .ZN(n14072) );
  AOI22_X1 U15186 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9767), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U15187 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15188 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15189 ( .A1(n11305), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12077) );
  NAND4_X1 U15190 ( .A1(n12080), .A2(n12079), .A3(n12078), .A4(n12077), .ZN(
        n12086) );
  AOI22_X1 U15191 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U15192 ( .A1(n11318), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15193 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11381), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15194 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12081) );
  NAND4_X1 U15195 ( .A1(n12084), .A2(n12083), .A3(n12082), .A4(n12081), .ZN(
        n12085) );
  NOR2_X1 U15196 ( .A1(n12086), .A2(n12085), .ZN(n12091) );
  INV_X1 U15197 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12088) );
  NAND2_X1 U15198 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12087) );
  OAI211_X1 U15199 ( .C1(n12300), .C2(n12088), .A(n13633), .B(n12087), .ZN(
        n12089) );
  INV_X1 U15200 ( .A(n12089), .ZN(n12090) );
  OAI21_X1 U15201 ( .B1(n12234), .B2(n12091), .A(n12090), .ZN(n12095) );
  OAI21_X1 U15202 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12093), .A(
        n12092), .ZN(n15749) );
  OR2_X1 U15203 ( .A1(n13633), .A2(n15749), .ZN(n12094) );
  NAND2_X1 U15204 ( .A1(n12095), .A2(n12094), .ZN(n14650) );
  XNOR2_X1 U15205 ( .A(n12097), .B(n12096), .ZN(n14856) );
  AOI22_X1 U15206 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U15207 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U15208 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11318), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12099) );
  AOI22_X1 U15209 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12098) );
  NAND4_X1 U15210 ( .A1(n12101), .A2(n12100), .A3(n12099), .A4(n12098), .ZN(
        n12107) );
  AOI22_X1 U15211 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U15212 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U15213 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U15214 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9746), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12102) );
  NAND4_X1 U15215 ( .A1(n12105), .A2(n12104), .A3(n12103), .A4(n12102), .ZN(
        n12106) );
  NOR2_X1 U15216 ( .A1(n12107), .A2(n12106), .ZN(n12110) );
  NAND2_X1 U15217 ( .A1(n12892), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12109) );
  NAND2_X1 U15218 ( .A1(n12891), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12108) );
  OAI211_X1 U15219 ( .C1(n12126), .C2(n12110), .A(n12109), .B(n12108), .ZN(
        n12111) );
  AOI21_X1 U15220 ( .B1(n14856), .B2(n12303), .A(n12111), .ZN(n14589) );
  OR2_X1 U15221 ( .A1(n14650), .A2(n14589), .ZN(n12129) );
  XOR2_X1 U15222 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n12112), .Z(
        n15754) );
  INV_X1 U15223 ( .A(n15754), .ZN(n12128) );
  AOI22_X1 U15224 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11376), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U15225 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11318), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U15226 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12114) );
  AOI22_X1 U15227 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9746), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12113) );
  NAND4_X1 U15228 ( .A1(n12116), .A2(n12115), .A3(n12114), .A4(n12113), .ZN(
        n12122) );
  AOI22_X1 U15229 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12120) );
  AOI22_X1 U15230 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15231 ( .A1(n13548), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12118) );
  AOI22_X1 U15232 ( .A1(n12216), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12117) );
  NAND4_X1 U15233 ( .A1(n12120), .A2(n12119), .A3(n12118), .A4(n12117), .ZN(
        n12121) );
  NOR2_X1 U15234 ( .A1(n12122), .A2(n12121), .ZN(n12125) );
  NAND2_X1 U15235 ( .A1(n12892), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12124) );
  NAND2_X1 U15236 ( .A1(n12891), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12123) );
  OAI211_X1 U15237 ( .C1(n12126), .C2(n12125), .A(n12124), .B(n12123), .ZN(
        n12127) );
  AOI21_X1 U15238 ( .B1(n12128), .B2(n12303), .A(n12127), .ZN(n14663) );
  NOR2_X1 U15239 ( .A1(n12129), .A2(n14663), .ZN(n14069) );
  AOI22_X1 U15240 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12214), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15241 ( .A1(n12168), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15242 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n9746), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12132) );
  AOI22_X1 U15243 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12131) );
  NAND4_X1 U15244 ( .A1(n12134), .A2(n12133), .A3(n12132), .A4(n12131), .ZN(
        n12141) );
  AOI22_X1 U15245 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U15246 ( .A1(n11376), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15247 ( .A1(n13548), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U15248 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12136) );
  NAND4_X1 U15249 ( .A1(n12139), .A2(n12138), .A3(n12137), .A4(n12136), .ZN(
        n12140) );
  NOR2_X1 U15250 ( .A1(n12141), .A2(n12140), .ZN(n12145) );
  INV_X1 U15251 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14729) );
  NAND2_X1 U15252 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12142) );
  OAI211_X1 U15253 ( .C1(n12300), .C2(n14729), .A(n13633), .B(n12142), .ZN(
        n12143) );
  INV_X1 U15254 ( .A(n12143), .ZN(n12144) );
  OAI21_X1 U15255 ( .B1(n12234), .B2(n12145), .A(n12144), .ZN(n12148) );
  OAI21_X1 U15256 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12146), .A(
        n12165), .ZN(n15667) );
  OR2_X1 U15257 ( .A1(n13633), .A2(n15667), .ZN(n12147) );
  NAND2_X1 U15258 ( .A1(n12148), .A2(n12147), .ZN(n14643) );
  NAND2_X1 U15259 ( .A1(n12150), .A2(n12149), .ZN(n14573) );
  AOI22_X1 U15260 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U15261 ( .A1(n12168), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U15262 ( .A1(n13548), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15263 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12151) );
  NAND4_X1 U15264 ( .A1(n12154), .A2(n12153), .A3(n12152), .A4(n12151), .ZN(
        n12161) );
  AOI22_X1 U15265 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15266 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15267 ( .A1(n12155), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U15268 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n9747), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12156) );
  NAND4_X1 U15269 ( .A1(n12159), .A2(n12158), .A3(n12157), .A4(n12156), .ZN(
        n12160) );
  NOR2_X1 U15270 ( .A1(n12161), .A2(n12160), .ZN(n12164) );
  AOI21_X1 U15271 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14822), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12162) );
  AOI21_X1 U15272 ( .B1(n12892), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12162), .ZN(
        n12163) );
  OAI21_X1 U15273 ( .B1(n12234), .B2(n12164), .A(n12163), .ZN(n12167) );
  XNOR2_X1 U15274 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n12165), .ZN(
        n14824) );
  NAND2_X1 U15275 ( .A1(n12303), .A2(n14824), .ZN(n12166) );
  NAND2_X1 U15276 ( .A1(n12167), .A2(n12166), .ZN(n14572) );
  AOI22_X1 U15277 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12214), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15278 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U15279 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n9747), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U15280 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12168), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12169) );
  NAND4_X1 U15281 ( .A1(n12172), .A2(n12171), .A3(n12170), .A4(n12169), .ZN(
        n12179) );
  AOI22_X1 U15282 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n9767), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U15283 ( .A1(n13548), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U15284 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12175) );
  AOI22_X1 U15285 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12135), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12174) );
  NAND4_X1 U15286 ( .A1(n12177), .A2(n12176), .A3(n12175), .A4(n12174), .ZN(
        n12178) );
  NOR2_X1 U15287 ( .A1(n12179), .A2(n12178), .ZN(n12184) );
  INV_X1 U15288 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n12181) );
  NAND2_X1 U15289 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12180) );
  OAI211_X1 U15290 ( .C1(n12300), .C2(n12181), .A(n13633), .B(n12180), .ZN(
        n12182) );
  INV_X1 U15291 ( .A(n12182), .ZN(n12183) );
  OAI21_X1 U15292 ( .B1(n12234), .B2(n12184), .A(n12183), .ZN(n12187) );
  OAI21_X1 U15293 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12185), .A(
        n12203), .ZN(n15744) );
  OR2_X1 U15294 ( .A1(n13633), .A2(n15744), .ZN(n12186) );
  AND2_X2 U15295 ( .A1(n14574), .A2(n14637), .ZN(n14630) );
  AOI22_X1 U15296 ( .A1(n13548), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15297 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15298 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15299 ( .A1(n11336), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12215), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12188) );
  NAND4_X1 U15300 ( .A1(n12191), .A2(n12190), .A3(n12189), .A4(n12188), .ZN(
        n12198) );
  AOI22_X1 U15301 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U15302 ( .A1(n12168), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15303 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12216), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15304 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11381), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12193) );
  NAND4_X1 U15305 ( .A1(n12196), .A2(n12195), .A3(n12194), .A4(n12193), .ZN(
        n12197) );
  NOR2_X1 U15306 ( .A1(n12198), .A2(n12197), .ZN(n12202) );
  OAI21_X1 U15307 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n12199), .A(n13633), 
        .ZN(n12200) );
  AOI21_X1 U15308 ( .B1(n12892), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12200), .ZN(
        n12201) );
  OAI21_X1 U15309 ( .B1(n12234), .B2(n12202), .A(n12201), .ZN(n12205) );
  XNOR2_X1 U15310 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12203), .ZN(
        n15734) );
  NAND2_X1 U15311 ( .A1(n12303), .A2(n15734), .ZN(n12204) );
  AOI22_X1 U15312 ( .A1(n11875), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15313 ( .A1(n11318), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12155), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U15314 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15315 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11381), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12209) );
  NAND4_X1 U15316 ( .A1(n12212), .A2(n12211), .A3(n12210), .A4(n12209), .ZN(
        n12222) );
  AOI22_X1 U15317 ( .A1(n12168), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9767), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15318 ( .A1(n12213), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11305), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12219) );
  AOI22_X1 U15319 ( .A1(n12214), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15320 ( .A1(n12216), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9739), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12217) );
  NAND4_X1 U15321 ( .A1(n12220), .A2(n12219), .A3(n12218), .A4(n12217), .ZN(
        n12221) );
  NOR2_X1 U15322 ( .A1(n12222), .A2(n12221), .ZN(n12227) );
  INV_X1 U15323 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14717) );
  NAND2_X1 U15324 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12223) );
  OAI211_X1 U15325 ( .C1(n12300), .C2(n14717), .A(n12224), .B(n12223), .ZN(
        n12225) );
  INV_X1 U15326 ( .A(n12225), .ZN(n12226) );
  OAI21_X1 U15327 ( .B1(n12234), .B2(n12227), .A(n12226), .ZN(n12230) );
  OAI21_X1 U15328 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12228), .A(
        n12239), .ZN(n15733) );
  OR2_X1 U15329 ( .A1(n13633), .A2(n15733), .ZN(n12229) );
  NAND2_X1 U15330 ( .A1(n12230), .A2(n12229), .ZN(n14620) );
  XOR2_X1 U15331 ( .A(n12233), .B(n12232), .Z(n12235) );
  NAND2_X1 U15332 ( .A1(n12235), .A2(n12297), .ZN(n12238) );
  INV_X1 U15333 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15634) );
  OAI21_X1 U15334 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15634), .A(n13633), 
        .ZN(n12236) );
  AOI21_X1 U15335 ( .B1(n12892), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12236), .ZN(
        n12237) );
  NAND2_X1 U15336 ( .A1(n12238), .A2(n12237), .ZN(n12241) );
  XNOR2_X1 U15337 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n12239), .ZN(
        n15624) );
  NAND2_X1 U15338 ( .A1(n12303), .A2(n15624), .ZN(n12240) );
  NAND2_X1 U15339 ( .A1(n12241), .A2(n12240), .ZN(n14614) );
  INV_X1 U15340 ( .A(n12242), .ZN(n12243) );
  XNOR2_X1 U15341 ( .A(n12244), .B(n12243), .ZN(n12245) );
  NAND2_X1 U15342 ( .A1(n12245), .A2(n12297), .ZN(n12253) );
  INV_X1 U15343 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14710) );
  NAND2_X1 U15344 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12246) );
  OAI211_X1 U15345 ( .C1(n12300), .C2(n14710), .A(n13633), .B(n12246), .ZN(
        n12247) );
  INV_X1 U15346 ( .A(n12247), .ZN(n12252) );
  INV_X1 U15347 ( .A(n12248), .ZN(n12249) );
  INV_X1 U15348 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14809) );
  NAND2_X1 U15349 ( .A1(n12249), .A2(n14809), .ZN(n12250) );
  NAND2_X1 U15350 ( .A1(n12258), .A2(n12250), .ZN(n15623) );
  NOR2_X1 U15351 ( .A1(n15623), .A2(n13633), .ZN(n12251) );
  AOI21_X1 U15352 ( .B1(n12253), .B2(n12252), .A(n12251), .ZN(n14605) );
  XOR2_X1 U15353 ( .A(n12255), .B(n12254), .Z(n12256) );
  NAND2_X1 U15354 ( .A1(n12256), .A2(n12297), .ZN(n12261) );
  OAI21_X1 U15355 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14796), .A(n13633), 
        .ZN(n12257) );
  AOI21_X1 U15356 ( .B1(n12892), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12257), .ZN(
        n12260) );
  XNOR2_X1 U15357 ( .A(n12258), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14800) );
  INV_X1 U15358 ( .A(n12262), .ZN(n12263) );
  XNOR2_X1 U15359 ( .A(n12264), .B(n12263), .ZN(n12267) );
  INV_X1 U15360 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14701) );
  NAND2_X1 U15361 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12265) );
  OAI211_X1 U15362 ( .C1(n12300), .C2(n14701), .A(n13633), .B(n12265), .ZN(
        n12266) );
  AOI21_X1 U15363 ( .B1(n12267), .B2(n12297), .A(n12266), .ZN(n12272) );
  INV_X1 U15364 ( .A(n12268), .ZN(n12269) );
  INV_X1 U15365 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14788) );
  NAND2_X1 U15366 ( .A1(n12269), .A2(n14788), .ZN(n12270) );
  NAND2_X1 U15367 ( .A1(n12280), .A2(n12270), .ZN(n14551) );
  NOR2_X1 U15368 ( .A1(n14551), .A2(n13633), .ZN(n12271) );
  XOR2_X1 U15369 ( .A(n12274), .B(n12273), .Z(n12275) );
  NAND2_X1 U15370 ( .A1(n12275), .A2(n12297), .ZN(n12279) );
  INV_X1 U15371 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14696) );
  NAND2_X1 U15372 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12276) );
  OAI211_X1 U15373 ( .C1(n12300), .C2(n14696), .A(n13633), .B(n12276), .ZN(
        n12277) );
  INV_X1 U15374 ( .A(n12277), .ZN(n12278) );
  NAND2_X1 U15375 ( .A1(n12279), .A2(n12278), .ZN(n12282) );
  XNOR2_X1 U15376 ( .A(n12280), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14777) );
  NAND2_X1 U15377 ( .A1(n14777), .A2(n12303), .ZN(n12281) );
  NAND2_X1 U15378 ( .A1(n12282), .A2(n12281), .ZN(n14534) );
  INV_X1 U15379 ( .A(n12284), .ZN(n12285) );
  XNOR2_X1 U15380 ( .A(n12286), .B(n12285), .ZN(n12289) );
  INV_X1 U15381 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14691) );
  NAND2_X1 U15382 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12287) );
  OAI211_X1 U15383 ( .C1(n12300), .C2(n14691), .A(n13633), .B(n12287), .ZN(
        n12288) );
  AOI21_X1 U15384 ( .B1(n12289), .B2(n12297), .A(n12288), .ZN(n12294) );
  INV_X1 U15385 ( .A(n12290), .ZN(n12291) );
  INV_X1 U15386 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14768) );
  NAND2_X1 U15387 ( .A1(n12291), .A2(n14768), .ZN(n12292) );
  NAND2_X1 U15388 ( .A1(n12302), .A2(n12292), .ZN(n14522) );
  NOR2_X1 U15389 ( .A1(n14522), .A2(n13633), .ZN(n12293) );
  XOR2_X1 U15390 ( .A(n12296), .B(n12295), .Z(n12298) );
  NAND2_X1 U15391 ( .A1(n12298), .A2(n12297), .ZN(n12306) );
  INV_X1 U15392 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14487) );
  OAI21_X1 U15393 ( .B1(n20516), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n20244), .ZN(n12299) );
  OAI21_X1 U15394 ( .B1(n12300), .B2(n14487), .A(n12299), .ZN(n12301) );
  INV_X1 U15395 ( .A(n12301), .ZN(n12305) );
  XNOR2_X1 U15396 ( .A(n12302), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14479) );
  INV_X1 U15397 ( .A(n14754), .ZN(n14690) );
  INV_X1 U15398 ( .A(n11785), .ZN(n12309) );
  NAND2_X1 U15399 ( .A1(n12310), .A2(n12309), .ZN(n13284) );
  INV_X1 U15400 ( .A(n12311), .ZN(n12312) );
  NAND4_X1 U15401 ( .A1(n12312), .A2(n13268), .A3(n13073), .A4(n12903), .ZN(
        n12899) );
  INV_X1 U15402 ( .A(n12899), .ZN(n12313) );
  NAND2_X1 U15403 ( .A1(n12313), .A2(n13244), .ZN(n12314) );
  INV_X1 U15404 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n12316) );
  INV_X1 U15405 ( .A(n12317), .ZN(n12318) );
  INV_X1 U15406 ( .A(n15366), .ZN(n15248) );
  OR2_X1 U15407 ( .A1(n20857), .A2(n15344), .ZN(n12319) );
  NOR2_X1 U15408 ( .A1(n15337), .A2(n12319), .ZN(n12320) );
  NOR2_X1 U15409 ( .A1(n12947), .A2(n19074), .ZN(n12347) );
  INV_X1 U15410 ( .A(n15396), .ZN(n16029) );
  INV_X1 U15411 ( .A(n16028), .ZN(n12321) );
  NAND2_X1 U15412 ( .A1(n12325), .A2(n15399), .ZN(n15374) );
  INV_X1 U15413 ( .A(n15371), .ZN(n12326) );
  INV_X1 U15414 ( .A(n15355), .ZN(n12327) );
  INV_X1 U15415 ( .A(n12328), .ZN(n15242) );
  NAND2_X1 U15416 ( .A1(n15230), .A2(n12331), .ZN(n12723) );
  NAND2_X1 U15417 ( .A1(n12722), .A2(n12332), .ZN(n12333) );
  XNOR2_X1 U15418 ( .A(n12723), .B(n12333), .ZN(n12952) );
  OR2_X1 U15419 ( .A1(n13951), .A2(n12335), .ZN(n12336) );
  NAND2_X1 U15420 ( .A1(n12334), .A2(n12336), .ZN(n15991) );
  OAI21_X1 U15421 ( .B1(n12337), .B2(n15285), .A(n15364), .ZN(n12726) );
  NOR2_X1 U15422 ( .A1(n18814), .A2(n19646), .ZN(n12948) );
  NOR3_X1 U15423 ( .A1(n15358), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n12338), .ZN(n12727) );
  AOI211_X1 U15424 ( .C1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n12726), .A(
        n12948), .B(n12727), .ZN(n12339) );
  OAI21_X1 U15425 ( .B1(n19072), .B2(n15991), .A(n12339), .ZN(n12344) );
  INV_X1 U15426 ( .A(n12340), .ZN(n12343) );
  INV_X1 U15427 ( .A(n12341), .ZN(n12342) );
  OAI21_X1 U15428 ( .B1(n12343), .B2(n12342), .A(n12733), .ZN(n18813) );
  INV_X1 U15429 ( .A(n18813), .ZN(n13997) );
  INV_X1 U15430 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16378) );
  INV_X1 U15431 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17672) );
  NOR2_X1 U15432 ( .A1(n17672), .A2(n17695), .ZN(n12348) );
  NAND2_X1 U15433 ( .A1(n17660), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17631) );
  NAND4_X1 U15434 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16518) );
  NOR2_X2 U15435 ( .A1(n17631), .A2(n16518), .ZN(n17592) );
  NAND2_X1 U15436 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17592), .ZN(
        n17571) );
  NAND2_X1 U15437 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17573) );
  NOR3_X2 U15438 ( .A1(n17571), .A2(n17573), .A3(n17553), .ZN(n17524) );
  NAND3_X1 U15439 ( .A1(n17524), .A2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17512) );
  INV_X1 U15440 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17513) );
  NOR2_X2 U15441 ( .A1(n17512), .A2(n17513), .ZN(n17487) );
  NAND3_X1 U15442 ( .A1(n17487), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17475) );
  INV_X1 U15443 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17474) );
  NOR2_X2 U15444 ( .A1(n17475), .A2(n17474), .ZN(n17447) );
  NAND2_X1 U15445 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17402) );
  NAND2_X1 U15446 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17370) );
  NOR2_X2 U15447 ( .A1(n12349), .A2(n17370), .ZN(n16236) );
  NAND2_X1 U15448 ( .A1(n16236), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12877) );
  INV_X1 U15449 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17727) );
  NOR2_X2 U15450 ( .A1(n12877), .A2(n17727), .ZN(n12357) );
  XNOR2_X1 U15451 ( .A(n16378), .B(n12357), .ZN(n16377) );
  INV_X1 U15452 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16388) );
  NAND2_X1 U15453 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16236), .ZN(
        n12350) );
  AOI21_X1 U15454 ( .B1(n16388), .B2(n12350), .A(n12357), .ZN(n16387) );
  INV_X1 U15455 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n20864) );
  NOR2_X1 U15456 ( .A1(n17727), .A2(n12349), .ZN(n12352) );
  NAND2_X1 U15457 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n12352), .ZN(
        n12351) );
  INV_X1 U15458 ( .A(n12350), .ZN(n12879) );
  AOI21_X1 U15459 ( .B1(n20864), .B2(n12351), .A(n12879), .ZN(n17360) );
  OAI21_X1 U15460 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n12352), .A(
        n12351), .ZN(n17375) );
  INV_X1 U15461 ( .A(n17375), .ZN(n16409) );
  INV_X1 U15462 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12353) );
  NAND2_X1 U15463 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17390), .ZN(
        n12354) );
  AOI21_X1 U15464 ( .B1(n12353), .B2(n12354), .A(n12352), .ZN(n17391) );
  INV_X1 U15465 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n20851) );
  INV_X1 U15466 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17422) );
  INV_X1 U15467 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17458) );
  NAND2_X1 U15468 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17488) );
  INV_X1 U15469 ( .A(n17487), .ZN(n17485) );
  NOR2_X1 U15470 ( .A1(n17727), .A2(n17485), .ZN(n17486) );
  INV_X1 U15471 ( .A(n17486), .ZN(n16519) );
  NOR2_X1 U15472 ( .A1(n17488), .A2(n16519), .ZN(n16494) );
  NAND2_X1 U15473 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16494), .ZN(
        n12356) );
  NOR2_X1 U15474 ( .A1(n17458), .A2(n12356), .ZN(n12359) );
  NAND2_X1 U15475 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n12359), .ZN(
        n12360) );
  NOR2_X1 U15476 ( .A1(n17422), .A2(n12360), .ZN(n17400) );
  INV_X1 U15477 ( .A(n17400), .ZN(n12364) );
  NOR2_X1 U15478 ( .A1(n20851), .A2(n12364), .ZN(n12355) );
  OAI21_X1 U15479 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n12355), .A(
        n12354), .ZN(n17405) );
  INV_X1 U15480 ( .A(n17405), .ZN(n16430) );
  AOI21_X1 U15481 ( .B1(n17422), .B2(n12360), .A(n17400), .ZN(n17427) );
  AOI21_X1 U15482 ( .B1(n17458), .B2(n12356), .A(n12359), .ZN(n17461) );
  OAI21_X1 U15483 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n16494), .A(
        n12356), .ZN(n17477) );
  INV_X1 U15484 ( .A(n17477), .ZN(n16485) );
  INV_X1 U15485 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16506) );
  NOR2_X1 U15486 ( .A1(n17727), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16714) );
  INV_X1 U15487 ( .A(n16714), .ZN(n16674) );
  NOR2_X1 U15488 ( .A1(n17512), .A2(n16674), .ZN(n16517) );
  NAND2_X1 U15489 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16517), .ZN(
        n16507) );
  NOR2_X1 U15490 ( .A1(n16506), .A2(n16507), .ZN(n16496) );
  NAND2_X1 U15491 ( .A1(n12357), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12358) );
  INV_X1 U15492 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12880) );
  INV_X4 U15493 ( .A(n9710), .ZN(n16688) );
  NOR2_X1 U15494 ( .A1(n16485), .A2(n16484), .ZN(n16483) );
  NOR2_X1 U15495 ( .A1(n16483), .A2(n16688), .ZN(n16475) );
  NOR2_X1 U15496 ( .A1(n17461), .A2(n16475), .ZN(n16474) );
  NOR2_X1 U15497 ( .A1(n16474), .A2(n16688), .ZN(n16465) );
  INV_X1 U15498 ( .A(n16465), .ZN(n12363) );
  INV_X1 U15499 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n21049) );
  INV_X1 U15500 ( .A(n12359), .ZN(n12361) );
  INV_X1 U15501 ( .A(n12360), .ZN(n17424) );
  AOI21_X1 U15502 ( .B1(n21049), .B2(n12361), .A(n17424), .ZN(n17455) );
  INV_X1 U15503 ( .A(n17455), .ZN(n12362) );
  NAND2_X1 U15504 ( .A1(n12363), .A2(n12362), .ZN(n16463) );
  AND2_X2 U15505 ( .A1(n16463), .A2(n9710), .ZN(n16452) );
  NOR2_X1 U15506 ( .A1(n17427), .A2(n16452), .ZN(n16451) );
  NOR2_X1 U15507 ( .A1(n16451), .A2(n16688), .ZN(n16444) );
  INV_X1 U15508 ( .A(n16444), .ZN(n12366) );
  OAI22_X1 U15509 ( .A1(n20851), .A2(n17400), .B1(n12364), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17413) );
  NAND2_X1 U15510 ( .A1(n12366), .A2(n12365), .ZN(n16442) );
  NOR2_X1 U15511 ( .A1(n16430), .A2(n16429), .ZN(n16428) );
  NOR2_X1 U15512 ( .A1(n16428), .A2(n16688), .ZN(n16421) );
  NOR2_X1 U15513 ( .A1(n17391), .A2(n16421), .ZN(n16420) );
  NOR2_X1 U15514 ( .A1(n16420), .A2(n16688), .ZN(n16408) );
  NOR2_X1 U15515 ( .A1(n16409), .A2(n16408), .ZN(n16407) );
  NOR2_X1 U15516 ( .A1(n16407), .A2(n16688), .ZN(n16402) );
  NOR2_X1 U15517 ( .A1(n17360), .A2(n16402), .ZN(n16401) );
  NOR2_X1 U15518 ( .A1(n16401), .A2(n16688), .ZN(n16386) );
  NOR2_X1 U15519 ( .A1(n16387), .A2(n16386), .ZN(n16385) );
  NOR2_X1 U15520 ( .A1(n16385), .A2(n16688), .ZN(n16376) );
  INV_X1 U15521 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18729) );
  INV_X1 U15522 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16356) );
  NAND4_X1 U15523 ( .A1(n18729), .A2(n18732), .A3(n16356), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n18588) );
  NOR2_X1 U15524 ( .A1(n16688), .A2(n18588), .ZN(n16724) );
  INV_X1 U15525 ( .A(n16724), .ZN(n12367) );
  NOR3_X1 U15526 ( .A1(n16377), .A2(n16376), .A3(n12367), .ZN(n12497) );
  NOR2_X1 U15527 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18706) );
  NAND2_X1 U15528 ( .A1(n18729), .A2(n18706), .ZN(n18742) );
  INV_X2 U15529 ( .A(n18527), .ZN(n18535) );
  AOI22_X1 U15530 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(n9716), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U15531 ( .A1(n16755), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17043), .ZN(n12381) );
  INV_X1 U15532 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n20866) );
  AOI22_X1 U15533 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17048), .ZN(n12368) );
  OAI21_X1 U15534 ( .B1(n20866), .B2(n12402), .A(n12368), .ZN(n12379) );
  NOR2_X2 U15535 ( .A1(n12369), .A2(n18535), .ZN(n12585) );
  AOI22_X1 U15536 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12570), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12377) );
  INV_X4 U15537 ( .A(n12560), .ZN(n17044) );
  AOI22_X1 U15538 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n17045), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17044), .ZN(n12376) );
  NOR2_X2 U15539 ( .A1(n12373), .A2(n18538), .ZN(n12542) );
  AOI22_X1 U15540 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17051), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17049), .ZN(n12375) );
  AOI22_X1 U15541 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10056), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12374) );
  NAND4_X1 U15542 ( .A1(n12377), .A2(n12376), .A3(n12375), .A4(n12374), .ZN(
        n12378) );
  NAND3_X2 U15543 ( .A1(n12382), .A2(n12381), .A3(n12380), .ZN(n18119) );
  AOI22_X1 U15544 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12391) );
  AOI22_X1 U15545 ( .A1(n17026), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12390) );
  AOI22_X1 U15546 ( .A1(n9740), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17033), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12383) );
  OAI21_X1 U15547 ( .B1(n12560), .B2(n18087), .A(n12383), .ZN(n12389) );
  AOI22_X1 U15548 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n9717), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12387) );
  AOI22_X1 U15549 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U15550 ( .A1(n16755), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12385) );
  AOI22_X1 U15551 ( .A1(n17048), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10056), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12384) );
  NAND4_X1 U15552 ( .A1(n12387), .A2(n12386), .A3(n12385), .A4(n12384), .ZN(
        n12388) );
  AOI22_X1 U15553 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12401) );
  AOI22_X1 U15554 ( .A1(n9715), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12400) );
  AOI22_X1 U15555 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12392) );
  OAI21_X1 U15556 ( .B1(n12560), .B2(n18107), .A(n12392), .ZN(n12398) );
  INV_X2 U15557 ( .A(n12402), .ZN(n16802) );
  AOI22_X1 U15558 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12396) );
  AOI22_X1 U15559 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12585), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12395) );
  AOI22_X1 U15560 ( .A1(n17026), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10056), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12394) );
  AOI22_X1 U15561 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12393) );
  NAND4_X1 U15562 ( .A1(n12396), .A2(n12395), .A3(n12394), .A4(n12393), .ZN(
        n12397) );
  AOI211_X1 U15563 ( .C1(n9718), .C2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n12398), .B(n12397), .ZN(n12399) );
  AOI22_X1 U15564 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9711), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U15565 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12412) );
  INV_X1 U15566 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18102) );
  AOI22_X1 U15567 ( .A1(n16755), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12404) );
  OAI21_X1 U15568 ( .B1(n12560), .B2(n18102), .A(n12404), .ZN(n12410) );
  AOI22_X1 U15569 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15570 ( .A1(n17026), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12407) );
  AOI22_X1 U15571 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12570), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12406) );
  AOI22_X1 U15572 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10056), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12405) );
  NAND4_X1 U15573 ( .A1(n12408), .A2(n12407), .A3(n12406), .A4(n12405), .ZN(
        n12409) );
  AOI211_X1 U15574 ( .C1(n9718), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n12410), .B(n12409), .ZN(n12411) );
  NAND3_X1 U15575 ( .A1(n12413), .A2(n12412), .A3(n12411), .ZN(n12466) );
  INV_X1 U15576 ( .A(n12466), .ZN(n18099) );
  AOI22_X1 U15577 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U15578 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U15579 ( .A1(n9740), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12542), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U15580 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10056), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12414) );
  NAND4_X1 U15581 ( .A1(n12417), .A2(n12416), .A3(n12415), .A4(n12414), .ZN(
        n12423) );
  AOI22_X1 U15582 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15583 ( .A1(n9716), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12420) );
  AOI22_X1 U15584 ( .A1(n17026), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12419) );
  AOI22_X1 U15585 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12544), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12418) );
  NAND4_X1 U15586 ( .A1(n12421), .A2(n12420), .A3(n12419), .A4(n12418), .ZN(
        n12422) );
  AOI22_X1 U15587 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12433) );
  AOI22_X1 U15588 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12432) );
  INV_X2 U15589 ( .A(n12519), .ZN(n17033) );
  AOI22_X1 U15590 ( .A1(n12585), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17033), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12424) );
  OAI21_X1 U15591 ( .B1(n12560), .B2(n20853), .A(n12424), .ZN(n12430) );
  AOI22_X1 U15592 ( .A1(n9715), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12428) );
  AOI22_X1 U15593 ( .A1(n17026), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12542), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12427) );
  AOI22_X1 U15594 ( .A1(n16686), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U15595 ( .A1(n16755), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10056), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12425) );
  NAND4_X1 U15596 ( .A1(n12428), .A2(n12427), .A3(n12426), .A4(n12425), .ZN(
        n12429) );
  NOR2_X1 U15597 ( .A1(n18109), .A2(n18115), .ZN(n12459) );
  NAND4_X1 U15598 ( .A1(n18084), .A2(n18104), .A3(n18099), .A4(n12459), .ZN(
        n12434) );
  AOI22_X1 U15599 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U15600 ( .A1(n17026), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12542), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12443) );
  AOI22_X1 U15601 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12435) );
  OAI21_X1 U15602 ( .B1(n12451), .B2(n20819), .A(n12435), .ZN(n12441) );
  AOI22_X1 U15603 ( .A1(n9716), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12439) );
  AOI22_X1 U15604 ( .A1(n12585), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15605 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10056), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U15606 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12436) );
  NAND4_X1 U15607 ( .A1(n12439), .A2(n12438), .A3(n12437), .A4(n12436), .ZN(
        n12440) );
  NAND3_X1 U15608 ( .A1(n18094), .A2(n18104), .A3(n18115), .ZN(n12464) );
  INV_X1 U15609 ( .A(n12464), .ZN(n12445) );
  NAND2_X1 U15610 ( .A1(n12661), .A2(n17098), .ZN(n12659) );
  AOI22_X1 U15611 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17017), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12449) );
  AOI22_X1 U15612 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n9740), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U15613 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12447) );
  AOI22_X1 U15614 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10056), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12446) );
  NAND4_X1 U15615 ( .A1(n12449), .A2(n12448), .A3(n12447), .A4(n12446), .ZN(
        n12457) );
  AOI22_X1 U15616 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U15617 ( .A1(n17026), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U15618 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17033), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12453) );
  INV_X1 U15619 ( .A(n12530), .ZN(n16870) );
  AOI22_X1 U15620 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12452) );
  NAND3_X1 U15621 ( .A1(n12455), .A2(n12454), .A3(n10079), .ZN(n12456) );
  NOR2_X1 U15622 ( .A1(n18090), .A2(n16678), .ZN(n12458) );
  NOR3_X1 U15623 ( .A1(n12458), .A2(n12471), .A3(n12466), .ZN(n12462) );
  NOR2_X1 U15624 ( .A1(n17097), .A2(n12459), .ZN(n12460) );
  NOR2_X1 U15625 ( .A1(n12458), .A2(n12640), .ZN(n12643) );
  OAI22_X1 U15626 ( .A1(n18104), .A2(n12460), .B1(n12459), .B2(n12643), .ZN(
        n12461) );
  OAI221_X1 U15627 ( .B1(n16678), .B2(n12464), .C1(n16678), .C2(n12659), .A(
        n12463), .ZN(n12648) );
  NOR2_X1 U15628 ( .A1(n17097), .A2(n18548), .ZN(n15611) );
  NOR2_X1 U15629 ( .A1(n18728), .A2(n18084), .ZN(n17306) );
  INV_X1 U15630 ( .A(n17306), .ZN(n12465) );
  AOI211_X1 U15631 ( .C1(n12466), .C2(n12467), .A(n12648), .B(n12647), .ZN(
        n12699) );
  NAND2_X1 U15632 ( .A1(n12468), .A2(n12699), .ZN(n12696) );
  NAND2_X1 U15633 ( .A1(n18119), .A2(n12466), .ZN(n12642) );
  NAND2_X1 U15634 ( .A1(n17305), .A2(n16678), .ZN(n12469) );
  NAND2_X1 U15635 ( .A1(n12468), .A2(n12640), .ZN(n12650) );
  NAND2_X1 U15636 ( .A1(n12469), .A2(n12650), .ZN(n16358) );
  INV_X1 U15637 ( .A(n12469), .ZN(n12470) );
  XNOR2_X1 U15638 ( .A(n18728), .B(n18094), .ZN(n12660) );
  INV_X1 U15639 ( .A(n12700), .ZN(n12472) );
  NOR2_X1 U15640 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18732), .ZN(n18584) );
  NAND2_X1 U15641 ( .A1(n18584), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18579) );
  AOI22_X1 U15642 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18555), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18703), .ZN(n12654) );
  XOR2_X1 U15643 ( .A(n12654), .B(n12652), .Z(n12484) );
  OAI22_X1 U15644 ( .A1(n18540), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18560), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12479) );
  OAI21_X1 U15645 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18697), .A(
        n12475), .ZN(n12476) );
  OAI22_X1 U15646 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18564), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12476), .ZN(n12482) );
  NOR2_X1 U15647 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18564), .ZN(
        n12477) );
  NAND2_X1 U15648 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12476), .ZN(
        n12481) );
  AOI22_X1 U15649 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12482), .B1(
        n12477), .B2(n12481), .ZN(n12658) );
  OAI21_X1 U15650 ( .B1(n12480), .B2(n12479), .A(n12658), .ZN(n12478) );
  AND2_X1 U15651 ( .A1(n12481), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12483) );
  OAI22_X1 U15652 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18525), .B1(
        n12483), .B2(n12482), .ZN(n12655) );
  INV_X1 U15653 ( .A(n18745), .ZN(n16677) );
  NAND2_X1 U15654 ( .A1(n18729), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18582) );
  INV_X1 U15655 ( .A(n18582), .ZN(n18421) );
  NAND2_X1 U15656 ( .A1(n18584), .A2(n18421), .ZN(n18577) );
  INV_X1 U15657 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18604) );
  INV_X1 U15658 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n16350) );
  NAND2_X2 U15659 ( .A1(n18719), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18666) );
  NOR2_X1 U15660 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16355) );
  INV_X1 U15661 ( .A(n16355), .ZN(n18593) );
  NAND3_X1 U15662 ( .A1(n18604), .A2(n18666), .A3(n18593), .ZN(n15509) );
  NAND2_X1 U15663 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18723) );
  INV_X1 U15664 ( .A(n18723), .ZN(n18730) );
  AOI211_X1 U15665 ( .C1(n18090), .C2(n15509), .A(n18730), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n12488) );
  INV_X1 U15666 ( .A(n12488), .ZN(n18573) );
  NOR2_X1 U15667 ( .A1(n16720), .A2(n16723), .ZN(n16560) );
  INV_X1 U15668 ( .A(n16560), .ZN(n16730) );
  NAND3_X1 U15669 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n12485) );
  INV_X1 U15670 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18650) );
  INV_X1 U15671 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18646) );
  INV_X1 U15672 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20847) );
  INV_X1 U15673 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18637) );
  INV_X1 U15674 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18634) );
  INV_X1 U15675 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18628) );
  INV_X1 U15676 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18624) );
  INV_X1 U15677 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18621) );
  INV_X1 U15678 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18619) );
  INV_X1 U15679 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18617) );
  INV_X1 U15680 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18613) );
  NAND3_X1 U15681 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16683) );
  NOR2_X1 U15682 ( .A1(n18613), .A2(n16683), .ZN(n16661) );
  NAND2_X1 U15683 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16661), .ZN(n16638) );
  NOR4_X1 U15684 ( .A1(n18621), .A2(n18619), .A3(n18617), .A4(n16638), .ZN(
        n16608) );
  NAND2_X1 U15685 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16608), .ZN(n16605) );
  NOR2_X1 U15686 ( .A1(n18624), .A2(n16605), .ZN(n16598) );
  NAND2_X1 U15687 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16598), .ZN(n16567) );
  NOR2_X1 U15688 ( .A1(n18628), .A2(n16567), .ZN(n16568) );
  NAND3_X1 U15689 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n16568), .ZN(n16558) );
  NOR2_X1 U15690 ( .A1(n18634), .A2(n16558), .ZN(n16538) );
  NAND2_X1 U15691 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n16538), .ZN(n16523) );
  NOR2_X1 U15692 ( .A1(n18637), .A2(n16523), .ZN(n16499) );
  NAND3_X1 U15693 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(n16499), .ZN(n16487) );
  NOR2_X1 U15694 ( .A1(n20847), .A2(n16487), .ZN(n16469) );
  NAND2_X1 U15695 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16469), .ZN(n16466) );
  NOR2_X1 U15696 ( .A1(n18646), .A2(n16466), .ZN(n16450) );
  NAND2_X1 U15697 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16450), .ZN(n16438) );
  NOR2_X1 U15698 ( .A1(n18650), .A2(n16438), .ZN(n16418) );
  NAND3_X1 U15699 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n16418), .ZN(n12486) );
  NOR2_X1 U15700 ( .A1(n16720), .A2(n12486), .ZN(n16399) );
  NOR2_X1 U15701 ( .A1(n16560), .A2(n16399), .ZN(n16425) );
  AOI21_X1 U15702 ( .B1(n16730), .B2(n12485), .A(n16425), .ZN(n16397) );
  NOR2_X1 U15703 ( .A1(n16704), .A2(n12486), .ZN(n16411) );
  NAND4_X1 U15704 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16411), .ZN(n12489) );
  NOR2_X1 U15705 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n12489), .ZN(n16380) );
  INV_X1 U15706 ( .A(n16380), .ZN(n12487) );
  INV_X1 U15707 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18663) );
  AOI21_X1 U15708 ( .B1(n16397), .B2(n12487), .A(n18663), .ZN(n12496) );
  INV_X1 U15709 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18665) );
  NOR3_X1 U15710 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18665), .A3(n12489), 
        .ZN(n12490) );
  AOI21_X1 U15711 ( .B1(n16721), .B2(P3_EBX_REG_31__SCAN_IN), .A(n12490), .ZN(
        n12494) );
  NAND2_X1 U15712 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18728), .ZN(n12491) );
  AOI211_X4 U15713 ( .C1(n16356), .C2(n18723), .A(n12492), .B(n12491), .ZN(
        n16731) );
  NOR3_X1 U15714 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16707) );
  INV_X1 U15715 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17075) );
  NAND2_X1 U15716 ( .A1(n16707), .A2(n17075), .ZN(n16696) );
  NOR2_X1 U15717 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16696), .ZN(n16671) );
  INV_X1 U15718 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17067) );
  NAND2_X1 U15719 ( .A1(n16671), .A2(n17067), .ZN(n16665) );
  INV_X1 U15720 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17064) );
  NAND2_X1 U15721 ( .A1(n16650), .A2(n17064), .ZN(n16642) );
  INV_X1 U15722 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20822) );
  NAND2_X1 U15723 ( .A1(n16628), .A2(n20822), .ZN(n16620) );
  INV_X1 U15724 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20970) );
  NAND2_X1 U15725 ( .A1(n16609), .A2(n20970), .ZN(n16593) );
  INV_X1 U15726 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20869) );
  NAND2_X1 U15727 ( .A1(n16580), .A2(n20869), .ZN(n16576) );
  INV_X1 U15728 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16550) );
  NAND2_X1 U15729 ( .A1(n16566), .A2(n16550), .ZN(n16549) );
  INV_X1 U15730 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16527) );
  NAND2_X1 U15731 ( .A1(n16530), .A2(n16527), .ZN(n16526) );
  INV_X1 U15732 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n20935) );
  NAND2_X1 U15733 ( .A1(n16509), .A2(n20935), .ZN(n16501) );
  INV_X1 U15734 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16883) );
  NAND2_X1 U15735 ( .A1(n16488), .A2(n16883), .ZN(n16480) );
  NOR2_X1 U15736 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16480), .ZN(n16461) );
  INV_X1 U15737 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16456) );
  NAND2_X1 U15738 ( .A1(n16461), .A2(n16456), .ZN(n16455) );
  NOR2_X1 U15739 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16455), .ZN(n16441) );
  INV_X1 U15740 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n20821) );
  NAND2_X1 U15741 ( .A1(n16441), .A2(n20821), .ZN(n16434) );
  NOR2_X1 U15742 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16434), .ZN(n16419) );
  INV_X1 U15743 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16414) );
  NAND2_X1 U15744 ( .A1(n16419), .A2(n16414), .ZN(n16413) );
  NOR2_X1 U15745 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16413), .ZN(n16400) );
  INV_X1 U15746 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16394) );
  NAND2_X1 U15747 ( .A1(n16400), .A2(n16394), .ZN(n16375) );
  NOR2_X1 U15748 ( .A1(n16706), .A2(n16375), .ZN(n16382) );
  INV_X1 U15749 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16738) );
  NAND2_X1 U15750 ( .A1(n16382), .A2(n16738), .ZN(n12493) );
  NAND3_X1 U15751 ( .A1(n12494), .A2(n12493), .A3(n10067), .ZN(n12495) );
  INV_X1 U15752 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16234) );
  NAND2_X1 U15753 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16234), .ZN(
        n12707) );
  AOI22_X1 U15754 ( .A1(n16755), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12507) );
  AOI22_X1 U15755 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U15756 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9711), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12498) );
  OAI21_X1 U15757 ( .B1(n9719), .B2(n20853), .A(n12498), .ZN(n12504) );
  INV_X1 U15758 ( .A(n12519), .ZN(n17045) );
  AOI22_X1 U15759 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U15760 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12501) );
  AOI22_X1 U15761 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U15762 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12499) );
  NAND4_X1 U15763 ( .A1(n12502), .A2(n12501), .A3(n12500), .A4(n12499), .ZN(
        n12503) );
  AOI211_X1 U15764 ( .C1(n12590), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n12504), .B(n12503), .ZN(n12505) );
  NAND3_X1 U15765 ( .A1(n12507), .A2(n12506), .A3(n12505), .ZN(n17217) );
  AOI22_X1 U15766 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12542), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12511) );
  AOI22_X1 U15767 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9718), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12510) );
  AOI22_X1 U15768 ( .A1(n9740), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12509) );
  AOI22_X1 U15769 ( .A1(n16755), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12508) );
  NAND4_X1 U15770 ( .A1(n12511), .A2(n12510), .A3(n12509), .A4(n12508), .ZN(
        n12518) );
  AOI22_X1 U15771 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9711), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12516) );
  AOI22_X1 U15772 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12515) );
  AOI22_X1 U15773 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12514) );
  AOI22_X1 U15774 ( .A1(n17033), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12513) );
  NAND4_X1 U15775 ( .A1(n12516), .A2(n12515), .A3(n12514), .A4(n12513), .ZN(
        n12517) );
  AOI22_X1 U15776 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12542), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12523) );
  AOI22_X1 U15777 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9718), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12522) );
  AOI22_X1 U15778 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10056), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12521) );
  AOI22_X1 U15779 ( .A1(n9740), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17033), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12520) );
  NAND4_X1 U15780 ( .A1(n12523), .A2(n12522), .A3(n12521), .A4(n12520), .ZN(
        n12529) );
  AOI22_X1 U15781 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12527) );
  AOI22_X1 U15782 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12526) );
  AOI22_X1 U15783 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12525) );
  AOI22_X1 U15784 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9711), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12524) );
  NAND4_X1 U15785 ( .A1(n12527), .A2(n12526), .A3(n12525), .A4(n12524), .ZN(
        n12528) );
  AOI22_X1 U15786 ( .A1(n12544), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12546), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12534) );
  AOI22_X1 U15787 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n16755), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12533) );
  AOI22_X1 U15788 ( .A1(n17026), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9711), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12532) );
  AOI22_X1 U15789 ( .A1(n12530), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10056), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12531) );
  AOI22_X1 U15790 ( .A1(n12542), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12535), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12539) );
  AOI22_X1 U15791 ( .A1(n16686), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12538) );
  AOI22_X1 U15792 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12585), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12537) );
  AOI22_X1 U15793 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9709), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12536) );
  INV_X1 U15794 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12552) );
  AOI22_X1 U15795 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10056), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12540) );
  OAI21_X1 U15796 ( .B1(n12560), .B2(n20819), .A(n12540), .ZN(n12541) );
  INV_X1 U15797 ( .A(n12541), .ZN(n12551) );
  AOI22_X1 U15798 ( .A1(n16755), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12542), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12550) );
  AOI22_X1 U15799 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9709), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12549) );
  AOI22_X1 U15800 ( .A1(n9715), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12544), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U15801 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12546), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12547) );
  INV_X1 U15802 ( .A(n12554), .ZN(n12558) );
  AOI22_X1 U15803 ( .A1(n17026), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12585), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12556) );
  AOI22_X1 U15804 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9711), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12555) );
  AND2_X1 U15805 ( .A1(n12556), .A2(n12555), .ZN(n12557) );
  NAND2_X1 U15806 ( .A1(n12558), .A2(n12557), .ZN(n17235) );
  NAND2_X1 U15807 ( .A1(n12678), .A2(n17235), .ZN(n12584) );
  AOI22_X1 U15808 ( .A1(n9716), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(n9717), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U15809 ( .A1(n16755), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12568) );
  AOI22_X1 U15810 ( .A1(n17033), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12559) );
  OAI21_X1 U15811 ( .B1(n9719), .B2(n18107), .A(n12559), .ZN(n12566) );
  AOI22_X1 U15812 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9711), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U15813 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17044), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U15814 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12562) );
  AOI22_X1 U15815 ( .A1(n17026), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10056), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12561) );
  NAND4_X1 U15816 ( .A1(n12564), .A2(n12563), .A3(n12562), .A4(n12561), .ZN(
        n12565) );
  AOI211_X1 U15817 ( .C1(n9718), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n12566), .B(n12565), .ZN(n12567) );
  NAND3_X1 U15818 ( .A1(n12569), .A2(n12568), .A3(n12567), .ZN(n17225) );
  NAND2_X1 U15819 ( .A1(n12602), .A2(n17225), .ZN(n12607) );
  AOI22_X1 U15820 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17044), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12575) );
  AOI22_X1 U15821 ( .A1(n9740), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17045), .ZN(n12574) );
  AOI22_X1 U15822 ( .A1(n17048), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n12571), .ZN(n12573) );
  AOI22_X1 U15823 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12572) );
  NAND4_X1 U15824 ( .A1(n12575), .A2(n12574), .A3(n12573), .A4(n12572), .ZN(
        n12581) );
  AOI22_X1 U15825 ( .A1(n9716), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(n9717), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U15826 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9718), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12578) );
  AOI22_X1 U15827 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12577) );
  AOI22_X1 U15828 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n16755), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17051), .ZN(n12576) );
  NAND4_X1 U15829 ( .A1(n12579), .A2(n12578), .A3(n12577), .A4(n12576), .ZN(
        n12580) );
  NOR2_X4 U15830 ( .A1(n16260), .A2(n17215), .ZN(n17638) );
  INV_X1 U15831 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17763) );
  INV_X1 U15832 ( .A(n16260), .ZN(n12582) );
  XOR2_X1 U15833 ( .A(n12583), .B(n17217), .Z(n12609) );
  INV_X1 U15834 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18019) );
  XNOR2_X1 U15835 ( .A(n12584), .B(n17230), .ZN(n12600) );
  INV_X1 U15836 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18043) );
  NOR2_X1 U15837 ( .A1(n18043), .A2(n12598), .ZN(n12599) );
  INV_X1 U15838 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18687) );
  NOR2_X1 U15839 ( .A1(n12678), .A2(n18687), .ZN(n12597) );
  AOI22_X1 U15840 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12570), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U15841 ( .A1(n9716), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12588) );
  AOI22_X1 U15842 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12587) );
  AOI22_X1 U15843 ( .A1(n12546), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10056), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12586) );
  NAND4_X1 U15844 ( .A1(n12589), .A2(n12588), .A3(n12587), .A4(n12586), .ZN(
        n12596) );
  AOI22_X1 U15845 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12594) );
  AOI22_X1 U15846 ( .A1(n12542), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12593) );
  AOI22_X1 U15847 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12592) );
  AOI22_X1 U15848 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12591) );
  NAND4_X1 U15849 ( .A1(n12594), .A2(n12593), .A3(n12592), .A4(n12591), .ZN(
        n12595) );
  NAND2_X1 U15850 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17730), .ZN(
        n17729) );
  NOR2_X1 U15851 ( .A1(n17729), .A2(n17722), .ZN(n17721) );
  NOR2_X1 U15852 ( .A1(n12597), .A2(n17721), .ZN(n17710) );
  NOR2_X1 U15853 ( .A1(n17710), .A2(n17709), .ZN(n17708) );
  XNOR2_X1 U15854 ( .A(n12600), .B(n12601), .ZN(n17700) );
  NOR2_X1 U15855 ( .A1(n12601), .A2(n12600), .ZN(n17688) );
  XOR2_X1 U15856 ( .A(n12602), .B(n17225), .Z(n12604) );
  INV_X1 U15857 ( .A(n12603), .ZN(n12605) );
  INV_X1 U15858 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18013) );
  XOR2_X1 U15859 ( .A(n18013), .B(n12604), .Z(n17690) );
  XNOR2_X1 U15860 ( .A(n12607), .B(n17222), .ZN(n17675) );
  NOR2_X1 U15861 ( .A1(n17674), .A2(n17675), .ZN(n12608) );
  NAND2_X1 U15862 ( .A1(n17674), .A2(n17675), .ZN(n17673) );
  OAI21_X1 U15863 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n12608), .A(
        n17673), .ZN(n17659) );
  INV_X1 U15864 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17972) );
  XOR2_X1 U15865 ( .A(n17972), .B(n12609), .Z(n17658) );
  NOR2_X1 U15866 ( .A1(n17659), .A2(n17658), .ZN(n17657) );
  NOR2_X2 U15867 ( .A1(n17657), .A2(n12610), .ZN(n12613) );
  XNOR2_X1 U15868 ( .A(n12612), .B(n12613), .ZN(n17653) );
  INV_X1 U15869 ( .A(n17653), .ZN(n12611) );
  INV_X1 U15870 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17988) );
  NAND2_X2 U15871 ( .A1(n12611), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17651) );
  INV_X1 U15872 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17953) );
  NAND2_X1 U15873 ( .A1(n17608), .A2(n17953), .ZN(n17596) );
  INV_X1 U15874 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17558) );
  NOR2_X1 U15875 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17878) );
  NAND2_X1 U15876 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17938) );
  INV_X1 U15877 ( .A(n17938), .ZN(n17599) );
  NAND2_X1 U15878 ( .A1(n17599), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17915) );
  INV_X1 U15879 ( .A(n17915), .ZN(n17942) );
  NAND2_X1 U15880 ( .A1(n17942), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17578) );
  INV_X1 U15881 ( .A(n17578), .ZN(n17893) );
  INV_X1 U15882 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17898) );
  NOR2_X1 U15883 ( .A1(n17558), .A2(n17898), .ZN(n17557) );
  NAND2_X1 U15884 ( .A1(n17893), .A2(n17557), .ZN(n17895) );
  INV_X1 U15885 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17880) );
  NOR2_X1 U15886 ( .A1(n17895), .A2(n17880), .ZN(n17842) );
  INV_X1 U15887 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17858) );
  INV_X1 U15888 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17849) );
  NAND2_X1 U15889 ( .A1(n17510), .A2(n17849), .ZN(n17509) );
  NAND2_X2 U15890 ( .A1(n17509), .A2(n17636), .ZN(n17428) );
  INV_X1 U15891 ( .A(n17521), .ZN(n12620) );
  INV_X1 U15892 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17782) );
  NOR2_X1 U15893 ( .A1(n17858), .A2(n17849), .ZN(n17502) );
  INV_X1 U15894 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17469) );
  INV_X1 U15895 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17837) );
  INV_X1 U15896 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17833) );
  NOR2_X1 U15897 ( .A1(n17837), .A2(n17833), .ZN(n17819) );
  INV_X1 U15898 ( .A(n17819), .ZN(n17466) );
  NOR2_X1 U15899 ( .A1(n17469), .A2(n17466), .ZN(n17439) );
  NAND3_X1 U15900 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17439), .A3(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12666) );
  INV_X1 U15901 ( .A(n12666), .ZN(n17758) );
  NAND2_X1 U15902 ( .A1(n17502), .A2(n17758), .ZN(n17759) );
  NOR2_X1 U15903 ( .A1(n17782), .A2(n17759), .ZN(n17777) );
  NOR2_X1 U15904 ( .A1(n17638), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17503) );
  NAND2_X1 U15905 ( .A1(n17503), .A2(n17837), .ZN(n12617) );
  NOR2_X1 U15906 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12617), .ZN(
        n17464) );
  NAND2_X1 U15907 ( .A1(n17464), .A2(n17469), .ZN(n17441) );
  NOR2_X2 U15908 ( .A1(n17417), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17416) );
  NAND2_X1 U15909 ( .A1(n17502), .A2(n12620), .ZN(n17462) );
  NAND2_X1 U15910 ( .A1(n17428), .A2(n17462), .ZN(n17463) );
  NAND2_X1 U15911 ( .A1(n17758), .A2(n17463), .ZN(n17429) );
  NOR3_X1 U15912 ( .A1(n17416), .A2(n17429), .A3(n17782), .ZN(n12622) );
  INV_X1 U15913 ( .A(n17416), .ZN(n17409) );
  NAND2_X1 U15914 ( .A1(n17636), .A2(n17409), .ZN(n12621) );
  NAND2_X1 U15915 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17739) );
  AND2_X1 U15916 ( .A1(n17638), .A2(n17739), .ZN(n12623) );
  NOR2_X1 U15917 ( .A1(n17638), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12625) );
  INV_X1 U15918 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16242) );
  NAND2_X1 U15919 ( .A1(n15533), .A2(n16242), .ZN(n12628) );
  INV_X1 U15920 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17366) );
  NAND2_X1 U15921 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15534), .ZN(
        n12629) );
  INV_X1 U15922 ( .A(n12629), .ZN(n12627) );
  AOI21_X2 U15923 ( .B1(n17636), .B2(n12628), .A(n12627), .ZN(n12636) );
  INV_X1 U15924 ( .A(n12636), .ZN(n12630) );
  NAND2_X1 U15925 ( .A1(n12629), .A2(n12628), .ZN(n15597) );
  NAND2_X1 U15926 ( .A1(n16234), .A2(n15597), .ZN(n15596) );
  AOI22_X1 U15927 ( .A1(n12707), .A2(n17636), .B1(n12630), .B2(n15596), .ZN(
        n12639) );
  NAND2_X1 U15928 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17638), .ZN(
        n12638) );
  INV_X1 U15929 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18688) );
  NAND2_X1 U15930 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18688), .ZN(
        n12635) );
  NAND2_X1 U15931 ( .A1(n17638), .A2(n18688), .ZN(n12631) );
  NAND2_X1 U15932 ( .A1(n12631), .A2(n12707), .ZN(n12632) );
  AOI21_X1 U15933 ( .B1(n12636), .B2(n12635), .A(n12634), .ZN(n12637) );
  AOI21_X1 U15934 ( .B1(n12639), .B2(n12638), .A(n12637), .ZN(n12876) );
  INV_X1 U15935 ( .A(n12876), .ZN(n12719) );
  NOR2_X1 U15936 ( .A1(n18090), .A2(n12640), .ZN(n12641) );
  NAND2_X1 U15937 ( .A1(n12641), .A2(n17098), .ZN(n12651) );
  INV_X1 U15938 ( .A(n12642), .ZN(n12697) );
  INV_X1 U15939 ( .A(n12643), .ZN(n12644) );
  NOR2_X1 U15940 ( .A1(n12645), .A2(n12644), .ZN(n12646) );
  OAI211_X1 U15941 ( .C1(n18104), .C2(n18548), .A(n12697), .B(n12646), .ZN(
        n12649) );
  INV_X1 U15942 ( .A(n16253), .ZN(n18521) );
  AOI211_X1 U15943 ( .C1(n12650), .C2(n12649), .A(n12648), .B(n12647), .ZN(
        n15515) );
  INV_X1 U15944 ( .A(n12651), .ZN(n12664) );
  AOI21_X1 U15945 ( .B1(n18709), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n12652), .ZN(n12653) );
  AOI21_X1 U15946 ( .B1(n12656), .B2(n12653), .A(n15508), .ZN(n18520) );
  AND2_X1 U15947 ( .A1(n12654), .A2(n12653), .ZN(n12657) );
  INV_X1 U15948 ( .A(n18516), .ZN(n15517) );
  AOI21_X1 U15949 ( .B1(n18104), .B2(n12659), .A(n15517), .ZN(n12663) );
  INV_X1 U15950 ( .A(n15509), .ZN(n18727) );
  OAI21_X1 U15951 ( .B1(n18727), .B2(n12660), .A(n18723), .ZN(n16357) );
  NOR3_X1 U15952 ( .A1(n12661), .A2(n15508), .A3(n16357), .ZN(n12662) );
  AOI211_X1 U15953 ( .C1(n12664), .C2(n18520), .A(n12663), .B(n12662), .ZN(
        n12665) );
  INV_X1 U15954 ( .A(n17502), .ZN(n17846) );
  INV_X1 U15955 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17751) );
  NAND2_X1 U15956 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17760) );
  NOR2_X1 U15957 ( .A1(n17763), .A2(n17760), .ZN(n17737) );
  INV_X1 U15958 ( .A(n17737), .ZN(n17364) );
  NOR2_X1 U15959 ( .A1(n17751), .A2(n17364), .ZN(n12704) );
  INV_X1 U15960 ( .A(n12704), .ZN(n17365) );
  NOR2_X1 U15961 ( .A1(n12666), .A2(n17365), .ZN(n12701) );
  NAND2_X1 U15962 ( .A1(n12701), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12702) );
  NOR2_X1 U15963 ( .A1(n17846), .A2(n12702), .ZN(n16261) );
  NAND2_X1 U15964 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16261), .ZN(
        n16225) );
  INV_X1 U15965 ( .A(n16225), .ZN(n12706) );
  INV_X1 U15966 ( .A(n17842), .ZN(n16223) );
  INV_X1 U15967 ( .A(n12678), .ZN(n17246) );
  NOR2_X1 U15968 ( .A1(n12674), .A2(n17235), .ZN(n12672) );
  NOR2_X1 U15969 ( .A1(n17230), .A2(n12672), .ZN(n12671) );
  NAND2_X1 U15970 ( .A1(n12671), .A2(n17225), .ZN(n12669) );
  NOR2_X1 U15971 ( .A1(n17222), .A2(n12669), .ZN(n12668) );
  NAND2_X1 U15972 ( .A1(n12668), .A2(n17217), .ZN(n12667) );
  NOR2_X1 U15973 ( .A1(n17215), .A2(n12667), .ZN(n12692) );
  XOR2_X1 U15974 ( .A(n17215), .B(n12667), .Z(n17644) );
  XOR2_X1 U15975 ( .A(n17217), .B(n12668), .Z(n12685) );
  XOR2_X1 U15976 ( .A(n17222), .B(n12669), .Z(n12670) );
  NAND2_X1 U15977 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12670), .ZN(
        n12684) );
  XOR2_X1 U15978 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n12670), .Z(
        n17670) );
  XOR2_X1 U15979 ( .A(n17225), .B(n12671), .Z(n12682) );
  XOR2_X1 U15980 ( .A(n17230), .B(n12672), .Z(n12673) );
  NAND2_X1 U15981 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12673), .ZN(
        n12680) );
  XOR2_X1 U15982 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n12673), .Z(
        n17698) );
  XOR2_X1 U15983 ( .A(n17235), .B(n12674), .Z(n12675) );
  OR2_X1 U15984 ( .A1(n18043), .A2(n12675), .ZN(n12679) );
  XOR2_X1 U15985 ( .A(n18043), .B(n12675), .Z(n17713) );
  AOI21_X1 U15986 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12678), .A(
        n17730), .ZN(n12677) );
  INV_X1 U15987 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21029) );
  NOR2_X1 U15988 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12678), .ZN(
        n12676) );
  AOI221_X1 U15989 ( .B1(n17730), .B2(n12678), .C1(n12677), .C2(n21029), .A(
        n12676), .ZN(n17712) );
  NAND2_X1 U15990 ( .A1(n17713), .A2(n17712), .ZN(n17711) );
  NAND2_X1 U15991 ( .A1(n12679), .A2(n17711), .ZN(n17697) );
  NAND2_X1 U15992 ( .A1(n17698), .A2(n17697), .ZN(n17696) );
  NAND2_X1 U15993 ( .A1(n12680), .A2(n17696), .ZN(n12681) );
  NAND2_X1 U15994 ( .A1(n12682), .A2(n12681), .ZN(n12683) );
  XOR2_X1 U15995 ( .A(n12682), .B(n12681), .Z(n17685) );
  NAND2_X1 U15996 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17685), .ZN(
        n17684) );
  NAND2_X1 U15997 ( .A1(n12683), .A2(n17684), .ZN(n17669) );
  NAND2_X1 U15998 ( .A1(n17670), .A2(n17669), .ZN(n17668) );
  NAND2_X1 U15999 ( .A1(n12684), .A2(n17668), .ZN(n12686) );
  NAND2_X1 U16000 ( .A1(n12685), .A2(n12686), .ZN(n12687) );
  XOR2_X1 U16001 ( .A(n12686), .B(n12685), .Z(n17662) );
  NAND2_X1 U16002 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17662), .ZN(
        n17661) );
  NAND2_X1 U16003 ( .A1(n12687), .A2(n17661), .ZN(n17645) );
  NOR2_X1 U16004 ( .A1(n17644), .A2(n17645), .ZN(n12688) );
  NOR2_X1 U16005 ( .A1(n12688), .A2(n17988), .ZN(n12689) );
  NAND2_X1 U16006 ( .A1(n12692), .A2(n12689), .ZN(n12693) );
  INV_X1 U16007 ( .A(n12689), .ZN(n12691) );
  NAND2_X1 U16008 ( .A1(n17644), .A2(n17645), .ZN(n17643) );
  NAND2_X1 U16009 ( .A1(n12692), .A2(n12691), .ZN(n12690) );
  OAI211_X1 U16010 ( .C1(n12692), .C2(n12691), .A(n17643), .B(n12690), .ZN(
        n17629) );
  NAND2_X1 U16011 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17629), .ZN(
        n17628) );
  NAND2_X1 U16012 ( .A1(n12706), .A2(n17799), .ZN(n16241) );
  NAND3_X1 U16013 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16256), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12694) );
  XNOR2_X1 U16014 ( .A(n18688), .B(n12694), .ZN(n12885) );
  NOR2_X1 U16015 ( .A1(n18104), .A2(n17098), .ZN(n18530) );
  NAND3_X1 U16016 ( .A1(n12642), .A2(n18728), .A3(n12700), .ZN(n12698) );
  NAND2_X1 U16017 ( .A1(n12699), .A2(n12698), .ZN(n18528) );
  NOR2_X1 U16018 ( .A1(n18037), .A2(n18050), .ZN(n18060) );
  NOR2_X1 U16019 ( .A1(n18663), .A2(n17892), .ZN(n12883) );
  INV_X2 U16020 ( .A(n18044), .ZN(n18061) );
  NOR2_X2 U16021 ( .A1(n18061), .A2(n18057), .ZN(n18052) );
  INV_X1 U16022 ( .A(n18052), .ZN(n18042) );
  NAND2_X1 U16023 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17968) );
  NAND3_X1 U16024 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17994) );
  INV_X1 U16025 ( .A(n17994), .ZN(n17970) );
  NAND2_X1 U16026 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17970), .ZN(
        n17987) );
  NOR2_X1 U16027 ( .A1(n17988), .A2(n17987), .ZN(n17977) );
  NAND2_X1 U16028 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17977), .ZN(
        n17910) );
  NOR2_X1 U16029 ( .A1(n17968), .A2(n17910), .ZN(n17868) );
  NAND2_X1 U16030 ( .A1(n17842), .A2(n17868), .ZN(n17844) );
  NOR2_X1 U16031 ( .A1(n17759), .A2(n17844), .ZN(n17738) );
  AOI21_X1 U16032 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17966) );
  NOR2_X1 U16033 ( .A1(n17966), .A2(n17910), .ZN(n17867) );
  NAND2_X1 U16034 ( .A1(n17842), .A2(n17867), .ZN(n17795) );
  NOR2_X1 U16035 ( .A1(n17846), .A2(n17795), .ZN(n17848) );
  AOI21_X1 U16036 ( .B1(n12701), .B2(n17848), .A(n17866), .ZN(n17745) );
  NAND2_X1 U16037 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17868), .ZN(
        n17957) );
  INV_X1 U16038 ( .A(n17957), .ZN(n17932) );
  NAND2_X1 U16039 ( .A1(n17842), .A2(n17932), .ZN(n17864) );
  INV_X1 U16040 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17850) );
  NOR2_X1 U16041 ( .A1(n17846), .A2(n17850), .ZN(n17471) );
  INV_X1 U16042 ( .A(n17471), .ZN(n17813) );
  OAI21_X1 U16043 ( .B1(n17864), .B2(n17813), .A(n18547), .ZN(n17817) );
  OAI21_X1 U16044 ( .B1(n17941), .B2(n17439), .A(n17817), .ZN(n17802) );
  AOI211_X1 U16045 ( .C1(n18547), .C2(n12702), .A(n17745), .B(n17802), .ZN(
        n12703) );
  OAI221_X1 U16046 ( .B1(n18549), .B2(n12704), .C1(n18549), .C2(n17738), .A(
        n12703), .ZN(n15529) );
  NAND3_X1 U16047 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12705) );
  INV_X1 U16048 ( .A(n17971), .ZN(n17973) );
  OAI211_X1 U16049 ( .C1(n15529), .C2(n12705), .A(n17973), .B(n18057), .ZN(
        n15598) );
  AOI21_X1 U16050 ( .B1(n18042), .B2(n15598), .A(n18688), .ZN(n12709) );
  NAND2_X1 U16051 ( .A1(n18057), .A2(n17973), .ZN(n18045) );
  NAND3_X1 U16052 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n18688), .ZN(n12713) );
  AOI21_X1 U16053 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18547), .A(
        n18534), .ZN(n18028) );
  OAI22_X1 U16054 ( .A1(n17866), .A2(n17795), .B1(n18028), .B2(n17844), .ZN(
        n17761) );
  NAND3_X1 U16055 ( .A1(n18057), .A2(n12706), .A3(n17761), .ZN(n15527) );
  OAI22_X1 U16056 ( .A1(n12707), .A2(n18045), .B1(n12713), .B2(n15527), .ZN(
        n12708) );
  NOR3_X1 U16057 ( .A1(n12883), .A2(n12709), .A3(n12708), .ZN(n12716) );
  NAND2_X1 U16058 ( .A1(n17981), .A2(n17636), .ZN(n12711) );
  INV_X1 U16059 ( .A(n16257), .ZN(n12714) );
  NAND2_X1 U16060 ( .A1(n16257), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16246) );
  OAI21_X1 U16061 ( .B1(n16234), .B2(n16246), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12712) );
  OAI21_X1 U16062 ( .B1(n12714), .B2(n12713), .A(n12712), .ZN(n12884) );
  NOR2_X1 U16063 ( .A1(n16252), .A2(n18521), .ZN(n17882) );
  NAND2_X1 U16064 ( .A1(n18057), .A2(n17882), .ZN(n17907) );
  INV_X1 U16065 ( .A(n12717), .ZN(n12718) );
  OAI21_X1 U16066 ( .B1(n12719), .B2(n17964), .A(n12718), .ZN(P3_U2831) );
  INV_X1 U16067 ( .A(n12332), .ZN(n12724) );
  NOR2_X1 U16068 ( .A1(n14207), .A2(n12724), .ZN(n12725) );
  NOR2_X1 U16069 ( .A1(n12727), .A2(n12726), .ZN(n15319) );
  INV_X1 U16070 ( .A(n12728), .ZN(n14095) );
  AOI21_X1 U16071 ( .B1(n12729), .B2(n12334), .A(n12728), .ZN(n18799) );
  NAND2_X1 U16072 ( .A1(n18799), .A2(n16143), .ZN(n12732) );
  INV_X1 U16073 ( .A(n12730), .ZN(n15323) );
  NOR2_X1 U16074 ( .A1(n18814), .A2(n19648), .ZN(n12738) );
  AOI21_X1 U16075 ( .B1(n15323), .B2(n15317), .A(n12738), .ZN(n12731) );
  OAI211_X1 U16076 ( .C1(n15319), .C2(n15317), .A(n12732), .B(n12731), .ZN(
        n12735) );
  AOI21_X1 U16077 ( .B1(n12734), .B2(n12733), .A(n14091), .ZN(n18800) );
  INV_X1 U16078 ( .A(n12737), .ZN(n12772) );
  AOI21_X1 U16079 ( .B1(n18795), .B2(n12772), .A(n12773), .ZN(n18794) );
  INV_X1 U16080 ( .A(n18794), .ZN(n12740) );
  AOI21_X1 U16081 ( .B1(n19055), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n12738), .ZN(n12739) );
  OAI21_X1 U16082 ( .B1(n12740), .B2(n19061), .A(n12739), .ZN(n12741) );
  INV_X1 U16083 ( .A(n12744), .ZN(n12745) );
  INV_X1 U16084 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15204) );
  INV_X1 U16085 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12871) );
  XNOR2_X1 U16086 ( .A(n12747), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15178) );
  INV_X1 U16087 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14139) );
  INV_X1 U16088 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15175) );
  XNOR2_X1 U16089 ( .A(n12746), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14244) );
  INV_X1 U16090 ( .A(n12747), .ZN(n12748) );
  AOI21_X1 U16091 ( .B1(n12749), .B2(n12871), .A(n12748), .ZN(n15001) );
  OAI21_X1 U16092 ( .B1(n9830), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n12749), .ZN(n15194) );
  INV_X1 U16093 ( .A(n15194), .ZN(n15007) );
  AOI21_X1 U16094 ( .B1(n15204), .B2(n12750), .A(n9830), .ZN(n15207) );
  INV_X1 U16095 ( .A(n12751), .ZN(n15951) );
  AOI21_X1 U16096 ( .B1(n12753), .B2(n15038), .A(n12752), .ZN(n15044) );
  OAI21_X1 U16097 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n11121), .A(
        n12753), .ZN(n12754) );
  INV_X1 U16098 ( .A(n12754), .ZN(n15969) );
  AOI21_X1 U16099 ( .B1(n18778), .B2(n12774), .A(n9820), .ZN(n18784) );
  AND2_X1 U16100 ( .A1(n12755), .A2(n15233), .ZN(n12757) );
  OR2_X1 U16101 ( .A1(n12757), .A2(n12756), .ZN(n18824) );
  INV_X1 U16102 ( .A(n18824), .ZN(n12771) );
  AOI21_X1 U16103 ( .B1(n10809), .B2(n12770), .A(n12758), .ZN(n18838) );
  AOI21_X1 U16104 ( .B1(n18853), .B2(n12759), .A(n12760), .ZN(n18859) );
  AOI21_X1 U16105 ( .B1(n10789), .B2(n12768), .A(n12769), .ZN(n16039) );
  AOI21_X1 U16106 ( .B1(n10781), .B2(n12767), .A(n12761), .ZN(n18872) );
  AOI21_X1 U16107 ( .B1(n14032), .B2(n12762), .A(n9777), .ZN(n18879) );
  AOI21_X1 U16108 ( .B1(n10763), .B2(n12765), .A(n12766), .ZN(n18915) );
  AOI21_X1 U16109 ( .B1(n16101), .B2(n12764), .A(n12763), .ZN(n16089) );
  OAI22_X1 U16110 ( .A1(n19727), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n15453) );
  OAI22_X1 U16111 ( .A1(n19727), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n10242), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15065) );
  AND2_X1 U16112 ( .A1(n15453), .A2(n15065), .ZN(n15049) );
  OAI21_X1 U16113 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12764), .ZN(n15051) );
  NAND2_X1 U16114 ( .A1(n15049), .A2(n15051), .ZN(n13618) );
  NOR2_X1 U16115 ( .A1(n16089), .A2(n13618), .ZN(n13814) );
  OAI21_X1 U16116 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12763), .A(
        n12765), .ZN(n19050) );
  NAND2_X1 U16117 ( .A1(n13814), .A2(n19050), .ZN(n18913) );
  NOR2_X1 U16118 ( .A1(n18915), .A2(n18913), .ZN(n18895) );
  OAI21_X1 U16119 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12766), .A(
        n12762), .ZN(n18898) );
  NAND2_X1 U16120 ( .A1(n18895), .A2(n18898), .ZN(n18878) );
  NOR2_X1 U16121 ( .A1(n18879), .A2(n18878), .ZN(n13791) );
  OAI21_X1 U16122 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n9777), .A(
        n12767), .ZN(n16081) );
  NAND2_X1 U16123 ( .A1(n13791), .A2(n16081), .ZN(n18869) );
  NOR2_X1 U16124 ( .A1(n18872), .A2(n18869), .ZN(n13776) );
  OAI21_X1 U16125 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12761), .A(
        n12768), .ZN(n16059) );
  NAND2_X1 U16126 ( .A1(n13776), .A2(n16059), .ZN(n12981) );
  NOR2_X1 U16127 ( .A1(n16039), .A2(n12981), .ZN(n13803) );
  OAI21_X1 U16128 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12769), .A(
        n12759), .ZN(n16038) );
  NAND2_X1 U16129 ( .A1(n13803), .A2(n16038), .ZN(n18857) );
  NOR2_X1 U16130 ( .A1(n18859), .A2(n18857), .ZN(n18843) );
  OAI21_X1 U16131 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12760), .A(
        n12770), .ZN(n18844) );
  NAND2_X1 U16132 ( .A1(n18843), .A2(n18844), .ZN(n18831) );
  NOR2_X1 U16133 ( .A1(n18838), .A2(n18831), .ZN(n18830) );
  OAI21_X1 U16134 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12758), .A(
        n12755), .ZN(n15244) );
  NAND2_X1 U16135 ( .A1(n18830), .A2(n15244), .ZN(n18822) );
  NOR2_X1 U16136 ( .A1(n12771), .A2(n18822), .ZN(n18807) );
  OAI21_X1 U16137 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12756), .A(
        n12772), .ZN(n18808) );
  NAND2_X1 U16138 ( .A1(n18807), .A2(n18808), .ZN(n18792) );
  NOR2_X1 U16139 ( .A1(n18794), .A2(n18792), .ZN(n14098) );
  OR2_X1 U16140 ( .A1(n12773), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12775) );
  NAND2_X1 U16141 ( .A1(n12775), .A2(n12774), .ZN(n15225) );
  NAND2_X1 U16142 ( .A1(n14098), .A2(n15225), .ZN(n18785) );
  OAI21_X1 U16143 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n9820), .A(
        n12776), .ZN(n16010) );
  NOR2_X1 U16144 ( .A1(n15969), .A2(n15968), .ZN(n15967) );
  NOR2_X1 U16145 ( .A1(n18896), .A2(n15967), .ZN(n15045) );
  NOR2_X1 U16146 ( .A1(n15044), .A2(n15045), .ZN(n15043) );
  NOR2_X1 U16147 ( .A1(n15951), .A2(n15950), .ZN(n15949) );
  NOR2_X1 U16148 ( .A1(n18896), .A2(n15949), .ZN(n15033) );
  NOR2_X1 U16149 ( .A1(n15207), .A2(n15033), .ZN(n15032) );
  NOR2_X1 U16150 ( .A1(n15178), .A2(n12778), .ZN(n14135) );
  INV_X1 U16151 ( .A(n14135), .ZN(n12780) );
  NAND4_X1 U16152 ( .A1(n19732), .A2(n19727), .A3(n19738), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19602) );
  AOI21_X1 U16153 ( .B1(n12778), .B2(n15178), .A(n19602), .ZN(n12779) );
  NAND2_X1 U16154 ( .A1(n12780), .A2(n12779), .ZN(n12831) );
  NAND2_X1 U16155 ( .A1(n9757), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12848) );
  INV_X1 U16156 ( .A(n12855), .ZN(n12781) );
  NAND2_X1 U16157 ( .A1(n9757), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12853) );
  NAND2_X1 U16158 ( .A1(n12781), .A2(n12853), .ZN(n12857) );
  NAND2_X1 U16159 ( .A1(n9757), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12860) );
  NAND2_X1 U16160 ( .A1(n12861), .A2(n12860), .ZN(n14136) );
  NAND2_X1 U16161 ( .A1(n9757), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12782) );
  XNOR2_X1 U16162 ( .A(n14136), .B(n12782), .ZN(n12921) );
  AND2_X1 U16163 ( .A1(n18753), .A2(n12783), .ZN(n12826) );
  INV_X1 U16164 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15975) );
  NAND2_X1 U16165 ( .A1(n19738), .A2(n19726), .ZN(n12827) );
  INV_X1 U16166 ( .A(n12827), .ZN(n12797) );
  NOR2_X1 U16167 ( .A1(n15975), .A2(n12797), .ZN(n12784) );
  NOR2_X1 U16168 ( .A1(n19546), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19477) );
  INV_X1 U16169 ( .A(n19477), .ZN(n12785) );
  NOR2_X1 U16170 ( .A1(n12786), .A2(n12785), .ZN(n16210) );
  INV_X1 U16171 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n12927) );
  INV_X1 U16172 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15128) );
  OAI22_X1 U16173 ( .A1(n14142), .A2(n15128), .B1(n14140), .B2(n12852), .ZN(
        n12787) );
  AOI21_X1 U16174 ( .B1(n14144), .B2(P2_REIP_REG_27__SCAN_IN), .A(n12787), 
        .ZN(n15025) );
  INV_X1 U16175 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n15122) );
  INV_X1 U16176 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15264) );
  OAI22_X1 U16177 ( .A1(n14142), .A2(n15122), .B1(n14140), .B2(n15264), .ZN(
        n12789) );
  AOI21_X1 U16178 ( .B1(n14144), .B2(P2_REIP_REG_28__SCAN_IN), .A(n12789), 
        .ZN(n15010) );
  INV_X1 U16179 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19667) );
  OR2_X1 U16180 ( .A1(n10908), .A2(n19667), .ZN(n12791) );
  AOI22_X1 U16181 ( .A1(n11131), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12790) );
  NAND2_X1 U16182 ( .A1(n12791), .A2(n12790), .ZN(n14994) );
  OR2_X1 U16183 ( .A1(n10908), .A2(n12927), .ZN(n12794) );
  AOI22_X1 U16184 ( .A1(n11131), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n10991), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12793) );
  NAND2_X1 U16185 ( .A1(n12794), .A2(n12793), .ZN(n12795) );
  NAND2_X1 U16186 ( .A1(n14996), .A2(n12795), .ZN(n14146) );
  OR2_X1 U16187 ( .A1(n14996), .A2(n12795), .ZN(n12796) );
  AND2_X1 U16188 ( .A1(n13014), .A2(n12797), .ZN(n12799) );
  AND2_X1 U16189 ( .A1(n12798), .A2(n12799), .ZN(n16206) );
  INV_X1 U16190 ( .A(n12798), .ZN(n13012) );
  NAND3_X1 U16191 ( .A1(n10216), .A2(n12827), .A3(n15975), .ZN(n12800) );
  AOI21_X1 U16192 ( .B1(n13012), .B2(n12800), .A(n12799), .ZN(n12801) );
  INV_X1 U16193 ( .A(n18922), .ZN(n18906) );
  INV_X1 U16194 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12818) );
  NAND2_X1 U16195 ( .A1(n18929), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18908) );
  NAND2_X1 U16196 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18939), .ZN(
        n12802) );
  OAI21_X1 U16197 ( .B1(n18906), .B2(n12818), .A(n12802), .ZN(n12803) );
  AOI21_X1 U16198 ( .B1(n14454), .B2(n18923), .A(n12803), .ZN(n12804) );
  OAI21_X1 U16199 ( .B1(n18929), .B2(n12927), .A(n12804), .ZN(n12805) );
  AOI21_X1 U16200 ( .B1(n12921), .B2(n18885), .A(n12805), .ZN(n12829) );
  NAND2_X1 U16201 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12809) );
  INV_X1 U16202 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n12806) );
  OAI22_X1 U16203 ( .A1(n12819), .A2(n12806), .B1(n19597), .B2(n15204), .ZN(
        n12807) );
  AOI21_X1 U16204 ( .B1(n14129), .B2(P2_REIP_REG_27__SCAN_IN), .A(n12807), 
        .ZN(n12808) );
  AND2_X1 U16205 ( .A1(n12809), .A2(n12808), .ZN(n15022) );
  NAND2_X1 U16206 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12813) );
  INV_X1 U16207 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n15014) );
  OAI22_X1 U16208 ( .A1(n12819), .A2(n15014), .B1(n19597), .B2(n9866), .ZN(
        n12811) );
  AOI21_X1 U16209 ( .B1(n14129), .B2(P2_REIP_REG_28__SCAN_IN), .A(n12811), 
        .ZN(n12812) );
  AND2_X1 U16210 ( .A1(n12813), .A2(n12812), .ZN(n15009) );
  NAND2_X1 U16211 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12817) );
  INV_X1 U16212 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12814) );
  OAI22_X1 U16213 ( .A1(n12819), .A2(n12814), .B1(n19597), .B2(n12871), .ZN(
        n12815) );
  AOI21_X1 U16214 ( .B1(n14129), .B2(P2_REIP_REG_29__SCAN_IN), .A(n12815), 
        .ZN(n12816) );
  NAND2_X1 U16215 ( .A1(n12817), .A2(n12816), .ZN(n12869) );
  NAND2_X1 U16216 ( .A1(n10254), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12822) );
  OAI22_X1 U16217 ( .A1(n12819), .A2(n12818), .B1(n19597), .B2(n15175), .ZN(
        n12820) );
  AOI21_X1 U16218 ( .B1(n14129), .B2(P2_REIP_REG_30__SCAN_IN), .A(n12820), 
        .ZN(n12821) );
  NAND2_X1 U16219 ( .A1(n12822), .A2(n12821), .ZN(n12824) );
  NOR2_X1 U16220 ( .A1(n12823), .A2(n12824), .ZN(n12825) );
  INV_X1 U16221 ( .A(n12826), .ZN(n12828) );
  NAND2_X1 U16222 ( .A1(n12831), .A2(n12830), .ZN(P2_U2825) );
  AND2_X1 U16223 ( .A1(n15766), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12833) );
  NOR2_X1 U16224 ( .A1(n12935), .A2(n12833), .ZN(n12834) );
  XNOR2_X1 U16225 ( .A(n12936), .B(n12834), .ZN(n14887) );
  OR2_X1 U16226 ( .A1(n12897), .A2(n11273), .ZN(n15564) );
  NOR2_X1 U16227 ( .A1(n15564), .A2(n19751), .ZN(n12835) );
  NAND3_X1 U16228 ( .A1(n15945), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15939) );
  INV_X1 U16229 ( .A(n15939), .ZN(n12839) );
  NOR2_X1 U16230 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20128) );
  AND2_X1 U16231 ( .A1(n12839), .A2(n20128), .ZN(n12940) );
  OR2_X1 U16232 ( .A1(n12840), .A2(n20128), .ZN(n20759) );
  AND2_X1 U16233 ( .A1(n20759), .A2(n15945), .ZN(n12841) );
  NAND2_X1 U16234 ( .A1(n15945), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15569) );
  NAND2_X1 U16235 ( .A1(n20516), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12842) );
  NAND2_X1 U16236 ( .A1(n15569), .A2(n12842), .ZN(n19935) );
  NAND2_X1 U16237 ( .A1(n19939), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14882) );
  OAI21_X1 U16238 ( .B1(n15795), .B2(n12843), .A(n14882), .ZN(n12844) );
  AOI21_X1 U16239 ( .B1(n15791), .B2(n14479), .A(n12844), .ZN(n12845) );
  INV_X1 U16240 ( .A(n12848), .ZN(n12849) );
  NAND2_X1 U16241 ( .A1(n12849), .A2(n9704), .ZN(n12850) );
  NAND2_X1 U16242 ( .A1(n12855), .A2(n12850), .ZN(n15028) );
  AND2_X1 U16243 ( .A1(n15188), .A2(n12852), .ZN(n12851) );
  INV_X1 U16244 ( .A(n12853), .ZN(n12854) );
  NAND2_X1 U16245 ( .A1(n12855), .A2(n12854), .ZN(n12856) );
  AND2_X1 U16246 ( .A1(n12857), .A2(n12856), .ZN(n15016) );
  NAND2_X1 U16247 ( .A1(n15016), .A2(n14238), .ZN(n15189) );
  INV_X1 U16248 ( .A(n15189), .ZN(n12858) );
  AOI21_X1 U16249 ( .B1(n12859), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14185), .ZN(n15185) );
  XNOR2_X1 U16250 ( .A(n12861), .B(n12860), .ZN(n12862) );
  INV_X1 U16251 ( .A(n12862), .ZN(n14997) );
  NAND3_X1 U16252 ( .A1(n14997), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14238), .ZN(n14234) );
  INV_X1 U16253 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14459) );
  OAI21_X1 U16254 ( .B1(n12862), .B2(n10934), .A(n14459), .ZN(n12919) );
  INV_X1 U16255 ( .A(n12863), .ZN(n12864) );
  NOR2_X1 U16256 ( .A1(n12852), .A2(n12864), .ZN(n12865) );
  AND2_X1 U16257 ( .A1(n12865), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12866) );
  NAND2_X1 U16258 ( .A1(n12867), .A2(n12866), .ZN(n12868) );
  AOI21_X1 U16259 ( .B1(n15197), .B2(n14459), .A(n14246), .ZN(n15257) );
  NOR2_X1 U16260 ( .A1(n15008), .A2(n12869), .ZN(n12870) );
  OR2_X1 U16261 ( .A1(n12823), .A2(n12870), .ZN(n15256) );
  NAND2_X1 U16262 ( .A1(n19044), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15252) );
  OAI21_X1 U16263 ( .B1(n16100), .B2(n12871), .A(n15252), .ZN(n12872) );
  AOI21_X1 U16264 ( .B1(n16090), .B2(n15001), .A(n12872), .ZN(n12873) );
  OAI21_X1 U16265 ( .B1(n15256), .B2(n16077), .A(n12873), .ZN(n12874) );
  AOI21_X1 U16266 ( .B1(n15257), .B2(n14248), .A(n12874), .ZN(n12875) );
  OAI21_X1 U16267 ( .B1(n15258), .B2(n16084), .A(n12875), .ZN(P2_U2985) );
  NAND2_X1 U16268 ( .A1(n12876), .A2(n17639), .ZN(n12890) );
  NAND2_X1 U16269 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18066) );
  NAND2_X1 U16270 ( .A1(n18678), .A2(n18066), .ZN(n18725) );
  INV_X1 U16271 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18689) );
  NOR2_X1 U16272 ( .A1(n18689), .A2(n16356), .ZN(n17705) );
  NAND2_X1 U16273 ( .A1(n18732), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18592) );
  NAND2_X1 U16274 ( .A1(n18525), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18691) );
  INV_X1 U16275 ( .A(n18691), .ZN(n18704) );
  NOR2_X1 U16276 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18735) );
  AOI21_X1 U16277 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n18735), .ZN(n18589) );
  NOR2_X1 U16278 ( .A1(n18704), .A2(n18589), .ZN(n18082) );
  NAND3_X1 U16279 ( .A1(n18729), .A2(n18678), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18423) );
  NOR2_X1 U16280 ( .A1(n18189), .A2(n18423), .ZN(n16237) );
  OR2_X1 U16281 ( .A1(n12877), .A2(n17572), .ZN(n16228) );
  XNOR2_X1 U16282 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12881) );
  NOR2_X1 U16283 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17508), .ZN(
        n16247) );
  NAND2_X1 U16284 ( .A1(n18460), .A2(n12877), .ZN(n12878) );
  OAI211_X1 U16285 ( .C1(n12879), .C2(n18592), .A(n17731), .B(n12878), .ZN(
        n16240) );
  NOR2_X1 U16286 ( .A1(n16247), .A2(n16240), .ZN(n16227) );
  OAI22_X1 U16287 ( .A1(n16228), .A2(n12881), .B1(n16227), .B2(n12880), .ZN(
        n12882) );
  AOI211_X1 U16288 ( .C1(n17530), .C2(n9710), .A(n12883), .B(n12882), .ZN(
        n12889) );
  NAND2_X1 U16289 ( .A1(n17640), .A2(n12884), .ZN(n12888) );
  INV_X1 U16290 ( .A(n12885), .ZN(n12886) );
  NAND2_X1 U16291 ( .A1(n12886), .A2(n17537), .ZN(n12887) );
  NAND2_X1 U16292 ( .A1(n12890), .A2(n10084), .ZN(P3_U2799) );
  AOI22_X1 U16293 ( .A1(n12892), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12891), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12893) );
  NAND2_X1 U16294 ( .A1(n13077), .A2(n20760), .ZN(n12898) );
  OR2_X1 U16295 ( .A1(n12897), .A2(n13638), .ZN(n13271) );
  OAI22_X1 U16296 ( .A1(n12896), .A2(n12898), .B1(n13280), .B2(n13271), .ZN(
        n13287) );
  OR2_X1 U16297 ( .A1(n13288), .A2(n20662), .ZN(n12900) );
  OAI22_X1 U16298 ( .A1(n13280), .A2(n12900), .B1(n13638), .B2(n12899), .ZN(
        n12901) );
  NAND2_X1 U16299 ( .A1(n14500), .A2(n10068), .ZN(n12918) );
  NOR4_X1 U16300 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12907) );
  NOR4_X1 U16301 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12906) );
  NOR4_X1 U16302 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12905) );
  NOR4_X1 U16303 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12904) );
  AND4_X1 U16304 ( .A1(n12907), .A2(n12906), .A3(n12905), .A4(n12904), .ZN(
        n12912) );
  NOR4_X1 U16305 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n12910) );
  NOR4_X1 U16306 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12909) );
  NOR4_X1 U16307 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12908) );
  INV_X1 U16308 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20674) );
  AND4_X1 U16309 ( .A1(n12910), .A2(n12909), .A3(n12908), .A4(n20674), .ZN(
        n12911) );
  NAND2_X1 U16310 ( .A1(n12912), .A2(n12911), .ZN(n12913) );
  INV_X1 U16311 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19124) );
  NOR2_X1 U16312 ( .A1(n15723), .A2(n19124), .ZN(n12916) );
  NOR2_X2 U16313 ( .A1(n13439), .A2(n19976), .ZN(n15720) );
  AOI22_X1 U16314 ( .A1(n15720), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15717), .ZN(n12914) );
  INV_X1 U16315 ( .A(n12914), .ZN(n12915) );
  NOR2_X1 U16316 ( .A1(n12916), .A2(n12915), .ZN(n12917) );
  NAND2_X1 U16317 ( .A1(n12918), .A2(n12917), .ZN(P1_U2873) );
  NAND2_X1 U16318 ( .A1(n12920), .A2(n12919), .ZN(n14237) );
  NAND2_X1 U16319 ( .A1(n14237), .A2(n14234), .ZN(n12925) );
  AOI21_X1 U16320 ( .B1(n12921), .B2(n14238), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14236) );
  INV_X1 U16321 ( .A(n12921), .ZN(n12922) );
  INV_X1 U16322 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14458) );
  OR3_X2 U16323 ( .A1(n12922), .A2(n10934), .A3(n14458), .ZN(n14235) );
  INV_X1 U16324 ( .A(n14235), .ZN(n12923) );
  NOR2_X1 U16325 ( .A1(n14236), .A2(n12923), .ZN(n12924) );
  XNOR2_X1 U16326 ( .A(n12925), .B(n12924), .ZN(n15184) );
  XOR2_X1 U16327 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n14246), .Z(
        n15182) );
  OAI21_X1 U16328 ( .B1(n12928), .B2(n15285), .A(n14197), .ZN(n15281) );
  AND2_X1 U16329 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12929) );
  AOI21_X1 U16330 ( .B1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n12929), .A(
        n15285), .ZN(n12926) );
  NOR2_X1 U16331 ( .A1(n15281), .A2(n12926), .ZN(n14461) );
  NOR2_X1 U16332 ( .A1(n18814), .A2(n12927), .ZN(n15177) );
  NAND2_X1 U16333 ( .A1(n14194), .A2(n12928), .ZN(n15259) );
  INV_X1 U16334 ( .A(n12929), .ZN(n12930) );
  OR2_X1 U16335 ( .A1(n15259), .A2(n12930), .ZN(n15251) );
  NOR3_X1 U16336 ( .A1(n15251), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14459), .ZN(n12931) );
  AOI211_X1 U16337 ( .C1(n14454), .C2(n19067), .A(n15177), .B(n12931), .ZN(
        n12932) );
  OAI21_X1 U16338 ( .B1(n14461), .B2(n14458), .A(n12932), .ZN(n12933) );
  OAI211_X1 U16339 ( .C1(n15184), .C2(n16163), .A(n12934), .B(n10060), .ZN(
        P2_U3016) );
  XNOR2_X1 U16340 ( .A(n12939), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14876) );
  NAND2_X1 U16341 ( .A1(n14500), .A2(n12940), .ZN(n12946) );
  INV_X1 U16342 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14504) );
  NAND2_X1 U16343 ( .A1(n15791), .A2(n13644), .ZN(n12943) );
  NAND2_X1 U16344 ( .A1(n19939), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14869) );
  OAI211_X1 U16345 ( .C1(n15795), .C2(n14504), .A(n12943), .B(n14869), .ZN(
        n12944) );
  OAI211_X1 U16346 ( .C1(n14876), .C2(n19757), .A(n12946), .B(n12945), .ZN(
        P1_U2968) );
  INV_X1 U16347 ( .A(n15991), .ZN(n18809) );
  AOI21_X1 U16348 ( .B1(n19055), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n12948), .ZN(n12949) );
  OAI21_X1 U16349 ( .B1(n18808), .B2(n19061), .A(n12949), .ZN(n12950) );
  INV_X1 U16350 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n20920) );
  NOR3_X1 U16351 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20920), .ZN(n12955) );
  NOR4_X1 U16352 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12954) );
  NAND4_X1 U16353 ( .A1(n19976), .A2(P1_W_R_N_REG_SCAN_IN), .A3(n12955), .A4(
        n12954), .ZN(U214) );
  NOR4_X1 U16354 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12959) );
  NOR4_X1 U16355 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n12958) );
  NOR4_X1 U16356 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12957) );
  NOR4_X1 U16357 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n12956) );
  NAND4_X1 U16358 ( .A1(n12959), .A2(n12958), .A3(n12957), .A4(n12956), .ZN(
        n12964) );
  NOR4_X1 U16359 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12962) );
  NOR4_X1 U16360 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n12961) );
  NOR4_X1 U16361 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n12960) );
  INV_X1 U16362 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19623) );
  NAND4_X1 U16363 ( .A1(n12962), .A2(n12961), .A3(n12960), .A4(n19623), .ZN(
        n12963) );
  OAI21_X1 U16364 ( .B1(n12964), .B2(n12963), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12965) );
  INV_X2 U16365 ( .A(n13917), .ZN(n13913) );
  NOR2_X1 U16366 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12967) );
  NOR4_X1 U16367 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12966) );
  NAND4_X1 U16368 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12967), .A4(n12966), .ZN(n12968) );
  NOR2_X1 U16369 ( .A1(n13913), .A2(n12968), .ZN(n16268) );
  NAND2_X1 U16370 ( .A1(n16268), .A2(U214), .ZN(U212) );
  NOR2_X1 U16371 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12968), .ZN(n16336)
         );
  AOI211_X1 U16372 ( .C1(n12971), .C2(n12970), .A(n12969), .B(n19602), .ZN(
        n12980) );
  AOI22_X1 U16373 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n18922), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n18912), .ZN(n12972) );
  INV_X1 U16374 ( .A(n12972), .ZN(n12979) );
  OAI22_X1 U16375 ( .A1(n12974), .A2(n18927), .B1(n18908), .B2(n12973), .ZN(
        n12978) );
  INV_X1 U16376 ( .A(n15111), .ZN(n12976) );
  INV_X1 U16377 ( .A(n15160), .ZN(n12975) );
  OAI22_X1 U16378 ( .A1(n12976), .A2(n18900), .B1(n18921), .B2(n12975), .ZN(
        n12977) );
  OR4_X1 U16379 ( .A1(n12980), .A2(n12979), .A3(n12978), .A4(n12977), .ZN(
        P2_U2832) );
  NAND2_X1 U16380 ( .A1(n18870), .A2(n18917), .ZN(n18829) );
  AOI211_X1 U16381 ( .C1(n16039), .C2(n12981), .A(n13803), .B(n18829), .ZN(
        n12995) );
  AOI22_X1 U16382 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18939), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n18912), .ZN(n12982) );
  OAI211_X1 U16383 ( .C1(n13541), .C2(n18906), .A(n12982), .B(n11123), .ZN(
        n12994) );
  OR2_X1 U16384 ( .A1(n12984), .A2(n12983), .ZN(n12986) );
  NAND2_X1 U16385 ( .A1(n12986), .A2(n12985), .ZN(n15432) );
  OAI22_X1 U16386 ( .A1(n12987), .A2(n18927), .B1(n18921), .B2(n15432), .ZN(
        n12993) );
  OAI21_X1 U16387 ( .B1(n12988), .B2(n12990), .A(n12989), .ZN(n13538) );
  NOR2_X1 U16388 ( .A1(n18870), .A2(n19602), .ZN(n18938) );
  INV_X1 U16389 ( .A(n18938), .ZN(n18816) );
  INV_X1 U16390 ( .A(n16039), .ZN(n12991) );
  OAI22_X1 U16391 ( .A1(n13538), .A2(n18900), .B1(n18816), .B2(n12991), .ZN(
        n12992) );
  OR4_X1 U16392 ( .A1(n12995), .A2(n12994), .A3(n12993), .A4(n12992), .ZN(
        P2_U2844) );
  INV_X1 U16393 ( .A(n12997), .ZN(n12996) );
  OR2_X1 U16394 ( .A1(n13491), .A2(n12996), .ZN(n15063) );
  INV_X1 U16395 ( .A(n15063), .ZN(n18936) );
  INV_X1 U16396 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13000) );
  NAND2_X1 U16397 ( .A1(n16207), .A2(n12997), .ZN(n13037) );
  INV_X1 U16398 ( .A(n13037), .ZN(n12998) );
  INV_X1 U16399 ( .A(n18751), .ZN(n13001) );
  AOI21_X1 U16400 ( .B1(n12998), .B2(n10216), .A(n13001), .ZN(n12999) );
  OAI21_X1 U16401 ( .B1(n18936), .B2(n13000), .A(n12999), .ZN(P2_U2814) );
  INV_X1 U16402 ( .A(n13135), .ZN(n16190) );
  INV_X1 U16403 ( .A(n18753), .ZN(n19729) );
  OAI21_X1 U16404 ( .B1(n13001), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n19729), 
        .ZN(n13002) );
  OAI21_X1 U16405 ( .B1(n16190), .B2(n19729), .A(n13002), .ZN(P2_U3612) );
  NAND2_X1 U16406 ( .A1(n10193), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13003) );
  AOI22_X1 U16407 ( .A1(n13306), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19697), .B2(n19715), .ZN(n13004) );
  INV_X1 U16408 ( .A(n13212), .ZN(n15454) );
  NOR2_X1 U16409 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13006) );
  NOR2_X1 U16410 ( .A1(n10193), .A2(n19727), .ZN(n13210) );
  OAI21_X1 U16411 ( .B1(n13007), .B2(n13006), .A(n13210), .ZN(n13008) );
  NOR2_X1 U16412 ( .A1(n16187), .A2(n16181), .ZN(n13498) );
  AND2_X1 U16413 ( .A1(n15461), .A2(n13009), .ZN(n13501) );
  MUX2_X1 U16414 ( .A(n10224), .B(n13005), .S(n18965), .Z(n13011) );
  OAI21_X1 U16415 ( .B1(n19710), .B2(n18951), .A(n13011), .ZN(P2_U2887) );
  INV_X1 U16416 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13958) );
  INV_X1 U16417 ( .A(n19731), .ZN(n18755) );
  OR2_X1 U16418 ( .A1(n13491), .A2(n18755), .ZN(n13013) );
  OAI21_X1 U16419 ( .B1(n13495), .B2(n13013), .A(n13133), .ZN(n13015) );
  NAND2_X1 U16420 ( .A1(n19029), .A2(n9776), .ZN(n19006) );
  NOR2_X1 U16421 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13490), .ZN(n19026) );
  INV_X1 U16422 ( .A(n19026), .ZN(n19031) );
  INV_X1 U16423 ( .A(n19031), .ZN(n19041) );
  AOI22_X1 U16424 ( .A1(n19026), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13016) );
  OAI21_X1 U16425 ( .B1(n13958), .B2(n19006), .A(n13016), .ZN(P2_U2934) );
  AOI22_X1 U16426 ( .A1(n19041), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13017) );
  OAI21_X1 U16427 ( .B1(n15128), .B2(n19006), .A(n13017), .ZN(P2_U2924) );
  INV_X1 U16428 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13916) );
  AOI22_X1 U16429 ( .A1(n19041), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13018) );
  OAI21_X1 U16430 ( .B1(n13916), .B2(n19006), .A(n13018), .ZN(P2_U2932) );
  AOI22_X1 U16431 ( .A1(n19041), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13019) );
  OAI21_X1 U16432 ( .B1(n11132), .B2(n19006), .A(n13019), .ZN(P2_U2927) );
  AOI22_X1 U16433 ( .A1(n19041), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13020) );
  OAI21_X1 U16434 ( .B1(n15122), .B2(n19006), .A(n13020), .ZN(P2_U2923) );
  INV_X1 U16435 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15116) );
  AOI22_X1 U16436 ( .A1(n19041), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13021) );
  OAI21_X1 U16437 ( .B1(n15116), .B2(n19006), .A(n13021), .ZN(P2_U2922) );
  INV_X1 U16438 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13120) );
  AOI22_X1 U16439 ( .A1(n19041), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13022) );
  OAI21_X1 U16440 ( .B1(n13120), .B2(n19006), .A(n13022), .ZN(P2_U2921) );
  INV_X1 U16441 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13111) );
  AOI22_X1 U16442 ( .A1(n19041), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13023) );
  OAI21_X1 U16443 ( .B1(n13111), .B2(n19006), .A(n13023), .ZN(P2_U2935) );
  INV_X1 U16444 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14041) );
  AOI22_X1 U16445 ( .A1(n19041), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13024) );
  OAI21_X1 U16446 ( .B1(n14041), .B2(n19006), .A(n13024), .ZN(P2_U2930) );
  INV_X1 U16447 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13998) );
  AOI22_X1 U16448 ( .A1(n19026), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13025) );
  OAI21_X1 U16449 ( .B1(n13998), .B2(n19006), .A(n13025), .ZN(P2_U2933) );
  INV_X1 U16450 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15158) );
  AOI22_X1 U16451 ( .A1(n19041), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13026) );
  OAI21_X1 U16452 ( .B1(n15158), .B2(n19006), .A(n13026), .ZN(P2_U2928) );
  INV_X1 U16453 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n15167) );
  AOI22_X1 U16454 ( .A1(n19041), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13027) );
  OAI21_X1 U16455 ( .B1(n15167), .B2(n19006), .A(n13027), .ZN(P2_U2929) );
  AOI22_X1 U16456 ( .A1(n19041), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13028) );
  OAI21_X1 U16457 ( .B1(n15139), .B2(n19006), .A(n13028), .ZN(P2_U2926) );
  INV_X1 U16458 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13129) );
  AOI22_X1 U16459 ( .A1(n19041), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13029) );
  OAI21_X1 U16460 ( .B1(n13129), .B2(n19006), .A(n13029), .ZN(P2_U2925) );
  INV_X1 U16461 ( .A(n20128), .ZN(n20743) );
  INV_X1 U16462 ( .A(n20743), .ZN(n20580) );
  NAND2_X1 U16463 ( .A1(n20580), .A2(n20957), .ZN(n19754) );
  INV_X1 U16464 ( .A(n19754), .ZN(n13030) );
  NOR2_X1 U16465 ( .A1(n13030), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13035)
         );
  AND2_X1 U16466 ( .A1(n13079), .A2(n13077), .ZN(n13068) );
  NAND2_X1 U16467 ( .A1(n13068), .A2(n13183), .ZN(n14491) );
  NOR2_X1 U16468 ( .A1(n13065), .A2(n19751), .ZN(n13031) );
  INV_X1 U16469 ( .A(n13638), .ZN(n13032) );
  OAI21_X1 U16470 ( .B1(n13033), .B2(n13032), .A(n20758), .ZN(n13034) );
  OAI21_X1 U16471 ( .B1(n13035), .B2(n20758), .A(n13034), .ZN(P1_U3487) );
  NAND2_X1 U16472 ( .A1(n10216), .A2(n19726), .ZN(n13036) );
  NOR2_X1 U16473 ( .A1(n13037), .A2(n13036), .ZN(n13038) );
  AOI22_X1 U16474 ( .A1(n13060), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n13107), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13041) );
  INV_X1 U16475 ( .A(n13038), .ZN(n13039) );
  NOR2_X2 U16476 ( .A1(n13039), .A2(n19737), .ZN(n13125) );
  AOI22_X1 U16477 ( .A1(n13917), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13913), .ZN(n19116) );
  INV_X1 U16478 ( .A(n19116), .ZN(n13040) );
  NAND2_X1 U16479 ( .A1(n13125), .A2(n13040), .ZN(n13087) );
  NAND2_X1 U16480 ( .A1(n13041), .A2(n13087), .ZN(P2_U2973) );
  AOI22_X1 U16481 ( .A1(n13060), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n13107), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13042) );
  AOI22_X1 U16482 ( .A1(n13917), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13913), .ZN(n19111) );
  INV_X1 U16483 ( .A(n19111), .ZN(n18996) );
  NAND2_X1 U16484 ( .A1(n13125), .A2(n18996), .ZN(n13105) );
  NAND2_X1 U16485 ( .A1(n13042), .A2(n13105), .ZN(P2_U2972) );
  AOI22_X1 U16486 ( .A1(n13060), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n13107), .ZN(n13043) );
  OAI22_X1 U16487 ( .A1(n13913), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13917), .ZN(n19106) );
  INV_X1 U16488 ( .A(n19106), .ZN(n15992) );
  NAND2_X1 U16489 ( .A1(n13125), .A2(n15992), .ZN(n13093) );
  NAND2_X1 U16490 ( .A1(n13043), .A2(n13093), .ZN(P2_U2971) );
  AOI22_X1 U16491 ( .A1(n13060), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n13107), .ZN(n13044) );
  AOI22_X1 U16492 ( .A1(n13917), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13913), .ZN(n13999) );
  INV_X1 U16493 ( .A(n13999), .ZN(n13478) );
  NAND2_X1 U16494 ( .A1(n13125), .A2(n13478), .ZN(n13091) );
  NAND2_X1 U16495 ( .A1(n13044), .A2(n13091), .ZN(P2_U2969) );
  AOI22_X1 U16496 ( .A1(n13060), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_1__SCAN_IN), .B2(n13107), .ZN(n13045) );
  AOI22_X1 U16497 ( .A1(n13917), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13913), .ZN(n13959) );
  INV_X1 U16498 ( .A(n13959), .ZN(n13328) );
  NAND2_X1 U16499 ( .A1(n13125), .A2(n13328), .ZN(n13049) );
  NAND2_X1 U16500 ( .A1(n13045), .A2(n13049), .ZN(P2_U2968) );
  AOI22_X1 U16501 ( .A1(n13060), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n13107), .ZN(n13048) );
  INV_X1 U16502 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13369) );
  OR2_X1 U16503 ( .A1(n13913), .A2(n13369), .ZN(n13047) );
  NAND2_X1 U16504 ( .A1(n13913), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13046) );
  NAND2_X1 U16505 ( .A1(n13047), .A2(n13046), .ZN(n15118) );
  NAND2_X1 U16506 ( .A1(n13125), .A2(n15118), .ZN(n13099) );
  NAND2_X1 U16507 ( .A1(n13048), .A2(n13099), .ZN(P2_U2980) );
  AOI22_X1 U16508 ( .A1(n13060), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n13107), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13050) );
  NAND2_X1 U16509 ( .A1(n13050), .A2(n13049), .ZN(P2_U2953) );
  AOI22_X1 U16510 ( .A1(n13060), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n13107), .ZN(n13053) );
  INV_X1 U16511 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n14017) );
  OR2_X1 U16512 ( .A1(n13913), .A2(n14017), .ZN(n13052) );
  NAND2_X1 U16513 ( .A1(n13913), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13051) );
  NAND2_X1 U16514 ( .A1(n13052), .A2(n13051), .ZN(n15130) );
  NAND2_X1 U16515 ( .A1(n13125), .A2(n15130), .ZN(n13101) );
  NAND2_X1 U16516 ( .A1(n13053), .A2(n13101), .ZN(P2_U2978) );
  AOI22_X1 U16517 ( .A1(n13060), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n13107), .ZN(n13056) );
  INV_X1 U16518 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13865) );
  OR2_X1 U16519 ( .A1(n13913), .A2(n13865), .ZN(n13055) );
  NAND2_X1 U16520 ( .A1(n13913), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13054) );
  NAND2_X1 U16521 ( .A1(n13055), .A2(n13054), .ZN(n15142) );
  NAND2_X1 U16522 ( .A1(n13125), .A2(n15142), .ZN(n13097) );
  NAND2_X1 U16523 ( .A1(n13056), .A2(n13097), .ZN(P2_U2976) );
  AOI22_X1 U16524 ( .A1(n13060), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n13107), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13058) );
  AOI22_X1 U16525 ( .A1(n13917), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13913), .ZN(n19127) );
  INV_X1 U16526 ( .A(n19127), .ZN(n13057) );
  NAND2_X1 U16527 ( .A1(n13125), .A2(n13057), .ZN(n13103) );
  NAND2_X1 U16528 ( .A1(n13058), .A2(n13103), .ZN(P2_U2974) );
  AOI22_X1 U16529 ( .A1(n13060), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n13107), .ZN(n13059) );
  AOI22_X1 U16530 ( .A1(n13917), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13913), .ZN(n19101) );
  INV_X1 U16531 ( .A(n19101), .ZN(n13594) );
  NAND2_X1 U16532 ( .A1(n13125), .A2(n13594), .ZN(n13089) );
  NAND2_X1 U16533 ( .A1(n13059), .A2(n13089), .ZN(P2_U2970) );
  INV_X1 U16534 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13062) );
  INV_X1 U16535 ( .A(n13125), .ZN(n13110) );
  AOI22_X1 U16536 ( .A1(n13917), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13913), .ZN(n13631) );
  INV_X1 U16537 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13061) );
  OAI222_X1 U16538 ( .A1(n13062), .A2(n13133), .B1(n13110), .B2(n13631), .C1(
        n13061), .C2(n13112), .ZN(P2_U2982) );
  INV_X1 U16539 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13064) );
  OAI22_X1 U16540 ( .A1(n13913), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13917), .ZN(n18973) );
  INV_X1 U16541 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13063) );
  OAI222_X1 U16542 ( .A1(n13064), .A2(n13112), .B1(n13110), .B2(n18973), .C1(
        n13063), .C2(n13133), .ZN(P2_U2967) );
  INV_X1 U16543 ( .A(n13065), .ZN(n13067) );
  NAND2_X1 U16544 ( .A1(n13280), .A2(n13638), .ZN(n13066) );
  OAI21_X1 U16545 ( .B1(n13068), .B2(n13067), .A(n13066), .ZN(n19752) );
  NAND3_X1 U16546 ( .A1(n13069), .A2(n13638), .A3(n15604), .ZN(n13070) );
  AND2_X1 U16547 ( .A1(n13070), .A2(n20760), .ZN(n20762) );
  NOR2_X1 U16548 ( .A1(n19752), .A2(n20762), .ZN(n15561) );
  OR2_X1 U16549 ( .A1(n15561), .A2(n19751), .ZN(n13084) );
  INV_X1 U16550 ( .A(n13084), .ZN(n19759) );
  INV_X1 U16551 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13086) );
  INV_X1 U16552 ( .A(n13273), .ZN(n13082) );
  NAND4_X1 U16553 ( .A1(n19978), .A2(n13073), .A3(n13072), .A4(n13071), .ZN(
        n13075) );
  OAI21_X1 U16554 ( .B1(n13076), .B2(n13075), .A(n13074), .ZN(n13080) );
  INV_X1 U16555 ( .A(n13077), .ZN(n13078) );
  AOI22_X1 U16556 ( .A1(n13080), .A2(n13280), .B1(n13079), .B2(n13078), .ZN(
        n13081) );
  OAI21_X1 U16557 ( .B1(n13082), .B2(n13280), .A(n13081), .ZN(n13083) );
  NAND2_X1 U16558 ( .A1(n13083), .A2(n20013), .ZN(n15562) );
  OR2_X1 U16559 ( .A1(n13084), .A2(n15562), .ZN(n13085) );
  OAI21_X1 U16560 ( .B1(n19759), .B2(n13086), .A(n13085), .ZN(P1_U3484) );
  AOI22_X1 U16561 ( .A1(n13130), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n13107), .ZN(n13088) );
  NAND2_X1 U16562 ( .A1(n13088), .A2(n13087), .ZN(P2_U2958) );
  AOI22_X1 U16563 ( .A1(n13130), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n13107), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13090) );
  NAND2_X1 U16564 ( .A1(n13090), .A2(n13089), .ZN(P2_U2955) );
  AOI22_X1 U16565 ( .A1(n13130), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n13107), .ZN(n13092) );
  NAND2_X1 U16566 ( .A1(n13092), .A2(n13091), .ZN(P2_U2954) );
  AOI22_X1 U16567 ( .A1(n13130), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n13107), .ZN(n13094) );
  NAND2_X1 U16568 ( .A1(n13094), .A2(n13093), .ZN(P2_U2956) );
  AOI22_X1 U16569 ( .A1(n13130), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n13107), .ZN(n13096) );
  AOI22_X1 U16570 ( .A1(n13917), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n13913), .ZN(n15153) );
  INV_X1 U16571 ( .A(n15153), .ZN(n13095) );
  NAND2_X1 U16572 ( .A1(n13125), .A2(n13095), .ZN(n13108) );
  NAND2_X1 U16573 ( .A1(n13096), .A2(n13108), .ZN(P2_U2960) );
  AOI22_X1 U16574 ( .A1(n13130), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n13107), .ZN(n13098) );
  NAND2_X1 U16575 ( .A1(n13098), .A2(n13097), .ZN(P2_U2961) );
  AOI22_X1 U16576 ( .A1(n13130), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n13107), .ZN(n13100) );
  NAND2_X1 U16577 ( .A1(n13100), .A2(n13099), .ZN(P2_U2965) );
  AOI22_X1 U16578 ( .A1(n13130), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n13107), .ZN(n13102) );
  NAND2_X1 U16579 ( .A1(n13102), .A2(n13101), .ZN(P2_U2963) );
  AOI22_X1 U16580 ( .A1(n13130), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n13107), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13104) );
  NAND2_X1 U16581 ( .A1(n13104), .A2(n13103), .ZN(P2_U2959) );
  AOI22_X1 U16582 ( .A1(n13130), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n13107), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13106) );
  NAND2_X1 U16583 ( .A1(n13106), .A2(n13105), .ZN(P2_U2957) );
  AOI22_X1 U16584 ( .A1(n13130), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_8__SCAN_IN), .B2(n13107), .ZN(n13109) );
  NAND2_X1 U16585 ( .A1(n13109), .A2(n13108), .ZN(P2_U2975) );
  INV_X1 U16586 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13113) );
  OAI222_X1 U16587 ( .A1(n13113), .A2(n13112), .B1(n13133), .B2(n13111), .C1(
        n13110), .C2(n18973), .ZN(P2_U2952) );
  INV_X1 U16588 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19019) );
  NAND2_X1 U16589 ( .A1(n13130), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13116) );
  INV_X1 U16590 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16297) );
  OR2_X1 U16591 ( .A1(n13913), .A2(n16297), .ZN(n13115) );
  NAND2_X1 U16592 ( .A1(n13913), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13114) );
  NAND2_X1 U16593 ( .A1(n13115), .A2(n13114), .ZN(n18992) );
  NAND2_X1 U16594 ( .A1(n13125), .A2(n18992), .ZN(n13127) );
  OAI211_X1 U16595 ( .C1(n19019), .C2(n13133), .A(n13116), .B(n13127), .ZN(
        P2_U2977) );
  NAND2_X1 U16596 ( .A1(n13130), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13119) );
  INV_X1 U16597 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14685) );
  OR2_X1 U16598 ( .A1(n13913), .A2(n14685), .ZN(n13118) );
  NAND2_X1 U16599 ( .A1(n13913), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13117) );
  AND2_X1 U16600 ( .A1(n13118), .A2(n13117), .ZN(n14452) );
  INV_X1 U16601 ( .A(n14452), .ZN(n18985) );
  NAND2_X1 U16602 ( .A1(n13125), .A2(n18985), .ZN(n13121) );
  OAI211_X1 U16603 ( .C1(n13120), .C2(n13133), .A(n13119), .B(n13121), .ZN(
        P2_U2966) );
  INV_X1 U16604 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19011) );
  NAND2_X1 U16605 ( .A1(n13130), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13122) );
  OAI211_X1 U16606 ( .C1(n19011), .C2(n13133), .A(n13122), .B(n13121), .ZN(
        P2_U2981) );
  INV_X1 U16607 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19014) );
  NAND2_X1 U16608 ( .A1(n13130), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13126) );
  INV_X1 U16609 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16294) );
  OR2_X1 U16610 ( .A1(n13913), .A2(n16294), .ZN(n13124) );
  NAND2_X1 U16611 ( .A1(n13913), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13123) );
  AND2_X1 U16612 ( .A1(n13124), .A2(n13123), .ZN(n15123) );
  INV_X1 U16613 ( .A(n15123), .ZN(n18988) );
  NAND2_X1 U16614 ( .A1(n13125), .A2(n18988), .ZN(n13131) );
  OAI211_X1 U16615 ( .C1(n19014), .C2(n13133), .A(n13126), .B(n13131), .ZN(
        P2_U2979) );
  NAND2_X1 U16616 ( .A1(n13130), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13128) );
  OAI211_X1 U16617 ( .C1(n13129), .C2(n13133), .A(n13128), .B(n13127), .ZN(
        P2_U2962) );
  NAND2_X1 U16618 ( .A1(n13130), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13132) );
  OAI211_X1 U16619 ( .C1(n15122), .C2(n13133), .A(n13132), .B(n13131), .ZN(
        P2_U2964) );
  NAND2_X1 U16620 ( .A1(n16187), .A2(n13134), .ZN(n13137) );
  NAND4_X1 U16621 ( .A1(n13135), .A2(n16183), .A3(n9729), .A4(n19726), .ZN(
        n13136) );
  NAND2_X1 U16622 ( .A1(n13137), .A2(n13136), .ZN(n13497) );
  INV_X1 U16623 ( .A(n13497), .ZN(n13139) );
  NAND2_X1 U16624 ( .A1(n13139), .A2(n13138), .ZN(n13140) );
  NAND2_X1 U16625 ( .A1(n15168), .A2(n13141), .ZN(n13632) );
  XNOR2_X1 U16626 ( .A(n13143), .B(n13142), .ZN(n13981) );
  INV_X1 U16627 ( .A(n13981), .ZN(n18901) );
  INV_X1 U16628 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19028) );
  OAI222_X1 U16629 ( .A1(n13632), .A2(n19116), .B1(n18901), .B2(n19004), .C1(
        n19028), .C2(n15168), .ZN(P2_U2913) );
  INV_X1 U16630 ( .A(n13145), .ZN(n13146) );
  OAI21_X1 U16631 ( .B1(n13148), .B2(n13147), .A(n13146), .ZN(n16160) );
  INV_X1 U16632 ( .A(n16160), .ZN(n18924) );
  NOR2_X1 U16633 ( .A1(n19710), .A2(n16160), .ZN(n13327) );
  INV_X1 U16634 ( .A(n13327), .ZN(n13149) );
  INV_X1 U16635 ( .A(n18998), .ZN(n15147) );
  OAI211_X1 U16636 ( .C1(n18937), .C2(n18924), .A(n13149), .B(n15147), .ZN(
        n13151) );
  AOI22_X1 U16637 ( .A1(n18924), .A2(n18980), .B1(n18995), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n13150) );
  OAI211_X1 U16638 ( .C1(n13632), .C2(n18973), .A(n13151), .B(n13150), .ZN(
        P2_U2919) );
  AOI21_X1 U16639 ( .B1(n13154), .B2(n13153), .A(n13152), .ZN(n15058) );
  INV_X1 U16640 ( .A(n15058), .ZN(n19690) );
  NAND2_X1 U16641 ( .A1(n16143), .A2(n9761), .ZN(n13159) );
  AOI221_X1 U16642 ( .B1(n13156), .B2(n13155), .C1(n13172), .C2(n13155), .A(
        n19079), .ZN(n13157) );
  INV_X1 U16643 ( .A(n13157), .ZN(n13158) );
  OR2_X1 U16644 ( .A1(n11123), .A2(n19624), .ZN(n13174) );
  NAND4_X1 U16645 ( .A1(n13160), .A2(n13159), .A3(n13158), .A4(n13174), .ZN(
        n13169) );
  AOI21_X1 U16646 ( .B1(n13163), .B2(n13162), .A(n13161), .ZN(n13173) );
  INV_X1 U16647 ( .A(n13173), .ZN(n13167) );
  NAND2_X1 U16648 ( .A1(n13165), .A2(n13164), .ZN(n13177) );
  NAND3_X1 U16649 ( .A1(n13178), .A2(n19069), .A3(n13177), .ZN(n13166) );
  OAI21_X1 U16650 ( .B1(n13167), .B2(n19074), .A(n13166), .ZN(n13168) );
  AOI211_X1 U16651 ( .C1(n19690), .C2(n19067), .A(n13169), .B(n13168), .ZN(
        n13170) );
  OAI21_X1 U16652 ( .B1(n13172), .B2(n13171), .A(n13170), .ZN(P2_U3044) );
  INV_X1 U16653 ( .A(n15051), .ZN(n15052) );
  NAND2_X1 U16654 ( .A1(n13173), .A2(n14248), .ZN(n13175) );
  OAI211_X1 U16655 ( .C1(n16100), .C2(n15057), .A(n13175), .B(n13174), .ZN(
        n13176) );
  AOI21_X1 U16656 ( .B1(n16090), .B2(n15052), .A(n13176), .ZN(n13180) );
  NAND3_X1 U16657 ( .A1(n13178), .A2(n19056), .A3(n13177), .ZN(n13179) );
  OAI211_X1 U16658 ( .C1(n13226), .C2(n16077), .A(n13180), .B(n13179), .ZN(
        P2_U3012) );
  INV_X1 U16659 ( .A(n15548), .ZN(n13182) );
  NAND2_X1 U16660 ( .A1(n13182), .A2(n13181), .ZN(n13186) );
  INV_X1 U16661 ( .A(n15604), .ZN(n15571) );
  NAND2_X1 U16662 ( .A1(n15571), .A2(n13183), .ZN(n13184) );
  NOR2_X1 U16663 ( .A1(n13280), .A2(n13184), .ZN(n13185) );
  NAND2_X1 U16664 ( .A1(n19897), .A2(n19978), .ZN(n19872) );
  NOR2_X1 U16665 ( .A1(n20957), .A2(n20244), .ZN(n15941) );
  NAND2_X1 U16666 ( .A1(n15945), .A2(n15941), .ZN(n19889) );
  AOI22_X1 U16667 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13188) );
  OAI21_X1 U16668 ( .B1(n14710), .B2(n19872), .A(n13188), .ZN(P1_U2912) );
  AOI22_X1 U16669 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13189) );
  OAI21_X1 U16670 ( .B1(n14691), .B2(n19872), .A(n13189), .ZN(P1_U2908) );
  AOI22_X1 U16671 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13190) );
  OAI21_X1 U16672 ( .B1(n14701), .B2(n19872), .A(n13190), .ZN(P1_U2910) );
  INV_X1 U16673 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13192) );
  AOI22_X1 U16674 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13191) );
  OAI21_X1 U16675 ( .B1(n13192), .B2(n19872), .A(n13191), .ZN(P1_U2917) );
  INV_X1 U16676 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13194) );
  AOI22_X1 U16677 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13193) );
  OAI21_X1 U16678 ( .B1(n13194), .B2(n19872), .A(n13193), .ZN(P1_U2906) );
  INV_X1 U16679 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13196) );
  AOI22_X1 U16680 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13195) );
  OAI21_X1 U16681 ( .B1(n13196), .B2(n19872), .A(n13195), .ZN(P1_U2913) );
  INV_X1 U16682 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13198) );
  AOI22_X1 U16683 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13197) );
  OAI21_X1 U16684 ( .B1(n13198), .B2(n19872), .A(n13197), .ZN(P1_U2919) );
  AOI22_X1 U16685 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13199) );
  OAI21_X1 U16686 ( .B1(n14696), .B2(n19872), .A(n13199), .ZN(P1_U2909) );
  AOI22_X1 U16687 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13200) );
  OAI21_X1 U16688 ( .B1(n12088), .B2(n19872), .A(n13200), .ZN(P1_U2920) );
  AOI22_X1 U16689 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13201) );
  OAI21_X1 U16690 ( .B1(n12181), .B2(n19872), .A(n13201), .ZN(P1_U2916) );
  AOI22_X1 U16691 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13202) );
  OAI21_X1 U16692 ( .B1(n14729), .B2(n19872), .A(n13202), .ZN(P1_U2918) );
  OR2_X1 U16693 ( .A1(n13204), .A2(n13203), .ZN(n13205) );
  AND2_X1 U16694 ( .A1(n13205), .A2(n13228), .ZN(n18890) );
  INV_X1 U16695 ( .A(n18890), .ZN(n16139) );
  INV_X1 U16696 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19025) );
  OAI222_X1 U16697 ( .A1(n13632), .A2(n19127), .B1(n16139), .B2(n19004), .C1(
        n19025), .C2(n15168), .ZN(P2_U2912) );
  NAND2_X1 U16698 ( .A1(n19708), .A2(n19715), .ZN(n19442) );
  INV_X1 U16699 ( .A(n19442), .ZN(n13207) );
  NOR2_X1 U16700 ( .A1(n19407), .A2(n13207), .ZN(n19284) );
  AND2_X1 U16701 ( .A1(n19284), .A2(n19697), .ZN(n19376) );
  AOI21_X1 U16702 ( .B1(n13306), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19376), .ZN(n13208) );
  NAND2_X1 U16703 ( .A1(n13234), .A2(n13235), .ZN(n13233) );
  NAND2_X1 U16704 ( .A1(n15454), .A2(n13213), .ZN(n13214) );
  INV_X1 U16705 ( .A(n13308), .ZN(n13215) );
  NOR2_X1 U16706 ( .A1(n19407), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13217) );
  NOR2_X1 U16707 ( .A1(n13303), .A2(n13217), .ZN(n19215) );
  AOI22_X1 U16708 ( .A1(n13306), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19697), .B2(n19215), .ZN(n13218) );
  INV_X1 U16709 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13220) );
  INV_X2 U16710 ( .A(n18965), .ZN(n13516) );
  MUX2_X1 U16711 ( .A(n13226), .B(n13225), .S(n13516), .Z(n13227) );
  OAI21_X1 U16712 ( .B1(n15488), .B2(n18951), .A(n13227), .ZN(P2_U2885) );
  NAND2_X1 U16713 ( .A1(n13229), .A2(n13228), .ZN(n13232) );
  INV_X1 U16714 ( .A(n13230), .ZN(n13231) );
  NAND2_X1 U16715 ( .A1(n13232), .A2(n13231), .ZN(n16123) );
  INV_X1 U16716 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19023) );
  OAI222_X1 U16717 ( .A1(n13632), .A2(n15153), .B1(n16123), .B2(n19004), .C1(
        n19023), .C2(n15168), .ZN(P2_U2911) );
  MUX2_X1 U16718 ( .A(n13236), .B(n13206), .S(n18965), .Z(n13237) );
  OAI21_X1 U16719 ( .B1(n19698), .B2(n18951), .A(n13237), .ZN(P2_U2886) );
  INV_X1 U16720 ( .A(n15142), .ZN(n13241) );
  OR2_X1 U16721 ( .A1(n13238), .A2(n13230), .ZN(n13240) );
  NAND2_X1 U16722 ( .A1(n13240), .A2(n13239), .ZN(n18877) );
  INV_X1 U16723 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19021) );
  OAI222_X1 U16724 ( .A1(n13632), .A2(n13241), .B1(n18877), .B2(n19004), .C1(
        n19021), .C2(n15168), .ZN(P2_U2910) );
  OAI21_X1 U16725 ( .B1(n13243), .B2(n13242), .A(n13414), .ZN(n13665) );
  OR2_X1 U16726 ( .A1(n13245), .A2(n13244), .ZN(n13246) );
  NAND2_X1 U16727 ( .A1(n13247), .A2(n13246), .ZN(n13656) );
  AOI22_X1 U16728 ( .A1(n14670), .A2(n13656), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14669), .ZN(n13248) );
  OAI21_X1 U16729 ( .B1(n13665), .B2(n14672), .A(n13248), .ZN(P1_U2871) );
  XNOR2_X1 U16730 ( .A(n13249), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13359) );
  OAI21_X1 U16731 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n15865), .A(
        n15881), .ZN(n19968) );
  INV_X1 U16732 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20748) );
  NOR2_X1 U16733 ( .A1(n15908), .A2(n20748), .ZN(n13354) );
  INV_X1 U16734 ( .A(n13656), .ZN(n13250) );
  NOR2_X1 U16735 ( .A1(n15909), .A2(n13250), .ZN(n13251) );
  AOI211_X1 U16736 ( .C1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n19968), .A(
        n13354), .B(n13251), .ZN(n13254) );
  NAND3_X1 U16737 ( .A1(n15907), .A2(n13252), .A3(n11656), .ZN(n13253) );
  OAI211_X1 U16738 ( .C1(n13359), .C2(n15872), .A(n13254), .B(n13253), .ZN(
        P1_U3030) );
  AND2_X1 U16739 ( .A1(n20763), .A2(n20662), .ZN(n13255) );
  OR2_X1 U16740 ( .A1(n19928), .A2(n19992), .ZN(n13441) );
  INV_X1 U16741 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13261) );
  NOR2_X2 U16742 ( .A1(n19928), .A2(n13256), .ZN(n19915) );
  INV_X1 U16743 ( .A(n19915), .ZN(n13260) );
  INV_X1 U16744 ( .A(DATAI_15_), .ZN(n13258) );
  INV_X1 U16745 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13257) );
  MUX2_X1 U16746 ( .A(n13258), .B(n13257), .S(n19976), .Z(n14739) );
  INV_X1 U16747 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13259) );
  OAI222_X1 U16748 ( .A1(n13441), .A2(n13261), .B1(n13260), .B2(n14739), .C1(
        n13259), .C2(n13360), .ZN(P1_U2967) );
  NOR2_X1 U16749 ( .A1(n11626), .A2(n13263), .ZN(n13264) );
  AND2_X1 U16750 ( .A1(n13265), .A2(n13264), .ZN(n13266) );
  NAND3_X1 U16751 ( .A1(n13267), .A2(n13266), .A3(n12896), .ZN(n13549) );
  INV_X1 U16752 ( .A(n13549), .ZN(n14982) );
  INV_X1 U16753 ( .A(n13268), .ZN(n13269) );
  OR2_X1 U16754 ( .A1(n13549), .A2(n13269), .ZN(n13558) );
  XNOR2_X1 U16755 ( .A(n14984), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13279) );
  INV_X1 U16756 ( .A(n13271), .ZN(n13272) );
  OR2_X1 U16757 ( .A1(n13273), .A2(n13272), .ZN(n13555) );
  XNOR2_X1 U16758 ( .A(n13274), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13275) );
  AOI22_X1 U16759 ( .A1(n13555), .A2(n13279), .B1(n15548), .B2(n13275), .ZN(
        n13276) );
  OAI21_X1 U16760 ( .B1(n13558), .B2(n13279), .A(n13276), .ZN(n13277) );
  INV_X1 U16761 ( .A(n13277), .ZN(n13278) );
  OAI21_X1 U16762 ( .B1(n13262), .B2(n14982), .A(n13278), .ZN(n13559) );
  NOR2_X1 U16763 ( .A1(n20957), .A2(n19933), .ZN(n14987) );
  INV_X1 U16764 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n20933) );
  OAI22_X1 U16765 ( .A1(n20933), .A2(n11656), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14988) );
  INV_X1 U16766 ( .A(n14988), .ZN(n13282) );
  INV_X1 U16767 ( .A(n13279), .ZN(n13281) );
  AOI222_X1 U16768 ( .A1(n13559), .A2(n14983), .B1(n14987), .B2(n13282), .C1(
        n13281), .C2(n15582), .ZN(n13296) );
  INV_X1 U16769 ( .A(n13283), .ZN(n13285) );
  OAI211_X1 U16770 ( .C1(n13640), .C2(n19996), .A(n13285), .B(n13284), .ZN(
        n13286) );
  INV_X1 U16771 ( .A(n13286), .ZN(n13294) );
  INV_X1 U16772 ( .A(n13287), .ZN(n13293) );
  OAI21_X1 U16773 ( .B1(n15548), .B2(n11626), .A(n15571), .ZN(n13289) );
  NAND2_X1 U16774 ( .A1(n13289), .A2(n13288), .ZN(n13291) );
  NAND3_X1 U16775 ( .A1(n13291), .A2(n20760), .A3(n13290), .ZN(n13292) );
  INV_X1 U16776 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19758) );
  NAND2_X1 U16777 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15941), .ZN(n15947) );
  OAI22_X1 U16778 ( .A1(n13562), .A2(n19751), .B1(n19758), .B2(n15947), .ZN(
        n13316) );
  AOI21_X1 U16779 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n15945), .A(n13316), 
        .ZN(n14991) );
  NAND2_X1 U16780 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n14991), .ZN(
        n13295) );
  OAI21_X1 U16781 ( .B1(n13296), .B2(n14991), .A(n13295), .ZN(P1_U3472) );
  INV_X1 U16782 ( .A(n13297), .ZN(n13298) );
  NAND2_X1 U16783 ( .A1(n13299), .A2(n13298), .ZN(n13300) );
  OAI21_X1 U16784 ( .B1(n13303), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19697), .ZN(n13304) );
  NOR2_X1 U16785 ( .A1(n19585), .A2(n13304), .ZN(n13305) );
  AOI21_X1 U16786 ( .B1(n13306), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13305), .ZN(n13307) );
  INV_X1 U16787 ( .A(n13335), .ZN(n13310) );
  AND2_X1 U16788 ( .A1(n14392), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13311) );
  INV_X1 U16789 ( .A(n13311), .ZN(n13309) );
  NAND2_X1 U16790 ( .A1(n13310), .A2(n13309), .ZN(n13312) );
  NAND2_X1 U16791 ( .A1(n13335), .A2(n13311), .ZN(n13700) );
  MUX2_X1 U16792 ( .A(n10598), .B(n16148), .S(n18965), .Z(n13313) );
  OAI21_X1 U16793 ( .B1(n19479), .B2(n18951), .A(n13313), .ZN(P2_U2884) );
  INV_X1 U16794 ( .A(n20127), .ZN(n20443) );
  NOR2_X1 U16795 ( .A1(n13314), .A2(n20443), .ZN(n13315) );
  XNOR2_X1 U16796 ( .A(n13315), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19841) );
  INV_X1 U16797 ( .A(n12896), .ZN(n13317) );
  NAND3_X1 U16798 ( .A1(n13317), .A2(n14983), .A3(n13316), .ZN(n13319) );
  INV_X1 U16799 ( .A(n14991), .ZN(n20730) );
  OAI22_X1 U16800 ( .A1(n19841), .A2(n13319), .B1(n13318), .B2(n20730), .ZN(
        P1_U3468) );
  INV_X1 U16801 ( .A(n20089), .ZN(n13570) );
  OAI22_X1 U16802 ( .A1(n13570), .A2(n14982), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14978), .ZN(n15547) );
  OAI22_X1 U16803 ( .A1(n20957), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20726), .ZN(n13320) );
  AOI21_X1 U16804 ( .B1(n15547), .B2(n14983), .A(n13320), .ZN(n13322) );
  AOI21_X1 U16805 ( .B1(n15548), .B2(n14983), .A(n14991), .ZN(n13321) );
  OAI22_X1 U16806 ( .A1(n13322), .A2(n14991), .B1(n13321), .B2(n11930), .ZN(
        P1_U3474) );
  XNOR2_X1 U16807 ( .A(n13324), .B(n13323), .ZN(n19706) );
  OR2_X1 U16808 ( .A1(n19702), .A2(n19706), .ZN(n13473) );
  NAND2_X1 U16809 ( .A1(n19702), .A2(n19706), .ZN(n13325) );
  NAND2_X1 U16810 ( .A1(n13473), .A2(n13325), .ZN(n13326) );
  NOR2_X1 U16811 ( .A1(n13326), .A2(n13327), .ZN(n13475) );
  AOI21_X1 U16812 ( .B1(n13327), .B2(n13326), .A(n13475), .ZN(n13331) );
  AOI22_X1 U16813 ( .A1(n18997), .A2(n13328), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n18995), .ZN(n13330) );
  NAND2_X1 U16814 ( .A1(n18980), .A2(n19706), .ZN(n13329) );
  OAI211_X1 U16815 ( .C1(n13331), .C2(n18998), .A(n13330), .B(n13329), .ZN(
        P2_U2918) );
  AND2_X1 U16816 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n10193), .ZN(
        n13332) );
  AOI21_X1 U16817 ( .B1(n13334), .B2(n13333), .A(n13332), .ZN(n13697) );
  NAND2_X1 U16818 ( .A1(n13335), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13336) );
  AND2_X1 U16819 ( .A1(n14392), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13698) );
  XOR2_X1 U16820 ( .A(n13345), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13343)
         );
  NAND2_X1 U16821 ( .A1(n13516), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n13342) );
  INV_X1 U16822 ( .A(n13338), .ZN(n13339) );
  AOI21_X1 U16823 ( .B1(n13340), .B2(n13749), .A(n13339), .ZN(n18916) );
  NAND2_X1 U16824 ( .A1(n18916), .A2(n18965), .ZN(n13341) );
  OAI211_X1 U16825 ( .C1(n13343), .C2(n18951), .A(n13342), .B(n13341), .ZN(
        P2_U2882) );
  INV_X1 U16826 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13344) );
  NOR2_X1 U16827 ( .A1(n13345), .A2(n13344), .ZN(n13346) );
  OAI211_X1 U16828 ( .C1(n13346), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n18966), .B(n13423), .ZN(n13352) );
  AND2_X1 U16829 ( .A1(n13338), .A2(n13347), .ZN(n13349) );
  OR2_X1 U16830 ( .A1(n13349), .A2(n13348), .ZN(n18899) );
  INV_X1 U16831 ( .A(n18899), .ZN(n13350) );
  NAND2_X1 U16832 ( .A1(n13350), .A2(n18965), .ZN(n13351) );
  OAI211_X1 U16833 ( .C1(n18965), .C2(n10769), .A(n13352), .B(n13351), .ZN(
        P2_U2881) );
  INV_X1 U16834 ( .A(n15130), .ZN(n13353) );
  INV_X1 U16835 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19017) );
  OAI222_X1 U16836 ( .A1(n13632), .A2(n13353), .B1(n15432), .B2(n19004), .C1(
        n19017), .C2(n15168), .ZN(P2_U2908) );
  INV_X1 U16837 ( .A(n13354), .ZN(n13355) );
  OAI21_X1 U16838 ( .B1(n15795), .B2(n13660), .A(n13355), .ZN(n13357) );
  NOR2_X1 U16839 ( .A1(n13665), .A2(n19975), .ZN(n13356) );
  AOI211_X1 U16840 ( .C1(n15791), .C2(n13660), .A(n13357), .B(n13356), .ZN(
        n13358) );
  OAI21_X1 U16841 ( .B1(n13359), .B2(n19757), .A(n13358), .ZN(P1_U2998) );
  INV_X2 U16842 ( .A(n13441), .ZN(n19923) );
  AOI22_X1 U16843 ( .A1(n19923), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n13470), .ZN(n13364) );
  NAND2_X1 U16844 ( .A1(n19974), .A2(DATAI_3_), .ZN(n13362) );
  NAND2_X1 U16845 ( .A1(n19976), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13361) );
  AND2_X1 U16846 ( .A1(n13362), .A2(n13361), .ZN(n20000) );
  INV_X1 U16847 ( .A(n20000), .ZN(n13363) );
  NAND2_X1 U16848 ( .A1(n19915), .A2(n13363), .ZN(n13442) );
  NAND2_X1 U16849 ( .A1(n13364), .A2(n13442), .ZN(P1_U2955) );
  AOI22_X1 U16850 ( .A1(n19923), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n13470), .ZN(n13368) );
  NAND2_X1 U16851 ( .A1(n19974), .A2(DATAI_7_), .ZN(n13366) );
  NAND2_X1 U16852 ( .A1(n19976), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13365) );
  AND2_X1 U16853 ( .A1(n13366), .A2(n13365), .ZN(n20017) );
  INV_X1 U16854 ( .A(n20017), .ZN(n13367) );
  NAND2_X1 U16855 ( .A1(n19915), .A2(n13367), .ZN(n13464) );
  NAND2_X1 U16856 ( .A1(n13368), .A2(n13464), .ZN(P1_U2959) );
  AOI22_X1 U16857 ( .A1(n19923), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n13470), .ZN(n13372) );
  INV_X1 U16858 ( .A(DATAI_13_), .ZN(n13370) );
  MUX2_X1 U16859 ( .A(n13370), .B(n13369), .S(n19976), .Z(n14745) );
  INV_X1 U16860 ( .A(n14745), .ZN(n13371) );
  NAND2_X1 U16861 ( .A1(n19915), .A2(n13371), .ZN(n13462) );
  NAND2_X1 U16862 ( .A1(n13372), .A2(n13462), .ZN(P1_U2965) );
  AOI22_X1 U16863 ( .A1(n19923), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n13470), .ZN(n13376) );
  NAND2_X1 U16864 ( .A1(n19974), .A2(DATAI_5_), .ZN(n13374) );
  NAND2_X1 U16865 ( .A1(n19976), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13373) );
  AND2_X1 U16866 ( .A1(n13374), .A2(n13373), .ZN(n20007) );
  INV_X1 U16867 ( .A(n20007), .ZN(n13375) );
  NAND2_X1 U16868 ( .A1(n19915), .A2(n13375), .ZN(n13460) );
  NAND2_X1 U16869 ( .A1(n13376), .A2(n13460), .ZN(P1_U2957) );
  AOI22_X1 U16870 ( .A1(n19923), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n13470), .ZN(n13379) );
  NAND2_X1 U16871 ( .A1(n19974), .A2(DATAI_4_), .ZN(n13378) );
  NAND2_X1 U16872 ( .A1(n19976), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13377) );
  AND2_X1 U16873 ( .A1(n13378), .A2(n13377), .ZN(n20003) );
  INV_X1 U16874 ( .A(n20003), .ZN(n15718) );
  NAND2_X1 U16875 ( .A1(n19915), .A2(n15718), .ZN(n13468) );
  NAND2_X1 U16876 ( .A1(n13379), .A2(n13468), .ZN(P1_U2956) );
  AOI22_X1 U16877 ( .A1(n19923), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n13470), .ZN(n13383) );
  NAND2_X1 U16878 ( .A1(n19974), .A2(DATAI_6_), .ZN(n13381) );
  NAND2_X1 U16879 ( .A1(n19976), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13380) );
  AND2_X1 U16880 ( .A1(n13381), .A2(n13380), .ZN(n20010) );
  INV_X1 U16881 ( .A(n20010), .ZN(n13382) );
  NAND2_X1 U16882 ( .A1(n19915), .A2(n13382), .ZN(n13450) );
  NAND2_X1 U16883 ( .A1(n13383), .A2(n13450), .ZN(P1_U2958) );
  XOR2_X1 U16884 ( .A(n13384), .B(n13385), .Z(n13417) );
  NOR2_X1 U16885 ( .A1(n19933), .A2(n11656), .ZN(n13386) );
  AOI21_X1 U16886 ( .B1(n13386), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n19944), .ZN(n13395) );
  AOI21_X1 U16887 ( .B1(n13389), .B2(n13388), .A(n13387), .ZN(n13669) );
  NAND2_X1 U16888 ( .A1(n13669), .A2(n19964), .ZN(n13394) );
  INV_X1 U16889 ( .A(n15902), .ZN(n14964) );
  OAI21_X1 U16890 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14964), .A(
        n15881), .ZN(n13392) );
  AND2_X1 U16891 ( .A1(n19953), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n13391) );
  NOR3_X1 U16892 ( .A1(n11656), .A2(n15900), .A3(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13390) );
  AOI211_X1 U16893 ( .C1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n13392), .A(
        n13391), .B(n13390), .ZN(n13393) );
  OAI211_X1 U16894 ( .C1(n13395), .C2(n15865), .A(n13394), .B(n13393), .ZN(
        n13396) );
  AOI21_X1 U16895 ( .B1(n13417), .B2(n19965), .A(n13396), .ZN(n13397) );
  INV_X1 U16896 ( .A(n13397), .ZN(P1_U3029) );
  INV_X1 U16897 ( .A(n13398), .ZN(n13399) );
  AOI21_X1 U16898 ( .B1(n13400), .B2(n19933), .A(n13399), .ZN(n19963) );
  INV_X1 U16899 ( .A(n19963), .ZN(n13405) );
  INV_X1 U16900 ( .A(n13401), .ZN(n13404) );
  OAI21_X1 U16901 ( .B1(n13404), .B2(n13403), .A(n13402), .ZN(n19941) );
  OAI222_X1 U16902 ( .A1(n13405), .A2(n14684), .B1(n11660), .B2(n14682), .C1(
        n19941), .C2(n14672), .ZN(P1_U2872) );
  XOR2_X1 U16903 ( .A(n13423), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13411)
         );
  OR2_X1 U16904 ( .A1(n13348), .A2(n13407), .ZN(n13408) );
  AND2_X1 U16905 ( .A1(n13406), .A2(n13408), .ZN(n18881) );
  INV_X1 U16906 ( .A(n18881), .ZN(n14035) );
  MUX2_X1 U16907 ( .A(n14035), .B(n13409), .S(n13516), .Z(n13410) );
  OAI21_X1 U16908 ( .B1(n13411), .B2(n18951), .A(n13410), .ZN(P2_U2880) );
  INV_X1 U16909 ( .A(n13412), .ZN(n13413) );
  AOI21_X1 U16910 ( .B1(n13415), .B2(n13414), .A(n13413), .ZN(n13420) );
  INV_X1 U16911 ( .A(n13420), .ZN(n13677) );
  AOI22_X1 U16912 ( .A1(n13669), .A2(n14670), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n14669), .ZN(n13416) );
  OAI21_X1 U16913 ( .B1(n13677), .B2(n14672), .A(n13416), .ZN(P1_U2870) );
  INV_X1 U16914 ( .A(n13417), .ZN(n13422) );
  AOI22_X1 U16915 ( .A1(n19936), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n19953), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13418) );
  OAI21_X1 U16916 ( .B1(n15787), .B2(n13667), .A(n13418), .ZN(n13419) );
  AOI21_X1 U16917 ( .B1(n13420), .B2(n12940), .A(n13419), .ZN(n13421) );
  OAI21_X1 U16918 ( .B1(n13422), .B2(n19757), .A(n13421), .ZN(P1_U2997) );
  XNOR2_X1 U16919 ( .A(n13520), .B(n13518), .ZN(n13428) );
  NAND2_X1 U16920 ( .A1(n13406), .A2(n13424), .ZN(n13425) );
  NAND2_X1 U16921 ( .A1(n13513), .A2(n13425), .ZN(n16126) );
  MUX2_X1 U16922 ( .A(n16126), .B(n13426), .S(n13516), .Z(n13427) );
  OAI21_X1 U16923 ( .B1(n13428), .B2(n18951), .A(n13427), .ZN(P2_U2879) );
  OR2_X1 U16924 ( .A1(n13431), .A2(n13430), .ZN(n13432) );
  NAND2_X1 U16925 ( .A1(n13429), .A2(n13432), .ZN(n19864) );
  INV_X1 U16926 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n19855) );
  OR2_X1 U16927 ( .A1(n13387), .A2(n13433), .ZN(n13434) );
  AND2_X1 U16928 ( .A1(n13580), .A2(n13434), .ZN(n19954) );
  INV_X1 U16929 ( .A(n19954), .ZN(n13435) );
  OAI222_X1 U16930 ( .A1(n19864), .A2(n14672), .B1(n14682), .B2(n19855), .C1(
        n13435), .C2(n14684), .ZN(P1_U2869) );
  NOR2_X1 U16931 ( .A1(n13438), .A2(n13436), .ZN(n13437) );
  NAND2_X1 U16932 ( .A1(n15728), .A2(n13438), .ZN(n15716) );
  NAND2_X1 U16933 ( .A1(n15716), .A2(n13439), .ZN(n15725) );
  OAI222_X1 U16934 ( .A1(n19864), .A2(n14740), .B1(n20000), .B2(n14744), .C1(
        n13440), .C2(n15728), .ZN(P1_U2901) );
  AOI22_X1 U16935 ( .A1(n19923), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n13470), .ZN(n13443) );
  NAND2_X1 U16936 ( .A1(n13443), .A2(n13442), .ZN(P1_U2940) );
  AOI22_X1 U16937 ( .A1(n19923), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n13470), .ZN(n13447) );
  NAND2_X1 U16938 ( .A1(n19974), .A2(DATAI_2_), .ZN(n13445) );
  NAND2_X1 U16939 ( .A1(n19976), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13444) );
  AND2_X1 U16940 ( .A1(n13445), .A2(n13444), .ZN(n19997) );
  INV_X1 U16941 ( .A(n19997), .ZN(n13446) );
  NAND2_X1 U16942 ( .A1(n19915), .A2(n13446), .ZN(n13448) );
  NAND2_X1 U16943 ( .A1(n13447), .A2(n13448), .ZN(P1_U2939) );
  AOI22_X1 U16944 ( .A1(n19923), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n13470), .ZN(n13449) );
  NAND2_X1 U16945 ( .A1(n13449), .A2(n13448), .ZN(P1_U2954) );
  AOI22_X1 U16946 ( .A1(n19923), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n13470), .ZN(n13451) );
  NAND2_X1 U16947 ( .A1(n13451), .A2(n13450), .ZN(P1_U2943) );
  AOI22_X1 U16948 ( .A1(n19923), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n13470), .ZN(n13455) );
  NAND2_X1 U16949 ( .A1(n19974), .A2(DATAI_0_), .ZN(n13453) );
  NAND2_X1 U16950 ( .A1(n19976), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13452) );
  AND2_X1 U16951 ( .A1(n13453), .A2(n13452), .ZN(n19985) );
  INV_X1 U16952 ( .A(n19985), .ZN(n13454) );
  NAND2_X1 U16953 ( .A1(n19915), .A2(n13454), .ZN(n13471) );
  NAND2_X1 U16954 ( .A1(n13455), .A2(n13471), .ZN(P1_U2952) );
  AOI22_X1 U16955 ( .A1(n19923), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n13470), .ZN(n13459) );
  NAND2_X1 U16956 ( .A1(n19974), .A2(DATAI_1_), .ZN(n13457) );
  NAND2_X1 U16957 ( .A1(n19976), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13456) );
  AND2_X1 U16958 ( .A1(n13457), .A2(n13456), .ZN(n19993) );
  INV_X1 U16959 ( .A(n19993), .ZN(n13458) );
  NAND2_X1 U16960 ( .A1(n19915), .A2(n13458), .ZN(n13466) );
  NAND2_X1 U16961 ( .A1(n13459), .A2(n13466), .ZN(P1_U2953) );
  AOI22_X1 U16962 ( .A1(n19923), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n13470), .ZN(n13461) );
  NAND2_X1 U16963 ( .A1(n13461), .A2(n13460), .ZN(P1_U2942) );
  AOI22_X1 U16964 ( .A1(n19923), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n13470), .ZN(n13463) );
  NAND2_X1 U16965 ( .A1(n13463), .A2(n13462), .ZN(P1_U2950) );
  AOI22_X1 U16966 ( .A1(n19923), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n13470), .ZN(n13465) );
  NAND2_X1 U16967 ( .A1(n13465), .A2(n13464), .ZN(P1_U2944) );
  AOI22_X1 U16968 ( .A1(n19923), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n13470), .ZN(n13467) );
  NAND2_X1 U16969 ( .A1(n13467), .A2(n13466), .ZN(P1_U2938) );
  AOI22_X1 U16970 ( .A1(n19923), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n13470), .ZN(n13469) );
  NAND2_X1 U16971 ( .A1(n13469), .A2(n13468), .ZN(P1_U2941) );
  AOI22_X1 U16972 ( .A1(n19923), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n13470), .ZN(n13472) );
  NAND2_X1 U16973 ( .A1(n13472), .A2(n13471), .ZN(P1_U2937) );
  INV_X1 U16974 ( .A(n13473), .ZN(n13474) );
  NOR2_X1 U16975 ( .A1(n13475), .A2(n13474), .ZN(n13477) );
  NAND2_X1 U16976 ( .A1(n15488), .A2(n15058), .ZN(n13589) );
  OAI21_X1 U16977 ( .B1(n15488), .B2(n15058), .A(n13589), .ZN(n13476) );
  NOR2_X1 U16978 ( .A1(n13477), .A2(n13476), .ZN(n13591) );
  AOI21_X1 U16979 ( .B1(n13477), .B2(n13476), .A(n13591), .ZN(n13481) );
  AOI22_X1 U16980 ( .A1(n18997), .A2(n13478), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n18995), .ZN(n13480) );
  NAND2_X1 U16981 ( .A1(n19690), .A2(n18980), .ZN(n13479) );
  OAI211_X1 U16982 ( .C1(n13481), .C2(n18998), .A(n13480), .B(n13479), .ZN(
        P2_U2917) );
  INV_X1 U16983 ( .A(n13483), .ZN(n13484) );
  XNOR2_X1 U16984 ( .A(n13482), .B(n13484), .ZN(n19955) );
  NAND2_X1 U16985 ( .A1(n19955), .A2(n19938), .ZN(n13489) );
  INV_X1 U16986 ( .A(n13485), .ZN(n19866) );
  INV_X1 U16987 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13486) );
  OAI22_X1 U16988 ( .A1(n15795), .A2(n20835), .B1(n15908), .B2(n13486), .ZN(
        n13487) );
  AOI21_X1 U16989 ( .B1(n19866), .B2(n15791), .A(n13487), .ZN(n13488) );
  OAI211_X1 U16990 ( .C1(n19975), .C2(n19864), .A(n13489), .B(n13488), .ZN(
        P1_U2996) );
  NOR2_X1 U16991 ( .A1(n19727), .A2(n13490), .ZN(n16219) );
  NOR2_X1 U16992 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19546), .ZN(n16220) );
  INV_X1 U16993 ( .A(n13491), .ZN(n16194) );
  NAND2_X1 U16994 ( .A1(n16194), .A2(n13492), .ZN(n13494) );
  OAI21_X1 U16995 ( .B1(n13495), .B2(n13494), .A(n13493), .ZN(n13496) );
  NOR3_X1 U16996 ( .A1(n13498), .A2(n13497), .A3(n13496), .ZN(n16170) );
  NOR2_X1 U16997 ( .A1(n16170), .A2(n18755), .ZN(n13499) );
  AOI211_X2 U16998 ( .C1(P2_FLUSH_REG_SCAN_IN), .C2(n16219), .A(n16220), .B(
        n13499), .ZN(n15524) );
  NAND2_X1 U16999 ( .A1(n16186), .A2(n16181), .ZN(n15471) );
  NOR2_X1 U17000 ( .A1(n13500), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15472) );
  INV_X1 U17001 ( .A(n15472), .ZN(n15479) );
  AOI22_X1 U17002 ( .A1(n15471), .A2(n15479), .B1(n10575), .B2(n9728), .ZN(
        n13507) );
  INV_X1 U17003 ( .A(n13501), .ZN(n13502) );
  NAND2_X1 U17004 ( .A1(n13502), .A2(n10846), .ZN(n13504) );
  AND2_X1 U17005 ( .A1(n13504), .A2(n13503), .ZN(n15480) );
  INV_X1 U17006 ( .A(n15475), .ZN(n15450) );
  NOR2_X1 U17007 ( .A1(n15450), .A2(n10575), .ZN(n13505) );
  NOR3_X1 U17008 ( .A1(n15480), .A2(n15472), .A3(n13505), .ZN(n13506) );
  MUX2_X1 U17009 ( .A(n13507), .B(n13506), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13509) );
  INV_X1 U17010 ( .A(n14294), .ZN(n13508) );
  OAI211_X1 U17011 ( .C1(n16148), .C2(n15461), .A(n13509), .B(n13508), .ZN(
        n16169) );
  AOI22_X1 U17012 ( .A1(n19681), .A2(n16214), .B1(n19596), .B2(n16169), .ZN(
        n13511) );
  NAND2_X1 U17013 ( .A1(n15524), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13510) );
  OAI21_X1 U17014 ( .B1(n15524), .B2(n13511), .A(n13510), .ZN(P2_U3596) );
  AND2_X1 U17015 ( .A1(n13513), .A2(n13512), .ZN(n13515) );
  OR2_X1 U17016 ( .A1(n13515), .A2(n13514), .ZN(n15442) );
  AND2_X1 U17017 ( .A1(n13518), .A2(n13517), .ZN(n13519) );
  INV_X1 U17018 ( .A(n13536), .ZN(n13532) );
  INV_X1 U17019 ( .A(n13520), .ZN(n13523) );
  OAI21_X1 U17020 ( .B1(n13523), .B2(n13522), .A(n13521), .ZN(n13524) );
  NAND3_X1 U17021 ( .A1(n13532), .A2(n18966), .A3(n13524), .ZN(n13526) );
  NAND2_X1 U17022 ( .A1(n13516), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n13525) );
  OAI211_X1 U17023 ( .C1(n15442), .C2(n13516), .A(n13526), .B(n13525), .ZN(
        P2_U2878) );
  AOI21_X1 U17024 ( .B1(n13529), .B2(n13429), .A(n13528), .ZN(n19848) );
  INV_X1 U17025 ( .A(n19848), .ZN(n13574) );
  XOR2_X1 U17026 ( .A(n13579), .B(n13580), .Z(n19946) );
  AOI22_X1 U17027 ( .A1(n19946), .A2(n14670), .B1(P1_EBX_REG_4__SCAN_IN), .B2(
        n14669), .ZN(n13530) );
  OAI21_X1 U17028 ( .B1(n13574), .B2(n14672), .A(n13530), .ZN(P1_U2868) );
  OAI21_X1 U17029 ( .B1(n13532), .B2(n18960), .A(n13531), .ZN(n13537) );
  AND2_X1 U17030 ( .A1(n13534), .A2(n13533), .ZN(n13535) );
  NAND3_X1 U17031 ( .A1(n13537), .A2(n18966), .A3(n13611), .ZN(n13540) );
  INV_X1 U17032 ( .A(n13538), .ZN(n16044) );
  NAND2_X1 U17033 ( .A1(n16044), .A2(n18965), .ZN(n13539) );
  OAI211_X1 U17034 ( .C1(n18965), .C2(n13541), .A(n13540), .B(n13539), .ZN(
        P2_U2876) );
  INV_X1 U17035 ( .A(n15118), .ZN(n13545) );
  OAI21_X1 U17036 ( .B1(n13544), .B2(n13542), .A(n13543), .ZN(n18864) );
  INV_X1 U17037 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n20918) );
  OAI222_X1 U17038 ( .A1(n13632), .A2(n13545), .B1(n18864), .B2(n19004), .C1(
        n20918), .C2(n15168), .ZN(P2_U2906) );
  OAI222_X1 U17039 ( .A1(n14747), .A2(n13677), .B1(n19997), .B2(n14744), .C1(
        n15728), .C2(n11917), .ZN(P1_U2902) );
  OAI222_X1 U17040 ( .A1(n14747), .A2(n13665), .B1(n19993), .B2(n14744), .C1(
        n15728), .C2(n11923), .ZN(P1_U2903) );
  INV_X1 U17041 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n13546) );
  OAI222_X1 U17042 ( .A1(n14747), .A2(n19941), .B1(n19985), .B2(n14744), .C1(
        n15728), .C2(n13546), .ZN(P1_U2904) );
  AOI21_X1 U17043 ( .B1(n14984), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11150), .ZN(n13547) );
  NOR2_X1 U17044 ( .A1(n13548), .A2(n13547), .ZN(n20727) );
  NAND2_X1 U17045 ( .A1(n20736), .A2(n13549), .ZN(n13557) );
  MUX2_X1 U17046 ( .A(n11158), .B(n20732), .S(n14984), .Z(n13551) );
  NOR2_X1 U17047 ( .A1(n13551), .A2(n13550), .ZN(n13554) );
  XNOR2_X1 U17048 ( .A(n13552), .B(n11150), .ZN(n13553) );
  AOI22_X1 U17049 ( .A1(n13555), .A2(n13554), .B1(n15548), .B2(n13553), .ZN(
        n13556) );
  OAI211_X1 U17050 ( .C1(n20727), .C2(n13558), .A(n13557), .B(n13556), .ZN(
        n20725) );
  MUX2_X1 U17051 ( .A(n20725), .B(n20732), .S(n13562), .Z(n15557) );
  NOR2_X1 U17052 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20957), .ZN(n13563) );
  AOI22_X1 U17053 ( .A1(n15557), .A2(n20957), .B1(n20732), .B2(n13563), .ZN(
        n13561) );
  INV_X1 U17054 ( .A(n13562), .ZN(n15549) );
  MUX2_X1 U17055 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13559), .S(
        n15549), .Z(n15555) );
  AOI22_X1 U17056 ( .A1(n13563), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15555), .B2(n20957), .ZN(n13560) );
  NOR2_X1 U17057 ( .A1(n13561), .A2(n13560), .ZN(n15567) );
  INV_X1 U17058 ( .A(n15567), .ZN(n13566) );
  OAI21_X1 U17059 ( .B1(n19841), .B2(n12896), .A(n15549), .ZN(n13565) );
  AOI21_X1 U17060 ( .B1(n13562), .B2(n13318), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n13564) );
  AOI22_X1 U17061 ( .A1(n13565), .A2(n13564), .B1(n13563), .B2(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15565) );
  OAI21_X1 U17062 ( .B1(n13566), .B2(n14985), .A(n15565), .ZN(n13568) );
  NOR2_X1 U17063 ( .A1(n13568), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n13567) );
  NOR2_X1 U17064 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20764) );
  INV_X1 U17065 ( .A(n13568), .ZN(n13569) );
  NAND2_X1 U17066 ( .A1(n13569), .A2(n15941), .ZN(n15577) );
  INV_X1 U17067 ( .A(n15577), .ZN(n13572) );
  NAND2_X1 U17068 ( .A1(n20446), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20737) );
  INV_X1 U17069 ( .A(n20737), .ZN(n14975) );
  OAI22_X1 U17070 ( .A1(n20438), .A2(n20743), .B1(n13570), .B2(n14975), .ZN(
        n13571) );
  OAI21_X1 U17071 ( .B1(n13572), .B2(n13571), .A(n20747), .ZN(n13573) );
  OAI21_X1 U17072 ( .B1(n20747), .B2(n20471), .A(n13573), .ZN(P1_U3478) );
  INV_X1 U17073 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19891) );
  OAI222_X1 U17074 ( .A1(n14747), .A2(n13574), .B1(n14744), .B2(n20003), .C1(
        n19891), .C2(n15728), .ZN(P1_U2900) );
  OR2_X1 U17075 ( .A1(n13528), .A2(n13576), .ZN(n13577) );
  AND2_X1 U17076 ( .A1(n13575), .A2(n13577), .ZN(n19832) );
  INV_X1 U17077 ( .A(n19832), .ZN(n13584) );
  OAI21_X1 U17078 ( .B1(n13580), .B2(n13579), .A(n13578), .ZN(n13581) );
  AND2_X1 U17079 ( .A1(n13581), .A2(n13711), .ZN(n19827) );
  AOI22_X1 U17080 ( .A1(n19827), .A2(n14670), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14669), .ZN(n13582) );
  OAI21_X1 U17081 ( .B1(n13584), .B2(n14672), .A(n13582), .ZN(P1_U2867) );
  INV_X1 U17082 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13583) );
  OAI222_X1 U17083 ( .A1(n13584), .A2(n14747), .B1(n20007), .B2(n14744), .C1(
        n13583), .C2(n15728), .ZN(P1_U2899) );
  OR2_X1 U17084 ( .A1(n13586), .A2(n13585), .ZN(n13588) );
  NAND2_X1 U17085 ( .A1(n13588), .A2(n13587), .ZN(n16151) );
  XNOR2_X1 U17086 ( .A(n19479), .B(n16151), .ZN(n13593) );
  INV_X1 U17087 ( .A(n13589), .ZN(n13590) );
  NOR2_X1 U17088 ( .A1(n13591), .A2(n13590), .ZN(n13592) );
  NOR2_X1 U17089 ( .A1(n13592), .A2(n13593), .ZN(n13692) );
  AOI21_X1 U17090 ( .B1(n13593), .B2(n13592), .A(n13692), .ZN(n13597) );
  AOI22_X1 U17091 ( .A1(n18997), .A2(n13594), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n18995), .ZN(n13596) );
  INV_X1 U17092 ( .A(n16151), .ZN(n19682) );
  NAND2_X1 U17093 ( .A1(n19682), .A2(n18980), .ZN(n13595) );
  OAI211_X1 U17094 ( .C1(n13597), .C2(n18998), .A(n13596), .B(n13595), .ZN(
        P2_U2916) );
  XOR2_X1 U17095 ( .A(n13598), .B(n13599), .Z(n19950) );
  INV_X1 U17096 ( .A(n19950), .ZN(n13603) );
  NAND2_X1 U17097 ( .A1(n19936), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13600) );
  NAND2_X1 U17098 ( .A1(n19939), .A2(P1_REIP_REG_4__SCAN_IN), .ZN(n19947) );
  OAI211_X1 U17099 ( .C1(n15787), .C2(n19852), .A(n13600), .B(n19947), .ZN(
        n13601) );
  AOI21_X1 U17100 ( .B1(n19848), .B2(n12940), .A(n13601), .ZN(n13602) );
  OAI21_X1 U17101 ( .B1(n13603), .B2(n19757), .A(n13602), .ZN(P1_U2995) );
  INV_X1 U17102 ( .A(n13604), .ZN(n13707) );
  NAND2_X1 U17103 ( .A1(n13575), .A2(n13605), .ZN(n13606) );
  AND2_X1 U17104 ( .A1(n13707), .A2(n13606), .ZN(n19822) );
  INV_X1 U17105 ( .A(n19822), .ZN(n13608) );
  XNOR2_X1 U17106 ( .A(n13711), .B(n13713), .ZN(n19814) );
  AOI22_X1 U17107 ( .A1(n19814), .A2(n14670), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14669), .ZN(n13607) );
  OAI21_X1 U17108 ( .B1(n13608), .B2(n14672), .A(n13607), .ZN(P1_U2866) );
  OAI222_X1 U17109 ( .A1(n14747), .A2(n13608), .B1(n20010), .B2(n14744), .C1(
        n15728), .C2(n11962), .ZN(P1_U2898) );
  INV_X1 U17110 ( .A(n15384), .ZN(n13609) );
  AOI21_X1 U17111 ( .B1(n13610), .B2(n13802), .A(n13609), .ZN(n18860) );
  NAND2_X1 U17112 ( .A1(n18860), .A2(n18965), .ZN(n13617) );
  OAI21_X1 U17113 ( .B1(n13611), .B2(n13613), .A(n13612), .ZN(n13615) );
  NAND3_X1 U17114 ( .A1(n13615), .A2(n18966), .A3(n13731), .ZN(n13616) );
  OAI211_X1 U17115 ( .C1(n18965), .C2(n10799), .A(n13617), .B(n13616), .ZN(
        P2_U2874) );
  NAND2_X1 U17116 ( .A1(n18870), .A2(n13618), .ZN(n13619) );
  XNOR2_X1 U17117 ( .A(n16089), .B(n13619), .ZN(n13620) );
  NAND2_X1 U17118 ( .A1(n13620), .A2(n18917), .ZN(n13627) );
  OAI22_X1 U17119 ( .A1(n10598), .A2(n18906), .B1(n10914), .B2(n18929), .ZN(
        n13621) );
  AOI21_X1 U17120 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18939), .A(
        n13621), .ZN(n13622) );
  OAI21_X1 U17121 ( .B1(n18927), .B2(n13623), .A(n13622), .ZN(n13625) );
  NOR2_X1 U17122 ( .A1(n16151), .A2(n18921), .ZN(n13624) );
  AOI211_X1 U17123 ( .C1(n18933), .C2(n10278), .A(n13625), .B(n13624), .ZN(
        n13626) );
  OAI211_X1 U17124 ( .C1(n19479), .C2(n15063), .A(n13627), .B(n13626), .ZN(
        P2_U2852) );
  OAI21_X1 U17125 ( .B1(n13628), .B2(n13630), .A(n13629), .ZN(n18842) );
  OAI222_X1 U17126 ( .A1(n13632), .A2(n13631), .B1(n18842), .B2(n19004), .C1(
        n13062), .C2(n15168), .ZN(P2_U2904) );
  INV_X1 U17127 ( .A(n20764), .ZN(n15943) );
  NOR3_X1 U17128 ( .A1(n15945), .A2(n20446), .A3(n15943), .ZN(n15576) );
  NOR3_X1 U17129 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20957), .A3(n13633), 
        .ZN(n13634) );
  OR2_X1 U17130 ( .A1(n19953), .A2(n13634), .ZN(n13635) );
  OR2_X1 U17131 ( .A1(n13638), .A2(n13642), .ZN(n13639) );
  NAND2_X1 U17132 ( .A1(n15629), .A2(n13639), .ZN(n19867) );
  INV_X1 U17133 ( .A(n19867), .ZN(n13676) );
  NOR2_X1 U17134 ( .A1(n13640), .A2(n13642), .ZN(n13674) );
  AND2_X1 U17135 ( .A1(n20760), .A2(n20516), .ZN(n15570) );
  AND2_X1 U17136 ( .A1(n13641), .A2(n15570), .ZN(n13647) );
  NAND2_X1 U17137 ( .A1(n19773), .A2(n19845), .ZN(n19816) );
  INV_X1 U17138 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20754) );
  NOR2_X1 U17139 ( .A1(n13644), .A2(n20957), .ZN(n13645) );
  OAI21_X1 U17140 ( .B1(n19858), .B2(n19865), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13653) );
  NAND2_X1 U17141 ( .A1(n19992), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13648) );
  NOR2_X1 U17142 ( .A1(n13648), .A2(n15570), .ZN(n13646) );
  INV_X1 U17143 ( .A(n13647), .ZN(n13651) );
  AND2_X1 U17144 ( .A1(n13649), .A2(n13648), .ZN(n13650) );
  AND2_X2 U17145 ( .A1(n13651), .A2(n13650), .ZN(n19837) );
  AOI22_X1 U17146 ( .A1(n19963), .A2(n19863), .B1(P1_EBX_REG_0__SCAN_IN), .B2(
        n19837), .ZN(n13652) );
  OAI211_X1 U17147 ( .C1(n15641), .C2(n20754), .A(n13653), .B(n13652), .ZN(
        n13654) );
  AOI21_X1 U17148 ( .B1(n20089), .B2(n13674), .A(n13654), .ZN(n13655) );
  OAI21_X1 U17149 ( .B1(n19941), .B2(n13676), .A(n13655), .ZN(P1_U2840) );
  INV_X1 U17150 ( .A(n13674), .ZN(n19860) );
  AOI22_X1 U17151 ( .A1(n19837), .A2(P1_EBX_REG_1__SCAN_IN), .B1(n19853), .B2(
        n20748), .ZN(n13658) );
  NAND2_X1 U17152 ( .A1(n13656), .A2(n19863), .ZN(n13657) );
  OAI211_X1 U17153 ( .C1(n19773), .C2(n20748), .A(n13658), .B(n13657), .ZN(
        n13659) );
  AOI21_X1 U17154 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19858), .A(
        n13659), .ZN(n13662) );
  NAND2_X1 U17155 ( .A1(n19865), .A2(n13660), .ZN(n13661) );
  OAI211_X1 U17156 ( .C1(n20508), .C2(n19860), .A(n13662), .B(n13661), .ZN(
        n13663) );
  INV_X1 U17157 ( .A(n13663), .ZN(n13664) );
  OAI21_X1 U17158 ( .B1(n13665), .B2(n13676), .A(n13664), .ZN(P1_U2839) );
  INV_X1 U17159 ( .A(n13262), .ZN(n19982) );
  AOI21_X1 U17160 ( .B1(n19853), .B2(P1_REIP_REG_1__SCAN_IN), .A(
        P1_REIP_REG_2__SCAN_IN), .ZN(n13672) );
  NAND2_X1 U17161 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n13666) );
  OAI21_X1 U17162 ( .B1(n19803), .B2(n13666), .A(n19816), .ZN(n19871) );
  INV_X1 U17163 ( .A(n13667), .ZN(n13668) );
  AOI22_X1 U17164 ( .A1(n13669), .A2(n19863), .B1(n13668), .B2(n19865), .ZN(
        n13671) );
  AOI22_X1 U17165 ( .A1(n19858), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n19837), .B2(P1_EBX_REG_2__SCAN_IN), .ZN(n13670) );
  OAI211_X1 U17166 ( .C1(n13672), .C2(n19871), .A(n13671), .B(n13670), .ZN(
        n13673) );
  AOI21_X1 U17167 ( .B1(n19982), .B2(n13674), .A(n13673), .ZN(n13675) );
  OAI21_X1 U17168 ( .B1(n13677), .B2(n13676), .A(n13675), .ZN(P1_U2838) );
  NAND2_X1 U17169 ( .A1(n19689), .A2(n19696), .ZN(n19163) );
  INV_X1 U17170 ( .A(n19163), .ZN(n19164) );
  AND2_X1 U17171 ( .A1(n19407), .A2(n19164), .ZN(n19206) );
  AOI21_X1 U17172 ( .B1(n13678), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13681) );
  OR2_X1 U17173 ( .A1(n19708), .A2(n19163), .ZN(n13683) );
  NAND2_X1 U17174 ( .A1(n13682), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19680) );
  NOR2_X1 U17175 ( .A1(n19681), .A2(n19680), .ZN(n13684) );
  INV_X1 U17176 ( .A(n13684), .ZN(n13679) );
  NAND2_X1 U17177 ( .A1(n13683), .A2(n13679), .ZN(n13680) );
  OAI211_X1 U17178 ( .C1(n19206), .C2(n13681), .A(n13680), .B(n19545), .ZN(
        n19208) );
  INV_X1 U17179 ( .A(n19208), .ZN(n13691) );
  INV_X1 U17180 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13690) );
  INV_X1 U17181 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16276) );
  INV_X1 U17182 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18080) );
  OAI22_X2 U17183 ( .A1(n16276), .A2(n19123), .B1(n18080), .B2(n19121), .ZN(
        n19547) );
  NOR2_X2 U17184 ( .A1(n18973), .A2(n19447), .ZN(n19540) );
  INV_X1 U17185 ( .A(n19697), .ZN(n19685) );
  OR3_X1 U17186 ( .A1(n13684), .A2(n13683), .A3(n19685), .ZN(n13686) );
  OAI21_X1 U17187 ( .B1(n10432), .B2(n19206), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13685) );
  NAND2_X1 U17188 ( .A1(n13686), .A2(n13685), .ZN(n19207) );
  AOI22_X1 U17189 ( .A1(n19547), .A2(n19201), .B1(n19540), .B2(n19207), .ZN(
        n13689) );
  AOI22_X1 U17190 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19120), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19119), .ZN(n19550) );
  INV_X1 U17191 ( .A(n19550), .ZN(n19508) );
  NOR2_X2 U17192 ( .A1(n19125), .A2(n10528), .ZN(n19539) );
  AOI22_X1 U17193 ( .A1(n19508), .A2(n19245), .B1(n19206), .B2(n19539), .ZN(
        n13688) );
  OAI211_X1 U17194 ( .C1(n13691), .C2(n13690), .A(n13689), .B(n13688), .ZN(
        P2_U3072) );
  AOI21_X1 U17195 ( .B1(n19479), .B2(n16151), .A(n13692), .ZN(n13696) );
  NAND2_X1 U17196 ( .A1(n13693), .A2(n13587), .ZN(n13695) );
  NAND2_X1 U17197 ( .A1(n13695), .A2(n9925), .ZN(n13819) );
  INV_X1 U17198 ( .A(n13819), .ZN(n13751) );
  NOR2_X1 U17199 ( .A1(n13696), .A2(n13751), .ZN(n19000) );
  INV_X1 U17200 ( .A(n13698), .ZN(n13699) );
  NAND3_X1 U17201 ( .A1(n13697), .A2(n13700), .A3(n13699), .ZN(n13701) );
  NAND2_X1 U17202 ( .A1(n13345), .A2(n13701), .ZN(n18999) );
  XNOR2_X1 U17203 ( .A(n19000), .B(n18999), .ZN(n13704) );
  AOI22_X1 U17204 ( .A1(n18997), .A2(n15992), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n18995), .ZN(n13703) );
  NAND2_X1 U17205 ( .A1(n18980), .A2(n13751), .ZN(n13702) );
  OAI211_X1 U17206 ( .C1(n13704), .C2(n18998), .A(n13703), .B(n13702), .ZN(
        P2_U2915) );
  NAND2_X1 U17207 ( .A1(n13707), .A2(n13706), .ZN(n13708) );
  AND2_X1 U17208 ( .A1(n13705), .A2(n13708), .ZN(n19809) );
  INV_X1 U17209 ( .A(n19809), .ZN(n13710) );
  OAI222_X1 U17210 ( .A1(n13710), .A2(n14747), .B1(n20017), .B2(n14744), .C1(
        n13709), .C2(n15728), .ZN(P1_U2897) );
  INV_X1 U17211 ( .A(n14672), .ZN(n14660) );
  INV_X1 U17212 ( .A(n13711), .ZN(n13714) );
  AOI21_X1 U17213 ( .B1(n13714), .B2(n13713), .A(n13712), .ZN(n13715) );
  OR2_X1 U17214 ( .A1(n13715), .A2(n13838), .ZN(n15916) );
  OAI22_X1 U17215 ( .A1(n15916), .A2(n14684), .B1(n13716), .B2(n14682), .ZN(
        n13717) );
  AOI21_X1 U17216 ( .B1(n19809), .B2(n14660), .A(n13717), .ZN(n13718) );
  INV_X1 U17217 ( .A(n13718), .ZN(P1_U2865) );
  AND2_X1 U17218 ( .A1(n13725), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19541) );
  NAND2_X1 U17219 ( .A1(n19541), .A2(n19479), .ZN(n19686) );
  NAND2_X1 U17220 ( .A1(n19689), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19251) );
  INV_X1 U17221 ( .A(n19251), .ZN(n19283) );
  NAND2_X1 U17222 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19283), .ZN(
        n19276) );
  NAND2_X1 U17223 ( .A1(n19686), .A2(n19276), .ZN(n13721) );
  NAND2_X1 U17224 ( .A1(n19407), .A2(n19283), .ZN(n19330) );
  INV_X1 U17225 ( .A(n19330), .ZN(n19333) );
  OAI211_X1 U17226 ( .C1(n19333), .C2(n19546), .A(n19545), .B(n13723), .ZN(
        n13719) );
  INV_X1 U17227 ( .A(n13719), .ZN(n13720) );
  NAND2_X1 U17228 ( .A1(n13721), .A2(n13720), .ZN(n19324) );
  INV_X1 U17229 ( .A(n19324), .ZN(n19313) );
  INV_X1 U17230 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13730) );
  NOR2_X2 U17231 ( .A1(n13999), .A2(n19447), .ZN(n19557) );
  OAI21_X1 U17232 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19276), .A(n19732), 
        .ZN(n13722) );
  NOR2_X2 U17233 ( .A1(n19125), .A2(n13724), .ZN(n19556) );
  INV_X1 U17234 ( .A(n19556), .ZN(n13727) );
  AOI22_X1 U17235 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19120), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19119), .ZN(n19458) );
  INV_X1 U17236 ( .A(n19458), .ZN(n19558) );
  NAND2_X1 U17237 ( .A1(n13725), .A2(n19212), .ZN(n19327) );
  AOI22_X1 U17238 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19119), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19120), .ZN(n19561) );
  AOI22_X1 U17239 ( .A1(n19347), .A2(n19558), .B1(n19318), .B2(n19455), .ZN(
        n13726) );
  OAI21_X1 U17240 ( .B1(n13727), .B2(n19330), .A(n13726), .ZN(n13728) );
  AOI21_X1 U17241 ( .B1(n19557), .B2(n19323), .A(n13728), .ZN(n13729) );
  OAI21_X1 U17242 ( .B1(n19313), .B2(n13730), .A(n13729), .ZN(P2_U3106) );
  XNOR2_X1 U17243 ( .A(n9778), .B(n13868), .ZN(n13738) );
  OR2_X1 U17244 ( .A1(n13732), .A2(n13733), .ZN(n13735) );
  AND2_X1 U17245 ( .A1(n13735), .A2(n13734), .ZN(n18839) );
  NOR2_X1 U17246 ( .A1(n18965), .A2(n10810), .ZN(n13736) );
  AOI21_X1 U17247 ( .B1(n18839), .B2(n18965), .A(n13736), .ZN(n13737) );
  OAI21_X1 U17248 ( .B1(n13738), .B2(n18951), .A(n13737), .ZN(P2_U2872) );
  XOR2_X1 U17249 ( .A(n13739), .B(n13740), .Z(n19047) );
  INV_X1 U17250 ( .A(n19047), .ZN(n13756) );
  XNOR2_X1 U17251 ( .A(n13741), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13742) );
  XNOR2_X1 U17252 ( .A(n13743), .B(n13742), .ZN(n19045) );
  NAND2_X1 U17253 ( .A1(n13745), .A2(n13744), .ZN(n13747) );
  NAND2_X1 U17254 ( .A1(n13747), .A2(n13746), .ZN(n13748) );
  NAND2_X1 U17255 ( .A1(n13749), .A2(n13748), .ZN(n18969) );
  INV_X1 U17256 ( .A(n16156), .ZN(n13977) );
  AOI21_X1 U17257 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13977), .A(
        n13976), .ZN(n13947) );
  NAND2_X1 U17258 ( .A1(n13947), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13753) );
  INV_X1 U17259 ( .A(n16132), .ZN(n16155) );
  NAND2_X1 U17260 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16155), .ZN(
        n13934) );
  OAI22_X1 U17261 ( .A1(n11123), .A2(n10920), .B1(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13934), .ZN(n13750) );
  AOI21_X1 U17262 ( .B1(n19067), .B2(n13751), .A(n13750), .ZN(n13752) );
  OAI211_X1 U17263 ( .C1(n18969), .C2(n19072), .A(n13753), .B(n13752), .ZN(
        n13754) );
  AOI21_X1 U17264 ( .B1(n19045), .B2(n16153), .A(n13754), .ZN(n13755) );
  OAI21_X1 U17265 ( .B1(n13756), .B2(n16163), .A(n13755), .ZN(P2_U3042) );
  NOR2_X1 U17266 ( .A1(n19132), .A2(n19738), .ZN(n19136) );
  NAND2_X1 U17267 ( .A1(n19681), .A2(n19136), .ZN(n13757) );
  NOR2_X1 U17268 ( .A1(n19689), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19406) );
  NAND2_X1 U17269 ( .A1(n19406), .A2(n19708), .ZN(n13762) );
  NAND2_X1 U17270 ( .A1(n13757), .A2(n13762), .ZN(n13761) );
  OAI21_X1 U17271 ( .B1(n10433), .B2(n19732), .A(n19546), .ZN(n13759) );
  INV_X1 U17272 ( .A(n19406), .ZN(n19409) );
  NOR3_X2 U17273 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19715), .A3(
        n19409), .ZN(n19379) );
  INV_X1 U17274 ( .A(n19379), .ZN(n13758) );
  AOI21_X1 U17275 ( .B1(n13759), .B2(n13758), .A(n19447), .ZN(n13760) );
  NAND2_X1 U17276 ( .A1(n13761), .A2(n13760), .ZN(n19372) );
  INV_X1 U17277 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13768) );
  AOI22_X1 U17278 ( .A1(n19558), .A2(n19400), .B1(n19556), .B2(n19379), .ZN(
        n13767) );
  INV_X1 U17279 ( .A(n13762), .ZN(n13763) );
  NAND2_X1 U17280 ( .A1(n13763), .A2(n19697), .ZN(n13765) );
  OAI21_X1 U17281 ( .B1(n10433), .B2(n19379), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13764) );
  NAND2_X1 U17282 ( .A1(n13765), .A2(n13764), .ZN(n19371) );
  AOI22_X1 U17283 ( .A1(n19455), .A2(n19370), .B1(n19557), .B2(n19371), .ZN(
        n13766) );
  OAI211_X1 U17284 ( .C1(n19364), .C2(n13768), .A(n13767), .B(n13766), .ZN(
        P2_U3122) );
  AOI22_X1 U17285 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19120), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19119), .ZN(n19488) );
  AOI22_X1 U17286 ( .A1(n19552), .A2(n19400), .B1(n19379), .B2(n13769), .ZN(
        n13771) );
  AOI22_X1 U17287 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19120), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19119), .ZN(n19555) );
  NOR2_X2 U17288 ( .A1(n13959), .A2(n19447), .ZN(n19551) );
  AOI22_X1 U17289 ( .A1(n19512), .A2(n19370), .B1(n19551), .B2(n19371), .ZN(
        n13770) );
  OAI211_X1 U17290 ( .C1(n19364), .C2(n13772), .A(n13771), .B(n13770), .ZN(
        P2_U3121) );
  INV_X1 U17291 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13775) );
  AOI22_X1 U17292 ( .A1(n19547), .A2(n19370), .B1(n19540), .B2(n19371), .ZN(
        n13774) );
  AOI22_X1 U17293 ( .A1(n19508), .A2(n19400), .B1(n19539), .B2(n19379), .ZN(
        n13773) );
  OAI211_X1 U17294 ( .C1(n19364), .C2(n13775), .A(n13774), .B(n13773), .ZN(
        P2_U3120) );
  NOR2_X1 U17295 ( .A1(n18896), .A2(n13776), .ZN(n13777) );
  XNOR2_X1 U17296 ( .A(n13777), .B(n16059), .ZN(n13789) );
  NOR2_X1 U17297 ( .A1(n13514), .A2(n13778), .ZN(n13779) );
  OR2_X1 U17298 ( .A1(n12988), .A2(n13779), .ZN(n16117) );
  OAI22_X1 U17299 ( .A1(n13781), .A2(n18927), .B1(n18908), .B2(n13780), .ZN(
        n13782) );
  INV_X1 U17300 ( .A(n13782), .ZN(n13783) );
  OAI211_X1 U17301 ( .C1(n18964), .C2(n18906), .A(n13783), .B(n11123), .ZN(
        n13784) );
  AOI21_X1 U17302 ( .B1(P2_REIP_REG_10__SCAN_IN), .B2(n18912), .A(n13784), 
        .ZN(n13787) );
  AOI21_X1 U17303 ( .B1(n13785), .B2(n13239), .A(n12983), .ZN(n18991) );
  NAND2_X1 U17304 ( .A1(n18923), .A2(n18991), .ZN(n13786) );
  OAI211_X1 U17305 ( .C1(n16117), .C2(n18900), .A(n13787), .B(n13786), .ZN(
        n13788) );
  AOI21_X1 U17306 ( .B1(n13789), .B2(n18917), .A(n13788), .ZN(n13790) );
  INV_X1 U17307 ( .A(n13790), .ZN(P2_U2845) );
  NOR2_X1 U17308 ( .A1(n18896), .A2(n13791), .ZN(n13792) );
  XNOR2_X1 U17309 ( .A(n13792), .B(n16081), .ZN(n13793) );
  NAND2_X1 U17310 ( .A1(n13793), .A2(n18917), .ZN(n13799) );
  AOI22_X1 U17311 ( .A1(n18922), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18939), .ZN(n13794) );
  OAI21_X1 U17312 ( .B1(n18921), .B2(n16123), .A(n13794), .ZN(n13796) );
  OAI21_X1 U17313 ( .B1(n10939), .B2(n18929), .A(n11123), .ZN(n13795) );
  AOI211_X1 U17314 ( .C1(n18885), .C2(n13797), .A(n13796), .B(n13795), .ZN(
        n13798) );
  OAI211_X1 U17315 ( .C1(n16126), .C2(n18900), .A(n13799), .B(n13798), .ZN(
        P2_U2847) );
  NAND2_X1 U17316 ( .A1(n12989), .A2(n13800), .ZN(n13801) );
  NAND2_X1 U17317 ( .A1(n13802), .A2(n13801), .ZN(n18959) );
  NOR2_X1 U17318 ( .A1(n18896), .A2(n13803), .ZN(n13804) );
  XNOR2_X1 U17319 ( .A(n13804), .B(n16038), .ZN(n13805) );
  NAND2_X1 U17320 ( .A1(n13805), .A2(n18917), .ZN(n13813) );
  AOI21_X1 U17321 ( .B1(n13806), .B2(n12985), .A(n13542), .ZN(n13807) );
  INV_X1 U17322 ( .A(n13807), .ZN(n18990) );
  AOI22_X1 U17323 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18939), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n18912), .ZN(n13808) );
  OAI211_X1 U17324 ( .C1(n18921), .C2(n18990), .A(n13808), .B(n18814), .ZN(
        n13811) );
  NOR2_X1 U17325 ( .A1(n13809), .A2(n18927), .ZN(n13810) );
  AOI211_X1 U17326 ( .C1(n18922), .C2(P2_EBX_REG_12__SCAN_IN), .A(n13811), .B(
        n13810), .ZN(n13812) );
  OAI211_X1 U17327 ( .C1(n18959), .C2(n18900), .A(n13813), .B(n13812), .ZN(
        P2_U2843) );
  INV_X1 U17328 ( .A(n19050), .ZN(n13817) );
  NOR2_X1 U17329 ( .A1(n18896), .A2(n13814), .ZN(n13816) );
  AOI21_X1 U17330 ( .B1(n13817), .B2(n13816), .A(n19602), .ZN(n13815) );
  OAI21_X1 U17331 ( .B1(n13817), .B2(n13816), .A(n13815), .ZN(n13825) );
  INV_X1 U17332 ( .A(n18969), .ZN(n19046) );
  AOI22_X1 U17333 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n18922), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18939), .ZN(n13818) );
  INV_X1 U17334 ( .A(n19044), .ZN(n18814) );
  OAI211_X1 U17335 ( .C1(n18921), .C2(n13819), .A(n13818), .B(n18814), .ZN(
        n13820) );
  AOI21_X1 U17336 ( .B1(n13821), .B2(n18885), .A(n13820), .ZN(n13822) );
  OAI21_X1 U17337 ( .B1(n18929), .B2(n10920), .A(n13822), .ZN(n13823) );
  AOI21_X1 U17338 ( .B1(n18933), .B2(n19046), .A(n13823), .ZN(n13824) );
  OAI211_X1 U17339 ( .C1(n18999), .C2(n15063), .A(n13825), .B(n13824), .ZN(
        P2_U2851) );
  NOR2_X1 U17340 ( .A1(n13827), .A2(n13828), .ZN(n13829) );
  OR2_X1 U17341 ( .A1(n13826), .A2(n13829), .ZN(n19782) );
  INV_X1 U17342 ( .A(n13836), .ZN(n13832) );
  INV_X1 U17343 ( .A(n13830), .ZN(n13831) );
  OAI21_X1 U17344 ( .B1(n13832), .B2(n13831), .A(n13927), .ZN(n15894) );
  INV_X1 U17345 ( .A(n15894), .ZN(n19776) );
  AOI22_X1 U17346 ( .A1(n19776), .A2(n14670), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n14669), .ZN(n13833) );
  OAI21_X1 U17347 ( .B1(n19782), .B2(n14672), .A(n13833), .ZN(P1_U2863) );
  AND2_X1 U17348 ( .A1(n13705), .A2(n13834), .ZN(n13835) );
  NOR2_X1 U17349 ( .A1(n13827), .A2(n13835), .ZN(n19795) );
  INV_X1 U17350 ( .A(n19795), .ZN(n13843) );
  INV_X1 U17351 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13839) );
  OAI21_X1 U17352 ( .B1(n13838), .B2(n13837), .A(n13836), .ZN(n19790) );
  OAI222_X1 U17353 ( .A1(n13843), .A2(n14672), .B1(n14682), .B2(n13839), .C1(
        n19790), .C2(n14684), .ZN(P1_U2864) );
  INV_X1 U17354 ( .A(DATAI_8_), .ZN(n13841) );
  INV_X1 U17355 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n13840) );
  MUX2_X1 U17356 ( .A(n13841), .B(n13840), .S(n19976), .Z(n19899) );
  OAI222_X1 U17357 ( .A1(n13843), .A2(n14747), .B1(n19899), .B2(n14744), .C1(
        n13842), .C2(n15728), .ZN(P1_U2896) );
  XOR2_X1 U17358 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n13844), .Z(
        n13845) );
  XNOR2_X1 U17359 ( .A(n13846), .B(n13845), .ZN(n15911) );
  INV_X1 U17360 ( .A(n15911), .ZN(n13850) );
  AOI22_X1 U17361 ( .A1(n19936), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19953), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13847) );
  OAI21_X1 U17362 ( .B1(n15787), .B2(n19793), .A(n13847), .ZN(n13848) );
  AOI21_X1 U17363 ( .B1(n19795), .B2(n12940), .A(n13848), .ZN(n13849) );
  OAI21_X1 U17364 ( .B1(n13850), .B2(n19757), .A(n13849), .ZN(P1_U2991) );
  AND2_X1 U17365 ( .A1(n13629), .A2(n13852), .ZN(n13853) );
  NOR2_X1 U17366 ( .A1(n13851), .A2(n13853), .ZN(n18981) );
  INV_X1 U17367 ( .A(n18981), .ZN(n13864) );
  NAND2_X1 U17368 ( .A1(n13734), .A2(n13854), .ZN(n13855) );
  NAND2_X1 U17369 ( .A1(n13950), .A2(n13855), .ZN(n18950) );
  INV_X1 U17370 ( .A(n18950), .ZN(n15247) );
  NOR2_X1 U17371 ( .A1(n13856), .A2(n18927), .ZN(n13859) );
  AOI22_X1 U17372 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18939), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n18912), .ZN(n13857) );
  OAI211_X1 U17373 ( .C1(n18906), .C2(n18947), .A(n13857), .B(n18814), .ZN(
        n13858) );
  AOI211_X1 U17374 ( .C1(n15247), .C2(n18933), .A(n13859), .B(n13858), .ZN(
        n13863) );
  NOR2_X1 U17375 ( .A1(n18896), .A2(n18830), .ZN(n13860) );
  XNOR2_X1 U17376 ( .A(n13860), .B(n15244), .ZN(n13861) );
  NAND2_X1 U17377 ( .A1(n13861), .A2(n18917), .ZN(n13862) );
  OAI211_X1 U17378 ( .C1(n13864), .C2(n18921), .A(n13863), .B(n13862), .ZN(
        P2_U2839) );
  INV_X1 U17379 ( .A(DATAI_9_), .ZN(n13866) );
  MUX2_X1 U17380 ( .A(n13866), .B(n13865), .S(n19976), .Z(n19902) );
  INV_X1 U17381 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13867) );
  OAI222_X1 U17382 ( .A1(n19782), .A2(n14747), .B1(n19902), .B2(n14744), .C1(
        n13867), .C2(n15728), .ZN(P1_U2895) );
  AOI22_X1 U17383 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13872) );
  AOI22_X1 U17384 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13871) );
  AOI22_X1 U17385 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13870) );
  AOI22_X1 U17386 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10407), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13869) );
  NAND4_X1 U17387 ( .A1(n13872), .A2(n13871), .A3(n13870), .A4(n13869), .ZN(
        n13878) );
  AOI22_X1 U17388 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13876) );
  AOI22_X1 U17389 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13875) );
  AOI22_X1 U17390 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13874) );
  AOI22_X1 U17391 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13873) );
  NAND4_X1 U17392 ( .A1(n13876), .A2(n13875), .A3(n13874), .A4(n13873), .ZN(
        n13877) );
  OR2_X1 U17393 ( .A1(n13878), .A2(n13877), .ZN(n13993) );
  INV_X1 U17394 ( .A(n13993), .ZN(n13889) );
  AOI22_X1 U17395 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10382), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13882) );
  AOI22_X1 U17396 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10406), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13881) );
  AOI22_X1 U17397 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13880) );
  AOI22_X1 U17398 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10407), .B1(
        n14294), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13879) );
  NAND4_X1 U17399 ( .A1(n13882), .A2(n13881), .A3(n13880), .A4(n13879), .ZN(
        n13888) );
  AOI22_X1 U17400 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10372), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13886) );
  AOI22_X1 U17401 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9707), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13885) );
  AOI22_X1 U17402 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10373), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13884) );
  AOI22_X1 U17403 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10360), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13883) );
  NAND4_X1 U17404 ( .A1(n13886), .A2(n13885), .A3(n13884), .A4(n13883), .ZN(
        n13887) );
  NOR2_X1 U17405 ( .A1(n13888), .A2(n13887), .ZN(n13953) );
  OR2_X1 U17406 ( .A1(n13889), .A2(n13953), .ZN(n13900) );
  AOI22_X1 U17407 ( .A1(n14293), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13893) );
  AOI22_X1 U17408 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13892) );
  AOI22_X1 U17409 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13891) );
  AOI22_X1 U17410 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10407), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13890) );
  NAND4_X1 U17411 ( .A1(n13893), .A2(n13892), .A3(n13891), .A4(n13890), .ZN(
        n13899) );
  AOI22_X1 U17412 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13897) );
  AOI22_X1 U17413 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13896) );
  AOI22_X1 U17414 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13895) );
  AOI22_X1 U17415 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13894) );
  NAND4_X1 U17416 ( .A1(n13897), .A2(n13896), .A3(n13895), .A4(n13894), .ZN(
        n13898) );
  NOR2_X1 U17417 ( .A1(n13899), .A2(n13898), .ZN(n18943) );
  NOR2_X1 U17418 ( .A1(n13900), .A2(n18943), .ZN(n13911) );
  AND2_X1 U17419 ( .A1(n14276), .A2(n13911), .ZN(n13996) );
  AOI22_X1 U17420 ( .A1(n14293), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13904) );
  AOI22_X1 U17421 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13903) );
  AOI22_X1 U17422 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13902) );
  AOI22_X1 U17423 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10407), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13901) );
  NAND4_X1 U17424 ( .A1(n13904), .A2(n13903), .A3(n13902), .A4(n13901), .ZN(
        n13910) );
  AOI22_X1 U17425 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13908) );
  AOI22_X1 U17426 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13907) );
  AOI22_X1 U17427 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13906) );
  AOI22_X1 U17428 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13905) );
  NAND4_X1 U17429 ( .A1(n13908), .A2(n13907), .A3(n13906), .A4(n13905), .ZN(
        n13909) );
  OR2_X1 U17430 ( .A1(n13910), .A2(n13909), .ZN(n13912) );
  AND2_X1 U17431 ( .A1(n13912), .A2(n13911), .ZN(n14273) );
  NAND2_X1 U17432 ( .A1(n14276), .A2(n14273), .ZN(n15980) );
  OAI21_X1 U17433 ( .B1(n13996), .B2(n13912), .A(n15980), .ZN(n13992) );
  NAND2_X1 U17434 ( .A1(n18800), .A2(n18980), .ZN(n13923) );
  NAND3_X1 U17435 ( .A1(n15168), .A2(n10203), .A3(n10193), .ZN(n13918) );
  NOR2_X2 U17436 ( .A1(n13918), .A2(n13913), .ZN(n18977) );
  INV_X1 U17437 ( .A(n13914), .ZN(n13915) );
  OAI22_X1 U17438 ( .A1(n19101), .A2(n15169), .B1(n15168), .B2(n13916), .ZN(
        n13921) );
  NOR2_X2 U17439 ( .A1(n13918), .A2(n13917), .ZN(n18976) );
  INV_X1 U17440 ( .A(n18976), .ZN(n14043) );
  INV_X1 U17441 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n13919) );
  NOR2_X1 U17442 ( .A1(n14043), .A2(n13919), .ZN(n13920) );
  AOI211_X1 U17443 ( .C1(BUF1_REG_19__SCAN_IN), .C2(n18977), .A(n13921), .B(
        n13920), .ZN(n13922) );
  OAI211_X1 U17444 ( .C1(n18998), .C2(n13992), .A(n13923), .B(n13922), .ZN(
        P2_U2900) );
  AOI21_X1 U17445 ( .B1(n12012), .B2(n12024), .A(n13925), .ZN(n15711) );
  INV_X1 U17446 ( .A(n15711), .ZN(n13975) );
  INV_X1 U17447 ( .A(n14014), .ZN(n13926) );
  AOI21_X1 U17448 ( .B1(n13928), .B2(n13927), .A(n13926), .ZN(n15706) );
  AOI22_X1 U17449 ( .A1(n15706), .A2(n14670), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14669), .ZN(n13929) );
  OAI21_X1 U17450 ( .B1(n13975), .B2(n14672), .A(n13929), .ZN(P1_U2862) );
  XNOR2_X1 U17451 ( .A(n13931), .B(n13930), .ZN(n16085) );
  OAI21_X1 U17452 ( .B1(n13694), .B2(n13933), .A(n13932), .ZN(n19003) );
  AOI221_X1 U17453 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n13936), .C2(n13935), .A(
        n13934), .ZN(n13937) );
  AOI21_X1 U17454 ( .B1(n19044), .B2(P2_REIP_REG_5__SCAN_IN), .A(n13937), .ZN(
        n13939) );
  NAND2_X1 U17455 ( .A1(n18916), .A2(n16143), .ZN(n13938) );
  OAI211_X1 U17456 ( .C1(n19003), .C2(n16161), .A(n13939), .B(n13938), .ZN(
        n13946) );
  OAI21_X1 U17457 ( .B1(n13943), .B2(n13941), .A(n13940), .ZN(n13942) );
  OAI21_X1 U17458 ( .B1(n13944), .B2(n13943), .A(n13942), .ZN(n16082) );
  NOR2_X1 U17459 ( .A1(n16082), .A2(n19074), .ZN(n13945) );
  AOI211_X1 U17460 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n13947), .A(
        n13946), .B(n13945), .ZN(n13948) );
  OAI21_X1 U17461 ( .B1(n16163), .B2(n16085), .A(n13948), .ZN(P2_U3041) );
  AND2_X1 U17462 ( .A1(n13950), .A2(n13949), .ZN(n13952) );
  OR2_X1 U17463 ( .A1(n13952), .A2(n13951), .ZN(n15334) );
  INV_X1 U17464 ( .A(n14276), .ZN(n18944) );
  NOR2_X1 U17465 ( .A1(n18946), .A2(n13953), .ZN(n13994) );
  AOI21_X1 U17466 ( .B1(n13953), .B2(n18946), .A(n13994), .ZN(n13962) );
  NAND2_X1 U17467 ( .A1(n13962), .A2(n18966), .ZN(n13955) );
  NAND2_X1 U17468 ( .A1(n13516), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13954) );
  OAI211_X1 U17469 ( .C1(n15334), .C2(n13516), .A(n13955), .B(n13954), .ZN(
        P2_U2870) );
  OR2_X1 U17470 ( .A1(n13851), .A2(n13956), .ZN(n13957) );
  NAND2_X1 U17471 ( .A1(n12340), .A2(n13957), .ZN(n18828) );
  OAI22_X1 U17472 ( .A1(n13959), .A2(n15169), .B1(n15168), .B2(n13958), .ZN(
        n13961) );
  NOR2_X1 U17473 ( .A1(n14043), .A2(n18088), .ZN(n13960) );
  AOI211_X1 U17474 ( .C1(BUF1_REG_17__SCAN_IN), .C2(n18977), .A(n13961), .B(
        n13960), .ZN(n13964) );
  NAND2_X1 U17475 ( .A1(n13962), .A2(n15147), .ZN(n13963) );
  OAI211_X1 U17476 ( .C1(n18828), .C2(n15994), .A(n13964), .B(n13963), .ZN(
        P2_U2902) );
  XNOR2_X1 U17477 ( .A(n13965), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13989) );
  XOR2_X1 U17478 ( .A(n13966), .B(n13967), .Z(n13987) );
  OAI22_X1 U17479 ( .A1(n19630), .A2(n18814), .B1(n19061), .B2(n18898), .ZN(
        n13969) );
  NOR2_X1 U17480 ( .A1(n16100), .A2(n9871), .ZN(n13968) );
  NOR2_X1 U17481 ( .A1(n13969), .A2(n13968), .ZN(n13970) );
  OAI21_X1 U17482 ( .B1(n18899), .B2(n16077), .A(n13970), .ZN(n13971) );
  AOI21_X1 U17483 ( .B1(n13987), .B2(n19056), .A(n13971), .ZN(n13972) );
  OAI21_X1 U17484 ( .B1(n13989), .B2(n16083), .A(n13972), .ZN(P2_U3008) );
  INV_X1 U17485 ( .A(DATAI_10_), .ZN(n13973) );
  MUX2_X1 U17486 ( .A(n13973), .B(n16297), .S(n19976), .Z(n19905) );
  INV_X1 U17487 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13974) );
  OAI222_X1 U17488 ( .A1(n14747), .A2(n13975), .B1(n19905), .B2(n14744), .C1(
        n13974), .C2(n15728), .ZN(P1_U2894) );
  AOI211_X1 U17489 ( .C1(n13977), .C2(n13979), .A(n13976), .B(n13978), .ZN(
        n13986) );
  NAND3_X1 U17490 ( .A1(n13979), .A2(n16155), .A3(n13978), .ZN(n13984) );
  OAI22_X1 U17491 ( .A1(n18899), .A2(n19072), .B1(n19630), .B2(n18814), .ZN(
        n13980) );
  INV_X1 U17492 ( .A(n13980), .ZN(n13983) );
  NAND2_X1 U17493 ( .A1(n13981), .A2(n19067), .ZN(n13982) );
  NAND3_X1 U17494 ( .A1(n13984), .A2(n13983), .A3(n13982), .ZN(n13985) );
  AOI211_X1 U17495 ( .C1(n13987), .C2(n19069), .A(n13986), .B(n13985), .ZN(
        n13988) );
  OAI21_X1 U17496 ( .B1(n13989), .B2(n19074), .A(n13988), .ZN(P2_U3040) );
  NAND2_X1 U17497 ( .A1(n18799), .A2(n18965), .ZN(n13991) );
  NAND2_X1 U17498 ( .A1(n13516), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n13990) );
  OAI211_X1 U17499 ( .C1(n13992), .C2(n18951), .A(n13991), .B(n13990), .ZN(
        P2_U2868) );
  NOR2_X1 U17500 ( .A1(n13994), .A2(n13993), .ZN(n13995) );
  NAND2_X1 U17501 ( .A1(n13997), .A2(n18980), .ZN(n14004) );
  OAI22_X1 U17502 ( .A1(n13999), .A2(n15169), .B1(n15168), .B2(n13998), .ZN(
        n14002) );
  INV_X1 U17503 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n14000) );
  NOR2_X1 U17504 ( .A1(n14043), .A2(n14000), .ZN(n14001) );
  AOI211_X1 U17505 ( .C1(BUF1_REG_18__SCAN_IN), .C2(n18977), .A(n14002), .B(
        n14001), .ZN(n14003) );
  OAI211_X1 U17506 ( .C1(n18998), .C2(n15988), .A(n14004), .B(n14003), .ZN(
        P2_U2901) );
  MUX2_X1 U17507 ( .A(n14006), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .S(
        n15766), .Z(n14007) );
  XNOR2_X1 U17508 ( .A(n14005), .B(n14007), .ZN(n15892) );
  INV_X1 U17509 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n14008) );
  OAI22_X1 U17510 ( .A1(n15795), .A2(n19779), .B1(n15908), .B2(n14008), .ZN(
        n14010) );
  NOR2_X1 U17511 ( .A1(n19782), .A2(n19975), .ZN(n14009) );
  AOI211_X1 U17512 ( .C1(n15791), .C2(n19783), .A(n14010), .B(n14009), .ZN(
        n14011) );
  OAI21_X1 U17513 ( .B1(n19757), .B2(n15892), .A(n14011), .ZN(P1_U2990) );
  OR2_X1 U17514 ( .A1(n13925), .A2(n14012), .ZN(n14013) );
  NAND2_X1 U17515 ( .A1(n14153), .A2(n14013), .ZN(n14155) );
  XNOR2_X1 U17516 ( .A(n14155), .B(n14152), .ZN(n15770) );
  INV_X1 U17517 ( .A(n15770), .ZN(n14020) );
  AOI21_X1 U17518 ( .B1(n14015), .B2(n14014), .A(n14674), .ZN(n15874) );
  AOI22_X1 U17519 ( .A1(n15874), .A2(n14670), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14669), .ZN(n14016) );
  OAI21_X1 U17520 ( .B1(n14020), .B2(n14672), .A(n14016), .ZN(P1_U2861) );
  INV_X1 U17521 ( .A(DATAI_11_), .ZN(n14018) );
  MUX2_X1 U17522 ( .A(n14018), .B(n14017), .S(n19976), .Z(n19908) );
  OAI222_X1 U17523 ( .A1(n14020), .A2(n14747), .B1(n19908), .B2(n14744), .C1(
        n14019), .C2(n15728), .ZN(P1_U2893) );
  XNOR2_X1 U17524 ( .A(n14022), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14023) );
  XNOR2_X1 U17525 ( .A(n14021), .B(n14023), .ZN(n16147) );
  INV_X1 U17526 ( .A(n16069), .ZN(n14031) );
  NAND2_X1 U17527 ( .A1(n14024), .A2(n14027), .ZN(n14028) );
  OAI21_X1 U17528 ( .B1(n14029), .B2(n14031), .A(n14028), .ZN(n14030) );
  OAI21_X1 U17529 ( .B1(n14026), .B2(n14031), .A(n14030), .ZN(n16144) );
  OAI22_X1 U17530 ( .A1(n16100), .A2(n14032), .B1(n19632), .B2(n18814), .ZN(
        n14033) );
  AOI21_X1 U17531 ( .B1(n16090), .B2(n18879), .A(n14033), .ZN(n14034) );
  OAI21_X1 U17532 ( .B1(n14035), .B2(n16077), .A(n14034), .ZN(n14036) );
  AOI21_X1 U17533 ( .B1(n16144), .B2(n19056), .A(n14036), .ZN(n14037) );
  OAI21_X1 U17534 ( .B1(n16083), .B2(n16147), .A(n14037), .ZN(P2_U3007) );
  OR2_X1 U17535 ( .A1(n14093), .A2(n14038), .ZN(n14040) );
  NAND2_X1 U17536 ( .A1(n14040), .A2(n14039), .ZN(n18791) );
  OAI22_X1 U17537 ( .A1(n19111), .A2(n15169), .B1(n15168), .B2(n14041), .ZN(
        n14045) );
  INV_X1 U17538 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n14042) );
  NOR2_X1 U17539 ( .A1(n14043), .A2(n14042), .ZN(n14044) );
  AOI211_X1 U17540 ( .C1(BUF1_REG_21__SCAN_IN), .C2(n18977), .A(n14045), .B(
        n14044), .ZN(n14068) );
  AOI22_X1 U17541 ( .A1(n14293), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14049) );
  AOI22_X1 U17542 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14048) );
  AOI22_X1 U17543 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14047) );
  AOI22_X1 U17544 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10407), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14046) );
  NAND4_X1 U17545 ( .A1(n14049), .A2(n14048), .A3(n14047), .A4(n14046), .ZN(
        n14055) );
  AOI22_X1 U17546 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14053) );
  AOI22_X1 U17547 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14052) );
  AOI22_X1 U17548 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14051) );
  AOI22_X1 U17549 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14050) );
  NAND4_X1 U17550 ( .A1(n14053), .A2(n14052), .A3(n14051), .A4(n14050), .ZN(
        n14054) );
  NOR2_X1 U17551 ( .A1(n14055), .A2(n14054), .ZN(n14271) );
  AOI22_X1 U17552 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n14293), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14059) );
  AOI22_X1 U17553 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14058) );
  AOI22_X1 U17554 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14057) );
  AOI22_X1 U17555 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10407), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14056) );
  NAND4_X1 U17556 ( .A1(n14059), .A2(n14058), .A3(n14057), .A4(n14056), .ZN(
        n14065) );
  AOI22_X1 U17557 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14063) );
  AOI22_X1 U17558 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n9708), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14062) );
  AOI22_X1 U17559 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10373), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14061) );
  AOI22_X1 U17560 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10360), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14060) );
  NAND4_X1 U17561 ( .A1(n14063), .A2(n14062), .A3(n14061), .A4(n14060), .ZN(
        n14064) );
  NOR2_X1 U17562 ( .A1(n14065), .A2(n14064), .ZN(n15979) );
  INV_X1 U17563 ( .A(n15164), .ZN(n14066) );
  AOI21_X1 U17564 ( .B1(n14271), .B2(n15982), .A(n14066), .ZN(n14087) );
  NAND2_X1 U17565 ( .A1(n14087), .A2(n15147), .ZN(n14067) );
  OAI211_X1 U17566 ( .C1(n18791), .C2(n15994), .A(n14068), .B(n14067), .ZN(
        P2_U2898) );
  AND2_X1 U17567 ( .A1(n14070), .A2(n14069), .ZN(n14653) );
  OAI21_X1 U17568 ( .B1(n14653), .B2(n14072), .A(n14071), .ZN(n14842) );
  OR2_X1 U17569 ( .A1(n14656), .A2(n14073), .ZN(n14074) );
  AND2_X1 U17570 ( .A1(n14645), .A2(n14074), .ZN(n15819) );
  AOI22_X1 U17571 ( .A1(n15819), .A2(n14670), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14669), .ZN(n14075) );
  OAI21_X1 U17572 ( .B1(n14842), .B2(n14672), .A(n14075), .ZN(P1_U2855) );
  OAI22_X1 U17573 ( .A1(n15716), .A2(n19993), .B1(n15728), .B2(n13198), .ZN(
        n14076) );
  AOI21_X1 U17574 ( .B1(n15720), .B2(DATAI_17_), .A(n14076), .ZN(n14078) );
  NAND2_X1 U17575 ( .A1(n14731), .A2(BUF1_REG_17__SCAN_IN), .ZN(n14077) );
  OAI211_X1 U17576 ( .C1(n14842), .C2(n14747), .A(n14078), .B(n14077), .ZN(
        P1_U2887) );
  INV_X1 U17577 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20692) );
  INV_X1 U17578 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n14593) );
  NOR2_X1 U17579 ( .A1(n20692), .A2(n14593), .ZN(n15674) );
  INV_X1 U17580 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20673) );
  NAND3_X1 U17581 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19844) );
  NOR2_X1 U17582 ( .A1(n20673), .A2(n19844), .ZN(n19774) );
  NAND4_X1 U17583 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n19775)
         );
  NOR2_X1 U17584 ( .A1(n14008), .A2(n19775), .ZN(n15705) );
  NAND3_X1 U17585 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n19774), .A3(n15705), 
        .ZN(n15700) );
  NAND2_X1 U17586 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14079) );
  NOR3_X1 U17587 ( .A1(n19845), .A2(n15700), .A3(n14079), .ZN(n15685) );
  NAND3_X1 U17588 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n15685), .ZN(n14577) );
  INV_X1 U17589 ( .A(n14577), .ZN(n15673) );
  NOR2_X1 U17590 ( .A1(n15700), .A2(n14079), .ZN(n14178) );
  NAND3_X1 U17591 ( .A1(n14178), .A2(P1_REIP_REG_14__SCAN_IN), .A3(
        P1_REIP_REG_13__SCAN_IN), .ZN(n14590) );
  NAND3_X1 U17592 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14578) );
  NOR3_X1 U17593 ( .A1(n19803), .A2(n14590), .A3(n14578), .ZN(n15643) );
  NOR2_X1 U17594 ( .A1(n15641), .A2(n15643), .ZN(n15665) );
  OAI221_X1 U17595 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n15674), .C1(
        P1_REIP_REG_17__SCAN_IN), .C2(n15673), .A(n15665), .ZN(n14083) );
  AOI22_X1 U17596 ( .A1(P1_EBX_REG_17__SCAN_IN), .A2(n19837), .B1(n19865), 
        .B2(n14845), .ZN(n14080) );
  INV_X1 U17597 ( .A(n19836), .ZN(n19777) );
  OAI211_X1 U17598 ( .C1(n19840), .C2(n14841), .A(n14080), .B(n19777), .ZN(
        n14081) );
  AOI21_X1 U17599 ( .B1(n15819), .B2(n19863), .A(n14081), .ZN(n14082) );
  OAI211_X1 U17600 ( .C1(n14842), .C2(n15629), .A(n14083), .B(n14082), .ZN(
        P1_U2823) );
  NOR2_X1 U17601 ( .A1(n14096), .A2(n14085), .ZN(n14086) );
  OR2_X1 U17602 ( .A1(n14084), .A2(n14086), .ZN(n18777) );
  NAND2_X1 U17603 ( .A1(n14087), .A2(n18966), .ZN(n14089) );
  NAND2_X1 U17604 ( .A1(n13516), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n14088) );
  OAI211_X1 U17605 ( .C1(n18777), .C2(n13516), .A(n14089), .B(n14088), .ZN(
        P2_U2866) );
  NOR2_X1 U17606 ( .A1(n14091), .A2(n14090), .ZN(n14092) );
  OR2_X1 U17607 ( .A1(n14093), .A2(n14092), .ZN(n15995) );
  AND2_X1 U17608 ( .A1(n14095), .A2(n14094), .ZN(n14097) );
  OR2_X1 U17609 ( .A1(n14097), .A2(n14096), .ZN(n15986) );
  INV_X1 U17610 ( .A(n15986), .ZN(n14104) );
  AOI22_X1 U17611 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18939), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18912), .ZN(n14100) );
  INV_X1 U17612 ( .A(n18829), .ZN(n18934) );
  OAI211_X1 U17613 ( .C1(n14098), .C2(n15225), .A(n18934), .B(n18785), .ZN(
        n14099) );
  OAI211_X1 U17614 ( .C1(n18906), .C2(n15983), .A(n14100), .B(n14099), .ZN(
        n14103) );
  OAI22_X1 U17615 ( .A1(n14101), .A2(n18927), .B1(n15225), .B2(n18816), .ZN(
        n14102) );
  AOI211_X1 U17616 ( .C1(n14104), .C2(n18933), .A(n14103), .B(n14102), .ZN(
        n14105) );
  OAI21_X1 U17617 ( .B1(n15995), .B2(n18921), .A(n14105), .ZN(P2_U2835) );
  INV_X1 U17618 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n16632) );
  NAND3_X1 U17619 ( .A1(n18104), .A2(n17097), .A3(n14106), .ZN(n14107) );
  INV_X1 U17620 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n20840) );
  INV_X1 U17621 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n14109) );
  NOR2_X1 U17622 ( .A1(n20840), .A2(n14109), .ZN(n17082) );
  NAND4_X1 U17623 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .A4(n17082), .ZN(n17074) );
  AND2_X2 U17624 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17012), .ZN(n17025) );
  INV_X1 U17625 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16971) );
  NOR3_X1 U17626 ( .A1(n16550), .A2(n16971), .A3(n20869), .ZN(n15503) );
  AND3_X1 U17627 ( .A1(n17097), .A2(n16985), .A3(n15503), .ZN(n16948) );
  NOR2_X1 U17628 ( .A1(n16971), .A2(n20869), .ZN(n14110) );
  AOI21_X1 U17629 ( .B1(n16985), .B2(n14110), .A(P3_EBX_REG_15__SCAN_IN), .ZN(
        n14111) );
  NOR2_X1 U17630 ( .A1(n16948), .A2(n14111), .ZN(n14123) );
  AOI22_X1 U17631 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n9714), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17044), .ZN(n14115) );
  INV_X1 U17632 ( .A(n9719), .ZN(n17046) );
  AOI22_X1 U17633 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14114) );
  AOI22_X1 U17634 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14113) );
  AOI22_X1 U17635 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12571), .B1(
        n17033), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14112) );
  NAND4_X1 U17636 ( .A1(n14115), .A2(n14114), .A3(n14113), .A4(n14112), .ZN(
        n14121) );
  AOI22_X1 U17637 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n9709), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n17017), .ZN(n14119) );
  AOI22_X1 U17638 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14118) );
  AOI22_X1 U17639 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n16755), .ZN(n14117) );
  AOI22_X1 U17640 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17050), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17048), .ZN(n14116) );
  NAND4_X1 U17641 ( .A1(n14119), .A2(n14118), .A3(n14117), .A4(n14116), .ZN(
        n14120) );
  NOR2_X1 U17642 ( .A1(n14121), .A2(n14120), .ZN(n17181) );
  INV_X1 U17643 ( .A(n17181), .ZN(n14122) );
  NOR2_X2 U17644 ( .A1(n17085), .A2(n17097), .ZN(n17089) );
  MUX2_X1 U17645 ( .A(n14123), .B(n14122), .S(n17089), .Z(P3_U2688) );
  OAI211_X1 U17646 ( .C1(n18686), .C2(n18535), .A(n16870), .B(n18525), .ZN(
        n18067) );
  NOR2_X1 U17647 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18067), .ZN(n14124) );
  NAND3_X1 U17648 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18676)
         );
  OAI21_X1 U17649 ( .B1(n14124), .B2(n18676), .A(n18189), .ZN(n18078) );
  INV_X1 U17650 ( .A(n18078), .ZN(n14125) );
  NOR2_X1 U17651 ( .A1(n17705), .A2(n18725), .ZN(n18071) );
  AOI21_X1 U17652 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18071), .ZN(n18072) );
  NOR2_X1 U17653 ( .A1(n14125), .A2(n18072), .ZN(n14127) );
  INV_X1 U17654 ( .A(n18423), .ZN(n18073) );
  NOR2_X1 U17655 ( .A1(n18678), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18126) );
  OR2_X1 U17656 ( .A1(n18126), .A2(n14125), .ZN(n18070) );
  OR2_X1 U17657 ( .A1(n18073), .A2(n18070), .ZN(n14126) );
  MUX2_X1 U17658 ( .A(n14127), .B(n14126), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  AOI22_X1 U17659 ( .A1(n14128), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14131) );
  NAND2_X1 U17660 ( .A1(n14129), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14130) );
  OAI211_X1 U17661 ( .C1(n14132), .C2(n14139), .A(n14131), .B(n14130), .ZN(
        n14133) );
  NAND2_X1 U17662 ( .A1(n14135), .A2(n18934), .ZN(n14151) );
  INV_X1 U17663 ( .A(n15953), .ZN(n14138) );
  NOR2_X1 U17664 ( .A1(n14136), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14137) );
  MUX2_X1 U17665 ( .A(n14138), .B(n14137), .S(n9757), .Z(n14239) );
  INV_X1 U17666 ( .A(P2_EAX_REG_31__SCAN_IN), .ZN(n14141) );
  OAI22_X1 U17667 ( .A1(n14142), .A2(n14141), .B1(n14140), .B2(n14139), .ZN(
        n14143) );
  AOI21_X1 U17668 ( .B1(n14144), .B2(P2_REIP_REG_31__SCAN_IN), .A(n14143), 
        .ZN(n14145) );
  XNOR2_X2 U17669 ( .A(n14146), .B(n14145), .ZN(n14467) );
  NAND2_X1 U17670 ( .A1(n18912), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14148) );
  AOI22_X1 U17671 ( .A1(n18922), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n18939), .ZN(n14147) );
  OAI211_X1 U17672 ( .C1(n14467), .C2(n18921), .A(n14148), .B(n14147), .ZN(
        n14149) );
  AOI21_X1 U17673 ( .B1(n14239), .B2(n18885), .A(n14149), .ZN(n14150) );
  OAI211_X1 U17674 ( .C1(n15976), .C2(n18900), .A(n14151), .B(n14150), .ZN(
        P2_U2824) );
  INV_X1 U17675 ( .A(n14152), .ZN(n14154) );
  OAI21_X1 U17676 ( .B1(n14155), .B2(n14154), .A(n14153), .ZN(n14676) );
  NAND2_X1 U17677 ( .A1(n14157), .A2(n14156), .ZN(n14664) );
  OAI21_X1 U17678 ( .B1(n14678), .B2(n14158), .A(n14664), .ZN(n14746) );
  OAI22_X1 U17679 ( .A1(n15765), .A2(n14161), .B1(n14160), .B2(n9736), .ZN(
        n15760) );
  NOR2_X1 U17680 ( .A1(n15766), .A2(n14162), .ZN(n14163) );
  NOR2_X1 U17681 ( .A1(n15760), .A2(n15759), .ZN(n15758) );
  NOR2_X1 U17682 ( .A1(n15758), .A2(n14164), .ZN(n14166) );
  XNOR2_X1 U17683 ( .A(n14166), .B(n14165), .ZN(n15855) );
  NAND2_X1 U17684 ( .A1(n15855), .A2(n19938), .ZN(n14170) );
  INV_X1 U17685 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n14167) );
  OAI22_X1 U17686 ( .A1(n15795), .A2(n14177), .B1(n15908), .B2(n14167), .ZN(
        n14168) );
  AOI21_X1 U17687 ( .B1(n15791), .B2(n14183), .A(n14168), .ZN(n14169) );
  OAI211_X1 U17688 ( .C1(n19975), .C2(n14746), .A(n14170), .B(n14169), .ZN(
        P1_U2986) );
  OR2_X1 U17689 ( .A1(n14172), .A2(n14173), .ZN(n14174) );
  AND2_X1 U17690 ( .A1(n14171), .A2(n14174), .ZN(n15854) );
  AOI22_X1 U17691 ( .A1(n15854), .A2(n14670), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14669), .ZN(n14175) );
  OAI21_X1 U17692 ( .B1(n14746), .B2(n14672), .A(n14175), .ZN(P1_U2859) );
  AOI22_X1 U17693 ( .A1(n15854), .A2(n19863), .B1(n19837), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14176) );
  OAI211_X1 U17694 ( .C1(n19840), .C2(n14177), .A(n14176), .B(n19777), .ZN(
        n14182) );
  OAI21_X1 U17695 ( .B1(n19845), .B2(n14178), .A(n19773), .ZN(n14179) );
  INV_X1 U17696 ( .A(n14179), .ZN(n15697) );
  INV_X1 U17697 ( .A(n15685), .ZN(n14180) );
  AOI22_X1 U17698 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n15697), .B1(n14180), 
        .B2(n14167), .ZN(n14181) );
  AOI211_X1 U17699 ( .C1(n19865), .C2(n14183), .A(n14182), .B(n14181), .ZN(
        n14184) );
  OAI21_X1 U17700 ( .B1(n14746), .B2(n15629), .A(n14184), .ZN(P1_U2827) );
  NOR2_X1 U17701 ( .A1(n14186), .A2(n14185), .ZN(n14189) );
  XOR2_X1 U17702 ( .A(n14189), .B(n14188), .Z(n14233) );
  AOI21_X1 U17703 ( .B1(n14190), .B2(n10025), .A(n10083), .ZN(n15097) );
  AOI21_X1 U17704 ( .B1(n14192), .B2(n15150), .A(n14191), .ZN(n15040) );
  INV_X1 U17705 ( .A(n15040), .ZN(n15140) );
  NAND2_X1 U17706 ( .A1(n16060), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n14226) );
  OAI21_X1 U17707 ( .B1(n16161), .B2(n15140), .A(n14226), .ZN(n14193) );
  AOI21_X1 U17708 ( .B1(n14194), .B2(n14196), .A(n14193), .ZN(n14195) );
  OAI21_X1 U17709 ( .B1(n14197), .B2(n14196), .A(n14195), .ZN(n14200) );
  NOR3_X1 U17710 ( .A1(n14229), .A2(n14228), .A3(n19074), .ZN(n14199) );
  AOI211_X1 U17711 ( .C1(n15097), .C2(n16143), .A(n14200), .B(n14199), .ZN(
        n14201) );
  OAI21_X1 U17712 ( .B1(n14233), .B2(n16163), .A(n14201), .ZN(P2_U3021) );
  NAND2_X1 U17713 ( .A1(n14203), .A2(n14202), .ZN(n14211) );
  INV_X1 U17714 ( .A(n14204), .ZN(n14205) );
  NAND2_X1 U17715 ( .A1(n15222), .A2(n15221), .ZN(n15220) );
  NAND2_X1 U17716 ( .A1(n15220), .A2(n14209), .ZN(n14210) );
  XOR2_X1 U17717 ( .A(n14211), .B(n14210), .Z(n14225) );
  NOR2_X1 U17718 ( .A1(n15224), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14212) );
  NOR2_X1 U17719 ( .A1(n15303), .A2(n14212), .ZN(n14223) );
  NOR2_X1 U17720 ( .A1(n18791), .A2(n16161), .ZN(n14217) );
  NAND2_X1 U17721 ( .A1(n16060), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n14219) );
  OAI21_X1 U17722 ( .B1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n14214), .A(
        n14213), .ZN(n14215) );
  OAI211_X1 U17723 ( .C1(n18777), .C2(n19072), .A(n14219), .B(n14215), .ZN(
        n14216) );
  AOI211_X1 U17724 ( .C1(n14223), .C2(n16153), .A(n14217), .B(n14216), .ZN(
        n14218) );
  OAI21_X1 U17725 ( .B1(n14225), .B2(n16163), .A(n14218), .ZN(P2_U3025) );
  OAI21_X1 U17726 ( .B1(n16100), .B2(n18778), .A(n14219), .ZN(n14220) );
  AOI21_X1 U17727 ( .B1(n16090), .B2(n18784), .A(n14220), .ZN(n14221) );
  OAI21_X1 U17728 ( .B1(n18777), .B2(n16077), .A(n14221), .ZN(n14222) );
  AOI21_X1 U17729 ( .B1(n14223), .B2(n14248), .A(n14222), .ZN(n14224) );
  OAI21_X1 U17730 ( .B1(n14225), .B2(n16084), .A(n14224), .ZN(P2_U2993) );
  NAND2_X1 U17731 ( .A1(n16090), .A2(n15044), .ZN(n14227) );
  OAI211_X1 U17732 ( .C1(n15038), .C2(n16100), .A(n14227), .B(n14226), .ZN(
        n14231) );
  NOR3_X1 U17733 ( .A1(n14229), .A2(n14228), .A3(n16083), .ZN(n14230) );
  OAI21_X1 U17734 ( .B1(n14233), .B2(n16084), .A(n14232), .ZN(P2_U2989) );
  NAND2_X1 U17735 ( .A1(n14239), .A2(n14238), .ZN(n14240) );
  XNOR2_X1 U17736 ( .A(n14240), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14241) );
  XNOR2_X1 U17737 ( .A(n14242), .B(n14241), .ZN(n14473) );
  NAND2_X1 U17738 ( .A1(n19044), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14463) );
  NAND2_X1 U17739 ( .A1(n19055), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14243) );
  OAI211_X1 U17740 ( .C1(n19061), .C2(n14244), .A(n14463), .B(n14243), .ZN(
        n14245) );
  INV_X1 U17741 ( .A(n14245), .ZN(n14250) );
  NAND2_X1 U17742 ( .A1(n14246), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14247) );
  XNOR2_X2 U17743 ( .A(n14247), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14471) );
  NAND2_X1 U17744 ( .A1(n14471), .A2(n14248), .ZN(n14249) );
  OAI21_X1 U17745 ( .B1(n14473), .B2(n16084), .A(n9802), .ZN(P2_U2983) );
  NAND2_X1 U17746 ( .A1(n18926), .A2(n14251), .ZN(n14252) );
  NAND2_X1 U17747 ( .A1(n19052), .A2(n14252), .ZN(n16162) );
  INV_X1 U17748 ( .A(n16162), .ZN(n14256) );
  OAI21_X1 U17749 ( .B1(n14254), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14253), .ZN(n16168) );
  OR2_X1 U17750 ( .A1(n11123), .A2(n18928), .ZN(n16166) );
  OAI21_X1 U17751 ( .B1(n16083), .B2(n16168), .A(n16166), .ZN(n14255) );
  AOI21_X1 U17752 ( .B1(n19056), .B2(n14256), .A(n14255), .ZN(n14259) );
  OAI21_X1 U17753 ( .B1(n19055), .B2(n14257), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14258) );
  OAI211_X1 U17754 ( .C1(n16077), .C2(n13005), .A(n14259), .B(n14258), .ZN(
        P2_U3014) );
  AOI22_X1 U17755 ( .A1(n14293), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14263) );
  AOI22_X1 U17756 ( .A1(n10406), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14262) );
  AOI22_X1 U17757 ( .A1(n10355), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14261) );
  AOI22_X1 U17758 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10407), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14260) );
  NAND4_X1 U17759 ( .A1(n14263), .A2(n14262), .A3(n14261), .A4(n14260), .ZN(
        n14270) );
  AOI22_X1 U17760 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14268) );
  AOI22_X1 U17761 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14267) );
  AOI22_X1 U17762 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14266) );
  AOI22_X1 U17763 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14265) );
  NAND4_X1 U17764 ( .A1(n14268), .A2(n14267), .A3(n14266), .A4(n14265), .ZN(
        n14269) );
  NOR2_X1 U17765 ( .A1(n14270), .A2(n14269), .ZN(n15165) );
  OR2_X1 U17766 ( .A1(n15165), .A2(n14271), .ZN(n14272) );
  NOR2_X1 U17767 ( .A1(n14272), .A2(n15979), .ZN(n14274) );
  AND2_X1 U17768 ( .A1(n14274), .A2(n14273), .ZN(n14275) );
  INV_X1 U17769 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n19227) );
  AOI22_X1 U17770 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14313), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14284) );
  AOI22_X1 U17771 ( .A1(n9755), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(n9748), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14283) );
  AOI22_X1 U17772 ( .A1(n9742), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n9771), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14282) );
  NAND2_X1 U17773 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n14280) );
  NAND2_X1 U17774 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14279) );
  AND2_X1 U17775 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14278) );
  OR2_X1 U17776 ( .A1(n14278), .A2(n14277), .ZN(n14440) );
  AND3_X1 U17777 ( .A1(n14280), .A2(n14279), .A3(n14440), .ZN(n14281) );
  NAND4_X1 U17778 ( .A1(n14284), .A2(n14283), .A3(n14282), .A4(n14281), .ZN(
        n14292) );
  INV_X1 U17779 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n19511) );
  AOI22_X1 U17780 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14313), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14290) );
  INV_X1 U17781 ( .A(n14440), .ZN(n14415) );
  NAND2_X1 U17782 ( .A1(n14439), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n14286) );
  NAND2_X1 U17783 ( .A1(n9754), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n14285) );
  AND3_X1 U17784 ( .A1(n14415), .A2(n14286), .A3(n14285), .ZN(n14289) );
  AOI22_X1 U17785 ( .A1(n9742), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9749), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14288) );
  AOI22_X1 U17786 ( .A1(n10296), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9759), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14287) );
  NAND4_X1 U17787 ( .A1(n14290), .A2(n14289), .A3(n14288), .A4(n14287), .ZN(
        n14291) );
  NAND2_X1 U17788 ( .A1(n14292), .A2(n14291), .ZN(n14330) );
  NOR2_X1 U17789 ( .A1(n19737), .A2(n14330), .ZN(n14312) );
  AOI22_X1 U17790 ( .A1(n14293), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10406), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14298) );
  AOI22_X1 U17791 ( .A1(n10354), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10352), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14297) );
  AOI22_X1 U17792 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10355), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14296) );
  AOI22_X1 U17793 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14295) );
  NAND4_X1 U17794 ( .A1(n14298), .A2(n14297), .A3(n14296), .A4(n14295), .ZN(
        n14307) );
  AOI22_X1 U17795 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10372), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14305) );
  AOI22_X1 U17796 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14304) );
  AOI22_X1 U17797 ( .A1(n10373), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10374), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14303) );
  AOI22_X1 U17798 ( .A1(n10388), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14302) );
  NAND4_X1 U17799 ( .A1(n14305), .A2(n14304), .A3(n14303), .A4(n14302), .ZN(
        n14306) );
  NOR2_X1 U17800 ( .A1(n14307), .A2(n14306), .ZN(n14329) );
  XNOR2_X1 U17801 ( .A(n14312), .B(n14329), .ZN(n14310) );
  INV_X1 U17802 ( .A(n14330), .ZN(n14308) );
  NAND2_X1 U17803 ( .A1(n19737), .A2(n14308), .ZN(n15108) );
  INV_X1 U17804 ( .A(n14312), .ZN(n14328) );
  AOI22_X1 U17805 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14319) );
  AOI22_X1 U17806 ( .A1(n9742), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10297), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14318) );
  AOI22_X1 U17807 ( .A1(n14313), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9759), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14317) );
  NAND2_X1 U17808 ( .A1(n9771), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14315) );
  NAND2_X1 U17809 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14314) );
  AND3_X1 U17810 ( .A1(n14315), .A2(n14314), .A3(n14440), .ZN(n14316) );
  NAND4_X1 U17811 ( .A1(n14319), .A2(n14318), .A3(n14317), .A4(n14316), .ZN(
        n14327) );
  AOI22_X1 U17812 ( .A1(n9755), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14313), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14325) );
  NAND2_X1 U17813 ( .A1(n9771), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n14321) );
  NAND2_X1 U17814 ( .A1(n9754), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n14320) );
  AND3_X1 U17815 ( .A1(n14415), .A2(n14321), .A3(n14320), .ZN(n14324) );
  AOI22_X1 U17816 ( .A1(n10295), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9760), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14323) );
  AOI22_X1 U17817 ( .A1(n9742), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10297), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14322) );
  NAND4_X1 U17818 ( .A1(n14325), .A2(n14324), .A3(n14323), .A4(n14322), .ZN(
        n14326) );
  NAND2_X1 U17819 ( .A1(n14327), .A2(n14326), .ZN(n14333) );
  OAI21_X1 U17820 ( .B1(n14329), .B2(n14328), .A(n14333), .ZN(n14335) );
  INV_X1 U17821 ( .A(n14329), .ZN(n14332) );
  NOR2_X1 U17822 ( .A1(n14333), .A2(n14330), .ZN(n14331) );
  NAND2_X1 U17823 ( .A1(n14332), .A2(n14331), .ZN(n14350) );
  INV_X1 U17824 ( .A(n14333), .ZN(n14334) );
  AOI22_X1 U17825 ( .A1(n14335), .A2(n14350), .B1(n19737), .B2(n14334), .ZN(
        n15103) );
  AOI22_X1 U17826 ( .A1(n10296), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14313), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14341) );
  NAND2_X1 U17827 ( .A1(n9771), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n14337) );
  NAND2_X1 U17828 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n14336) );
  AND3_X1 U17829 ( .A1(n14415), .A2(n14337), .A3(n14336), .ZN(n14340) );
  AOI22_X1 U17830 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9760), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14339) );
  AOI22_X1 U17831 ( .A1(n9742), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9749), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14338) );
  NAND4_X1 U17832 ( .A1(n14341), .A2(n14340), .A3(n14339), .A4(n14338), .ZN(
        n14349) );
  AOI22_X1 U17833 ( .A1(n9755), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14313), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14347) );
  AOI22_X1 U17834 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n9759), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14346) );
  AOI22_X1 U17835 ( .A1(n9742), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n9748), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14345) );
  NAND2_X1 U17836 ( .A1(n9771), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n14343) );
  NAND2_X1 U17837 ( .A1(n9754), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14342) );
  AND3_X1 U17838 ( .A1(n14343), .A2(n14342), .A3(n14440), .ZN(n14344) );
  NAND4_X1 U17839 ( .A1(n14347), .A2(n14346), .A3(n14345), .A4(n14344), .ZN(
        n14348) );
  AND2_X1 U17840 ( .A1(n14349), .A2(n14348), .ZN(n14352) );
  INV_X1 U17841 ( .A(n14350), .ZN(n14351) );
  NAND2_X1 U17842 ( .A1(n14351), .A2(n14352), .ZN(n14377) );
  OAI211_X1 U17843 ( .C1(n14352), .C2(n14351), .A(n14392), .B(n14377), .ZN(
        n14355) );
  INV_X1 U17844 ( .A(n14352), .ZN(n14353) );
  NOR2_X1 U17845 ( .A1(n10215), .A2(n14353), .ZN(n15095) );
  INV_X1 U17846 ( .A(n14354), .ZN(n15148) );
  AOI22_X1 U17847 ( .A1(n10296), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14313), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14363) );
  NAND2_X1 U17848 ( .A1(n9771), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n14359) );
  NAND2_X1 U17849 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n14358) );
  AND3_X1 U17850 ( .A1(n14415), .A2(n14359), .A3(n14358), .ZN(n14362) );
  AOI22_X1 U17851 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9759), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14361) );
  AOI22_X1 U17852 ( .A1(n9742), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10297), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14360) );
  NAND4_X1 U17853 ( .A1(n14363), .A2(n14362), .A3(n14361), .A4(n14360), .ZN(
        n14371) );
  AOI22_X1 U17854 ( .A1(n9755), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14313), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14369) );
  AOI22_X1 U17855 ( .A1(n10295), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9760), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14368) );
  AOI22_X1 U17856 ( .A1(n9742), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n9748), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14367) );
  NAND2_X1 U17857 ( .A1(n9771), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n14365) );
  NAND2_X1 U17858 ( .A1(n9754), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14364) );
  AND3_X1 U17859 ( .A1(n14365), .A2(n14364), .A3(n14440), .ZN(n14366) );
  NAND4_X1 U17860 ( .A1(n14369), .A2(n14368), .A3(n14367), .A4(n14366), .ZN(
        n14370) );
  AND2_X1 U17861 ( .A1(n14371), .A2(n14370), .ZN(n14375) );
  XNOR2_X1 U17862 ( .A(n14377), .B(n14375), .ZN(n14372) );
  NAND2_X1 U17863 ( .A1(n19737), .A2(n14375), .ZN(n15090) );
  INV_X1 U17864 ( .A(n14375), .ZN(n14376) );
  NOR2_X1 U17865 ( .A1(n14377), .A2(n14376), .ZN(n14393) );
  INV_X1 U17866 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n20817) );
  AOI22_X1 U17867 ( .A1(n10295), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14313), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14383) );
  NAND2_X1 U17868 ( .A1(n9760), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14379) );
  NAND2_X1 U17869 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n14378) );
  AND3_X1 U17870 ( .A1(n14415), .A2(n14379), .A3(n14378), .ZN(n14382) );
  AOI22_X1 U17871 ( .A1(n10296), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10297), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14381) );
  INV_X1 U17872 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n21013) );
  AOI22_X1 U17873 ( .A1(n9742), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9771), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14380) );
  NAND4_X1 U17874 ( .A1(n14383), .A2(n14382), .A3(n14381), .A4(n14380), .ZN(
        n14391) );
  AOI22_X1 U17875 ( .A1(n9755), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n9742), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14389) );
  AOI22_X1 U17876 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n9749), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14388) );
  AOI22_X1 U17877 ( .A1(n14313), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9759), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14387) );
  NAND2_X1 U17878 ( .A1(n9771), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14385) );
  NAND2_X1 U17879 ( .A1(n9754), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14384) );
  AND3_X1 U17880 ( .A1(n14385), .A2(n14384), .A3(n14440), .ZN(n14386) );
  NAND4_X1 U17881 ( .A1(n14389), .A2(n14388), .A3(n14387), .A4(n14386), .ZN(
        n14390) );
  AND2_X1 U17882 ( .A1(n14391), .A2(n14390), .ZN(n14396) );
  NAND2_X1 U17883 ( .A1(n14393), .A2(n14396), .ZN(n15077) );
  OAI211_X1 U17884 ( .C1(n14393), .C2(n14396), .A(n14392), .B(n15077), .ZN(
        n14394) );
  INV_X1 U17885 ( .A(n14396), .ZN(n14397) );
  NOR2_X1 U17886 ( .A1(n10215), .A2(n14397), .ZN(n15085) );
  NAND2_X1 U17887 ( .A1(n15083), .A2(n15085), .ZN(n15084) );
  INV_X1 U17888 ( .A(n14398), .ZN(n15078) );
  AOI22_X1 U17889 ( .A1(n10296), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14313), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14404) );
  NAND2_X1 U17890 ( .A1(n9771), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n14400) );
  NAND2_X1 U17891 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n14399) );
  AND3_X1 U17892 ( .A1(n14415), .A2(n14400), .A3(n14399), .ZN(n14403) );
  AOI22_X1 U17893 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9760), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14402) );
  AOI22_X1 U17894 ( .A1(n9742), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9749), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14401) );
  NAND4_X1 U17895 ( .A1(n14404), .A2(n14403), .A3(n14402), .A4(n14401), .ZN(
        n14412) );
  AOI22_X1 U17896 ( .A1(n10296), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14313), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14410) );
  AOI22_X1 U17897 ( .A1(n10295), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9760), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14409) );
  AOI22_X1 U17898 ( .A1(n9742), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9749), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14408) );
  NAND2_X1 U17899 ( .A1(n9771), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14406) );
  NAND2_X1 U17900 ( .A1(n9754), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n14405) );
  AND3_X1 U17901 ( .A1(n14406), .A2(n14405), .A3(n14440), .ZN(n14407) );
  NAND4_X1 U17902 ( .A1(n14410), .A2(n14409), .A3(n14408), .A4(n14407), .ZN(
        n14411) );
  NAND2_X1 U17903 ( .A1(n14412), .A2(n14411), .ZN(n15080) );
  AOI21_X2 U17904 ( .B1(n15084), .B2(n15078), .A(n15080), .ZN(n15074) );
  AOI22_X1 U17905 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9742), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14419) );
  NAND2_X1 U17906 ( .A1(n9759), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14414) );
  NAND2_X1 U17907 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n14413) );
  AND3_X1 U17908 ( .A1(n14415), .A2(n14414), .A3(n14413), .ZN(n14418) );
  AOI22_X1 U17909 ( .A1(n9755), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10297), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14417) );
  AOI22_X1 U17910 ( .A1(n14313), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9771), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14416) );
  NAND4_X1 U17911 ( .A1(n14419), .A2(n14418), .A3(n14417), .A4(n14416), .ZN(
        n14427) );
  AOI22_X1 U17912 ( .A1(n10296), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9742), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14425) );
  AOI22_X1 U17913 ( .A1(n10295), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9748), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14424) );
  AOI22_X1 U17914 ( .A1(n14313), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9759), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14423) );
  NAND2_X1 U17915 ( .A1(n9771), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n14421) );
  NAND2_X1 U17916 ( .A1(n9754), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n14420) );
  AND3_X1 U17917 ( .A1(n14421), .A2(n14420), .A3(n14440), .ZN(n14422) );
  NAND4_X1 U17918 ( .A1(n14425), .A2(n14424), .A3(n14423), .A4(n14422), .ZN(
        n14426) );
  NAND2_X1 U17919 ( .A1(n14427), .A2(n14426), .ZN(n14429) );
  OR3_X1 U17920 ( .A1(n15077), .A2(n19737), .A3(n15080), .ZN(n14428) );
  NOR2_X1 U17921 ( .A1(n14428), .A2(n14429), .ZN(n14430) );
  AOI21_X1 U17922 ( .B1(n14429), .B2(n14428), .A(n14430), .ZN(n15073) );
  AND2_X2 U17923 ( .A1(n15074), .A2(n15073), .ZN(n15114) );
  NOR2_X1 U17924 ( .A1(n15114), .A2(n14430), .ZN(n14449) );
  AOI22_X1 U17925 ( .A1(n10296), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9742), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14432) );
  AOI22_X1 U17926 ( .A1(n14313), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9748), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14431) );
  NAND2_X1 U17927 ( .A1(n14432), .A2(n14431), .ZN(n14447) );
  INV_X1 U17928 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14436) );
  AOI22_X1 U17929 ( .A1(n9770), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9759), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14435) );
  AOI21_X1 U17930 ( .B1(n9754), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(n14440), .ZN(n14434) );
  OAI211_X1 U17931 ( .C1(n10298), .C2(n14436), .A(n14435), .B(n14434), .ZN(
        n14446) );
  AOI22_X1 U17932 ( .A1(n9769), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n9755), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14438) );
  AOI22_X1 U17933 ( .A1(n9742), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n9749), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14437) );
  NAND2_X1 U17934 ( .A1(n14438), .A2(n14437), .ZN(n14445) );
  AOI22_X1 U17935 ( .A1(n14313), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9759), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14443) );
  NAND2_X1 U17936 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14442) );
  NAND2_X1 U17937 ( .A1(n9771), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n14441) );
  NAND4_X1 U17938 ( .A1(n14443), .A2(n14442), .A3(n14441), .A4(n14440), .ZN(
        n14444) );
  OAI22_X1 U17939 ( .A1(n14447), .A2(n14446), .B1(n14445), .B2(n14444), .ZN(
        n14448) );
  XNOR2_X1 U17940 ( .A(n14449), .B(n14448), .ZN(n14457) );
  NOR2_X1 U17941 ( .A1(n15180), .A2(n13516), .ZN(n14450) );
  AOI21_X1 U17942 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n13516), .A(n14450), .ZN(
        n14451) );
  OAI21_X1 U17943 ( .B1(n14457), .B2(n18951), .A(n14451), .ZN(P2_U2857) );
  OAI22_X1 U17944 ( .A1(n14452), .A2(n15169), .B1(n15168), .B2(n13120), .ZN(
        n14453) );
  AOI21_X1 U17945 ( .B1(n14454), .B2(n18980), .A(n14453), .ZN(n14456) );
  AOI22_X1 U17946 ( .A1(n18976), .A2(BUF2_REG_30__SCAN_IN), .B1(n18977), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n14455) );
  OAI211_X1 U17947 ( .C1(n14457), .C2(n18998), .A(n14456), .B(n14455), .ZN(
        P2_U2889) );
  NOR4_X1 U17948 ( .A1(n15251), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14459), .A4(n14458), .ZN(n14460) );
  OAI21_X1 U17949 ( .B1(n15285), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14461), .ZN(n14462) );
  INV_X1 U17950 ( .A(n14462), .ZN(n14464) );
  INV_X1 U17951 ( .A(n14468), .ZN(n14469) );
  OAI21_X1 U17952 ( .B1(n15976), .B2(n19072), .A(n14469), .ZN(n14470) );
  OAI21_X1 U17953 ( .B1(n14473), .B2(n16163), .A(n14472), .ZN(P2_U3015) );
  NAND2_X1 U17954 ( .A1(n14521), .A2(n14476), .ZN(n14477) );
  AOI22_X1 U17955 ( .A1(n14878), .A2(n14670), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14669), .ZN(n14478) );
  OAI21_X1 U17956 ( .B1(n14474), .B2(n14672), .A(n14478), .ZN(P1_U2843) );
  INV_X1 U17957 ( .A(n14479), .ZN(n14481) );
  AOI22_X1 U17958 ( .A1(n19858), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        n19837), .B2(P1_EBX_REG_29__SCAN_IN), .ZN(n14480) );
  OAI21_X1 U17959 ( .B1(n19851), .B2(n14481), .A(n14480), .ZN(n14485) );
  INV_X1 U17960 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20702) );
  NAND3_X1 U17961 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_18__SCAN_IN), .ZN(n15645) );
  INV_X1 U17962 ( .A(n15645), .ZN(n15642) );
  NAND2_X1 U17963 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n15642), .ZN(n15625) );
  NOR3_X1 U17964 ( .A1(n14590), .A2(n14578), .A3(n15625), .ZN(n14482) );
  NAND3_X1 U17965 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(n14482), .ZN(n15614) );
  NOR2_X1 U17966 ( .A1(n20702), .A2(n15614), .ZN(n14560) );
  AND2_X1 U17967 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n14560), .ZN(n14547) );
  NAND2_X1 U17968 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n14547), .ZN(n14483) );
  NOR2_X1 U17969 ( .A1(n14483), .A2(n19845), .ZN(n14525) );
  NAND3_X1 U17970 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .A3(n14525), .ZN(n14508) );
  INV_X1 U17971 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14509) );
  AND2_X1 U17972 ( .A1(n14483), .A2(n19853), .ZN(n14546) );
  INV_X1 U17973 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20707) );
  INV_X1 U17974 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20708) );
  NOR2_X1 U17975 ( .A1(n20707), .A2(n20708), .ZN(n14526) );
  NOR2_X1 U17976 ( .A1(n19845), .A2(n14526), .ZN(n14529) );
  NOR3_X1 U17977 ( .A1(n10076), .A2(n14529), .A3(n14509), .ZN(n14501) );
  AOI21_X1 U17978 ( .B1(n14508), .B2(n14509), .A(n14501), .ZN(n14484) );
  AOI211_X1 U17979 ( .C1(n14878), .C2(n19863), .A(n14485), .B(n14484), .ZN(
        n14486) );
  OAI21_X1 U17980 ( .B1(n14474), .B2(n15629), .A(n14486), .ZN(P1_U2811) );
  OAI22_X1 U17981 ( .A1(n15716), .A2(n14745), .B1(n15728), .B2(n14487), .ZN(
        n14488) );
  AOI21_X1 U17982 ( .B1(n15720), .B2(DATAI_29_), .A(n14488), .ZN(n14490) );
  NAND2_X1 U17983 ( .A1(n14731), .A2(BUF1_REG_29__SCAN_IN), .ZN(n14489) );
  OAI211_X1 U17984 ( .C1(n14474), .C2(n14740), .A(n14490), .B(n14489), .ZN(
        P1_U2875) );
  NAND2_X1 U17985 ( .A1(n14491), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n14493)
         );
  NAND3_X1 U17986 ( .A1(n14493), .A2(n14492), .A3(n19754), .ZN(P1_U2801) );
  AOI22_X1 U17987 ( .A1(n14497), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13069), .ZN(n14498) );
  AOI21_X1 U17988 ( .B1(n14501), .B2(P1_REIP_REG_30__SCAN_IN), .A(n15641), 
        .ZN(n14513) );
  INV_X1 U17989 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14507) );
  NOR4_X1 U17990 ( .A1(n14509), .A2(n14507), .A3(P1_REIP_REG_31__SCAN_IN), 
        .A4(n14508), .ZN(n14502) );
  AOI21_X1 U17991 ( .B1(n19837), .B2(P1_EBX_REG_31__SCAN_IN), .A(n14502), .ZN(
        n14503) );
  OAI21_X1 U17992 ( .B1(n19840), .B2(n14504), .A(n14503), .ZN(n14505) );
  AOI21_X1 U17993 ( .B1(n14513), .B2(P1_REIP_REG_31__SCAN_IN), .A(n14505), 
        .ZN(n14506) );
  NAND2_X1 U17994 ( .A1(n14754), .A2(n19821), .ZN(n14515) );
  OAI21_X1 U17995 ( .B1(n14509), .B2(n14508), .A(n14507), .ZN(n14512) );
  AOI22_X1 U17996 ( .A1(n19858), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n19837), .ZN(n14510) );
  OAI21_X1 U17997 ( .B1(n19851), .B2(n14748), .A(n14510), .ZN(n14511) );
  AOI21_X1 U17998 ( .B1(n14513), .B2(n14512), .A(n14511), .ZN(n14514) );
  OAI211_X1 U17999 ( .C1(n19791), .C2(n14516), .A(n14515), .B(n14514), .ZN(
        P1_U2810) );
  AOI21_X1 U18000 ( .B1(n14517), .B2(n14518), .A(n12836), .ZN(n14770) );
  INV_X1 U18001 ( .A(n14770), .ZN(n14695) );
  OR2_X1 U18002 ( .A1(n14538), .A2(n14519), .ZN(n14520) );
  NAND2_X1 U18003 ( .A1(n14521), .A2(n14520), .ZN(n14893) );
  AOI22_X1 U18004 ( .A1(n19858), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n19837), .B2(P1_EBX_REG_28__SCAN_IN), .ZN(n14524) );
  INV_X1 U18005 ( .A(n14522), .ZN(n14766) );
  NAND2_X1 U18006 ( .A1(n19865), .A2(n14766), .ZN(n14523) );
  OAI211_X1 U18007 ( .C1(n14893), .C2(n19791), .A(n14524), .B(n14523), .ZN(
        n14528) );
  INV_X1 U18008 ( .A(n14525), .ZN(n14537) );
  NOR3_X1 U18009 ( .A1(n14537), .A2(n14526), .A3(n20708), .ZN(n14527) );
  NOR2_X1 U18010 ( .A1(n14528), .A2(n14527), .ZN(n14531) );
  OAI21_X1 U18011 ( .B1(n10076), .B2(n14529), .A(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14530) );
  OAI211_X1 U18012 ( .C1(n14695), .C2(n15629), .A(n14531), .B(n14530), .ZN(
        P1_U2812) );
  INV_X1 U18013 ( .A(n14517), .ZN(n14533) );
  AOI21_X1 U18014 ( .B1(n14534), .B2(n14544), .A(n14533), .ZN(n14781) );
  INV_X1 U18015 ( .A(n14781), .ZN(n14700) );
  NAND2_X1 U18016 ( .A1(n19858), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14536) );
  AOI22_X1 U18017 ( .A1(n19837), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_REIP_REG_27__SCAN_IN), .B2(n10076), .ZN(n14535) );
  OAI211_X1 U18018 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14537), .A(n14536), 
        .B(n14535), .ZN(n14541) );
  AOI21_X1 U18019 ( .B1(n14539), .B2(n14550), .A(n14538), .ZN(n14902) );
  INV_X1 U18020 ( .A(n14902), .ZN(n14600) );
  NOR2_X1 U18021 ( .A1(n14600), .A2(n19791), .ZN(n14540) );
  AOI211_X1 U18022 ( .C1(n19865), .C2(n14777), .A(n14541), .B(n14540), .ZN(
        n14542) );
  OAI21_X1 U18023 ( .B1(n14700), .B2(n15629), .A(n14542), .ZN(P1_U2813) );
  AOI21_X1 U18024 ( .B1(n14545), .B2(n14543), .A(n14532), .ZN(n14790) );
  INV_X1 U18025 ( .A(n14790), .ZN(n14705) );
  AOI22_X1 U18026 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n10076), .B1(n14547), 
        .B2(n14546), .ZN(n14556) );
  NAND2_X1 U18027 ( .A1(n14565), .A2(n14548), .ZN(n14549) );
  NAND2_X1 U18028 ( .A1(n14550), .A2(n14549), .ZN(n14909) );
  AOI22_X1 U18029 ( .A1(n19858), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n19837), .B2(P1_EBX_REG_26__SCAN_IN), .ZN(n14553) );
  INV_X1 U18030 ( .A(n14551), .ZN(n14786) );
  NAND2_X1 U18031 ( .A1(n19865), .A2(n14786), .ZN(n14552) );
  OAI211_X1 U18032 ( .C1(n14909), .C2(n19791), .A(n14553), .B(n14552), .ZN(
        n14554) );
  INV_X1 U18033 ( .A(n14554), .ZN(n14555) );
  OAI211_X1 U18034 ( .C1(n14705), .C2(n15629), .A(n14556), .B(n14555), .ZN(
        P1_U2814) );
  OAI21_X1 U18035 ( .B1(n14557), .B2(n14558), .A(n14543), .ZN(n14797) );
  INV_X1 U18036 ( .A(n14797), .ZN(n14570) );
  AOI22_X1 U18037 ( .A1(n19865), .A2(n14800), .B1(n19837), .B2(
        P1_EBX_REG_25__SCAN_IN), .ZN(n14562) );
  INV_X1 U18038 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14559) );
  NAND3_X1 U18039 ( .A1(n19853), .A2(n14560), .A3(n14559), .ZN(n14561) );
  OAI211_X1 U18040 ( .C1(n19840), .C2(n14796), .A(n14562), .B(n14561), .ZN(
        n14569) );
  OR2_X1 U18041 ( .A1(n14609), .A2(n14563), .ZN(n14564) );
  NAND2_X1 U18042 ( .A1(n14565), .A2(n14564), .ZN(n14920) );
  NAND2_X1 U18043 ( .A1(n19853), .A2(n15614), .ZN(n14566) );
  NAND2_X1 U18044 ( .A1(n19773), .A2(n14566), .ZN(n15626) );
  NOR2_X1 U18045 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n19845), .ZN(n15615) );
  OAI21_X1 U18046 ( .B1(n15626), .B2(n15615), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14567) );
  OAI21_X1 U18047 ( .B1(n14920), .B2(n19791), .A(n14567), .ZN(n14568) );
  AOI211_X1 U18048 ( .C1(n14570), .C2(n19821), .A(n14569), .B(n14568), .ZN(
        n14571) );
  INV_X1 U18049 ( .A(n14571), .ZN(P1_U2815) );
  INV_X1 U18050 ( .A(n14572), .ZN(n14575) );
  INV_X1 U18051 ( .A(n14573), .ZN(n14642) );
  INV_X1 U18052 ( .A(n14574), .ZN(n14638) );
  AOI21_X1 U18053 ( .B1(n14576), .B2(n14647), .A(n14634), .ZN(n15804) );
  INV_X1 U18054 ( .A(n19837), .ZN(n19856) );
  NAND2_X1 U18055 ( .A1(n19865), .A2(n14824), .ZN(n14582) );
  INV_X1 U18056 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14821) );
  NOR2_X1 U18057 ( .A1(n14578), .A2(n14577), .ZN(n15669) );
  NAND2_X1 U18058 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15669), .ZN(n15659) );
  INV_X1 U18059 ( .A(n15659), .ZN(n14580) );
  OAI21_X1 U18060 ( .B1(n19840), .B2(n14822), .A(n19777), .ZN(n14579) );
  AOI21_X1 U18061 ( .B1(n14821), .B2(n14580), .A(n14579), .ZN(n14581) );
  OAI211_X1 U18062 ( .C1(n14583), .C2(n19856), .A(n14582), .B(n14581), .ZN(
        n14584) );
  AOI21_X1 U18063 ( .B1(n15804), .B2(n19863), .A(n14584), .ZN(n14587) );
  INV_X1 U18064 ( .A(n15669), .ZN(n15644) );
  OAI22_X1 U18065 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15644), .B1(n15641), 
        .B2(n15643), .ZN(n14585) );
  NAND2_X1 U18066 ( .A1(n14585), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n14586) );
  OAI211_X1 U18067 ( .C1(n14827), .C2(n15629), .A(n14587), .B(n14586), .ZN(
        P1_U2821) );
  INV_X1 U18068 ( .A(n14651), .ZN(n14588) );
  AOI21_X1 U18069 ( .B1(n14589), .B2(n14666), .A(n14588), .ZN(n14858) );
  INV_X1 U18070 ( .A(n14858), .ZN(n14741) );
  AOI21_X1 U18071 ( .B1(n19853), .B2(n14590), .A(n19803), .ZN(n15690) );
  AOI22_X1 U18072 ( .A1(n19858), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n19837), .B2(P1_EBX_REG_15__SCAN_IN), .ZN(n14591) );
  OAI211_X1 U18073 ( .C1(n14593), .C2(n15690), .A(n14591), .B(n19777), .ZN(
        n14592) );
  AOI21_X1 U18074 ( .B1(n15673), .B2(n14593), .A(n14592), .ZN(n14598) );
  OAI21_X1 U18075 ( .B1(n14171), .B2(n14667), .A(n14594), .ZN(n14595) );
  AND2_X1 U18076 ( .A1(n14595), .A2(n14655), .ZN(n15827) );
  INV_X1 U18077 ( .A(n14856), .ZN(n14596) );
  AOI22_X1 U18078 ( .A1(n15827), .A2(n19863), .B1(n19865), .B2(n14596), .ZN(
        n14597) );
  OAI211_X1 U18079 ( .C1(n14741), .C2(n15629), .A(n14598), .B(n14597), .ZN(
        P1_U2825) );
  INV_X1 U18080 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14599) );
  OAI22_X1 U18081 ( .A1(n14867), .A2(n14684), .B1(n14682), .B2(n14599), .ZN(
        P1_U2841) );
  INV_X1 U18082 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n21059) );
  OAI222_X1 U18083 ( .A1(n14672), .A2(n14695), .B1(n21059), .B2(n14682), .C1(
        n14893), .C2(n14684), .ZN(P1_U2844) );
  INV_X1 U18084 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14601) );
  OAI222_X1 U18085 ( .A1(n14672), .A2(n14700), .B1(n14682), .B2(n14601), .C1(
        n14600), .C2(n14684), .ZN(P1_U2845) );
  OAI222_X1 U18086 ( .A1(n14672), .A2(n14705), .B1(n14602), .B2(n14682), .C1(
        n14909), .C2(n14684), .ZN(P1_U2846) );
  INV_X1 U18087 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14603) );
  OAI222_X1 U18088 ( .A1(n14672), .A2(n14797), .B1(n14603), .B2(n14682), .C1(
        n14920), .C2(n14684), .ZN(P1_U2847) );
  NOR2_X1 U18089 ( .A1(n14604), .A2(n14605), .ZN(n14606) );
  OR2_X1 U18090 ( .A1(n14557), .A2(n14606), .ZN(n14806) );
  NOR2_X1 U18091 ( .A1(n14616), .A2(n14607), .ZN(n14608) );
  OR2_X1 U18092 ( .A1(n14609), .A2(n14608), .ZN(n15619) );
  OAI22_X1 U18093 ( .A1(n15619), .A2(n14684), .B1(n14610), .B2(n14682), .ZN(
        n14611) );
  INV_X1 U18094 ( .A(n14611), .ZN(n14612) );
  OAI21_X1 U18095 ( .B1(n14806), .B2(n14672), .A(n14612), .ZN(P1_U2848) );
  AOI21_X1 U18096 ( .B1(n14614), .B2(n14613), .A(n14604), .ZN(n14615) );
  INV_X1 U18097 ( .A(n14615), .ZN(n15630) );
  AOI21_X1 U18098 ( .B1(n14617), .B2(n14624), .A(n14616), .ZN(n15798) );
  AOI22_X1 U18099 ( .A1(n15798), .A2(n14670), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n14669), .ZN(n14618) );
  OAI21_X1 U18100 ( .B1(n15630), .B2(n14672), .A(n14618), .ZN(P1_U2849) );
  NAND2_X1 U18101 ( .A1(n14619), .A2(n14620), .ZN(n14621) );
  NAND2_X1 U18102 ( .A1(n14628), .A2(n14622), .ZN(n14623) );
  NAND2_X1 U18103 ( .A1(n14624), .A2(n14623), .ZN(n15648) );
  OAI22_X1 U18104 ( .A1(n15648), .A2(n14684), .B1(n14625), .B2(n14682), .ZN(
        n14626) );
  AOI21_X1 U18105 ( .B1(n15730), .B2(n14660), .A(n14626), .ZN(n14627) );
  INV_X1 U18106 ( .A(n14627), .ZN(P1_U2850) );
  OAI21_X1 U18107 ( .B1(n14636), .B2(n14629), .A(n14628), .ZN(n15592) );
  INV_X1 U18108 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14632) );
  OAI21_X1 U18109 ( .B1(n14630), .B2(n14631), .A(n14619), .ZN(n15649) );
  OAI222_X1 U18110 ( .A1(n15592), .A2(n14684), .B1(n14632), .B2(n14682), .C1(
        n15649), .C2(n14672), .ZN(P1_U2851) );
  NOR2_X1 U18111 ( .A1(n14634), .A2(n14633), .ZN(n14635) );
  OR2_X1 U18112 ( .A1(n14636), .A2(n14635), .ZN(n15664) );
  INV_X1 U18113 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15657) );
  INV_X1 U18114 ( .A(n14637), .ZN(n14639) );
  AOI21_X1 U18115 ( .B1(n14639), .B2(n14638), .A(n14630), .ZN(n15740) );
  INV_X1 U18116 ( .A(n15740), .ZN(n14640) );
  OAI222_X1 U18117 ( .A1(n14684), .A2(n15664), .B1(n15657), .B2(n14682), .C1(
        n14640), .C2(n14672), .ZN(P1_U2852) );
  AOI22_X1 U18118 ( .A1(n15804), .A2(n14670), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14669), .ZN(n14641) );
  OAI21_X1 U18119 ( .B1(n14827), .B2(n14672), .A(n14641), .ZN(P1_U2853) );
  AOI21_X1 U18120 ( .B1(n14643), .B2(n14071), .A(n14642), .ZN(n15670) );
  NAND2_X1 U18121 ( .A1(n14645), .A2(n14644), .ZN(n14646) );
  NAND2_X1 U18122 ( .A1(n14647), .A2(n14646), .ZN(n15811) );
  OAI22_X1 U18123 ( .A1(n15811), .A2(n14684), .B1(n20872), .B2(n14682), .ZN(
        n14648) );
  AOI21_X1 U18124 ( .B1(n15670), .B2(n14660), .A(n14648), .ZN(n14649) );
  INV_X1 U18125 ( .A(n14649), .ZN(P1_U2854) );
  AND2_X1 U18126 ( .A1(n14655), .A2(n14654), .ZN(n14657) );
  OR2_X1 U18127 ( .A1(n14657), .A2(n14656), .ZN(n15684) );
  OAI22_X1 U18128 ( .A1(n15684), .A2(n14684), .B1(n14658), .B2(n14682), .ZN(
        n14659) );
  AOI21_X1 U18129 ( .B1(n15745), .B2(n14660), .A(n14659), .ZN(n14661) );
  INV_X1 U18130 ( .A(n14661), .ZN(P1_U2856) );
  AOI22_X1 U18131 ( .A1(n15827), .A2(n14670), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14669), .ZN(n14662) );
  OAI21_X1 U18132 ( .B1(n14741), .B2(n14672), .A(n14662), .ZN(P1_U2857) );
  NAND2_X1 U18133 ( .A1(n14664), .A2(n14663), .ZN(n14665) );
  INV_X1 U18134 ( .A(n14667), .ZN(n14668) );
  XNOR2_X1 U18135 ( .A(n14171), .B(n14668), .ZN(n15834) );
  AOI22_X1 U18136 ( .A1(n15834), .A2(n14670), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n14669), .ZN(n14671) );
  OAI21_X1 U18137 ( .B1(n14743), .B2(n14672), .A(n14671), .ZN(P1_U2858) );
  NOR2_X1 U18138 ( .A1(n14674), .A2(n14673), .ZN(n14675) );
  OR2_X1 U18139 ( .A1(n14172), .A2(n14675), .ZN(n15860) );
  INV_X1 U18140 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14683) );
  INV_X1 U18141 ( .A(n14676), .ZN(n14680) );
  INV_X1 U18142 ( .A(n14677), .ZN(n14679) );
  INV_X1 U18143 ( .A(n15761), .ZN(n14681) );
  OAI222_X1 U18144 ( .A1(n15860), .A2(n14684), .B1(n14683), .B2(n14682), .C1(
        n14681), .C2(n14672), .ZN(P1_U2860) );
  INV_X1 U18145 ( .A(DATAI_14_), .ZN(n14686) );
  MUX2_X1 U18146 ( .A(n14686), .B(n14685), .S(n19976), .Z(n19913) );
  OAI22_X1 U18147 ( .A1(n15716), .A2(n19913), .B1(n15728), .B2(n13194), .ZN(
        n14687) );
  AOI21_X1 U18148 ( .B1(n15720), .B2(DATAI_30_), .A(n14687), .ZN(n14689) );
  NAND2_X1 U18149 ( .A1(n14731), .A2(BUF1_REG_30__SCAN_IN), .ZN(n14688) );
  OAI211_X1 U18150 ( .C1(n14690), .C2(n14740), .A(n14689), .B(n14688), .ZN(
        P1_U2874) );
  INV_X1 U18151 ( .A(DATAI_12_), .ZN(n20966) );
  MUX2_X1 U18152 ( .A(n20966), .B(n16294), .S(n19976), .Z(n15724) );
  OAI22_X1 U18153 ( .A1(n15716), .A2(n15724), .B1(n15728), .B2(n14691), .ZN(
        n14692) );
  AOI21_X1 U18154 ( .B1(n15720), .B2(DATAI_28_), .A(n14692), .ZN(n14694) );
  NAND2_X1 U18155 ( .A1(n14731), .A2(BUF1_REG_28__SCAN_IN), .ZN(n14693) );
  OAI211_X1 U18156 ( .C1(n14695), .C2(n14740), .A(n14694), .B(n14693), .ZN(
        P1_U2876) );
  OAI22_X1 U18157 ( .A1(n15716), .A2(n19908), .B1(n15728), .B2(n14696), .ZN(
        n14697) );
  AOI21_X1 U18158 ( .B1(n15720), .B2(DATAI_27_), .A(n14697), .ZN(n14699) );
  NAND2_X1 U18159 ( .A1(n14731), .A2(BUF1_REG_27__SCAN_IN), .ZN(n14698) );
  OAI211_X1 U18160 ( .C1(n14700), .C2(n14740), .A(n14699), .B(n14698), .ZN(
        P1_U2877) );
  OAI22_X1 U18161 ( .A1(n15716), .A2(n19905), .B1(n15728), .B2(n14701), .ZN(
        n14702) );
  AOI21_X1 U18162 ( .B1(n15720), .B2(DATAI_26_), .A(n14702), .ZN(n14704) );
  NAND2_X1 U18163 ( .A1(n14731), .A2(BUF1_REG_26__SCAN_IN), .ZN(n14703) );
  OAI211_X1 U18164 ( .C1(n14705), .C2(n14740), .A(n14704), .B(n14703), .ZN(
        P1_U2878) );
  INV_X1 U18165 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14706) );
  OAI22_X1 U18166 ( .A1(n15716), .A2(n19902), .B1(n15728), .B2(n14706), .ZN(
        n14707) );
  AOI21_X1 U18167 ( .B1(n15720), .B2(DATAI_25_), .A(n14707), .ZN(n14709) );
  NAND2_X1 U18168 ( .A1(n14731), .A2(BUF1_REG_25__SCAN_IN), .ZN(n14708) );
  OAI211_X1 U18169 ( .C1(n14797), .C2(n14740), .A(n14709), .B(n14708), .ZN(
        P1_U2879) );
  OAI22_X1 U18170 ( .A1(n15716), .A2(n19899), .B1(n15728), .B2(n14710), .ZN(
        n14711) );
  AOI21_X1 U18171 ( .B1(n15720), .B2(DATAI_24_), .A(n14711), .ZN(n14713) );
  NAND2_X1 U18172 ( .A1(n14731), .A2(BUF1_REG_24__SCAN_IN), .ZN(n14712) );
  OAI211_X1 U18173 ( .C1(n14806), .C2(n14740), .A(n14713), .B(n14712), .ZN(
        P1_U2880) );
  OAI22_X1 U18174 ( .A1(n15716), .A2(n20017), .B1(n15728), .B2(n13196), .ZN(
        n14714) );
  AOI21_X1 U18175 ( .B1(n15720), .B2(DATAI_23_), .A(n14714), .ZN(n14716) );
  NAND2_X1 U18176 ( .A1(n14731), .A2(BUF1_REG_23__SCAN_IN), .ZN(n14715) );
  OAI211_X1 U18177 ( .C1(n15630), .C2(n14740), .A(n14716), .B(n14715), .ZN(
        P1_U2881) );
  INV_X1 U18178 ( .A(n15730), .ZN(n14721) );
  OAI22_X1 U18179 ( .A1(n15716), .A2(n20010), .B1(n15728), .B2(n14717), .ZN(
        n14718) );
  AOI21_X1 U18180 ( .B1(n15720), .B2(DATAI_22_), .A(n14718), .ZN(n14720) );
  NAND2_X1 U18181 ( .A1(n14731), .A2(BUF1_REG_22__SCAN_IN), .ZN(n14719) );
  OAI211_X1 U18182 ( .C1(n14721), .C2(n14740), .A(n14720), .B(n14719), .ZN(
        P1_U2882) );
  INV_X1 U18183 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14722) );
  OAI22_X1 U18184 ( .A1(n15716), .A2(n20007), .B1(n15728), .B2(n14722), .ZN(
        n14723) );
  AOI21_X1 U18185 ( .B1(n15720), .B2(DATAI_21_), .A(n14723), .ZN(n14725) );
  NAND2_X1 U18186 ( .A1(n14731), .A2(BUF1_REG_21__SCAN_IN), .ZN(n14724) );
  OAI211_X1 U18187 ( .C1(n15649), .C2(n14740), .A(n14725), .B(n14724), .ZN(
        P1_U2883) );
  OAI22_X1 U18188 ( .A1(n15716), .A2(n20000), .B1(n15728), .B2(n13192), .ZN(
        n14726) );
  AOI21_X1 U18189 ( .B1(n15720), .B2(DATAI_19_), .A(n14726), .ZN(n14728) );
  NAND2_X1 U18190 ( .A1(n14731), .A2(BUF1_REG_19__SCAN_IN), .ZN(n14727) );
  OAI211_X1 U18191 ( .C1(n14827), .C2(n14740), .A(n14728), .B(n14727), .ZN(
        P1_U2885) );
  INV_X1 U18192 ( .A(n15670), .ZN(n14734) );
  OAI22_X1 U18193 ( .A1(n15716), .A2(n19997), .B1(n15728), .B2(n14729), .ZN(
        n14730) );
  AOI21_X1 U18194 ( .B1(n15720), .B2(DATAI_18_), .A(n14730), .ZN(n14733) );
  NAND2_X1 U18195 ( .A1(n14731), .A2(BUF1_REG_18__SCAN_IN), .ZN(n14732) );
  OAI211_X1 U18196 ( .C1(n14734), .C2(n14740), .A(n14733), .B(n14732), .ZN(
        P1_U2886) );
  INV_X1 U18197 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n14738) );
  NAND2_X1 U18198 ( .A1(n15745), .A2(n15726), .ZN(n14737) );
  OAI22_X1 U18199 ( .A1(n15716), .A2(n19985), .B1(n15728), .B2(n12088), .ZN(
        n14735) );
  AOI21_X1 U18200 ( .B1(n15720), .B2(DATAI_16_), .A(n14735), .ZN(n14736) );
  OAI211_X1 U18201 ( .C1(n15723), .C2(n14738), .A(n14737), .B(n14736), .ZN(
        P1_U2888) );
  OAI222_X1 U18202 ( .A1(n14741), .A2(n14740), .B1(n15728), .B2(n13261), .C1(
        n14744), .C2(n14739), .ZN(P1_U2889) );
  INV_X1 U18203 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14742) );
  OAI222_X1 U18204 ( .A1(n14743), .A2(n14747), .B1(n19913), .B2(n14744), .C1(
        n14742), .C2(n15728), .ZN(P1_U2890) );
  OAI222_X1 U18205 ( .A1(n14747), .A2(n14746), .B1(n14745), .B2(n14744), .C1(
        n15728), .C2(n12062), .ZN(P1_U2891) );
  INV_X1 U18206 ( .A(n14748), .ZN(n14749) );
  NAND2_X1 U18207 ( .A1(n15791), .A2(n14749), .ZN(n14751) );
  OAI211_X1 U18208 ( .C1(n14752), .C2(n15795), .A(n14751), .B(n14750), .ZN(
        n14753) );
  AOI21_X1 U18209 ( .B1(n14754), .B2(n12940), .A(n14753), .ZN(n14755) );
  OAI21_X1 U18210 ( .B1(n14756), .B2(n19757), .A(n14755), .ZN(P1_U2969) );
  NAND2_X1 U18211 ( .A1(n15766), .A2(n14907), .ZN(n14758) );
  NAND2_X1 U18212 ( .A1(n14757), .A2(n14758), .ZN(n14762) );
  NAND2_X1 U18213 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14759) );
  NOR2_X1 U18214 ( .A1(n14762), .A2(n14759), .ZN(n14764) );
  NOR4_X1 U18215 ( .A1(n14760), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14761) );
  AND2_X1 U18216 ( .A1(n14762), .A2(n14761), .ZN(n14763) );
  MUX2_X1 U18217 ( .A(n14764), .B(n14763), .S(n10088), .Z(n14765) );
  XNOR2_X1 U18218 ( .A(n14765), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14897) );
  NAND2_X1 U18219 ( .A1(n15791), .A2(n14766), .ZN(n14767) );
  NAND2_X1 U18220 ( .A1(n19939), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14892) );
  OAI211_X1 U18221 ( .C1(n14768), .C2(n15795), .A(n14767), .B(n14892), .ZN(
        n14769) );
  AOI21_X1 U18222 ( .B1(n14770), .B2(n12940), .A(n14769), .ZN(n14771) );
  OAI21_X1 U18223 ( .B1(n19757), .B2(n14897), .A(n14771), .ZN(P1_U2971) );
  NAND2_X1 U18224 ( .A1(n12832), .A2(n10088), .ZN(n14774) );
  NAND2_X1 U18225 ( .A1(n14772), .A2(n15766), .ZN(n14773) );
  XNOR2_X1 U18226 ( .A(n14776), .B(n14775), .ZN(n14905) );
  INV_X1 U18227 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14779) );
  NAND2_X1 U18228 ( .A1(n15791), .A2(n14777), .ZN(n14778) );
  NAND2_X1 U18229 ( .A1(n19939), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14899) );
  OAI211_X1 U18230 ( .C1(n14779), .C2(n15795), .A(n14778), .B(n14899), .ZN(
        n14780) );
  AOI21_X1 U18231 ( .B1(n14781), .B2(n12940), .A(n14780), .ZN(n14782) );
  OAI21_X1 U18232 ( .B1(n14905), .B2(n19757), .A(n14782), .ZN(P1_U2972) );
  INV_X1 U18233 ( .A(n14757), .ZN(n14802) );
  OAI21_X1 U18234 ( .B1(n14802), .B2(n14907), .A(n15766), .ZN(n14783) );
  NAND2_X1 U18235 ( .A1(n14784), .A2(n14783), .ZN(n14785) );
  XNOR2_X1 U18236 ( .A(n14785), .B(n14906), .ZN(n14914) );
  NAND2_X1 U18237 ( .A1(n15791), .A2(n14786), .ZN(n14787) );
  NAND2_X1 U18238 ( .A1(n19939), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14908) );
  OAI211_X1 U18239 ( .C1(n15795), .C2(n14788), .A(n14787), .B(n14908), .ZN(
        n14789) );
  AOI21_X1 U18240 ( .B1(n14790), .B2(n12940), .A(n14789), .ZN(n14791) );
  OAI21_X1 U18241 ( .B1(n19757), .B2(n14914), .A(n14791), .ZN(P1_U2973) );
  NAND2_X1 U18242 ( .A1(n14792), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14803) );
  MUX2_X1 U18243 ( .A(n14929), .B(n14793), .S(n10088), .Z(n14794) );
  AOI21_X1 U18244 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14803), .A(
        n14794), .ZN(n14795) );
  XNOR2_X1 U18245 ( .A(n14795), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14924) );
  NAND2_X1 U18246 ( .A1(n19939), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14919) );
  OAI21_X1 U18247 ( .B1(n15795), .B2(n14796), .A(n14919), .ZN(n14799) );
  NOR2_X1 U18248 ( .A1(n14797), .A2(n19975), .ZN(n14798) );
  AOI211_X1 U18249 ( .C1(n15791), .C2(n14800), .A(n14799), .B(n14798), .ZN(
        n14801) );
  OAI21_X1 U18250 ( .B1(n19757), .B2(n14924), .A(n14801), .ZN(P1_U2974) );
  NAND2_X1 U18251 ( .A1(n14802), .A2(n10088), .ZN(n14804) );
  MUX2_X1 U18252 ( .A(n10088), .B(n14804), .S(n14803), .Z(n14805) );
  XNOR2_X1 U18253 ( .A(n14805), .B(n14929), .ZN(n14934) );
  INV_X1 U18254 ( .A(n14806), .ZN(n15621) );
  INV_X1 U18255 ( .A(n15623), .ZN(n14807) );
  NAND2_X1 U18256 ( .A1(n15791), .A2(n14807), .ZN(n14808) );
  NAND2_X1 U18257 ( .A1(n19939), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14925) );
  OAI211_X1 U18258 ( .C1(n15795), .C2(n14809), .A(n14808), .B(n14925), .ZN(
        n14810) );
  AOI21_X1 U18259 ( .B1(n15621), .B2(n12940), .A(n14810), .ZN(n14811) );
  OAI21_X1 U18260 ( .B1(n14934), .B2(n19757), .A(n14811), .ZN(P1_U2975) );
  XNOR2_X1 U18261 ( .A(n15766), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14812) );
  XNOR2_X1 U18262 ( .A(n14757), .B(n14812), .ZN(n15797) );
  INV_X1 U18263 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14813) );
  OAI22_X1 U18264 ( .A1(n15795), .A2(n15634), .B1(n15908), .B2(n14813), .ZN(
        n14815) );
  NOR2_X1 U18265 ( .A1(n15630), .A2(n19975), .ZN(n14814) );
  AOI211_X1 U18266 ( .C1(n15791), .C2(n15624), .A(n14815), .B(n14814), .ZN(
        n14816) );
  OAI21_X1 U18267 ( .B1(n15797), .B2(n19757), .A(n14816), .ZN(P1_U2976) );
  MUX2_X1 U18268 ( .A(n11556), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .S(
        n9737), .Z(n14819) );
  NAND2_X1 U18269 ( .A1(n15766), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14946) );
  INV_X1 U18270 ( .A(n14817), .ZN(n14818) );
  AOI21_X1 U18271 ( .B1(n10088), .B2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n14818), .ZN(n15588) );
  MUX2_X1 U18272 ( .A(n14819), .B(n14946), .S(n15588), .Z(n14820) );
  NAND3_X1 U18273 ( .A1(n15588), .A2(n10088), .A3(n11556), .ZN(n15589) );
  NAND2_X1 U18274 ( .A1(n14820), .A2(n15589), .ZN(n15805) );
  NAND2_X1 U18275 ( .A1(n15805), .A2(n19938), .ZN(n14826) );
  OAI22_X1 U18276 ( .A1(n15795), .A2(n14822), .B1(n15908), .B2(n14821), .ZN(
        n14823) );
  AOI21_X1 U18277 ( .B1(n15791), .B2(n14824), .A(n14823), .ZN(n14825) );
  OAI211_X1 U18278 ( .C1(n19975), .C2(n14827), .A(n14826), .B(n14825), .ZN(
        P1_U2980) );
  OAI21_X1 U18279 ( .B1(n11555), .B2(n14828), .A(n14817), .ZN(n15812) );
  AOI22_X1 U18280 ( .A1(n19936), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n19953), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14829) );
  OAI21_X1 U18281 ( .B1(n15787), .B2(n15667), .A(n14829), .ZN(n14830) );
  AOI21_X1 U18282 ( .B1(n15670), .B2(n12940), .A(n14830), .ZN(n14831) );
  OAI21_X1 U18283 ( .B1(n19757), .B2(n15812), .A(n14831), .ZN(P1_U2981) );
  NAND2_X1 U18284 ( .A1(n10088), .A2(n14832), .ZN(n14837) );
  NOR2_X1 U18285 ( .A1(n10047), .A2(n14833), .ZN(n14848) );
  AOI21_X1 U18286 ( .B1(n14848), .B2(n14835), .A(n14834), .ZN(n14836) );
  MUX2_X1 U18287 ( .A(n14837), .B(n10088), .S(n14836), .Z(n14839) );
  INV_X1 U18288 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14838) );
  XNOR2_X1 U18289 ( .A(n14839), .B(n14838), .ZN(n15818) );
  INV_X1 U18290 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14840) );
  OAI22_X1 U18291 ( .A1(n15795), .A2(n14841), .B1(n15908), .B2(n14840), .ZN(
        n14844) );
  NOR2_X1 U18292 ( .A1(n14842), .A2(n19975), .ZN(n14843) );
  AOI211_X1 U18293 ( .C1(n15791), .C2(n14845), .A(n14844), .B(n14843), .ZN(
        n14846) );
  OAI21_X1 U18294 ( .B1(n19757), .B2(n15818), .A(n14846), .ZN(P1_U2982) );
  NOR2_X1 U18295 ( .A1(n15750), .A2(n14849), .ZN(n14958) );
  INV_X1 U18296 ( .A(n14958), .ZN(n14851) );
  NAND2_X1 U18297 ( .A1(n14851), .A2(n14850), .ZN(n14854) );
  NAND2_X1 U18298 ( .A1(n14852), .A2(n14957), .ZN(n14853) );
  XNOR2_X1 U18299 ( .A(n14854), .B(n14853), .ZN(n15828) );
  INV_X1 U18300 ( .A(n15828), .ZN(n14860) );
  AOI22_X1 U18301 ( .A1(n19936), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n19953), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n14855) );
  OAI21_X1 U18302 ( .B1(n15787), .B2(n14856), .A(n14855), .ZN(n14857) );
  AOI21_X1 U18303 ( .B1(n14858), .B2(n12940), .A(n14857), .ZN(n14859) );
  OAI21_X1 U18304 ( .B1(n14860), .B2(n19757), .A(n14859), .ZN(P1_U2984) );
  MUX2_X1 U18305 ( .A(n15765), .B(n14861), .S(n10088), .Z(n14862) );
  XOR2_X1 U18306 ( .A(n11696), .B(n14862), .Z(n15890) );
  INV_X1 U18307 ( .A(n15890), .ZN(n14866) );
  AOI22_X1 U18308 ( .A1(n19936), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n19939), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14863) );
  OAI21_X1 U18309 ( .B1(n15787), .B2(n15709), .A(n14863), .ZN(n14864) );
  AOI21_X1 U18310 ( .B1(n15711), .B2(n12940), .A(n14864), .ZN(n14865) );
  OAI21_X1 U18311 ( .B1(n14866), .B2(n19757), .A(n14865), .ZN(P1_U2989) );
  INV_X1 U18312 ( .A(n14867), .ZN(n14874) );
  NAND2_X1 U18313 ( .A1(n20933), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14871) );
  NAND3_X1 U18314 ( .A1(n14868), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15882), .ZN(n14870) );
  OAI211_X1 U18315 ( .C1(n14872), .C2(n14871), .A(n14870), .B(n14869), .ZN(
        n14873) );
  AOI21_X1 U18316 ( .B1(n14874), .B2(n19964), .A(n14873), .ZN(n14875) );
  OAI21_X1 U18317 ( .B1(n14876), .B2(n15872), .A(n14875), .ZN(P1_U3000) );
  INV_X1 U18318 ( .A(n14877), .ZN(n14885) );
  INV_X1 U18319 ( .A(n14878), .ZN(n14883) );
  NAND3_X1 U18320 ( .A1(n14898), .A2(n14880), .A3(n14879), .ZN(n14881) );
  OAI211_X1 U18321 ( .C1(n14883), .C2(n15909), .A(n14882), .B(n14881), .ZN(
        n14884) );
  AOI21_X1 U18322 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n14885), .A(
        n14884), .ZN(n14886) );
  OAI21_X1 U18323 ( .B1(n14887), .B2(n15872), .A(n14886), .ZN(P1_U3002) );
  INV_X1 U18324 ( .A(n14888), .ZN(n14890) );
  NAND3_X1 U18325 ( .A1(n14898), .A2(n14890), .A3(n14889), .ZN(n14891) );
  OAI211_X1 U18326 ( .C1(n14893), .C2(n15909), .A(n14892), .B(n14891), .ZN(
        n14894) );
  INV_X1 U18327 ( .A(n14894), .ZN(n14896) );
  NAND3_X1 U18328 ( .A1(n14912), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15882), .ZN(n14895) );
  OAI211_X1 U18329 ( .C1(n14897), .C2(n15872), .A(n14896), .B(n14895), .ZN(
        P1_U3003) );
  INV_X1 U18330 ( .A(n14898), .ZN(n14900) );
  OAI21_X1 U18331 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14900), .A(
        n14899), .ZN(n14901) );
  AOI21_X1 U18332 ( .B1(n14902), .B2(n19964), .A(n14901), .ZN(n14904) );
  NAND3_X1 U18333 ( .A1(n14912), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15882), .ZN(n14903) );
  OAI211_X1 U18334 ( .C1(n14905), .C2(n15872), .A(n14904), .B(n14903), .ZN(
        P1_U3004) );
  OAI21_X1 U18335 ( .B1(n14907), .B2(n15802), .A(n14906), .ZN(n14911) );
  OAI21_X1 U18336 ( .B1(n14909), .B2(n15909), .A(n14908), .ZN(n14910) );
  AOI21_X1 U18337 ( .B1(n14912), .B2(n14911), .A(n14910), .ZN(n14913) );
  OAI21_X1 U18338 ( .B1(n14914), .B2(n15872), .A(n14913), .ZN(P1_U3005) );
  INV_X1 U18339 ( .A(n14915), .ZN(n14922) );
  NOR2_X1 U18340 ( .A1(n14929), .A2(n11559), .ZN(n14928) );
  NAND3_X1 U18341 ( .A1(n14917), .A2(n14928), .A3(n14916), .ZN(n14918) );
  OAI211_X1 U18342 ( .C1(n14920), .C2(n15909), .A(n14919), .B(n14918), .ZN(
        n14921) );
  AOI21_X1 U18343 ( .B1(n14922), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n14921), .ZN(n14923) );
  OAI21_X1 U18344 ( .B1(n14924), .B2(n15872), .A(n14923), .ZN(P1_U3006) );
  INV_X1 U18345 ( .A(n15619), .ZN(n14927) );
  INV_X1 U18346 ( .A(n14925), .ZN(n14926) );
  AOI21_X1 U18347 ( .B1(n14927), .B2(n19964), .A(n14926), .ZN(n14933) );
  AOI21_X1 U18348 ( .B1(n15900), .B2(n15865), .A(n14928), .ZN(n14931) );
  OAI21_X1 U18349 ( .B1(n11559), .B2(n15802), .A(n14929), .ZN(n14930) );
  OAI21_X1 U18350 ( .B1(n15796), .B2(n14931), .A(n14930), .ZN(n14932) );
  OAI211_X1 U18351 ( .C1(n14934), .C2(n15872), .A(n14933), .B(n14932), .ZN(
        P1_U3007) );
  INV_X1 U18352 ( .A(n15591), .ZN(n14945) );
  NAND2_X1 U18353 ( .A1(n14936), .A2(n14935), .ZN(n14937) );
  XNOR2_X1 U18354 ( .A(n14937), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15729) );
  NAND2_X1 U18355 ( .A1(n15729), .A2(n19965), .ZN(n14943) );
  AOI21_X1 U18356 ( .B1(n11557), .B2(n14944), .A(n14938), .ZN(n14941) );
  INV_X1 U18357 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14939) );
  OAI22_X1 U18358 ( .A1(n15648), .A2(n15909), .B1(n15908), .B2(n14939), .ZN(
        n14940) );
  AOI21_X1 U18359 ( .B1(n15593), .B2(n14941), .A(n14940), .ZN(n14942) );
  OAI211_X1 U18360 ( .C1(n14945), .C2(n14944), .A(n14943), .B(n14942), .ZN(
        P1_U3009) );
  OAI21_X1 U18361 ( .B1(n14817), .B2(n14946), .A(n15589), .ZN(n14948) );
  XNOR2_X1 U18362 ( .A(n14948), .B(n14947), .ZN(n15741) );
  INV_X1 U18363 ( .A(n15741), .ZN(n14955) );
  AOI21_X1 U18364 ( .B1(n15848), .B2(n14949), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14950) );
  OAI21_X1 U18365 ( .B1(n14950), .B2(n15803), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14954) );
  INV_X1 U18366 ( .A(n15664), .ZN(n14952) );
  NOR3_X1 U18367 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11556), .A3(
        n15808), .ZN(n14951) );
  INV_X1 U18368 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20698) );
  NOR2_X1 U18369 ( .A1(n15908), .A2(n20698), .ZN(n15739) );
  AOI211_X1 U18370 ( .C1(n14952), .C2(n19964), .A(n14951), .B(n15739), .ZN(
        n14953) );
  OAI211_X1 U18371 ( .C1(n14955), .C2(n15872), .A(n14954), .B(n14953), .ZN(
        P1_U3011) );
  NAND2_X1 U18372 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14956), .ZN(
        n15825) );
  NOR2_X1 U18373 ( .A1(n15831), .A2(n15825), .ZN(n15817) );
  INV_X1 U18374 ( .A(n15817), .ZN(n14969) );
  OAI21_X1 U18375 ( .B1(n14958), .B2(n11550), .A(n14957), .ZN(n14960) );
  XNOR2_X1 U18376 ( .A(n14960), .B(n14959), .ZN(n15746) );
  NAND2_X1 U18377 ( .A1(n15746), .A2(n19965), .ZN(n14968) );
  INV_X1 U18378 ( .A(n14961), .ZN(n15849) );
  INV_X1 U18379 ( .A(n15865), .ZN(n19945) );
  INV_X1 U18380 ( .A(n15881), .ZN(n15842) );
  AOI21_X1 U18381 ( .B1(n19945), .B2(n14962), .A(n15842), .ZN(n15906) );
  OAI21_X1 U18382 ( .B1(n21043), .B2(n15833), .A(n15907), .ZN(n14963) );
  OAI211_X1 U18383 ( .C1(n14964), .C2(n15849), .A(n15906), .B(n14963), .ZN(
        n15809) );
  INV_X1 U18384 ( .A(n15809), .ZN(n15832) );
  OAI21_X1 U18385 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15825), .A(
        n15832), .ZN(n14966) );
  OAI22_X1 U18386 ( .A1(n15684), .A2(n15909), .B1(n15908), .B2(n20692), .ZN(
        n14965) );
  AOI21_X1 U18387 ( .B1(n14966), .B2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n14965), .ZN(n14967) );
  OAI211_X1 U18388 ( .C1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n14969), .A(
        n14968), .B(n14967), .ZN(P1_U3015) );
  NAND2_X1 U18389 ( .A1(n9766), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20587) );
  OAI211_X1 U18390 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n9766), .A(n20587), 
        .B(n20580), .ZN(n14971) );
  OAI21_X1 U18391 ( .B1(n14975), .B2(n20508), .A(n14971), .ZN(n14972) );
  MUX2_X1 U18392 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14972), .S(
        n20747), .Z(P1_U3477) );
  XNOR2_X1 U18393 ( .A(n14974), .B(n20587), .ZN(n14976) );
  OAI22_X1 U18394 ( .A1(n14976), .A2(n20743), .B1(n13262), .B2(n14975), .ZN(
        n14977) );
  MUX2_X1 U18395 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14977), .S(
        n20747), .Z(P1_U3476) );
  NOR2_X1 U18396 ( .A1(n14985), .A2(n14984), .ZN(n14980) );
  INV_X1 U18397 ( .A(n14978), .ZN(n14979) );
  AOI22_X1 U18398 ( .A1(n15548), .A2(n13274), .B1(n14980), .B2(n14979), .ZN(
        n14981) );
  OAI21_X1 U18399 ( .B1(n20508), .B2(n14982), .A(n14981), .ZN(n15550) );
  INV_X1 U18400 ( .A(n15550), .ZN(n14990) );
  INV_X1 U18401 ( .A(n14983), .ZN(n20728) );
  NOR3_X1 U18402 ( .A1(n14985), .A2(n14984), .A3(n20726), .ZN(n14986) );
  AOI21_X1 U18403 ( .B1(n14988), .B2(n14987), .A(n14986), .ZN(n14989) );
  OAI21_X1 U18404 ( .B1(n14990), .B2(n20728), .A(n14989), .ZN(n14992) );
  MUX2_X1 U18405 ( .A(n14992), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n14991), .Z(P1_U3473) );
  NOR2_X1 U18406 ( .A1(n14993), .A2(n14994), .ZN(n14995) );
  AOI22_X1 U18407 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n18922), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n18912), .ZN(n14999) );
  AOI22_X1 U18408 ( .A1(n14997), .A2(n18885), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18939), .ZN(n14998) );
  OAI211_X1 U18409 ( .C1(n15253), .C2(n18921), .A(n14999), .B(n14998), .ZN(
        n15003) );
  AOI211_X1 U18410 ( .C1(n15001), .C2(n9811), .A(n15000), .B(n19602), .ZN(
        n15002) );
  NOR2_X1 U18411 ( .A1(n15003), .A2(n15002), .ZN(n15004) );
  OAI21_X1 U18412 ( .B1(n15256), .B2(n18900), .A(n15004), .ZN(P2_U2826) );
  AOI211_X1 U18413 ( .C1(n15007), .C2(n15006), .A(n15005), .B(n19602), .ZN(
        n15021) );
  AOI21_X1 U18414 ( .B1(n15009), .B2(n15024), .A(n15008), .ZN(n15269) );
  INV_X1 U18415 ( .A(n15269), .ZN(n15019) );
  AND2_X1 U18416 ( .A1(n15027), .A2(n15010), .ZN(n15011) );
  NOR2_X1 U18417 ( .A1(n14993), .A2(n15011), .ZN(n15262) );
  NAND2_X1 U18418 ( .A1(n15262), .A2(n18923), .ZN(n15013) );
  NAND2_X1 U18419 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18939), .ZN(
        n15012) );
  OAI211_X1 U18420 ( .C1(n18906), .C2(n15014), .A(n15013), .B(n15012), .ZN(
        n15015) );
  AOI21_X1 U18421 ( .B1(n18912), .B2(P2_REIP_REG_28__SCAN_IN), .A(n15015), 
        .ZN(n15018) );
  NAND2_X1 U18422 ( .A1(n15016), .A2(n18885), .ZN(n15017) );
  OAI211_X1 U18423 ( .C1(n15019), .C2(n18900), .A(n15018), .B(n15017), .ZN(
        n15020) );
  OR2_X1 U18424 ( .A1(n15021), .A2(n15020), .ZN(P2_U2827) );
  NAND2_X1 U18425 ( .A1(n12810), .A2(n15022), .ZN(n15023) );
  NAND2_X1 U18426 ( .A1(n15024), .A2(n15023), .ZN(n15278) );
  NAND2_X1 U18427 ( .A1(n12788), .A2(n15025), .ZN(n15026) );
  NAND2_X1 U18428 ( .A1(n15027), .A2(n15026), .ZN(n15277) );
  AOI22_X1 U18429 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n18922), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n18912), .ZN(n15031) );
  OAI22_X1 U18430 ( .A1(n15028), .A2(n18927), .B1(n18908), .B2(n15204), .ZN(
        n15029) );
  INV_X1 U18431 ( .A(n15029), .ZN(n15030) );
  OAI211_X1 U18432 ( .C1(n15277), .C2(n18921), .A(n15031), .B(n15030), .ZN(
        n15035) );
  AOI211_X1 U18433 ( .C1(n15207), .C2(n15033), .A(n15032), .B(n19602), .ZN(
        n15034) );
  NOR2_X1 U18434 ( .A1(n15035), .A2(n15034), .ZN(n15036) );
  OAI21_X1 U18435 ( .B1(n15278), .B2(n18900), .A(n15036), .ZN(P2_U2828) );
  AOI22_X1 U18436 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n18922), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n18912), .ZN(n15037) );
  OAI21_X1 U18437 ( .B1(n15038), .B2(n18908), .A(n15037), .ZN(n15039) );
  AOI21_X1 U18438 ( .B1(n15040), .B2(n18923), .A(n15039), .ZN(n15041) );
  OAI21_X1 U18439 ( .B1(n15042), .B2(n18927), .A(n15041), .ZN(n15047) );
  AOI211_X1 U18440 ( .C1(n15045), .C2(n15044), .A(n15043), .B(n19602), .ZN(
        n15046) );
  AOI211_X1 U18441 ( .C1(n18933), .C2(n15097), .A(n15047), .B(n15046), .ZN(
        n15048) );
  INV_X1 U18442 ( .A(n15048), .ZN(P2_U2830) );
  INV_X1 U18443 ( .A(n15064), .ZN(n15050) );
  AOI221_X1 U18444 ( .B1(n15052), .B2(n15064), .C1(n15051), .C2(n15050), .A(
        n19602), .ZN(n15053) );
  INV_X1 U18445 ( .A(n15053), .ZN(n15062) );
  NAND2_X1 U18446 ( .A1(n18885), .A2(n15054), .ZN(n15056) );
  AOI22_X1 U18447 ( .A1(P2_EBX_REG_2__SCAN_IN), .A2(n18922), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n18912), .ZN(n15055) );
  OAI211_X1 U18448 ( .C1(n18908), .C2(n15057), .A(n15056), .B(n15055), .ZN(
        n15060) );
  NOR2_X1 U18449 ( .A1(n15058), .A2(n18921), .ZN(n15059) );
  AOI211_X1 U18450 ( .C1(n18933), .C2(n9761), .A(n15060), .B(n15059), .ZN(
        n15061) );
  OAI211_X1 U18451 ( .C1(n15488), .C2(n15063), .A(n15062), .B(n15061), .ZN(
        P2_U2853) );
  OAI21_X1 U18452 ( .B1(n15453), .B2(n15065), .A(n15064), .ZN(n15459) );
  AOI22_X1 U18453 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(n18922), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n18912), .ZN(n15066) );
  OAI21_X1 U18454 ( .B1(n10242), .B2(n18908), .A(n15066), .ZN(n15067) );
  AOI21_X1 U18455 ( .B1(n18938), .B2(n10242), .A(n15067), .ZN(n15068) );
  OAI21_X1 U18456 ( .B1(n18927), .B2(n19053), .A(n15068), .ZN(n15069) );
  AOI21_X1 U18457 ( .B1(n18923), .B2(n19706), .A(n15069), .ZN(n15070) );
  OAI21_X1 U18458 ( .B1(n13206), .B2(n18900), .A(n15070), .ZN(n15071) );
  AOI21_X1 U18459 ( .B1(n19702), .B2(n18936), .A(n15071), .ZN(n15072) );
  OAI21_X1 U18460 ( .B1(n15459), .B2(n19602), .A(n15072), .ZN(P2_U2854) );
  NOR2_X1 U18461 ( .A1(n15074), .A2(n15073), .ZN(n15115) );
  NAND2_X1 U18462 ( .A1(n13516), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15075) );
  OAI211_X1 U18463 ( .C1(n15256), .C2(n13516), .A(n15076), .B(n15075), .ZN(
        P2_U2858) );
  NAND2_X1 U18464 ( .A1(n15078), .A2(n15077), .ZN(n15079) );
  XOR2_X1 U18465 ( .A(n15080), .B(n15079), .Z(n15127) );
  NAND2_X1 U18466 ( .A1(n13516), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15082) );
  NAND2_X1 U18467 ( .A1(n15269), .A2(n18965), .ZN(n15081) );
  OAI211_X1 U18468 ( .C1(n15127), .C2(n18951), .A(n15082), .B(n15081), .ZN(
        P2_U2859) );
  OAI21_X1 U18469 ( .B1(n15083), .B2(n15085), .A(n15084), .ZN(n15133) );
  NOR2_X1 U18470 ( .A1(n15278), .A2(n13516), .ZN(n15086) );
  AOI21_X1 U18471 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n13516), .A(n15086), .ZN(
        n15087) );
  OAI21_X1 U18472 ( .B1(n15133), .B2(n18951), .A(n15087), .ZN(P2_U2860) );
  INV_X1 U18473 ( .A(n15088), .ZN(n15958) );
  AOI21_X1 U18474 ( .B1(n15091), .B2(n15090), .A(n15089), .ZN(n15134) );
  NAND2_X1 U18475 ( .A1(n15134), .A2(n18966), .ZN(n15093) );
  NAND2_X1 U18476 ( .A1(n13516), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15092) );
  OAI211_X1 U18477 ( .C1(n15958), .C2(n13516), .A(n15093), .B(n15092), .ZN(
        P2_U2861) );
  OAI21_X1 U18478 ( .B1(n15096), .B2(n15095), .A(n15094), .ZN(n15145) );
  NAND2_X1 U18479 ( .A1(n13516), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15099) );
  NAND2_X1 U18480 ( .A1(n15097), .A2(n18965), .ZN(n15098) );
  OAI211_X1 U18481 ( .C1(n15145), .C2(n18951), .A(n15099), .B(n15098), .ZN(
        P2_U2862) );
  NAND2_X1 U18482 ( .A1(n15101), .A2(n15100), .ZN(n15102) );
  NAND2_X1 U18483 ( .A1(n10025), .A2(n15102), .ZN(n15964) );
  NAND2_X1 U18484 ( .A1(n15104), .A2(n15103), .ZN(n15146) );
  NAND3_X1 U18485 ( .A1(n15148), .A2(n18966), .A3(n15146), .ZN(n15106) );
  NAND2_X1 U18486 ( .A1(n13516), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n15105) );
  OAI211_X1 U18487 ( .C1(n15964), .C2(n13516), .A(n15106), .B(n15105), .ZN(
        P2_U2863) );
  AOI21_X1 U18488 ( .B1(n15109), .B2(n15108), .A(n15107), .ZN(n15110) );
  INV_X1 U18489 ( .A(n15110), .ZN(n15163) );
  NAND2_X1 U18490 ( .A1(n13516), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15113) );
  NAND2_X1 U18491 ( .A1(n15111), .A2(n18965), .ZN(n15112) );
  OAI211_X1 U18492 ( .C1(n15163), .C2(n18951), .A(n15113), .B(n15112), .ZN(
        P2_U2864) );
  OR3_X1 U18493 ( .A1(n15115), .A2(n15114), .A3(n18998), .ZN(n15121) );
  OAI22_X1 U18494 ( .A1(n15253), .A2(n15994), .B1(n15168), .B2(n15116), .ZN(
        n15117) );
  AOI21_X1 U18495 ( .B1(n18974), .B2(n15118), .A(n15117), .ZN(n15120) );
  AOI22_X1 U18496 ( .A1(n18976), .A2(BUF2_REG_29__SCAN_IN), .B1(n18977), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15119) );
  NAND3_X1 U18497 ( .A1(n15121), .A2(n15120), .A3(n15119), .ZN(P2_U2890) );
  OAI22_X1 U18498 ( .A1(n15123), .A2(n15169), .B1(n15168), .B2(n15122), .ZN(
        n15124) );
  AOI21_X1 U18499 ( .B1(n15262), .B2(n18980), .A(n15124), .ZN(n15126) );
  AOI22_X1 U18500 ( .A1(n18976), .A2(BUF2_REG_28__SCAN_IN), .B1(n18977), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15125) );
  OAI211_X1 U18501 ( .C1(n15127), .C2(n18998), .A(n15126), .B(n15125), .ZN(
        P2_U2891) );
  OAI22_X1 U18502 ( .A1(n15994), .A2(n15277), .B1(n15168), .B2(n15128), .ZN(
        n15129) );
  AOI21_X1 U18503 ( .B1(n18974), .B2(n15130), .A(n15129), .ZN(n15132) );
  AOI22_X1 U18504 ( .A1(n18976), .A2(BUF2_REG_27__SCAN_IN), .B1(n18977), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15131) );
  OAI211_X1 U18505 ( .C1(n15133), .C2(n18998), .A(n15132), .B(n15131), .ZN(
        P2_U2892) );
  NAND2_X1 U18506 ( .A1(n15134), .A2(n15147), .ZN(n15138) );
  AOI22_X1 U18507 ( .A1(n18980), .A2(n15961), .B1(n18995), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15137) );
  AOI22_X1 U18508 ( .A1(n18976), .A2(BUF2_REG_26__SCAN_IN), .B1(n18977), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15136) );
  NAND2_X1 U18509 ( .A1(n18974), .A2(n18992), .ZN(n15135) );
  NAND4_X1 U18510 ( .A1(n15138), .A2(n15137), .A3(n15136), .A4(n15135), .ZN(
        P2_U2893) );
  OAI22_X1 U18511 ( .A1(n15994), .A2(n15140), .B1(n15168), .B2(n15139), .ZN(
        n15141) );
  AOI21_X1 U18512 ( .B1(n18974), .B2(n15142), .A(n15141), .ZN(n15144) );
  AOI22_X1 U18513 ( .A1(n18976), .A2(BUF2_REG_25__SCAN_IN), .B1(n18977), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15143) );
  OAI211_X1 U18514 ( .C1(n15145), .C2(n18998), .A(n15144), .B(n15143), .ZN(
        P2_U2894) );
  NAND3_X1 U18515 ( .A1(n15148), .A2(n15147), .A3(n15146), .ZN(n15157) );
  INV_X1 U18516 ( .A(n15149), .ZN(n15151) );
  OAI21_X1 U18517 ( .B1(n15152), .B2(n15151), .A(n15150), .ZN(n15290) );
  INV_X1 U18518 ( .A(n15290), .ZN(n15965) );
  OAI22_X1 U18519 ( .A1(n15153), .A2(n15169), .B1(n15168), .B2(n11132), .ZN(
        n15154) );
  AOI21_X1 U18520 ( .B1(n18980), .B2(n15965), .A(n15154), .ZN(n15156) );
  AOI22_X1 U18521 ( .A1(n18976), .A2(BUF2_REG_24__SCAN_IN), .B1(n18977), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15155) );
  NAND3_X1 U18522 ( .A1(n15157), .A2(n15156), .A3(n15155), .ZN(P2_U2895) );
  OAI22_X1 U18523 ( .A1(n19127), .A2(n15169), .B1(n15168), .B2(n15158), .ZN(
        n15159) );
  AOI21_X1 U18524 ( .B1(n18980), .B2(n15160), .A(n15159), .ZN(n15162) );
  AOI22_X1 U18525 ( .A1(n18976), .A2(BUF2_REG_23__SCAN_IN), .B1(n18977), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n15161) );
  OAI211_X1 U18526 ( .C1(n15163), .C2(n18998), .A(n15162), .B(n15161), .ZN(
        P2_U2896) );
  AOI21_X1 U18527 ( .B1(n15165), .B2(n15164), .A(n14309), .ZN(n15977) );
  INV_X1 U18528 ( .A(n15977), .ZN(n15174) );
  XNOR2_X1 U18529 ( .A(n15166), .B(n11065), .ZN(n15541) );
  INV_X1 U18530 ( .A(n15541), .ZN(n15171) );
  OAI22_X1 U18531 ( .A1(n19116), .A2(n15169), .B1(n15168), .B2(n15167), .ZN(
        n15170) );
  AOI21_X1 U18532 ( .B1(n18980), .B2(n15171), .A(n15170), .ZN(n15173) );
  AOI22_X1 U18533 ( .A1(n18976), .A2(BUF2_REG_22__SCAN_IN), .B1(n18977), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n15172) );
  OAI211_X1 U18534 ( .C1(n15174), .C2(n18998), .A(n15173), .B(n15172), .ZN(
        P2_U2897) );
  NOR2_X1 U18535 ( .A1(n16100), .A2(n15175), .ZN(n15176) );
  AOI211_X1 U18536 ( .C1(n15178), .C2(n16090), .A(n15177), .B(n15176), .ZN(
        n15179) );
  OAI21_X1 U18537 ( .B1(n15180), .B2(n16077), .A(n15179), .ZN(n15181) );
  AOI21_X1 U18538 ( .B1(n15182), .B2(n14248), .A(n15181), .ZN(n15183) );
  OAI21_X1 U18539 ( .B1(n15184), .B2(n16084), .A(n15183), .ZN(P2_U2984) );
  XNOR2_X1 U18540 ( .A(n15189), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15190) );
  XNOR2_X1 U18541 ( .A(n15191), .B(n15190), .ZN(n15271) );
  INV_X1 U18542 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n15192) );
  NOR2_X1 U18543 ( .A1(n18814), .A2(n15192), .ZN(n15261) );
  AOI21_X1 U18544 ( .B1(n19055), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15261), .ZN(n15193) );
  OAI21_X1 U18545 ( .B1(n19061), .B2(n15194), .A(n15193), .ZN(n15199) );
  INV_X1 U18546 ( .A(n15195), .ZN(n15196) );
  OAI21_X1 U18547 ( .B1(n15195), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15197), .ZN(n15266) );
  NOR2_X1 U18548 ( .A1(n15266), .A2(n16083), .ZN(n15198) );
  AOI211_X1 U18549 ( .C1(n19063), .C2(n15269), .A(n15199), .B(n15198), .ZN(
        n15200) );
  OAI21_X1 U18550 ( .B1(n15271), .B2(n16084), .A(n15200), .ZN(P2_U2986) );
  INV_X1 U18551 ( .A(n15201), .ZN(n15202) );
  OAI21_X1 U18552 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15202), .A(
        n15196), .ZN(n15284) );
  OR2_X1 U18553 ( .A1(n15203), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15273) );
  NAND3_X1 U18554 ( .A1(n15273), .A2(n15272), .A3(n19056), .ZN(n15209) );
  INV_X1 U18555 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19664) );
  OR2_X1 U18556 ( .A1(n18814), .A2(n19664), .ZN(n15275) );
  OAI21_X1 U18557 ( .B1(n16100), .B2(n15204), .A(n15275), .ZN(n15206) );
  NOR2_X1 U18558 ( .A1(n15278), .A2(n16077), .ZN(n15205) );
  AOI211_X1 U18559 ( .C1(n16090), .C2(n15207), .A(n15206), .B(n15205), .ZN(
        n15208) );
  OAI211_X1 U18560 ( .C1(n16083), .C2(n15284), .A(n15209), .B(n15208), .ZN(
        P2_U2987) );
  INV_X1 U18561 ( .A(n9788), .ZN(n15212) );
  XOR2_X1 U18562 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n15210), .Z(
        n15211) );
  XNOR2_X1 U18563 ( .A(n15212), .B(n15211), .ZN(n15297) );
  AOI21_X1 U18564 ( .B1(n15286), .B2(n15214), .A(n15213), .ZN(n15295) );
  INV_X1 U18565 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19657) );
  OR2_X1 U18566 ( .A1(n18814), .A2(n19657), .ZN(n15288) );
  OAI21_X1 U18567 ( .B1(n16100), .B2(n15215), .A(n15288), .ZN(n15216) );
  AOI21_X1 U18568 ( .B1(n16090), .B2(n15969), .A(n15216), .ZN(n15217) );
  OAI21_X1 U18569 ( .B1(n15964), .B2(n16077), .A(n15217), .ZN(n15218) );
  AOI21_X1 U18570 ( .B1(n15295), .B2(n14248), .A(n15218), .ZN(n15219) );
  OAI21_X1 U18571 ( .B1(n15297), .B2(n16084), .A(n15219), .ZN(P2_U2990) );
  OAI21_X1 U18572 ( .B1(n15222), .B2(n15221), .A(n15220), .ZN(n15329) );
  AOI21_X1 U18573 ( .B1(n15223), .B2(n15318), .A(n15224), .ZN(n15327) );
  NOR2_X1 U18574 ( .A1(n18814), .A2(n19650), .ZN(n15321) );
  NOR2_X1 U18575 ( .A1(n15225), .A2(n19061), .ZN(n15226) );
  AOI211_X1 U18576 ( .C1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n19055), .A(
        n15321), .B(n15226), .ZN(n15227) );
  OAI21_X1 U18577 ( .B1(n15986), .B2(n16077), .A(n15227), .ZN(n15228) );
  AOI21_X1 U18578 ( .B1(n15327), .B2(n14248), .A(n15228), .ZN(n15229) );
  OAI21_X1 U18579 ( .B1(n15329), .B2(n16084), .A(n15229), .ZN(P2_U2994) );
  OAI21_X1 U18580 ( .B1(n15232), .B2(n15231), .A(n15230), .ZN(n15341) );
  INV_X1 U18581 ( .A(n15341), .ZN(n15241) );
  INV_X1 U18582 ( .A(n15334), .ZN(n18821) );
  NOR2_X1 U18583 ( .A1(n19644), .A2(n11123), .ZN(n15235) );
  OAI22_X1 U18584 ( .A1(n16100), .A2(n15233), .B1(n19061), .B2(n18824), .ZN(
        n15234) );
  AOI211_X1 U18585 ( .C1(n18821), .C2(n19063), .A(n15235), .B(n15234), .ZN(
        n15240) );
  INV_X1 U18586 ( .A(n15330), .ZN(n15238) );
  INV_X1 U18587 ( .A(n15236), .ZN(n15237) );
  OAI211_X1 U18588 ( .C1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n15238), .A(
        n15237), .B(n14248), .ZN(n15239) );
  OAI211_X1 U18589 ( .C1(n15241), .C2(n16084), .A(n15240), .B(n15239), .ZN(
        P2_U2997) );
  XNOR2_X1 U18590 ( .A(n15243), .B(n15242), .ZN(n15353) );
  NOR2_X1 U18591 ( .A1(n19061), .A2(n15244), .ZN(n15246) );
  OAI22_X1 U18592 ( .A1(n16100), .A2(n10814), .B1(n15346), .B2(n18814), .ZN(
        n15245) );
  AOI211_X1 U18593 ( .C1(n15247), .C2(n19063), .A(n15246), .B(n15245), .ZN(
        n15250) );
  OAI211_X1 U18594 ( .C1(n15248), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n14248), .B(n15330), .ZN(n15249) );
  OAI211_X1 U18595 ( .C1(n15353), .C2(n16084), .A(n15250), .B(n15249), .ZN(
        P2_U2998) );
  NOR2_X1 U18596 ( .A1(n15259), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15274) );
  NOR2_X1 U18597 ( .A1(n15281), .A2(n15274), .ZN(n15265) );
  OAI21_X1 U18598 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n15259), .A(
        n15265), .ZN(n15255) );
  OAI21_X1 U18599 ( .B1(n15253), .B2(n16161), .A(n15252), .ZN(n15254) );
  NOR3_X1 U18600 ( .A1(n15259), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n12852), .ZN(n15260) );
  AOI211_X1 U18601 ( .C1(n19067), .C2(n15262), .A(n15261), .B(n15260), .ZN(
        n15263) );
  OAI21_X1 U18602 ( .B1(n15265), .B2(n15264), .A(n15263), .ZN(n15268) );
  NOR2_X1 U18603 ( .A1(n15266), .A2(n19074), .ZN(n15267) );
  AOI211_X1 U18604 ( .C1(n15269), .C2(n16143), .A(n15268), .B(n15267), .ZN(
        n15270) );
  OAI21_X1 U18605 ( .B1(n15271), .B2(n16163), .A(n15270), .ZN(P2_U3018) );
  NAND3_X1 U18606 ( .A1(n15273), .A2(n15272), .A3(n19069), .ZN(n15283) );
  INV_X1 U18607 ( .A(n15274), .ZN(n15276) );
  OAI211_X1 U18608 ( .C1(n16161), .C2(n15277), .A(n15276), .B(n15275), .ZN(
        n15280) );
  NOR2_X1 U18609 ( .A1(n15278), .A2(n19072), .ZN(n15279) );
  AOI211_X1 U18610 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15281), .A(
        n15280), .B(n15279), .ZN(n15282) );
  OAI211_X1 U18611 ( .C1(n15284), .C2(n19074), .A(n15283), .B(n15282), .ZN(
        P2_U3019) );
  OAI21_X1 U18612 ( .B1(n15287), .B2(n15285), .A(n15311), .ZN(n15292) );
  NAND3_X1 U18613 ( .A1(n15309), .A2(n15287), .A3(n15286), .ZN(n15289) );
  OAI211_X1 U18614 ( .C1(n16161), .C2(n15290), .A(n15289), .B(n15288), .ZN(
        n15291) );
  AOI21_X1 U18615 ( .B1(n15292), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15291), .ZN(n15293) );
  OAI21_X1 U18616 ( .B1(n15964), .B2(n19072), .A(n15293), .ZN(n15294) );
  AOI21_X1 U18617 ( .B1(n15295), .B2(n16153), .A(n15294), .ZN(n15296) );
  OAI21_X1 U18618 ( .B1(n15297), .B2(n16163), .A(n15296), .ZN(P2_U3022) );
  INV_X1 U18619 ( .A(n15299), .ZN(n15300) );
  NOR2_X1 U18620 ( .A1(n15301), .A2(n15300), .ZN(n15302) );
  XNOR2_X1 U18621 ( .A(n15298), .B(n15302), .ZN(n16002) );
  INV_X1 U18622 ( .A(n16002), .ZN(n15316) );
  INV_X1 U18623 ( .A(n16005), .ZN(n15304) );
  OR2_X1 U18624 ( .A1(n15303), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16000) );
  NAND3_X1 U18625 ( .A1(n15304), .A2(n16153), .A3(n16000), .ZN(n15315) );
  OR2_X1 U18626 ( .A1(n14084), .A2(n15305), .ZN(n15306) );
  NAND2_X1 U18627 ( .A1(n10843), .A2(n15306), .ZN(n16001) );
  INV_X1 U18628 ( .A(n16001), .ZN(n15313) );
  NOR2_X1 U18629 ( .A1(n16161), .A2(n15541), .ZN(n15308) );
  NOR2_X1 U18630 ( .A1(n11059), .A2(n11123), .ZN(n15307) );
  AOI211_X1 U18631 ( .C1(n15309), .C2(n20973), .A(n15308), .B(n15307), .ZN(
        n15310) );
  OAI21_X1 U18632 ( .B1(n15311), .B2(n20973), .A(n15310), .ZN(n15312) );
  AOI21_X1 U18633 ( .B1(n15313), .B2(n16143), .A(n15312), .ZN(n15314) );
  OAI211_X1 U18634 ( .C1(n15316), .C2(n16163), .A(n15315), .B(n15314), .ZN(
        P2_U3024) );
  NOR2_X1 U18635 ( .A1(n15995), .A2(n16161), .ZN(n15326) );
  XNOR2_X1 U18636 ( .A(n15317), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15322) );
  NOR2_X1 U18637 ( .A1(n15319), .A2(n15318), .ZN(n15320) );
  AOI211_X1 U18638 ( .C1(n15323), .C2(n15322), .A(n15321), .B(n15320), .ZN(
        n15324) );
  OAI21_X1 U18639 ( .B1(n19072), .B2(n15986), .A(n15324), .ZN(n15325) );
  AOI211_X1 U18640 ( .C1(n15327), .C2(n16153), .A(n15326), .B(n15325), .ZN(
        n15328) );
  OAI21_X1 U18641 ( .B1(n15329), .B2(n16163), .A(n15328), .ZN(P2_U3026) );
  OAI21_X1 U18642 ( .B1(n16153), .B2(n15331), .A(n15330), .ZN(n15332) );
  OAI211_X1 U18643 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15333), .A(
        n15332), .B(n15364), .ZN(n15351) );
  AOI21_X1 U18644 ( .B1(n15337), .B2(n19078), .A(n15351), .ZN(n15345) );
  INV_X1 U18645 ( .A(n18828), .ZN(n15340) );
  OAI22_X1 U18646 ( .A1(n15334), .A2(n19072), .B1(n19644), .B2(n18814), .ZN(
        n15339) );
  OAI21_X1 U18647 ( .B1(n15335), .B2(n19074), .A(n15358), .ZN(n15336) );
  NAND2_X1 U18648 ( .A1(n15336), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15349) );
  NOR3_X1 U18649 ( .A1(n15349), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15337), .ZN(n15338) );
  AOI211_X1 U18650 ( .C1(n19067), .C2(n15340), .A(n15339), .B(n15338), .ZN(
        n15343) );
  NAND2_X1 U18651 ( .A1(n15341), .A2(n19069), .ZN(n15342) );
  OAI211_X1 U18652 ( .C1(n15345), .C2(n15344), .A(n15343), .B(n15342), .ZN(
        P2_U3029) );
  OAI22_X1 U18653 ( .A1(n18950), .A2(n19072), .B1(n15346), .B2(n18814), .ZN(
        n15347) );
  AOI21_X1 U18654 ( .B1(n18981), .B2(n19067), .A(n15347), .ZN(n15348) );
  OAI21_X1 U18655 ( .B1(n15349), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15348), .ZN(n15350) );
  AOI21_X1 U18656 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15351), .A(
        n15350), .ZN(n15352) );
  OAI21_X1 U18657 ( .B1(n16163), .B2(n15353), .A(n15352), .ZN(P2_U3030) );
  NAND2_X1 U18658 ( .A1(n15355), .A2(n15354), .ZN(n15357) );
  XOR2_X1 U18659 ( .A(n15357), .B(n15356), .Z(n16012) );
  INV_X1 U18660 ( .A(n18842), .ZN(n15369) );
  INV_X1 U18661 ( .A(n15358), .ZN(n15360) );
  INV_X1 U18662 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19642) );
  NOR2_X1 U18663 ( .A1(n19642), .A2(n11123), .ZN(n15359) );
  AOI21_X1 U18664 ( .B1(n15360), .B2(n15363), .A(n15359), .ZN(n15362) );
  NAND2_X1 U18665 ( .A1(n18839), .A2(n16143), .ZN(n15361) );
  OAI211_X1 U18666 ( .C1(n15364), .C2(n15363), .A(n15362), .B(n15361), .ZN(
        n15368) );
  OAI21_X1 U18667 ( .B1(n15365), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15366), .ZN(n16011) );
  NOR2_X1 U18668 ( .A1(n16011), .A2(n19074), .ZN(n15367) );
  AOI211_X1 U18669 ( .C1(n19067), .C2(n15369), .A(n15368), .B(n15367), .ZN(
        n15370) );
  OAI21_X1 U18670 ( .B1(n16012), .B2(n16163), .A(n15370), .ZN(P2_U3031) );
  AND2_X1 U18671 ( .A1(n15372), .A2(n15371), .ZN(n15373) );
  XNOR2_X1 U18672 ( .A(n15374), .B(n15373), .ZN(n16016) );
  INV_X1 U18673 ( .A(n16016), .ZN(n15394) );
  AND2_X1 U18674 ( .A1(n15410), .A2(n15376), .ZN(n15377) );
  OR2_X1 U18675 ( .A1(n15377), .A2(n15365), .ZN(n16019) );
  NOR2_X1 U18676 ( .A1(n16019), .A2(n19074), .ZN(n15392) );
  INV_X1 U18677 ( .A(n15402), .ZN(n15378) );
  NOR2_X1 U18678 ( .A1(n15379), .A2(n15378), .ZN(n15382) );
  NAND2_X1 U18679 ( .A1(n15402), .A2(n10731), .ZN(n16103) );
  NAND2_X1 U18680 ( .A1(n16102), .A2(n16103), .ZN(n15406) );
  AOI21_X1 U18681 ( .B1(n15402), .B2(n15409), .A(n15406), .ZN(n15380) );
  INV_X1 U18682 ( .A(n15380), .ZN(n15381) );
  MUX2_X1 U18683 ( .A(n15382), .B(n15381), .S(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n15391) );
  INV_X1 U18684 ( .A(n13732), .ZN(n15386) );
  NAND2_X1 U18685 ( .A1(n15384), .A2(n15383), .ZN(n15385) );
  NAND2_X1 U18686 ( .A1(n15386), .A2(n15385), .ZN(n18955) );
  NOR2_X1 U18687 ( .A1(n18955), .A2(n19072), .ZN(n15390) );
  AOI21_X1 U18688 ( .B1(n15387), .B2(n13543), .A(n13628), .ZN(n15388) );
  INV_X1 U18689 ( .A(n15388), .ZN(n18987) );
  OAI22_X1 U18690 ( .A1(n16161), .A2(n18987), .B1(n11020), .B2(n18814), .ZN(
        n15389) );
  NOR4_X1 U18691 ( .A1(n15392), .A2(n15391), .A3(n15390), .A4(n15389), .ZN(
        n15393) );
  OAI21_X1 U18692 ( .B1(n16163), .B2(n15394), .A(n15393), .ZN(P2_U3032) );
  OR2_X1 U18693 ( .A1(n15395), .A2(n16028), .ZN(n15397) );
  NAND2_X1 U18694 ( .A1(n15397), .A2(n15396), .ZN(n15401) );
  NAND2_X1 U18695 ( .A1(n15399), .A2(n15398), .ZN(n15400) );
  XNOR2_X1 U18696 ( .A(n15401), .B(n15400), .ZN(n16024) );
  NAND2_X1 U18697 ( .A1(n15402), .A2(n15409), .ZN(n15403) );
  NOR2_X1 U18698 ( .A1(n10731), .A2(n15403), .ZN(n15405) );
  INV_X1 U18699 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19639) );
  NOR2_X1 U18700 ( .A1(n19639), .A2(n18814), .ZN(n15404) );
  AOI211_X1 U18701 ( .C1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n15406), .A(
        n15405), .B(n15404), .ZN(n15407) );
  OAI21_X1 U18702 ( .B1(n16161), .B2(n18864), .A(n15407), .ZN(n15413) );
  OR2_X1 U18703 ( .A1(n16031), .A2(n10731), .ZN(n16033) );
  NAND2_X1 U18704 ( .A1(n16033), .A2(n15409), .ZN(n15411) );
  NAND2_X1 U18705 ( .A1(n15411), .A2(n15410), .ZN(n16023) );
  NOR2_X1 U18706 ( .A1(n16023), .A2(n19074), .ZN(n15412) );
  AOI211_X1 U18707 ( .C1(n16143), .C2(n18860), .A(n15413), .B(n15412), .ZN(
        n15414) );
  OAI21_X1 U18708 ( .B1(n16163), .B2(n16024), .A(n15414), .ZN(P2_U3033) );
  NOR2_X1 U18709 ( .A1(n15415), .A2(n15416), .ZN(n15418) );
  NOR2_X1 U18710 ( .A1(n15418), .A2(n15417), .ZN(n15422) );
  NAND2_X1 U18711 ( .A1(n15420), .A2(n15419), .ZN(n15421) );
  XNOR2_X1 U18712 ( .A(n15422), .B(n15421), .ZN(n16041) );
  INV_X1 U18713 ( .A(n15423), .ZN(n15425) );
  INV_X1 U18714 ( .A(n16031), .ZN(n15424) );
  AOI21_X1 U18715 ( .B1(n15427), .B2(n15425), .A(n15424), .ZN(n16040) );
  INV_X1 U18716 ( .A(n16113), .ZN(n15441) );
  NOR2_X1 U18717 ( .A1(n10990), .A2(n18814), .ZN(n15429) );
  AOI211_X1 U18718 ( .C1(n16114), .C2(n15427), .A(n15426), .B(n16115), .ZN(
        n15428) );
  AOI211_X1 U18719 ( .C1(n15441), .C2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15429), .B(n15428), .ZN(n15431) );
  NAND2_X1 U18720 ( .A1(n16044), .A2(n16143), .ZN(n15430) );
  OAI211_X1 U18721 ( .C1(n16161), .C2(n15432), .A(n15431), .B(n15430), .ZN(
        n15433) );
  AOI21_X1 U18722 ( .B1(n16040), .B2(n16153), .A(n15433), .ZN(n15434) );
  OAI21_X1 U18723 ( .B1(n16041), .B2(n16163), .A(n15434), .ZN(P2_U3035) );
  INV_X1 U18724 ( .A(n16048), .ZN(n15435) );
  NOR2_X1 U18725 ( .A1(n15435), .A2(n16047), .ZN(n15436) );
  XOR2_X1 U18726 ( .A(n15436), .B(n15415), .Z(n16062) );
  OAI21_X1 U18727 ( .B1(n9727), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15437), .ZN(n16061) );
  INV_X1 U18728 ( .A(n16061), .ZN(n15446) );
  NOR2_X1 U18729 ( .A1(n10963), .A2(n18814), .ZN(n15439) );
  AOI221_X1 U18730 ( .B1(n15441), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n15440), .C2(n20889), .A(n15439), .ZN(n15444) );
  INV_X1 U18731 ( .A(n15442), .ZN(n18873) );
  NAND2_X1 U18732 ( .A1(n18873), .A2(n16143), .ZN(n15443) );
  OAI211_X1 U18733 ( .C1(n16161), .C2(n18877), .A(n15444), .B(n15443), .ZN(
        n15445) );
  AOI21_X1 U18734 ( .B1(n15446), .B2(n16153), .A(n15445), .ZN(n15447) );
  OAI21_X1 U18735 ( .B1(n16163), .B2(n16062), .A(n15447), .ZN(P2_U3037) );
  OR2_X1 U18736 ( .A1(n13005), .A2(n15461), .ZN(n15452) );
  INV_X1 U18737 ( .A(n10887), .ZN(n15449) );
  AND2_X1 U18738 ( .A1(n15449), .A2(n15448), .ZN(n15466) );
  MUX2_X1 U18739 ( .A(n15466), .B(n15450), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15451) );
  NAND2_X1 U18740 ( .A1(n15452), .A2(n15451), .ZN(n16172) );
  INV_X1 U18741 ( .A(n15453), .ZN(n18935) );
  AOI22_X1 U18742 ( .A1(n18896), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18935), .B2(n18870), .ZN(n15460) );
  AOI22_X1 U18743 ( .A1(n16172), .A2(n19596), .B1(P2_STATE2_REG_1__SCAN_IN), 
        .B2(n15460), .ZN(n15456) );
  NAND2_X1 U18744 ( .A1(n15454), .A2(n16214), .ZN(n15455) );
  AOI21_X1 U18745 ( .B1(n15456), .B2(n15455), .A(n15524), .ZN(n15457) );
  AOI21_X1 U18746 ( .B1(n15524), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n15457), .ZN(n15458) );
  INV_X1 U18747 ( .A(n15458), .ZN(P2_U3601) );
  OAI21_X1 U18748 ( .B1(n18870), .B2(n19059), .A(n15459), .ZN(n15484) );
  INV_X1 U18749 ( .A(n15484), .ZN(n15467) );
  NOR2_X1 U18750 ( .A1(n15460), .A2(n19597), .ZN(n15483) );
  NOR2_X1 U18751 ( .A1(n10303), .A2(n10304), .ZN(n15465) );
  INV_X1 U18752 ( .A(n15461), .ZN(n15470) );
  NAND2_X1 U18753 ( .A1(n19064), .A2(n15470), .ZN(n15464) );
  NAND2_X1 U18754 ( .A1(n9728), .A2(n15462), .ZN(n15463) );
  OAI211_X1 U18755 ( .C1(n15466), .C2(n15465), .A(n15464), .B(n15463), .ZN(
        n16173) );
  AOI222_X1 U18756 ( .A1(n15467), .A2(n15483), .B1(n16173), .B2(n19596), .C1(
        n19702), .C2(n16214), .ZN(n15469) );
  NAND2_X1 U18757 ( .A1(n15524), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15468) );
  OAI21_X1 U18758 ( .B1(n15524), .B2(n15469), .A(n15468), .ZN(P2_U3600) );
  INV_X1 U18759 ( .A(n16214), .ZN(n15486) );
  NAND2_X1 U18760 ( .A1(n9761), .A2(n15470), .ZN(n15482) );
  OAI21_X1 U18761 ( .B1(n9760), .B2(n15472), .A(n15471), .ZN(n15477) );
  NOR2_X1 U18762 ( .A1(n15473), .A2(n10575), .ZN(n15474) );
  NAND2_X1 U18763 ( .A1(n15475), .A2(n15474), .ZN(n15476) );
  NAND2_X1 U18764 ( .A1(n15477), .A2(n15476), .ZN(n15478) );
  AOI21_X1 U18765 ( .B1(n15480), .B2(n15479), .A(n15478), .ZN(n15481) );
  NAND2_X1 U18766 ( .A1(n15482), .A2(n15481), .ZN(n16171) );
  AOI22_X1 U18767 ( .A1(n16171), .A2(n19596), .B1(n15484), .B2(n15483), .ZN(
        n15485) );
  OAI21_X1 U18768 ( .B1(n15488), .B2(n15486), .A(n15485), .ZN(n15487) );
  MUX2_X1 U18769 ( .A(n15487), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15524), .Z(P2_U3599) );
  NAND2_X1 U18770 ( .A1(n19535), .A2(n19593), .ZN(n15489) );
  AOI21_X1 U18771 ( .B1(n15489), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19685), 
        .ZN(n15494) );
  NAND2_X1 U18772 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19441) );
  INV_X1 U18773 ( .A(n19441), .ZN(n19474) );
  NAND2_X1 U18774 ( .A1(n19284), .A2(n19474), .ZN(n15497) );
  NAND2_X1 U18775 ( .A1(n15494), .A2(n15497), .ZN(n15493) );
  NAND2_X1 U18776 ( .A1(n15495), .A2(n19546), .ZN(n15491) );
  NAND2_X1 U18777 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19474), .ZN(
        n19542) );
  NOR2_X1 U18778 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19542), .ZN(
        n19530) );
  NOR2_X1 U18779 ( .A1(n19697), .A2(n19530), .ZN(n15490) );
  AOI21_X1 U18780 ( .B1(n15491), .B2(n15490), .A(n19447), .ZN(n15492) );
  NAND2_X1 U18781 ( .A1(n15493), .A2(n15492), .ZN(n19532) );
  INV_X1 U18782 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15502) );
  INV_X1 U18783 ( .A(n15494), .ZN(n15498) );
  OAI21_X1 U18784 ( .B1(n15495), .B2(n19530), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15496) );
  AOI22_X1 U18785 ( .A1(n19558), .A2(n19574), .B1(n19556), .B2(n19530), .ZN(
        n15499) );
  OAI21_X1 U18786 ( .B1(n19535), .B2(n19561), .A(n15499), .ZN(n15500) );
  AOI21_X1 U18787 ( .B1(n19557), .B2(n19531), .A(n15500), .ZN(n15501) );
  OAI21_X1 U18788 ( .B1(n19529), .B2(n15502), .A(n15501), .ZN(P2_U3162) );
  INV_X1 U18789 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16837) );
  NAND4_X1 U18790 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(P3_EBX_REG_26__SCAN_IN), .A4(P3_EBX_REG_25__SCAN_IN), .ZN(n15504)
         );
  NOR3_X1 U18791 ( .A1(n16456), .A2(n16837), .A3(n15504), .ZN(n15505) );
  NAND4_X1 U18792 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(n16896), .A4(n15505), .ZN(n16737) );
  NOR2_X1 U18793 ( .A1(n16738), .A2(n16737), .ZN(n16836) );
  NAND2_X1 U18794 ( .A1(n17079), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n15507) );
  NAND2_X1 U18795 ( .A1(n16836), .A2(n17097), .ZN(n15506) );
  OAI22_X1 U18796 ( .A1(n16836), .A2(n15507), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n15506), .ZN(P3_U2672) );
  NOR2_X1 U18797 ( .A1(n18730), .A2(n15508), .ZN(n15513) );
  AOI21_X1 U18798 ( .B1(n15513), .B2(n17247), .A(n15610), .ZN(n15514) );
  OAI211_X1 U18799 ( .C1(n15517), .C2(n15516), .A(n15515), .B(n15514), .ZN(
        n18546) );
  INV_X1 U18800 ( .A(n18546), .ZN(n18558) );
  NAND2_X1 U18801 ( .A1(n18732), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18083) );
  INV_X1 U18802 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18068) );
  OR2_X1 U18803 ( .A1(n18068), .A2(n18676), .ZN(n15518) );
  OAI211_X1 U18804 ( .C1(n18579), .C2(n18558), .A(n18083), .B(n15518), .ZN(
        n18707) );
  AOI21_X1 U18805 ( .B1(n18527), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15521) );
  NOR2_X1 U18806 ( .A1(n15521), .A2(n15520), .ZN(n18570) );
  NAND3_X1 U18807 ( .A1(n18707), .A2(n18706), .A3(n18570), .ZN(n15522) );
  OAI21_X1 U18808 ( .B1(n18707), .B2(n18525), .A(n15522), .ZN(P3_U3284) );
  INV_X1 U18809 ( .A(n15524), .ZN(n15526) );
  NAND4_X1 U18810 ( .A1(n16194), .A2(n19737), .A3(n19596), .A4(n16193), .ZN(
        n15523) );
  OR2_X1 U18811 ( .A1(n15524), .A2(n15523), .ZN(n15525) );
  OAI21_X1 U18812 ( .B1(n15526), .B2(n16201), .A(n15525), .ZN(P2_U3595) );
  OAI21_X1 U18813 ( .B1(n18055), .B2(n16241), .A(n15527), .ZN(n15528) );
  AOI21_X1 U18814 ( .B1(n16257), .B2(n17980), .A(n15528), .ZN(n15602) );
  AOI21_X1 U18815 ( .B1(n17948), .B2(n9918), .A(n15529), .ZN(n16254) );
  OAI21_X1 U18816 ( .B1(n17971), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16254), .ZN(n15532) );
  AOI21_X1 U18817 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16256), .A(
        n18055), .ZN(n15530) );
  AOI211_X1 U18818 ( .C1(n17980), .C2(n16246), .A(n15530), .B(n18052), .ZN(
        n15599) );
  INV_X1 U18819 ( .A(n15599), .ZN(n15531) );
  AOI21_X1 U18820 ( .B1(n18057), .B2(n15532), .A(n15531), .ZN(n15537) );
  NOR2_X1 U18821 ( .A1(n15534), .A2(n15533), .ZN(n15535) );
  XOR2_X1 U18822 ( .A(n16242), .B(n15535), .Z(n16245) );
  AOI22_X1 U18823 ( .A1(n18061), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n17979), 
        .B2(n16245), .ZN(n15536) );
  OAI221_X1 U18824 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15602), 
        .C1(n16242), .C2(n15537), .A(n15536), .ZN(P3_U2833) );
  OAI21_X1 U18825 ( .B1(n15538), .B2(n16010), .A(n18917), .ZN(n15545) );
  AOI22_X1 U18826 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18939), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18912), .ZN(n15539) );
  OAI21_X1 U18827 ( .B1(n15540), .B2(n18927), .A(n15539), .ZN(n15543) );
  OAI22_X1 U18828 ( .A1(n16001), .A2(n18900), .B1(n18921), .B2(n15541), .ZN(
        n15542) );
  AOI211_X1 U18829 ( .C1(P2_EBX_REG_22__SCAN_IN), .C2(n18922), .A(n15543), .B(
        n15542), .ZN(n15544) );
  OAI21_X1 U18830 ( .B1(n15546), .B2(n15545), .A(n15544), .ZN(P2_U2833) );
  INV_X1 U18831 ( .A(n15557), .ZN(n15560) );
  AOI21_X1 U18832 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15548), .A(
        n15547), .ZN(n15554) );
  INV_X1 U18833 ( .A(n15554), .ZN(n15551) );
  OAI211_X1 U18834 ( .C1(n15552), .C2(n15551), .A(n15550), .B(n15549), .ZN(
        n15553) );
  OAI211_X1 U18835 ( .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n15554), .A(
        n15553), .B(n20439), .ZN(n15558) );
  AND2_X1 U18836 ( .A1(n20284), .A2(n15558), .ZN(n15556) );
  OAI222_X1 U18837 ( .A1(n20284), .A2(n15558), .B1(n20746), .B2(n15557), .C1(
        n15556), .C2(n15555), .ZN(n15559) );
  OAI21_X1 U18838 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15560), .A(
        n15559), .ZN(n15568) );
  OAI21_X1 U18839 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15561), .ZN(n15563) );
  NAND4_X1 U18840 ( .A1(n15565), .A2(n15564), .A3(n15563), .A4(n15562), .ZN(
        n15566) );
  AOI211_X1 U18841 ( .C1(n15568), .C2(n19973), .A(n15567), .B(n15566), .ZN(
        n15580) );
  INV_X1 U18842 ( .A(n15580), .ZN(n15575) );
  OAI21_X1 U18843 ( .B1(n15569), .B2(n20760), .A(n15579), .ZN(n15574) );
  NAND4_X1 U18844 ( .A1(n11626), .A2(n15572), .A3(n15571), .A4(n15570), .ZN(
        n15573) );
  NAND2_X1 U18845 ( .A1(n15574), .A2(n15573), .ZN(n15940) );
  AOI221_X1 U18846 ( .B1(n15945), .B2(n20957), .C1(n15575), .C2(n20957), .A(
        n15940), .ZN(n15946) );
  AOI21_X1 U18847 ( .B1(n20662), .B2(n20244), .A(n15576), .ZN(n15578) );
  OAI211_X1 U18848 ( .C1(n15580), .C2(n15579), .A(n15578), .B(n15577), .ZN(
        n15581) );
  NOR2_X1 U18849 ( .A1(n15946), .A2(n15581), .ZN(n15585) );
  NAND2_X1 U18850 ( .A1(n20764), .A2(n15582), .ZN(n15583) );
  NAND2_X1 U18851 ( .A1(n15945), .A2(n15583), .ZN(n15584) );
  OAI22_X1 U18852 ( .A1(n15585), .A2(n15945), .B1(n15946), .B2(n15584), .ZN(
        P1_U3161) );
  NAND2_X1 U18853 ( .A1(n15766), .A2(n15586), .ZN(n15587) );
  OAI22_X1 U18854 ( .A1(n15589), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n15588), .B2(n15587), .ZN(n15590) );
  XOR2_X1 U18855 ( .A(n11557), .B(n15590), .Z(n15738) );
  AOI22_X1 U18856 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15591), .B1(
        n19953), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15595) );
  INV_X1 U18857 ( .A(n15592), .ZN(n15650) );
  AOI22_X1 U18858 ( .A1(n15593), .A2(n11557), .B1(n19964), .B2(n15650), .ZN(
        n15594) );
  OAI211_X1 U18859 ( .C1(n15872), .C2(n15738), .A(n15595), .B(n15594), .ZN(
        P1_U3010) );
  NAND2_X1 U18860 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16234), .ZN(
        n16224) );
  OAI21_X1 U18861 ( .B1(n15597), .B2(n16234), .A(n15596), .ZN(n16231) );
  AOI21_X1 U18862 ( .B1(n15599), .B2(n15598), .A(n16234), .ZN(n15600) );
  AOI21_X1 U18863 ( .B1(n17979), .B2(n16231), .A(n15600), .ZN(n15601) );
  NAND2_X1 U18864 ( .A1(n18061), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16226) );
  OAI211_X1 U18865 ( .C1(n15602), .C2(n16224), .A(n15601), .B(n16226), .ZN(
        P3_U2832) );
  INV_X1 U18866 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20959) );
  OAI221_X1 U18867 ( .B1(n20662), .B2(HOLD), .C1(n20662), .C2(n20959), .A(
        P1_STATE_REG_1__SCAN_IN), .ZN(n15605) );
  INV_X1 U18868 ( .A(HOLD), .ZN(n20668) );
  OAI211_X1 U18869 ( .C1(n20959), .C2(n20668), .A(P1_STATE_REG_0__SCAN_IN), 
        .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n15603) );
  NAND3_X1 U18870 ( .A1(n15605), .A2(n15604), .A3(n15603), .ZN(P1_U3195) );
  INV_X1 U18871 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16346) );
  NOR2_X1 U18872 ( .A1(n19888), .A2(n16346), .ZN(P1_U2905) );
  NOR2_X1 U18873 ( .A1(n19733), .A2(n19727), .ZN(n19595) );
  NAND2_X1 U18874 ( .A1(n19595), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15607) );
  AND2_X1 U18875 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19699) );
  AOI21_X1 U18876 ( .B1(n19699), .B2(n19727), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15606) );
  AOI21_X1 U18877 ( .B1(n15607), .B2(n15606), .A(n16219), .ZN(P2_U3178) );
  INV_X1 U18878 ( .A(n16211), .ZN(n19718) );
  INV_X1 U18879 ( .A(n19713), .ZN(n19714) );
  NOR2_X1 U18880 ( .A1(n16204), .A2(n19714), .ZN(P2_U3047) );
  INV_X1 U18881 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17304) );
  NOR2_X2 U18882 ( .A1(n17096), .A2(n17304), .ZN(n17242) );
  INV_X1 U18883 ( .A(n17096), .ZN(n15612) );
  NAND2_X1 U18884 ( .A1(n17097), .A2(n15612), .ZN(n17182) );
  NAND2_X1 U18885 ( .A1(n15611), .A2(n15612), .ZN(n17239) );
  NAND2_X2 U18886 ( .A1(n18548), .A2(n15612), .ZN(n17231) );
  AOI22_X1 U18887 ( .A1(n17241), .A2(BUF2_REG_0__SCAN_IN), .B1(n17218), .B2(
        n17730), .ZN(n15613) );
  OAI221_X1 U18888 ( .B1(n17242), .B2(n17304), .C1(n17242), .C2(n17182), .A(
        n15613), .ZN(P3_U2735) );
  INV_X1 U18889 ( .A(n15614), .ZN(n15616) );
  AOI22_X1 U18890 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n15626), .B1(n15616), 
        .B2(n15615), .ZN(n15618) );
  AOI22_X1 U18891 ( .A1(n19858), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n19837), .B2(P1_EBX_REG_24__SCAN_IN), .ZN(n15617) );
  OAI211_X1 U18892 ( .C1(n15619), .C2(n19791), .A(n15618), .B(n15617), .ZN(
        n15620) );
  AOI21_X1 U18893 ( .B1(n15621), .B2(n19821), .A(n15620), .ZN(n15622) );
  OAI21_X1 U18894 ( .B1(n15623), .B2(n19851), .A(n15622), .ZN(P1_U2816) );
  AOI22_X1 U18895 ( .A1(n19865), .A2(n15624), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n19837), .ZN(n15633) );
  NOR2_X1 U18896 ( .A1(n15625), .A2(n15644), .ZN(n15635) );
  AOI21_X1 U18897 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n15635), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n15628) );
  INV_X1 U18898 ( .A(n15626), .ZN(n15627) );
  OAI22_X1 U18899 ( .A1(n15630), .A2(n15629), .B1(n15628), .B2(n15627), .ZN(
        n15631) );
  AOI21_X1 U18900 ( .B1(n19863), .B2(n15798), .A(n15631), .ZN(n15632) );
  OAI211_X1 U18901 ( .C1(n15634), .C2(n19840), .A(n15633), .B(n15632), .ZN(
        P1_U2817) );
  INV_X1 U18902 ( .A(n15635), .ZN(n15639) );
  INV_X1 U18903 ( .A(n15733), .ZN(n15636) );
  AOI22_X1 U18904 ( .A1(n19865), .A2(n15636), .B1(n19837), .B2(
        P1_EBX_REG_22__SCAN_IN), .ZN(n15638) );
  NAND2_X1 U18905 ( .A1(n19858), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15637) );
  OAI211_X1 U18906 ( .C1(n15639), .C2(P1_REIP_REG_22__SCAN_IN), .A(n15638), 
        .B(n15637), .ZN(n15640) );
  AOI21_X1 U18907 ( .B1(n15730), .B2(n19821), .A(n15640), .ZN(n15647) );
  AOI21_X1 U18908 ( .B1(n15643), .B2(n15642), .A(n15641), .ZN(n15661) );
  NOR3_X1 U18909 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n15645), .A3(n15644), 
        .ZN(n15651) );
  OAI21_X1 U18910 ( .B1(n15661), .B2(n15651), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15646) );
  OAI211_X1 U18911 ( .C1(n15648), .C2(n19791), .A(n15647), .B(n15646), .ZN(
        P1_U2818) );
  AOI22_X1 U18912 ( .A1(n19858), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n19837), .B2(P1_EBX_REG_21__SCAN_IN), .ZN(n15655) );
  AOI22_X1 U18913 ( .A1(n15734), .A2(n19865), .B1(P1_REIP_REG_21__SCAN_IN), 
        .B2(n15661), .ZN(n15654) );
  INV_X1 U18914 ( .A(n15649), .ZN(n15735) );
  AOI22_X1 U18915 ( .A1(n15735), .A2(n19821), .B1(n19863), .B2(n15650), .ZN(
        n15653) );
  INV_X1 U18916 ( .A(n15651), .ZN(n15652) );
  NAND4_X1 U18917 ( .A1(n15655), .A2(n15654), .A3(n15653), .A4(n15652), .ZN(
        P1_U2819) );
  INV_X1 U18918 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15656) );
  OAI222_X1 U18919 ( .A1(n15657), .A2(n19856), .B1(n19840), .B2(n15656), .C1(
        n15744), .C2(n19851), .ZN(n15658) );
  INV_X1 U18920 ( .A(n15658), .ZN(n15663) );
  OAI21_X1 U18921 ( .B1(n14821), .B2(n15659), .A(n20698), .ZN(n15660) );
  AOI22_X1 U18922 ( .A1(n15740), .A2(n19821), .B1(n15661), .B2(n15660), .ZN(
        n15662) );
  OAI211_X1 U18923 ( .C1(n19791), .C2(n15664), .A(n15663), .B(n15662), .ZN(
        P1_U2820) );
  AOI22_X1 U18924 ( .A1(n19837), .A2(P1_EBX_REG_18__SCAN_IN), .B1(n15665), 
        .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n15666) );
  OAI21_X1 U18925 ( .B1(n19851), .B2(n15667), .A(n15666), .ZN(n15668) );
  AOI211_X1 U18926 ( .C1(n19858), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n19836), .B(n15668), .ZN(n15672) );
  INV_X1 U18927 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20694) );
  AOI22_X1 U18928 ( .A1(n15670), .A2(n19821), .B1(n20694), .B2(n15669), .ZN(
        n15671) );
  OAI211_X1 U18929 ( .C1(n19791), .C2(n15811), .A(n15672), .B(n15671), .ZN(
        P1_U2822) );
  OAI21_X1 U18930 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n15673), .ZN(n15675) );
  NOR2_X1 U18931 ( .A1(n15675), .A2(n15674), .ZN(n15682) );
  NAND2_X1 U18932 ( .A1(n19837), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n15676) );
  NAND2_X1 U18933 ( .A1(n15676), .A2(n19777), .ZN(n15677) );
  AOI21_X1 U18934 ( .B1(n19858), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15677), .ZN(n15680) );
  INV_X1 U18935 ( .A(n15749), .ZN(n15678) );
  NAND2_X1 U18936 ( .A1(n19865), .A2(n15678), .ZN(n15679) );
  OAI211_X1 U18937 ( .C1(n15690), .C2(n20692), .A(n15680), .B(n15679), .ZN(
        n15681) );
  AOI211_X1 U18938 ( .C1(n15745), .C2(n19821), .A(n15682), .B(n15681), .ZN(
        n15683) );
  OAI21_X1 U18939 ( .B1(n19791), .B2(n15684), .A(n15683), .ZN(P1_U2824) );
  AOI21_X1 U18940 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15685), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15691) );
  AOI22_X1 U18941 ( .A1(n19858), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n19837), .B2(P1_EBX_REG_14__SCAN_IN), .ZN(n15686) );
  INV_X1 U18942 ( .A(n15686), .ZN(n15687) );
  AOI211_X1 U18943 ( .C1(n15834), .C2(n19863), .A(n19836), .B(n15687), .ZN(
        n15689) );
  AOI22_X1 U18944 ( .A1(n15755), .A2(n19821), .B1(n19865), .B2(n15754), .ZN(
        n15688) );
  OAI211_X1 U18945 ( .C1(n15691), .C2(n15690), .A(n15689), .B(n15688), .ZN(
        P1_U2826) );
  NOR2_X1 U18946 ( .A1(n19845), .A2(n15700), .ZN(n15699) );
  AOI21_X1 U18947 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15699), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15698) );
  AOI21_X1 U18948 ( .B1(n19837), .B2(P1_EBX_REG_12__SCAN_IN), .A(n19836), .ZN(
        n15693) );
  NAND2_X1 U18949 ( .A1(n19858), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15692) );
  OAI211_X1 U18950 ( .C1(n15860), .C2(n19791), .A(n15693), .B(n15692), .ZN(
        n15694) );
  INV_X1 U18951 ( .A(n15694), .ZN(n15696) );
  AOI22_X1 U18952 ( .A1(n15762), .A2(n19865), .B1(n19821), .B2(n15761), .ZN(
        n15695) );
  OAI211_X1 U18953 ( .C1(n15698), .C2(n15697), .A(n15696), .B(n15695), .ZN(
        P1_U2828) );
  INV_X1 U18954 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20686) );
  AOI22_X1 U18955 ( .A1(n19863), .A2(n15874), .B1(n15699), .B2(n20686), .ZN(
        n15704) );
  AOI21_X1 U18956 ( .B1(n19853), .B2(n15700), .A(n19803), .ZN(n15714) );
  AOI22_X1 U18957 ( .A1(n19858), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n19837), .B2(P1_EBX_REG_11__SCAN_IN), .ZN(n15701) );
  OAI211_X1 U18958 ( .C1(n20686), .C2(n15714), .A(n15701), .B(n19777), .ZN(
        n15702) );
  AOI21_X1 U18959 ( .B1(n19821), .B2(n15770), .A(n15702), .ZN(n15703) );
  OAI211_X1 U18960 ( .C1(n15773), .C2(n19851), .A(n15704), .B(n15703), .ZN(
        P1_U2829) );
  INV_X1 U18961 ( .A(n19774), .ZN(n19802) );
  NOR2_X1 U18962 ( .A1(n19845), .A2(n19802), .ZN(n19826) );
  AOI21_X1 U18963 ( .B1(n15705), .B2(n19826), .A(P1_REIP_REG_10__SCAN_IN), 
        .ZN(n15715) );
  INV_X1 U18964 ( .A(n15706), .ZN(n15887) );
  OAI22_X1 U18965 ( .A1(n15887), .A2(n19791), .B1(n15707), .B2(n19856), .ZN(
        n15708) );
  AOI211_X1 U18966 ( .C1(n19858), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19836), .B(n15708), .ZN(n15713) );
  INV_X1 U18967 ( .A(n15709), .ZN(n15710) );
  AOI22_X1 U18968 ( .A1(n15711), .A2(n19821), .B1(n15710), .B2(n19865), .ZN(
        n15712) );
  OAI211_X1 U18969 ( .C1(n15715), .C2(n15714), .A(n15713), .B(n15712), .ZN(
        P1_U2830) );
  INV_X1 U18970 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16283) );
  INV_X1 U18971 ( .A(n15716), .ZN(n15719) );
  AOI22_X1 U18972 ( .A1(n15719), .A2(n15718), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n15717), .ZN(n15722) );
  AOI22_X1 U18973 ( .A1(n15740), .A2(n15726), .B1(n15720), .B2(DATAI_20_), 
        .ZN(n15721) );
  OAI211_X1 U18974 ( .C1(n15723), .C2(n16283), .A(n15722), .B(n15721), .ZN(
        P1_U2884) );
  INV_X1 U18975 ( .A(n15724), .ZN(n19911) );
  AOI22_X1 U18976 ( .A1(n15761), .A2(n15726), .B1(n19911), .B2(n15725), .ZN(
        n15727) );
  OAI21_X1 U18977 ( .B1(n15728), .B2(n12045), .A(n15727), .ZN(P1_U2892) );
  AOI22_X1 U18978 ( .A1(n19936), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n19939), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15732) );
  AOI22_X1 U18979 ( .A1(n15730), .A2(n12940), .B1(n19938), .B2(n15729), .ZN(
        n15731) );
  OAI211_X1 U18980 ( .C1(n15787), .C2(n15733), .A(n15732), .B(n15731), .ZN(
        P1_U2977) );
  AOI22_X1 U18981 ( .A1(n19936), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n19939), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15737) );
  AOI22_X1 U18982 ( .A1(n15735), .A2(n12940), .B1(n15791), .B2(n15734), .ZN(
        n15736) );
  OAI211_X1 U18983 ( .C1(n19757), .C2(n15738), .A(n15737), .B(n15736), .ZN(
        P1_U2978) );
  AOI21_X1 U18984 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19936), .A(
        n15739), .ZN(n15743) );
  AOI22_X1 U18985 ( .A1(n15741), .A2(n19938), .B1(n15740), .B2(n12940), .ZN(
        n15742) );
  OAI211_X1 U18986 ( .C1(n15787), .C2(n15744), .A(n15743), .B(n15742), .ZN(
        P1_U2979) );
  AOI22_X1 U18987 ( .A1(n19936), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n19939), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15748) );
  AOI22_X1 U18988 ( .A1(n15746), .A2(n19938), .B1(n12940), .B2(n15745), .ZN(
        n15747) );
  OAI211_X1 U18989 ( .C1(n15787), .C2(n15749), .A(n15748), .B(n15747), .ZN(
        P1_U2983) );
  OAI21_X1 U18990 ( .B1(n15751), .B2(n15766), .A(n15750), .ZN(n15753) );
  XNOR2_X1 U18991 ( .A(n15766), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15752) );
  XNOR2_X1 U18992 ( .A(n15753), .B(n15752), .ZN(n15847) );
  AOI22_X1 U18993 ( .A1(n19936), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n19953), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15757) );
  AOI22_X1 U18994 ( .A1(n15755), .A2(n12940), .B1(n15791), .B2(n15754), .ZN(
        n15756) );
  OAI211_X1 U18995 ( .C1(n15847), .C2(n19757), .A(n15757), .B(n15756), .ZN(
        P1_U2985) );
  AOI21_X1 U18996 ( .B1(n15760), .B2(n15759), .A(n15758), .ZN(n15873) );
  AOI22_X1 U18997 ( .A1(n19936), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n19939), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15764) );
  AOI22_X1 U18998 ( .A1(n15791), .A2(n15762), .B1(n12940), .B2(n15761), .ZN(
        n15763) );
  OAI211_X1 U18999 ( .C1(n15873), .C2(n19757), .A(n15764), .B(n15763), .ZN(
        P1_U2987) );
  AOI22_X1 U19000 ( .A1(n19936), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n19953), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15772) );
  NOR2_X1 U19001 ( .A1(n14861), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15768) );
  NOR2_X1 U19002 ( .A1(n15765), .A2(n11696), .ZN(n15767) );
  MUX2_X1 U19003 ( .A(n15768), .B(n15767), .S(n9737), .Z(n15769) );
  XOR2_X1 U19004 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n15769), .Z(
        n15875) );
  AOI22_X1 U19005 ( .A1(n19938), .A2(n15875), .B1(n12940), .B2(n15770), .ZN(
        n15771) );
  OAI211_X1 U19006 ( .C1(n15787), .C2(n15773), .A(n15772), .B(n15771), .ZN(
        P1_U2988) );
  AOI22_X1 U19007 ( .A1(n19936), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n19953), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15779) );
  NAND2_X1 U19008 ( .A1(n15775), .A2(n15774), .ZN(n15776) );
  NAND2_X1 U19009 ( .A1(n15777), .A2(n15776), .ZN(n15918) );
  AOI22_X1 U19010 ( .A1(n15918), .A2(n19938), .B1(n12940), .B2(n19809), .ZN(
        n15778) );
  OAI211_X1 U19011 ( .C1(n15787), .C2(n19812), .A(n15779), .B(n15778), .ZN(
        P1_U2992) );
  INV_X1 U19012 ( .A(n15780), .ZN(n19825) );
  AOI22_X1 U19013 ( .A1(n19936), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n19953), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15786) );
  NAND2_X1 U19014 ( .A1(n15783), .A2(n15782), .ZN(n15784) );
  XNOR2_X1 U19015 ( .A(n15781), .B(n15784), .ZN(n15924) );
  AOI22_X1 U19016 ( .A1(n15924), .A2(n19938), .B1(n12940), .B2(n19822), .ZN(
        n15785) );
  OAI211_X1 U19017 ( .C1(n15787), .C2(n19825), .A(n15786), .B(n15785), .ZN(
        P1_U2993) );
  INV_X1 U19018 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19830) );
  INV_X1 U19019 ( .A(n15789), .ZN(n15790) );
  XNOR2_X1 U19020 ( .A(n15788), .B(n15790), .ZN(n15930) );
  INV_X1 U19021 ( .A(n19835), .ZN(n15792) );
  AOI222_X1 U19022 ( .A1(n15930), .A2(n19938), .B1(n12940), .B2(n19832), .C1(
        n15792), .C2(n15791), .ZN(n15794) );
  AND2_X1 U19023 ( .A1(n19953), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n15931) );
  INV_X1 U19024 ( .A(n15931), .ZN(n15793) );
  OAI211_X1 U19025 ( .C1(n19830), .C2(n15795), .A(n15794), .B(n15793), .ZN(
        P1_U2994) );
  AOI22_X1 U19026 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n15796), .B1(
        n19939), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n15801) );
  INV_X1 U19027 ( .A(n15797), .ZN(n15799) );
  AOI22_X1 U19028 ( .A1(n15799), .A2(n19965), .B1(n19964), .B2(n15798), .ZN(
        n15800) );
  OAI211_X1 U19029 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n15802), .A(
        n15801), .B(n15800), .ZN(P1_U3008) );
  AOI22_X1 U19030 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15803), .B1(
        n19953), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15807) );
  AOI22_X1 U19031 ( .A1(n15805), .A2(n19965), .B1(n19964), .B2(n15804), .ZN(
        n15806) );
  OAI211_X1 U19032 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15808), .A(
        n15807), .B(n15806), .ZN(P1_U3012) );
  AOI21_X1 U19033 ( .B1(n15907), .B2(n15810), .A(n15809), .ZN(n15824) );
  NOR3_X1 U19034 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15810), .A3(
        n15825), .ZN(n15814) );
  OAI22_X1 U19035 ( .A1(n15812), .A2(n15872), .B1(n15909), .B2(n15811), .ZN(
        n15813) );
  AOI211_X1 U19036 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n19939), .A(n15814), 
        .B(n15813), .ZN(n15815) );
  OAI21_X1 U19037 ( .B1(n15824), .B2(n15816), .A(n15815), .ZN(P1_U3013) );
  AOI21_X1 U19038 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15817), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15823) );
  INV_X1 U19039 ( .A(n15818), .ZN(n15820) );
  AOI22_X1 U19040 ( .A1(n15820), .A2(n19965), .B1(n19964), .B2(n15819), .ZN(
        n15822) );
  NAND2_X1 U19041 ( .A1(n19939), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15821) );
  OAI211_X1 U19042 ( .C1(n15824), .C2(n15823), .A(n15822), .B(n15821), .ZN(
        P1_U3014) );
  NOR2_X1 U19043 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15825), .ZN(
        n15826) );
  AOI21_X1 U19044 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n19939), .A(n15826), 
        .ZN(n15830) );
  AOI22_X1 U19045 ( .A1(n15828), .A2(n19965), .B1(n19964), .B2(n15827), .ZN(
        n15829) );
  OAI211_X1 U19046 ( .C1(n15832), .C2(n15831), .A(n15830), .B(n15829), .ZN(
        P1_U3016) );
  NAND2_X1 U19047 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15880) );
  OAI21_X1 U19048 ( .B1(n15880), .B2(n15900), .A(n15865), .ZN(n15928) );
  NAND2_X1 U19049 ( .A1(n15884), .A2(n15928), .ZN(n15927) );
  NOR3_X1 U19050 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15833), .A3(
        n15927), .ZN(n15838) );
  NAND2_X1 U19051 ( .A1(n15834), .A2(n19964), .ZN(n15836) );
  NAND2_X1 U19052 ( .A1(n19939), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n15835) );
  NAND2_X1 U19053 ( .A1(n15836), .A2(n15835), .ZN(n15837) );
  NOR2_X1 U19054 ( .A1(n15838), .A2(n15837), .ZN(n15846) );
  AND2_X1 U19055 ( .A1(n15751), .A2(n15839), .ZN(n15850) );
  OAI22_X1 U19056 ( .A1(n15849), .A2(n15848), .B1(n15840), .B2(n15853), .ZN(
        n15841) );
  AOI211_X1 U19057 ( .C1(n19945), .C2(n15843), .A(n15842), .B(n15841), .ZN(
        n15858) );
  INV_X1 U19058 ( .A(n15858), .ZN(n15844) );
  OAI21_X1 U19059 ( .B1(n15850), .B2(n15844), .A(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15845) );
  OAI211_X1 U19060 ( .C1(n15847), .C2(n15872), .A(n15846), .B(n15845), .ZN(
        P1_U3017) );
  NOR2_X1 U19061 ( .A1(n15849), .A2(n15848), .ZN(n15852) );
  NOR2_X1 U19062 ( .A1(n15908), .A2(n14167), .ZN(n15851) );
  AOI211_X1 U19063 ( .C1(n15853), .C2(n15852), .A(n15851), .B(n15850), .ZN(
        n15857) );
  AOI22_X1 U19064 ( .A1(n15855), .A2(n19965), .B1(n19964), .B2(n15854), .ZN(
        n15856) );
  OAI211_X1 U19065 ( .C1(n15858), .C2(n15751), .A(n15857), .B(n15856), .ZN(
        P1_U3018) );
  INV_X1 U19066 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15859) );
  OAI22_X1 U19067 ( .A1(n15860), .A2(n15909), .B1(n15908), .B2(n15859), .ZN(
        n15861) );
  INV_X1 U19068 ( .A(n15861), .ZN(n15871) );
  OR2_X1 U19069 ( .A1(n15863), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15879) );
  OAI21_X1 U19070 ( .B1(n15863), .B2(n15862), .A(n15902), .ZN(n15864) );
  OAI211_X1 U19071 ( .C1(n15868), .C2(n15865), .A(n15906), .B(n15864), .ZN(
        n15876) );
  INV_X1 U19072 ( .A(n15876), .ZN(n15866) );
  OAI21_X1 U19073 ( .B1(n15900), .B2(n15879), .A(n15866), .ZN(n15869) );
  NOR2_X1 U19074 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15927), .ZN(
        n15867) );
  AOI22_X1 U19075 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15869), .B1(
        n15868), .B2(n15867), .ZN(n15870) );
  OAI211_X1 U19076 ( .C1(n15873), .C2(n15872), .A(n15871), .B(n15870), .ZN(
        P1_U3019) );
  AOI22_X1 U19077 ( .A1(n15874), .A2(n19964), .B1(n19953), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n15878) );
  AOI22_X1 U19078 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15876), .B1(
        n19965), .B2(n15875), .ZN(n15877) );
  OAI211_X1 U19079 ( .C1(n15927), .C2(n15879), .A(n15878), .B(n15877), .ZN(
        P1_U3020) );
  NAND2_X1 U19080 ( .A1(n15884), .A2(n15885), .ZN(n15883) );
  NAND2_X1 U19081 ( .A1(n15902), .A2(n15880), .ZN(n15904) );
  NAND2_X1 U19082 ( .A1(n15881), .A2(n15904), .ZN(n19943) );
  OAI21_X1 U19083 ( .B1(n15883), .B2(n19943), .A(n15882), .ZN(n15899) );
  NAND3_X1 U19084 ( .A1(n15885), .A2(n15884), .A3(n15928), .ZN(n15893) );
  AOI221_X1 U19085 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n11696), .C2(n14006), .A(
        n15893), .ZN(n15889) );
  INV_X1 U19086 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n15886) );
  OAI22_X1 U19087 ( .A1(n15887), .A2(n15909), .B1(n15886), .B2(n15908), .ZN(
        n15888) );
  AOI211_X1 U19088 ( .C1(n15890), .C2(n19965), .A(n15889), .B(n15888), .ZN(
        n15891) );
  OAI21_X1 U19089 ( .B1(n11696), .B2(n15899), .A(n15891), .ZN(P1_U3021) );
  INV_X1 U19090 ( .A(n15892), .ZN(n15897) );
  NOR2_X1 U19091 ( .A1(n15893), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15896) );
  OAI22_X1 U19092 ( .A1(n15894), .A2(n15909), .B1(n14008), .B2(n15908), .ZN(
        n15895) );
  AOI211_X1 U19093 ( .C1(n15897), .C2(n19965), .A(n15896), .B(n15895), .ZN(
        n15898) );
  OAI21_X1 U19094 ( .B1(n14006), .B2(n15899), .A(n15898), .ZN(P1_U3022) );
  NAND2_X1 U19095 ( .A1(n15901), .A2(n11501), .ZN(n15937) );
  NAND2_X1 U19096 ( .A1(n15902), .A2(n19942), .ZN(n15903) );
  AND2_X1 U19097 ( .A1(n15904), .A2(n15903), .ZN(n15905) );
  AND2_X1 U19098 ( .A1(n15906), .A2(n15905), .ZN(n15934) );
  OAI21_X1 U19099 ( .B1(n15900), .B2(n15937), .A(n15934), .ZN(n15923) );
  AOI21_X1 U19100 ( .B1(n15912), .B2(n15907), .A(n15923), .ZN(n15922) );
  INV_X1 U19101 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20681) );
  OAI22_X1 U19102 ( .A1(n19790), .A2(n15909), .B1(n20681), .B2(n15908), .ZN(
        n15910) );
  AOI21_X1 U19103 ( .B1(n15911), .B2(n19965), .A(n15910), .ZN(n15914) );
  NOR2_X1 U19104 ( .A1(n15912), .A2(n15927), .ZN(n15917) );
  OAI221_X1 U19105 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n15915), .C2(n15921), .A(
        n15917), .ZN(n15913) );
  OAI211_X1 U19106 ( .C1(n15922), .C2(n15915), .A(n15914), .B(n15913), .ZN(
        P1_U3023) );
  INV_X1 U19107 ( .A(n15916), .ZN(n19801) );
  AOI22_X1 U19108 ( .A1(n19801), .A2(n19964), .B1(n19953), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n15920) );
  AOI22_X1 U19109 ( .A1(n15918), .A2(n19965), .B1(n15917), .B2(n15921), .ZN(
        n15919) );
  OAI211_X1 U19110 ( .C1(n15922), .C2(n15921), .A(n15920), .B(n15919), .ZN(
        P1_U3024) );
  AOI22_X1 U19111 ( .A1(n19814), .A2(n19964), .B1(n19953), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n15926) );
  AOI22_X1 U19112 ( .A1(n15924), .A2(n19965), .B1(n15923), .B2(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15925) );
  OAI211_X1 U19113 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n15927), .A(
        n15926), .B(n15925), .ZN(P1_U3025) );
  INV_X1 U19114 ( .A(n19944), .ZN(n15929) );
  NAND2_X1 U19115 ( .A1(n15929), .A2(n15928), .ZN(n19958) );
  NAND2_X1 U19116 ( .A1(n15930), .A2(n19965), .ZN(n15933) );
  AOI21_X1 U19117 ( .B1(n19827), .B2(n19964), .A(n15931), .ZN(n15932) );
  OAI211_X1 U19118 ( .C1(n11501), .C2(n15934), .A(n15933), .B(n15932), .ZN(
        n15935) );
  INV_X1 U19119 ( .A(n15935), .ZN(n15936) );
  OAI21_X1 U19120 ( .B1(n15937), .B2(n19958), .A(n15936), .ZN(P1_U3026) );
  NAND4_X1 U19121 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n20244), .A4(n20760), .ZN(n15938) );
  NAND2_X1 U19122 ( .A1(n15939), .A2(n15938), .ZN(n20650) );
  OAI21_X1 U19123 ( .B1(n15941), .B2(n20650), .A(n15940), .ZN(n15942) );
  OAI221_X1 U19124 ( .B1(n15943), .B2(n20446), .C1(n15943), .C2(n20760), .A(
        n15942), .ZN(n15944) );
  AOI221_X1 U19125 ( .B1(n15946), .B2(n20957), .C1(n15945), .C2(n20957), .A(
        n15944), .ZN(P1_U3162) );
  NOR2_X1 U19126 ( .A1(n15946), .A2(n15945), .ZN(n15948) );
  OAI21_X1 U19127 ( .B1(n15948), .B2(n20446), .A(n15947), .ZN(P1_U3466) );
  AOI211_X1 U19128 ( .C1(n15951), .C2(n15950), .A(n15949), .B(n19602), .ZN(
        n15960) );
  OAI22_X1 U19129 ( .A1(n18906), .A2(n15952), .B1(n18908), .B2(n9865), .ZN(
        n15956) );
  AOI211_X1 U19130 ( .C1(n15954), .C2(P2_EBX_REG_26__SCAN_IN), .A(n15953), .B(
        n18927), .ZN(n15955) );
  AOI211_X1 U19131 ( .C1(n18912), .C2(P2_REIP_REG_26__SCAN_IN), .A(n15956), 
        .B(n15955), .ZN(n15957) );
  OAI21_X1 U19132 ( .B1(n15958), .B2(n18900), .A(n15957), .ZN(n15959) );
  AOI211_X1 U19133 ( .C1(n18923), .C2(n15961), .A(n15960), .B(n15959), .ZN(
        n15962) );
  INV_X1 U19134 ( .A(n15962), .ZN(P2_U2829) );
  AOI22_X1 U19135 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n18922), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18912), .ZN(n15974) );
  AOI22_X1 U19136 ( .A1(n15963), .A2(n18885), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18939), .ZN(n15973) );
  INV_X1 U19137 ( .A(n15964), .ZN(n15966) );
  AOI22_X1 U19138 ( .A1(n15966), .A2(n18933), .B1(n15965), .B2(n18923), .ZN(
        n15972) );
  AOI21_X1 U19139 ( .B1(n15969), .B2(n15968), .A(n15967), .ZN(n15970) );
  NAND2_X1 U19140 ( .A1(n18917), .A2(n15970), .ZN(n15971) );
  NAND4_X1 U19141 ( .A1(n15974), .A2(n15973), .A3(n15972), .A4(n15971), .ZN(
        P2_U2831) );
  AOI22_X1 U19142 ( .A1(n18965), .A2(n15976), .B1(n15975), .B2(n13516), .ZN(
        P2_U2856) );
  AOI22_X1 U19143 ( .A1(n15977), .A2(n18966), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n13516), .ZN(n15978) );
  OAI21_X1 U19144 ( .B1(n13516), .B2(n16001), .A(n15978), .ZN(P2_U2865) );
  NAND2_X1 U19145 ( .A1(n15980), .A2(n15979), .ZN(n15981) );
  NAND2_X1 U19146 ( .A1(n15982), .A2(n15981), .ZN(n15993) );
  OAI22_X1 U19147 ( .A1(n15993), .A2(n18951), .B1(n18965), .B2(n15983), .ZN(
        n15984) );
  INV_X1 U19148 ( .A(n15984), .ZN(n15985) );
  OAI21_X1 U19149 ( .B1(n13516), .B2(n15986), .A(n15985), .ZN(P2_U2867) );
  OAI22_X1 U19150 ( .A1(n15988), .A2(n18951), .B1(n18965), .B2(n15987), .ZN(
        n15989) );
  INV_X1 U19151 ( .A(n15989), .ZN(n15990) );
  OAI21_X1 U19152 ( .B1(n13516), .B2(n15991), .A(n15990), .ZN(P2_U2869) );
  AOI22_X1 U19153 ( .A1(n15992), .A2(n18974), .B1(n18995), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n15999) );
  AOI22_X1 U19154 ( .A1(n18977), .A2(BUF1_REG_20__SCAN_IN), .B1(n18976), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n15998) );
  OAI22_X1 U19155 ( .A1(n15995), .A2(n15994), .B1(n18998), .B2(n15993), .ZN(
        n15996) );
  INV_X1 U19156 ( .A(n15996), .ZN(n15997) );
  NAND3_X1 U19157 ( .A1(n15999), .A2(n15998), .A3(n15997), .ZN(P2_U2899) );
  AOI22_X1 U19158 ( .A1(n19055), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19044), .ZN(n16009) );
  NAND2_X1 U19159 ( .A1(n16000), .A2(n14248), .ZN(n16006) );
  OR2_X1 U19160 ( .A1(n16001), .A2(n16077), .ZN(n16004) );
  NAND2_X1 U19161 ( .A1(n16002), .A2(n19056), .ZN(n16003) );
  OAI211_X1 U19162 ( .C1(n16006), .C2(n16005), .A(n16004), .B(n16003), .ZN(
        n16007) );
  INV_X1 U19163 ( .A(n16007), .ZN(n16008) );
  OAI211_X1 U19164 ( .C1(n19061), .C2(n16010), .A(n16009), .B(n16008), .ZN(
        P2_U2992) );
  AOI22_X1 U19165 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19044), .B1(n16090), 
        .B2(n18838), .ZN(n16015) );
  OAI22_X1 U19166 ( .A1(n16012), .A2(n16084), .B1(n16083), .B2(n16011), .ZN(
        n16013) );
  AOI21_X1 U19167 ( .B1(n19063), .B2(n18839), .A(n16013), .ZN(n16014) );
  OAI211_X1 U19168 ( .C1(n16100), .C2(n10809), .A(n16015), .B(n16014), .ZN(
        P2_U2999) );
  AOI22_X1 U19169 ( .A1(n19055), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19044), .ZN(n16022) );
  NAND2_X1 U19170 ( .A1(n16016), .A2(n19056), .ZN(n16018) );
  OR2_X1 U19171 ( .A1(n18955), .A2(n16077), .ZN(n16017) );
  OAI211_X1 U19172 ( .C1(n16019), .C2(n16083), .A(n16018), .B(n16017), .ZN(
        n16020) );
  INV_X1 U19173 ( .A(n16020), .ZN(n16021) );
  OAI211_X1 U19174 ( .C1(n19061), .C2(n18844), .A(n16022), .B(n16021), .ZN(
        P2_U3000) );
  AOI22_X1 U19175 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n16060), .B1(n16090), 
        .B2(n18859), .ZN(n16027) );
  OAI22_X1 U19176 ( .A1(n16024), .A2(n16084), .B1(n16083), .B2(n16023), .ZN(
        n16025) );
  AOI21_X1 U19177 ( .B1(n19063), .B2(n18860), .A(n16025), .ZN(n16026) );
  OAI211_X1 U19178 ( .C1(n16100), .C2(n18853), .A(n16027), .B(n16026), .ZN(
        P2_U3001) );
  AOI22_X1 U19179 ( .A1(n19055), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19044), .ZN(n16037) );
  NOR2_X1 U19180 ( .A1(n16029), .A2(n16028), .ZN(n16030) );
  XNOR2_X1 U19181 ( .A(n15395), .B(n16030), .ZN(n16111) );
  INV_X1 U19182 ( .A(n16111), .ZN(n16035) );
  INV_X1 U19183 ( .A(n18959), .ZN(n16034) );
  NAND2_X1 U19184 ( .A1(n16031), .A2(n10731), .ZN(n16032) );
  AOI222_X1 U19185 ( .A1(n16035), .A2(n19056), .B1(n19063), .B2(n16034), .C1(
        n14248), .C2(n16108), .ZN(n16036) );
  OAI211_X1 U19186 ( .C1(n19061), .C2(n16038), .A(n16037), .B(n16036), .ZN(
        P2_U3002) );
  AOI22_X1 U19187 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19044), .B1(n16090), 
        .B2(n16039), .ZN(n16046) );
  INV_X1 U19188 ( .A(n16040), .ZN(n16042) );
  OAI22_X1 U19189 ( .A1(n16042), .A2(n16083), .B1(n16041), .B2(n16084), .ZN(
        n16043) );
  AOI21_X1 U19190 ( .B1(n19063), .B2(n16044), .A(n16043), .ZN(n16045) );
  OAI211_X1 U19191 ( .C1(n16100), .C2(n10789), .A(n16046), .B(n16045), .ZN(
        P2_U3003) );
  AOI22_X1 U19192 ( .A1(n19055), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19044), .ZN(n16058) );
  OR2_X1 U19193 ( .A1(n15415), .A2(n16047), .ZN(n16049) );
  NAND2_X1 U19194 ( .A1(n16049), .A2(n16048), .ZN(n16054) );
  INV_X1 U19195 ( .A(n16050), .ZN(n16051) );
  NOR2_X1 U19196 ( .A1(n16052), .A2(n16051), .ZN(n16053) );
  XNOR2_X1 U19197 ( .A(n16054), .B(n16053), .ZN(n16122) );
  INV_X1 U19198 ( .A(n16122), .ZN(n16056) );
  INV_X1 U19199 ( .A(n16117), .ZN(n18961) );
  AND2_X1 U19200 ( .A1(n15437), .A2(n16114), .ZN(n16055) );
  NOR2_X1 U19201 ( .A1(n15423), .A2(n16055), .ZN(n16119) );
  AOI222_X1 U19202 ( .A1(n16056), .A2(n19056), .B1(n19063), .B2(n18961), .C1(
        n14248), .C2(n16119), .ZN(n16057) );
  OAI211_X1 U19203 ( .C1(n19061), .C2(n16059), .A(n16058), .B(n16057), .ZN(
        P2_U3004) );
  AOI22_X1 U19204 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n16060), .B1(n16090), 
        .B2(n18872), .ZN(n16065) );
  OAI22_X1 U19205 ( .A1(n16062), .A2(n16084), .B1(n16083), .B2(n16061), .ZN(
        n16063) );
  AOI21_X1 U19206 ( .B1(n19063), .B2(n18873), .A(n16063), .ZN(n16064) );
  OAI211_X1 U19207 ( .C1(n16100), .C2(n10781), .A(n16065), .B(n16064), .ZN(
        P2_U3005) );
  AOI22_X1 U19208 ( .A1(n19055), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19044), .ZN(n16080) );
  INV_X1 U19209 ( .A(n16067), .ZN(n16068) );
  XNOR2_X1 U19210 ( .A(n16066), .B(n16068), .ZN(n16125) );
  NAND2_X1 U19211 ( .A1(n16125), .A2(n14248), .ZN(n16076) );
  NAND2_X1 U19212 ( .A1(n14026), .A2(n16069), .ZN(n16074) );
  INV_X1 U19213 ( .A(n16070), .ZN(n16072) );
  NOR2_X1 U19214 ( .A1(n16072), .A2(n16071), .ZN(n16073) );
  XNOR2_X1 U19215 ( .A(n16074), .B(n16073), .ZN(n16129) );
  NAND2_X1 U19216 ( .A1(n16129), .A2(n19056), .ZN(n16075) );
  OAI211_X1 U19217 ( .C1(n16077), .C2(n16126), .A(n16076), .B(n16075), .ZN(
        n16078) );
  INV_X1 U19218 ( .A(n16078), .ZN(n16079) );
  OAI211_X1 U19219 ( .C1(n19061), .C2(n16081), .A(n16080), .B(n16079), .ZN(
        P2_U3006) );
  AOI22_X1 U19220 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19044), .B1(n16090), 
        .B2(n18915), .ZN(n16088) );
  OAI22_X1 U19221 ( .A1(n16085), .A2(n16084), .B1(n16083), .B2(n16082), .ZN(
        n16086) );
  AOI21_X1 U19222 ( .B1(n19063), .B2(n18916), .A(n16086), .ZN(n16087) );
  OAI211_X1 U19223 ( .C1(n16100), .C2(n10763), .A(n16088), .B(n16087), .ZN(
        P2_U3009) );
  AOI22_X1 U19224 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19044), .B1(n16090), 
        .B2(n16089), .ZN(n16099) );
  XNOR2_X1 U19225 ( .A(n16091), .B(n10262), .ZN(n16092) );
  XNOR2_X1 U19226 ( .A(n16093), .B(n16092), .ZN(n16159) );
  INV_X1 U19227 ( .A(n16159), .ZN(n16097) );
  NAND2_X1 U19228 ( .A1(n16094), .A2(n9825), .ZN(n16095) );
  AND2_X1 U19229 ( .A1(n16096), .A2(n16095), .ZN(n16154) );
  AOI222_X1 U19230 ( .A1(n16097), .A2(n19056), .B1(n10278), .B2(n19063), .C1(
        n14248), .C2(n16154), .ZN(n16098) );
  OAI211_X1 U19231 ( .C1(n16101), .C2(n16100), .A(n16099), .B(n16098), .ZN(
        P2_U3011) );
  INV_X1 U19232 ( .A(n16102), .ZN(n16106) );
  NAND2_X1 U19233 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19044), .ZN(n16104) );
  OAI211_X1 U19234 ( .C1(n16161), .C2(n18990), .A(n16104), .B(n16103), .ZN(
        n16105) );
  AOI21_X1 U19235 ( .B1(n16106), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n16105), .ZN(n16110) );
  NOR2_X1 U19236 ( .A1(n18959), .A2(n19072), .ZN(n16107) );
  AOI21_X1 U19237 ( .B1(n16108), .B2(n16153), .A(n16107), .ZN(n16109) );
  OAI211_X1 U19238 ( .C1(n16111), .C2(n16163), .A(n16110), .B(n16109), .ZN(
        P2_U3034) );
  NAND2_X1 U19239 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19044), .ZN(n16112) );
  OAI221_X1 U19240 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16115), 
        .C1(n16114), .C2(n16113), .A(n16112), .ZN(n16116) );
  AOI21_X1 U19241 ( .B1(n18991), .B2(n19067), .A(n16116), .ZN(n16121) );
  NOR2_X1 U19242 ( .A1(n16117), .A2(n19072), .ZN(n16118) );
  AOI21_X1 U19243 ( .B1(n16119), .B2(n16153), .A(n16118), .ZN(n16120) );
  OAI211_X1 U19244 ( .C1(n16122), .C2(n16163), .A(n16121), .B(n16120), .ZN(
        P2_U3036) );
  INV_X1 U19245 ( .A(n16123), .ZN(n16124) );
  AOI22_X1 U19246 ( .A1(n19067), .A2(n16124), .B1(P2_REIP_REG_8__SCAN_IN), 
        .B2(n19044), .ZN(n16138) );
  INV_X1 U19247 ( .A(n16125), .ZN(n16127) );
  OAI22_X1 U19248 ( .A1(n16127), .A2(n19074), .B1(n19072), .B2(n16126), .ZN(
        n16128) );
  AOI21_X1 U19249 ( .B1(n19069), .B2(n16129), .A(n16128), .ZN(n16137) );
  OAI21_X1 U19250 ( .B1(n16156), .B2(n16133), .A(n16130), .ZN(n16131) );
  INV_X1 U19251 ( .A(n16131), .ZN(n16142) );
  NOR3_X1 U19252 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n16133), .A3(
        n16132), .ZN(n16141) );
  OAI21_X1 U19253 ( .B1(n16142), .B2(n16141), .A(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16136) );
  NAND3_X1 U19254 ( .A1(n16134), .A2(n16155), .A3(n10643), .ZN(n16135) );
  NAND4_X1 U19255 ( .A1(n16138), .A2(n16137), .A3(n16136), .A4(n16135), .ZN(
        P2_U3038) );
  OAI22_X1 U19256 ( .A1(n16139), .A2(n16161), .B1(n19632), .B2(n18814), .ZN(
        n16140) );
  AOI211_X1 U19257 ( .C1(n16142), .C2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n16141), .B(n16140), .ZN(n16146) );
  AOI22_X1 U19258 ( .A1(n16144), .A2(n19069), .B1(n16143), .B2(n18881), .ZN(
        n16145) );
  OAI211_X1 U19259 ( .C1(n19074), .C2(n16147), .A(n16146), .B(n16145), .ZN(
        P2_U3039) );
  OAI22_X1 U19260 ( .A1(n16148), .A2(n19072), .B1(n10914), .B2(n18814), .ZN(
        n16149) );
  INV_X1 U19261 ( .A(n16149), .ZN(n16150) );
  OAI21_X1 U19262 ( .B1(n16151), .B2(n16161), .A(n16150), .ZN(n16152) );
  AOI21_X1 U19263 ( .B1(n16154), .B2(n16153), .A(n16152), .ZN(n16158) );
  AOI22_X1 U19264 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16156), .B1(
        n16155), .B2(n10262), .ZN(n16157) );
  OAI211_X1 U19265 ( .C1(n16159), .C2(n16163), .A(n16158), .B(n16157), .ZN(
        P2_U3043) );
  OAI22_X1 U19266 ( .A1(n14251), .A2(n19070), .B1(n19072), .B2(n13005), .ZN(
        n16165) );
  OAI22_X1 U19267 ( .A1(n16163), .A2(n16162), .B1(n16161), .B2(n16160), .ZN(
        n16164) );
  AOI211_X1 U19268 ( .C1(n14251), .C2(n19078), .A(n16165), .B(n16164), .ZN(
        n16167) );
  OAI211_X1 U19269 ( .C1(n19074), .C2(n16168), .A(n16167), .B(n16166), .ZN(
        P2_U3046) );
  INV_X1 U19270 ( .A(n16170), .ZN(n16200) );
  AOI22_X1 U19271 ( .A1(n16170), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n16169), .B2(n16200), .ZN(n16199) );
  OAI22_X1 U19272 ( .A1(n16200), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16171), .B2(n16170), .ZN(n16198) );
  INV_X1 U19273 ( .A(n16198), .ZN(n16177) );
  NAND2_X1 U19274 ( .A1(n16177), .A2(n19696), .ZN(n16178) );
  NAND2_X1 U19275 ( .A1(n16173), .A2(n19708), .ZN(n16175) );
  OAI22_X1 U19276 ( .A1(n16173), .A2(n19708), .B1(n19715), .B2(n16172), .ZN(
        n16174) );
  NAND2_X1 U19277 ( .A1(n16175), .A2(n16174), .ZN(n16176) );
  OAI211_X1 U19278 ( .C1(n16177), .C2(n19696), .A(n16176), .B(n16200), .ZN(
        n16179) );
  AND3_X1 U19279 ( .A1(n16199), .A2(n16178), .A3(n16179), .ZN(n16180) );
  OAI22_X1 U19280 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16180), .B1(
        n16199), .B2(n16179), .ZN(n16205) );
  INV_X1 U19281 ( .A(n16181), .ZN(n16182) );
  NAND2_X1 U19282 ( .A1(n16187), .A2(n16182), .ZN(n16185) );
  INV_X1 U19283 ( .A(n16183), .ZN(n16192) );
  NAND2_X1 U19284 ( .A1(n9729), .A2(n16192), .ZN(n16184) );
  OAI211_X1 U19285 ( .C1(n16187), .C2(n16186), .A(n16185), .B(n16184), .ZN(
        n16188) );
  INV_X1 U19286 ( .A(n16188), .ZN(n19723) );
  NAND2_X1 U19287 ( .A1(n16189), .A2(n10216), .ZN(n16197) );
  NAND2_X1 U19288 ( .A1(n16190), .A2(n19739), .ZN(n19734) );
  INV_X1 U19289 ( .A(n9729), .ZN(n16191) );
  AOI211_X1 U19290 ( .C1(n19726), .C2(n19734), .A(n16192), .B(n16191), .ZN(
        n18756) );
  OAI21_X1 U19291 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n18756), .ZN(n16196) );
  NAND3_X1 U19292 ( .A1(n16194), .A2(n19737), .A3(n16193), .ZN(n16195) );
  NAND4_X1 U19293 ( .A1(n19723), .A2(n16197), .A3(n16196), .A4(n16195), .ZN(
        n16203) );
  OAI22_X1 U19294 ( .A1(n16201), .A2(n16200), .B1(n16199), .B2(n16198), .ZN(
        n16202) );
  AOI211_X1 U19295 ( .C1(n16205), .C2(n16204), .A(n16203), .B(n16202), .ZN(
        n16218) );
  NAND2_X1 U19296 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19732), .ZN(n19599) );
  AOI21_X1 U19297 ( .B1(n16207), .B2(n16206), .A(n18755), .ZN(n16212) );
  INV_X1 U19298 ( .A(n16212), .ZN(n16208) );
  OAI21_X1 U19299 ( .B1(n19726), .B2(n19599), .A(n16208), .ZN(n16209) );
  AOI211_X1 U19300 ( .C1(n16219), .C2(n16211), .A(n16210), .B(n16209), .ZN(
        n16217) );
  NAND2_X1 U19301 ( .A1(n16218), .A2(n16212), .ZN(n16222) );
  NAND2_X1 U19302 ( .A1(n16222), .A2(n19031), .ZN(n19603) );
  INV_X1 U19303 ( .A(n19603), .ZN(n19598) );
  INV_X1 U19304 ( .A(n19742), .ZN(n16213) );
  OAI21_X1 U19305 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16214), .A(n16213), 
        .ZN(n16215) );
  OAI21_X1 U19306 ( .B1(n19598), .B2(n19726), .A(n16215), .ZN(n16216) );
  OAI211_X1 U19307 ( .C1(n16218), .C2(n18755), .A(n16217), .B(n16216), .ZN(
        P2_U3176) );
  INV_X1 U19308 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19546) );
  NOR2_X1 U19309 ( .A1(n16220), .A2(n16219), .ZN(n16221) );
  OAI21_X1 U19310 ( .B1(n19546), .B2(n16222), .A(n16221), .ZN(P2_U3593) );
  AOI21_X1 U19311 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16256), .A(
        n17735), .ZN(n16244) );
  AOI21_X1 U19312 ( .B1(n17640), .B2(n16246), .A(n16244), .ZN(n16235) );
  AOI22_X1 U19313 ( .A1(n17933), .A2(n17537), .B1(n17640), .B2(n17935), .ZN(
        n17598) );
  NOR3_X1 U19314 ( .A1(n16225), .A2(n16224), .A3(n17536), .ZN(n16230) );
  OAI221_X1 U19315 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16228), .C1(
        n16378), .C2(n16227), .A(n16226), .ZN(n16229) );
  AOI211_X1 U19316 ( .C1(n17530), .C2(n16377), .A(n16230), .B(n16229), .ZN(
        n16233) );
  NAND2_X1 U19317 ( .A1(n17639), .A2(n16231), .ZN(n16232) );
  OAI211_X1 U19318 ( .C1(n16235), .C2(n16234), .A(n16233), .B(n16232), .ZN(
        P3_U2800) );
  INV_X1 U19319 ( .A(n16236), .ZN(n16238) );
  OAI21_X1 U19320 ( .B1(n16238), .B2(n18190), .A(n16388), .ZN(n16239) );
  AOI22_X1 U19321 ( .A1(n18061), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n16240), 
        .B2(n16239), .ZN(n16251) );
  NAND2_X1 U19322 ( .A1(n16242), .A2(n16241), .ZN(n16243) );
  AOI22_X1 U19323 ( .A1(n17639), .A2(n16245), .B1(n16244), .B2(n16243), .ZN(
        n16250) );
  OAI211_X1 U19324 ( .C1(n16257), .C2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n17640), .B(n16246), .ZN(n16249) );
  OAI21_X1 U19325 ( .B1(n16247), .B2(n17530), .A(n16387), .ZN(n16248) );
  NAND4_X1 U19326 ( .A1(n16251), .A2(n16250), .A3(n16249), .A4(n16248), .ZN(
        P3_U2801) );
  NAND2_X1 U19327 ( .A1(n18061), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17372) );
  AOI21_X1 U19328 ( .B1(n17638), .B2(n17378), .A(n17377), .ZN(n17363) );
  AOI22_X1 U19329 ( .A1(n17638), .A2(n17366), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17636), .ZN(n17362) );
  NOR2_X1 U19330 ( .A1(n17363), .A2(n17362), .ZN(n17361) );
  OAI211_X1 U19331 ( .C1(n16260), .C2(n17378), .A(n16253), .B(n16252), .ZN(
        n16255) );
  OAI211_X1 U19332 ( .C1(n17361), .C2(n16255), .A(n16254), .B(n18042), .ZN(
        n16259) );
  INV_X1 U19333 ( .A(n17882), .ZN(n17934) );
  OAI22_X1 U19334 ( .A1(n16257), .A2(n17934), .B1(n16256), .B2(n18037), .ZN(
        n16258) );
  OAI211_X1 U19335 ( .C1(n16259), .C2(n16258), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17892), .ZN(n16265) );
  NOR3_X1 U19336 ( .A1(n17361), .A2(n17964), .A3(n16260), .ZN(n16262) );
  OAI22_X1 U19337 ( .A1(n18037), .A2(n17883), .B1(n17881), .B2(n17934), .ZN(
        n17843) );
  NOR2_X1 U19338 ( .A1(n17761), .A2(n17843), .ZN(n17806) );
  NOR2_X1 U19339 ( .A1(n17806), .A2(n18050), .ZN(n17773) );
  OAI211_X1 U19340 ( .C1(n16262), .C2(n17773), .A(n16261), .B(n17366), .ZN(
        n16264) );
  NAND3_X1 U19341 ( .A1(n17979), .A2(n17377), .A3(n17362), .ZN(n16263) );
  NAND4_X1 U19342 ( .A1(n17372), .A2(n16265), .A3(n16264), .A4(n16263), .ZN(
        P3_U2834) );
  NOR3_X1 U19343 ( .A1(P3_D_C_N_REG_SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), .A3(
        P3_BE_N_REG_0__SCAN_IN), .ZN(n16267) );
  NOR4_X1 U19344 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_2__SCAN_IN), 
        .A3(P3_BE_N_REG_3__SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16266) );
  NAND4_X1 U19345 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16267), .A3(n16266), .A4(
        U215), .ZN(U213) );
  INV_X1 U19346 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19005) );
  INV_X2 U19347 ( .A(U214), .ZN(n16309) );
  NOR2_X2 U19348 ( .A1(n16309), .A2(n16268), .ZN(n16310) );
  OAI222_X1 U19349 ( .A1(U212), .A2(n19005), .B1(n16313), .B2(n19124), .C1(
        U214), .C2(n16346), .ZN(U216) );
  INV_X1 U19350 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n19114) );
  AOI22_X1 U19351 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n16309), .ZN(n16269) );
  OAI21_X1 U19352 ( .B1(n19114), .B2(n16313), .A(n16269), .ZN(U217) );
  INV_X1 U19353 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n16343) );
  INV_X1 U19354 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n19109) );
  INV_X1 U19355 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n20987) );
  OAI222_X1 U19356 ( .A1(U212), .A2(n16343), .B1(n16313), .B2(n19109), .C1(
        U214), .C2(n20987), .ZN(U218) );
  INV_X1 U19357 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n19104) );
  AOI22_X1 U19358 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16309), .ZN(n16270) );
  OAI21_X1 U19359 ( .B1(n19104), .B2(n16313), .A(n16270), .ZN(U219) );
  INV_X1 U19360 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n19099) );
  AOI22_X1 U19361 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16309), .ZN(n16271) );
  OAI21_X1 U19362 ( .B1(n19099), .B2(n16313), .A(n16271), .ZN(U220) );
  INV_X1 U19363 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16273) );
  AOI22_X1 U19364 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16309), .ZN(n16272) );
  OAI21_X1 U19365 ( .B1(n16273), .B2(n16313), .A(n16272), .ZN(U221) );
  AOI222_X1 U19366 ( .A1(n16304), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(n16310), 
        .B2(BUF1_REG_25__SCAN_IN), .C1(n16309), .C2(P1_DATAO_REG_25__SCAN_IN), 
        .ZN(n16274) );
  INV_X1 U19367 ( .A(n16274), .ZN(U222) );
  AOI22_X1 U19368 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16309), .ZN(n16275) );
  OAI21_X1 U19369 ( .B1(n16276), .B2(n16313), .A(n16275), .ZN(U223) );
  INV_X1 U19370 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16278) );
  AOI22_X1 U19371 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16309), .ZN(n16277) );
  OAI21_X1 U19372 ( .B1(n16278), .B2(n16313), .A(n16277), .ZN(U224) );
  INV_X1 U19373 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16280) );
  AOI22_X1 U19374 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16309), .ZN(n16279) );
  OAI21_X1 U19375 ( .B1(n16280), .B2(n16313), .A(n16279), .ZN(U225) );
  AOI222_X1 U19376 ( .A1(n16304), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(n16310), 
        .B2(BUF1_REG_21__SCAN_IN), .C1(n16309), .C2(P1_DATAO_REG_21__SCAN_IN), 
        .ZN(n16281) );
  INV_X1 U19377 ( .A(n16281), .ZN(U226) );
  AOI22_X1 U19378 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16309), .ZN(n16282) );
  OAI21_X1 U19379 ( .B1(n16283), .B2(n16313), .A(n16282), .ZN(U227) );
  INV_X1 U19380 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20816) );
  AOI22_X1 U19381 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16309), .ZN(n16284) );
  OAI21_X1 U19382 ( .B1(n20816), .B2(n16313), .A(n16284), .ZN(U228) );
  INV_X1 U19383 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16286) );
  AOI22_X1 U19384 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16309), .ZN(n16285) );
  OAI21_X1 U19385 ( .B1(n16286), .B2(n16313), .A(n16285), .ZN(U229) );
  INV_X1 U19386 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16288) );
  AOI22_X1 U19387 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16309), .ZN(n16287) );
  OAI21_X1 U19388 ( .B1(n16288), .B2(n16313), .A(n16287), .ZN(U230) );
  AOI22_X1 U19389 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16309), .ZN(n16289) );
  OAI21_X1 U19390 ( .B1(n14738), .B2(n16313), .A(n16289), .ZN(U231) );
  AOI22_X1 U19391 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16309), .ZN(n16290) );
  OAI21_X1 U19392 ( .B1(n13257), .B2(n16313), .A(n16290), .ZN(U232) );
  AOI22_X1 U19393 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16309), .ZN(n16291) );
  OAI21_X1 U19394 ( .B1(n14685), .B2(n16313), .A(n16291), .ZN(U233) );
  INV_X1 U19395 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n20909) );
  AOI22_X1 U19396 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16310), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16304), .ZN(n16292) );
  OAI21_X1 U19397 ( .B1(n20909), .B2(U214), .A(n16292), .ZN(U234) );
  AOI22_X1 U19398 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16309), .ZN(n16293) );
  OAI21_X1 U19399 ( .B1(n16294), .B2(n16313), .A(n16293), .ZN(U235) );
  INV_X1 U19400 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n19015) );
  AOI22_X1 U19401 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16310), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16309), .ZN(n16295) );
  OAI21_X1 U19402 ( .B1(n19015), .B2(U212), .A(n16295), .ZN(U236) );
  AOI22_X1 U19403 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16309), .ZN(n16296) );
  OAI21_X1 U19404 ( .B1(n16297), .B2(n16313), .A(n16296), .ZN(U237) );
  INV_X1 U19405 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16323) );
  AOI22_X1 U19406 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16310), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16309), .ZN(n16298) );
  OAI21_X1 U19407 ( .B1(n16323), .B2(U212), .A(n16298), .ZN(U238) );
  INV_X1 U19408 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16300) );
  AOI22_X1 U19409 ( .A1(BUF1_REG_8__SCAN_IN), .A2(n16310), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16309), .ZN(n16299) );
  OAI21_X1 U19410 ( .B1(n16300), .B2(U212), .A(n16299), .ZN(U239) );
  INV_X1 U19411 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n21028) );
  AOI22_X1 U19412 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16310), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16304), .ZN(n16301) );
  OAI21_X1 U19413 ( .B1(n21028), .B2(U214), .A(n16301), .ZN(U240) );
  INV_X1 U19414 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16320) );
  AOI22_X1 U19415 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n16310), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16309), .ZN(n16302) );
  OAI21_X1 U19416 ( .B1(n16320), .B2(U212), .A(n16302), .ZN(U241) );
  INV_X1 U19417 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n20979) );
  AOI22_X1 U19418 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16310), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16304), .ZN(n16303) );
  OAI21_X1 U19419 ( .B1(n20979), .B2(U214), .A(n16303), .ZN(U242) );
  INV_X1 U19420 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16306) );
  AOI22_X1 U19421 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16304), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16309), .ZN(n16305) );
  OAI21_X1 U19422 ( .B1(n16306), .B2(n16313), .A(n16305), .ZN(U243) );
  INV_X1 U19423 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16317) );
  AOI22_X1 U19424 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16310), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16309), .ZN(n16307) );
  OAI21_X1 U19425 ( .B1(n16317), .B2(U212), .A(n16307), .ZN(U244) );
  INV_X1 U19426 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16316) );
  AOI22_X1 U19427 ( .A1(BUF1_REG_2__SCAN_IN), .A2(n16310), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16309), .ZN(n16308) );
  OAI21_X1 U19428 ( .B1(n16316), .B2(U212), .A(n16308), .ZN(U245) );
  INV_X1 U19429 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16315) );
  AOI22_X1 U19430 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16310), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16309), .ZN(n16311) );
  OAI21_X1 U19431 ( .B1(n16315), .B2(U212), .A(n16311), .ZN(U246) );
  INV_X1 U19432 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16314) );
  INV_X1 U19433 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16312) );
  INV_X1 U19434 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n20930) );
  OAI222_X1 U19435 ( .A1(U212), .A2(n16314), .B1(n16313), .B2(n16312), .C1(
        U214), .C2(n20930), .ZN(U247) );
  INV_X1 U19436 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18081) );
  AOI22_X1 U19437 ( .A1(n16345), .A2(n16314), .B1(n18081), .B2(U215), .ZN(U251) );
  INV_X1 U19438 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18089) );
  AOI22_X1 U19439 ( .A1(n16345), .A2(n16315), .B1(n18089), .B2(U215), .ZN(U252) );
  INV_X1 U19440 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18093) );
  AOI22_X1 U19441 ( .A1(n16345), .A2(n16316), .B1(n18093), .B2(U215), .ZN(U253) );
  INV_X1 U19442 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18098) );
  AOI22_X1 U19443 ( .A1(n16345), .A2(n16317), .B1(n18098), .B2(U215), .ZN(U254) );
  OAI22_X1 U19444 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16345), .ZN(n16318) );
  INV_X1 U19445 ( .A(n16318), .ZN(U255) );
  OAI22_X1 U19446 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16336), .ZN(n16319) );
  INV_X1 U19447 ( .A(n16319), .ZN(U256) );
  INV_X1 U19448 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18113) );
  AOI22_X1 U19449 ( .A1(n16345), .A2(n16320), .B1(n18113), .B2(U215), .ZN(U257) );
  OAI22_X1 U19450 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16336), .ZN(n16321) );
  INV_X1 U19451 ( .A(n16321), .ZN(U258) );
  OAI22_X1 U19452 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16336), .ZN(n16322) );
  INV_X1 U19453 ( .A(n16322), .ZN(U259) );
  INV_X1 U19454 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17341) );
  AOI22_X1 U19455 ( .A1(n16345), .A2(n16323), .B1(n17341), .B2(U215), .ZN(U260) );
  OAI22_X1 U19456 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16336), .ZN(n16324) );
  INV_X1 U19457 ( .A(n16324), .ZN(U261) );
  INV_X1 U19458 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17345) );
  AOI22_X1 U19459 ( .A1(n16345), .A2(n19015), .B1(n17345), .B2(U215), .ZN(U262) );
  OAI22_X1 U19460 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16336), .ZN(n16325) );
  INV_X1 U19461 ( .A(n16325), .ZN(U263) );
  OAI22_X1 U19462 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16336), .ZN(n16326) );
  INV_X1 U19463 ( .A(n16326), .ZN(U264) );
  OAI22_X1 U19464 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16336), .ZN(n16327) );
  INV_X1 U19465 ( .A(n16327), .ZN(U265) );
  OAI22_X1 U19466 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16345), .ZN(n16328) );
  INV_X1 U19467 ( .A(n16328), .ZN(U266) );
  OAI22_X1 U19468 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16336), .ZN(n16329) );
  INV_X1 U19469 ( .A(n16329), .ZN(U267) );
  OAI22_X1 U19470 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16345), .ZN(n16330) );
  INV_X1 U19471 ( .A(n16330), .ZN(U268) );
  OAI22_X1 U19472 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16336), .ZN(n16331) );
  INV_X1 U19473 ( .A(n16331), .ZN(U269) );
  OAI22_X1 U19474 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16345), .ZN(n16332) );
  INV_X1 U19475 ( .A(n16332), .ZN(U270) );
  OAI22_X1 U19476 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16345), .ZN(n16333) );
  INV_X1 U19477 ( .A(n16333), .ZN(U271) );
  INV_X1 U19478 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16334) );
  AOI22_X1 U19479 ( .A1(n16345), .A2(n16334), .B1(n14042), .B2(U215), .ZN(U272) );
  OAI22_X1 U19480 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16345), .ZN(n16335) );
  INV_X1 U19481 ( .A(n16335), .ZN(U273) );
  OAI22_X1 U19482 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16336), .ZN(n16337) );
  INV_X1 U19483 ( .A(n16337), .ZN(U274) );
  OAI22_X1 U19484 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16345), .ZN(n16338) );
  INV_X1 U19485 ( .A(n16338), .ZN(U275) );
  OAI22_X1 U19486 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16345), .ZN(n16339) );
  INV_X1 U19487 ( .A(n16339), .ZN(U276) );
  OAI22_X1 U19488 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16345), .ZN(n16340) );
  INV_X1 U19489 ( .A(n16340), .ZN(U277) );
  OAI22_X1 U19490 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16345), .ZN(n16341) );
  INV_X1 U19491 ( .A(n16341), .ZN(U278) );
  OAI22_X1 U19492 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16345), .ZN(n16342) );
  INV_X1 U19493 ( .A(n16342), .ZN(U279) );
  INV_X1 U19494 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n19110) );
  AOI22_X1 U19495 ( .A1(n16345), .A2(n16343), .B1(n19110), .B2(U215), .ZN(U280) );
  OAI22_X1 U19496 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16345), .ZN(n16344) );
  INV_X1 U19497 ( .A(n16344), .ZN(U281) );
  INV_X1 U19498 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19122) );
  AOI22_X1 U19499 ( .A1(n16345), .A2(n19005), .B1(n19122), .B2(U215), .ZN(U282) );
  INV_X1 U19500 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17249) );
  AOI222_X1 U19501 ( .A1(n19005), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16346), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n17249), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16347) );
  INV_X2 U19502 ( .A(n16349), .ZN(n16348) );
  INV_X1 U19503 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18625) );
  INV_X1 U19504 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19636) );
  AOI22_X1 U19505 ( .A1(n16348), .A2(n18625), .B1(n19636), .B2(n16349), .ZN(
        U347) );
  INV_X1 U19506 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n21056) );
  INV_X1 U19507 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19635) );
  AOI22_X1 U19508 ( .A1(n16348), .A2(n21056), .B1(n19635), .B2(n16349), .ZN(
        U348) );
  INV_X1 U19509 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18622) );
  INV_X1 U19510 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19634) );
  AOI22_X1 U19511 ( .A1(n16348), .A2(n18622), .B1(n19634), .B2(n16349), .ZN(
        U349) );
  INV_X1 U19512 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18620) );
  INV_X1 U19513 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19633) );
  AOI22_X1 U19514 ( .A1(n16348), .A2(n18620), .B1(n19633), .B2(n16349), .ZN(
        U350) );
  INV_X1 U19515 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18618) );
  INV_X1 U19516 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19631) );
  AOI22_X1 U19517 ( .A1(n16348), .A2(n18618), .B1(n19631), .B2(n16349), .ZN(
        U351) );
  INV_X1 U19518 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18616) );
  INV_X1 U19519 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19629) );
  AOI22_X1 U19520 ( .A1(n16348), .A2(n18616), .B1(n19629), .B2(n16349), .ZN(
        U352) );
  INV_X1 U19521 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18614) );
  INV_X1 U19522 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19627) );
  AOI22_X1 U19523 ( .A1(n16348), .A2(n18614), .B1(n19627), .B2(n16349), .ZN(
        U353) );
  INV_X1 U19524 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18612) );
  INV_X1 U19525 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19626) );
  AOI22_X1 U19526 ( .A1(n16348), .A2(n18612), .B1(n19626), .B2(n16349), .ZN(
        U354) );
  INV_X1 U19527 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18664) );
  INV_X1 U19528 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19670) );
  AOI22_X1 U19529 ( .A1(n16348), .A2(n18664), .B1(n19670), .B2(n16349), .ZN(
        U355) );
  INV_X1 U19530 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18662) );
  INV_X1 U19531 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19668) );
  AOI22_X1 U19532 ( .A1(n16348), .A2(n18662), .B1(n19668), .B2(n16349), .ZN(
        U356) );
  INV_X1 U19533 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18659) );
  INV_X1 U19534 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19666) );
  AOI22_X1 U19535 ( .A1(n16348), .A2(n18659), .B1(n19666), .B2(n16349), .ZN(
        U357) );
  INV_X1 U19536 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18657) );
  INV_X1 U19537 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19663) );
  AOI22_X1 U19538 ( .A1(n16348), .A2(n18657), .B1(n19663), .B2(n16349), .ZN(
        U358) );
  INV_X1 U19539 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18655) );
  INV_X1 U19540 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19662) );
  AOI22_X1 U19541 ( .A1(n16348), .A2(n18655), .B1(n19662), .B2(n16349), .ZN(
        U359) );
  INV_X1 U19542 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18653) );
  INV_X1 U19543 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19660) );
  AOI22_X1 U19544 ( .A1(n16348), .A2(n18653), .B1(n19660), .B2(n16349), .ZN(
        U360) );
  INV_X1 U19545 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18651) );
  INV_X1 U19546 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19658) );
  AOI22_X1 U19547 ( .A1(n16348), .A2(n18651), .B1(n19658), .B2(n16349), .ZN(
        U361) );
  INV_X1 U19548 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18648) );
  INV_X1 U19549 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19656) );
  AOI22_X1 U19550 ( .A1(n16348), .A2(n18648), .B1(n19656), .B2(n16349), .ZN(
        U362) );
  INV_X1 U19551 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18647) );
  INV_X1 U19552 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19654) );
  AOI22_X1 U19553 ( .A1(n16348), .A2(n18647), .B1(n19654), .B2(n16349), .ZN(
        U363) );
  INV_X1 U19554 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18644) );
  INV_X1 U19555 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19653) );
  AOI22_X1 U19556 ( .A1(n16348), .A2(n18644), .B1(n19653), .B2(n16349), .ZN(
        U364) );
  INV_X1 U19557 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18610) );
  INV_X1 U19558 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19625) );
  AOI22_X1 U19559 ( .A1(n16348), .A2(n18610), .B1(n19625), .B2(n16349), .ZN(
        U365) );
  INV_X1 U19560 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18643) );
  INV_X1 U19561 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19651) );
  AOI22_X1 U19562 ( .A1(n16348), .A2(n18643), .B1(n19651), .B2(n16349), .ZN(
        U366) );
  INV_X1 U19563 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18641) );
  INV_X1 U19564 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19649) );
  AOI22_X1 U19565 ( .A1(n16348), .A2(n18641), .B1(n19649), .B2(n16349), .ZN(
        U367) );
  INV_X1 U19566 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18640) );
  INV_X1 U19567 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19647) );
  AOI22_X1 U19568 ( .A1(n16348), .A2(n18640), .B1(n19647), .B2(n16349), .ZN(
        U368) );
  INV_X1 U19569 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18638) );
  INV_X1 U19570 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19645) );
  AOI22_X1 U19571 ( .A1(n16348), .A2(n18638), .B1(n19645), .B2(n16349), .ZN(
        U369) );
  INV_X1 U19572 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18636) );
  INV_X1 U19573 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n21063) );
  AOI22_X1 U19574 ( .A1(n16348), .A2(n18636), .B1(n21063), .B2(n16349), .ZN(
        U370) );
  INV_X1 U19575 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n20870) );
  INV_X1 U19576 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19643) );
  AOI22_X1 U19577 ( .A1(n16348), .A2(n20870), .B1(n19643), .B2(n16349), .ZN(
        U371) );
  INV_X1 U19578 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18633) );
  INV_X1 U19579 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19641) );
  AOI22_X1 U19580 ( .A1(n16348), .A2(n18633), .B1(n19641), .B2(n16349), .ZN(
        U372) );
  INV_X1 U19581 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18631) );
  INV_X1 U19582 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19640) );
  AOI22_X1 U19583 ( .A1(n16348), .A2(n18631), .B1(n19640), .B2(n16349), .ZN(
        U373) );
  INV_X1 U19584 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18629) );
  INV_X1 U19585 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19638) );
  AOI22_X1 U19586 ( .A1(n16348), .A2(n18629), .B1(n19638), .B2(n16349), .ZN(
        U374) );
  INV_X1 U19587 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18627) );
  INV_X1 U19588 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19637) );
  AOI22_X1 U19589 ( .A1(n16348), .A2(n18627), .B1(n19637), .B2(n16349), .ZN(
        U375) );
  INV_X1 U19590 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18608) );
  AOI22_X1 U19591 ( .A1(n16348), .A2(n18608), .B1(n19623), .B2(n16349), .ZN(
        U376) );
  INV_X1 U19592 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18607) );
  NAND2_X1 U19593 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18607), .ZN(n18599) );
  NAND2_X1 U19594 ( .A1(n18604), .A2(n16350), .ZN(n18594) );
  OAI21_X1 U19595 ( .B1(n18604), .B2(n18599), .A(n18594), .ZN(n18675) );
  AOI21_X1 U19596 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18675), .ZN(n16351) );
  INV_X1 U19597 ( .A(n16351), .ZN(P3_U2633) );
  INV_X1 U19598 ( .A(n16358), .ZN(n16352) );
  OAI21_X1 U19599 ( .B1(n16352), .B2(n17307), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16353) );
  OAI21_X1 U19600 ( .B1(n18742), .B2(n18732), .A(n16353), .ZN(P3_U2634) );
  INV_X1 U19601 ( .A(n18740), .ZN(n18739) );
  AOI21_X1 U19602 ( .B1(n18604), .B2(n18607), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16354) );
  AOI22_X1 U19603 ( .A1(n18739), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16354), 
        .B2(n18740), .ZN(P3_U2635) );
  OAI21_X1 U19604 ( .B1(n16355), .B2(BS16), .A(n18675), .ZN(n18673) );
  OAI21_X1 U19605 ( .B1(n18675), .B2(n16356), .A(n18673), .ZN(P3_U2636) );
  AND3_X1 U19606 ( .A1(n18519), .A2(n16358), .A3(n16357), .ZN(n18522) );
  NOR2_X1 U19607 ( .A1(n18522), .A2(n18579), .ZN(n18721) );
  OAI21_X1 U19608 ( .B1(n18721), .B2(n18068), .A(n16359), .ZN(P3_U2637) );
  NOR4_X1 U19609 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_20__SCAN_IN), .ZN(n16363) );
  NOR4_X1 U19610 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16362) );
  NOR4_X1 U19611 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n16361) );
  NOR4_X1 U19612 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16360) );
  NAND4_X1 U19613 ( .A1(n16363), .A2(n16362), .A3(n16361), .A4(n16360), .ZN(
        n16369) );
  NOR4_X1 U19614 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_31__SCAN_IN), .A3(P3_DATAWIDTH_REG_2__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16367) );
  AOI211_X1 U19615 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_19__SCAN_IN), .B(
        P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n16366) );
  NOR4_X1 U19616 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16365) );
  NOR4_X1 U19617 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16364) );
  NAND4_X1 U19618 ( .A1(n16367), .A2(n16366), .A3(n16365), .A4(n16364), .ZN(
        n16368) );
  NOR2_X1 U19619 ( .A1(n16369), .A2(n16368), .ZN(n18718) );
  INV_X1 U19620 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16371) );
  NOR3_X1 U19621 ( .A1(P3_DATAWIDTH_REG_0__SCAN_IN), .A2(
        P3_REIP_REG_0__SCAN_IN), .A3(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n16372)
         );
  OAI21_X1 U19622 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16372), .A(n18718), .ZN(
        n16370) );
  OAI21_X1 U19623 ( .B1(n18718), .B2(n16371), .A(n16370), .ZN(P3_U2638) );
  INV_X1 U19624 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18711) );
  INV_X1 U19625 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18674) );
  AOI21_X1 U19626 ( .B1(n18711), .B2(n18674), .A(n16372), .ZN(n16374) );
  INV_X1 U19627 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16373) );
  INV_X1 U19628 ( .A(n18718), .ZN(n18713) );
  AOI22_X1 U19629 ( .A1(n18718), .A2(n16374), .B1(n16373), .B2(n18713), .ZN(
        P3_U2639) );
  NAND2_X1 U19630 ( .A1(n16731), .A2(n16375), .ZN(n16392) );
  XOR2_X1 U19631 ( .A(n16377), .B(n16376), .Z(n16381) );
  INV_X1 U19632 ( .A(n18588), .ZN(n16713) );
  OAI22_X1 U19633 ( .A1(n16397), .A2(n18665), .B1(n16378), .B2(n16693), .ZN(
        n16379) );
  OAI21_X1 U19634 ( .B1(n16732), .B2(n16382), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16383) );
  OAI211_X1 U19635 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16392), .A(n16384), .B(
        n16383), .ZN(P3_U2641) );
  INV_X1 U19636 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18661) );
  AOI211_X1 U19637 ( .C1(n16387), .C2(n16386), .A(n16385), .B(n18588), .ZN(
        n16391) );
  NAND3_X1 U19638 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16411), .ZN(n16389) );
  OAI22_X1 U19639 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16389), .B1(n16388), 
        .B2(n16693), .ZN(n16390) );
  AOI211_X1 U19640 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16721), .A(n16391), .B(
        n16390), .ZN(n16396) );
  INV_X1 U19641 ( .A(n16392), .ZN(n16393) );
  OAI21_X1 U19642 ( .B1(n16400), .B2(n16394), .A(n16393), .ZN(n16395) );
  OAI211_X1 U19643 ( .C1(n16397), .C2(n18661), .A(n16396), .B(n16395), .ZN(
        P3_U2642) );
  INV_X1 U19644 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18656) );
  NOR2_X1 U19645 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18656), .ZN(n16398) );
  AOI22_X1 U19646 ( .A1(n16721), .A2(P3_EBX_REG_28__SCAN_IN), .B1(n16411), 
        .B2(n16398), .ZN(n16406) );
  AOI21_X1 U19647 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16399), .A(n16560), 
        .ZN(n16412) );
  AOI211_X1 U19648 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16413), .A(n16400), .B(
        n16706), .ZN(n16404) );
  AOI211_X1 U19649 ( .C1(n17360), .C2(n16402), .A(n16401), .B(n18588), .ZN(
        n16403) );
  AOI211_X1 U19650 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16412), .A(n16404), 
        .B(n16403), .ZN(n16405) );
  OAI211_X1 U19651 ( .C1(n20864), .C2(n16693), .A(n16406), .B(n16405), .ZN(
        P3_U2643) );
  AOI22_X1 U19652 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16725), .B1(
        n16721), .B2(P3_EBX_REG_27__SCAN_IN), .ZN(n16417) );
  AOI211_X1 U19653 ( .C1(n16409), .C2(n16408), .A(n16407), .B(n18588), .ZN(
        n16410) );
  AOI221_X1 U19654 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16412), .C1(n16411), 
        .C2(n16412), .A(n16410), .ZN(n16416) );
  OAI211_X1 U19655 ( .C1(n16419), .C2(n16414), .A(n16731), .B(n16413), .ZN(
        n16415) );
  NAND3_X1 U19656 ( .A1(n16417), .A2(n16416), .A3(n16415), .ZN(P3_U2644) );
  AOI22_X1 U19657 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16725), .B1(
        n16721), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16427) );
  INV_X1 U19658 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18652) );
  NAND2_X1 U19659 ( .A1(n16723), .A2(n16418), .ZN(n16431) );
  INV_X1 U19660 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18654) );
  OAI21_X1 U19661 ( .B1(n18652), .B2(n16431), .A(n18654), .ZN(n16424) );
  AOI211_X1 U19662 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16434), .A(n16419), .B(
        n16706), .ZN(n16423) );
  AOI211_X1 U19663 ( .C1(n17391), .C2(n16421), .A(n16420), .B(n18588), .ZN(
        n16422) );
  AOI211_X1 U19664 ( .C1(n16425), .C2(n16424), .A(n16423), .B(n16422), .ZN(
        n16426) );
  NAND2_X1 U19665 ( .A1(n16427), .A2(n16426), .ZN(P3_U2645) );
  AOI21_X1 U19666 ( .B1(n16438), .B2(n16723), .A(n16720), .ZN(n16459) );
  INV_X1 U19667 ( .A(n16459), .ZN(n16447) );
  AOI21_X1 U19668 ( .B1(n16723), .B2(n18650), .A(n16447), .ZN(n16437) );
  AOI211_X1 U19669 ( .C1(n16430), .C2(n16429), .A(n16428), .B(n18588), .ZN(
        n16433) );
  OAI22_X1 U19670 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16431), .B1(n20821), 
        .B2(n16692), .ZN(n16432) );
  AOI211_X1 U19671 ( .C1(n16725), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16433), .B(n16432), .ZN(n16436) );
  OAI211_X1 U19672 ( .C1(n16441), .C2(n20821), .A(n16731), .B(n16434), .ZN(
        n16435) );
  OAI211_X1 U19673 ( .C1(n16437), .C2(n18652), .A(n16436), .B(n16435), .ZN(
        P3_U2646) );
  INV_X1 U19674 ( .A(n16438), .ZN(n16440) );
  NOR2_X1 U19675 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16704), .ZN(n16439) );
  AOI22_X1 U19676 ( .A1(n16721), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16440), 
        .B2(n16439), .ZN(n16449) );
  AOI211_X1 U19677 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16455), .A(n16441), .B(
        n16706), .ZN(n16446) );
  INV_X1 U19678 ( .A(n16442), .ZN(n16443) );
  AOI211_X1 U19679 ( .C1(n17413), .C2(n16444), .A(n16443), .B(n18588), .ZN(
        n16445) );
  AOI211_X1 U19680 ( .C1(n16447), .C2(P3_REIP_REG_24__SCAN_IN), .A(n16446), 
        .B(n16445), .ZN(n16448) );
  OAI211_X1 U19681 ( .C1(n20851), .C2(n16693), .A(n16449), .B(n16448), .ZN(
        P3_U2647) );
  AOI21_X1 U19682 ( .B1(n16723), .B2(n16450), .A(P3_REIP_REG_23__SCAN_IN), 
        .ZN(n16460) );
  AOI211_X1 U19683 ( .C1(n17427), .C2(n16452), .A(n16451), .B(n18588), .ZN(
        n16454) );
  OAI22_X1 U19684 ( .A1(n17422), .A2(n16693), .B1(n16692), .B2(n16456), .ZN(
        n16453) );
  NOR2_X1 U19685 ( .A1(n16454), .A2(n16453), .ZN(n16458) );
  OAI211_X1 U19686 ( .C1(n16461), .C2(n16456), .A(n16731), .B(n16455), .ZN(
        n16457) );
  OAI211_X1 U19687 ( .C1(n16460), .C2(n16459), .A(n16458), .B(n16457), .ZN(
        P3_U2648) );
  AOI211_X1 U19688 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16480), .A(n16461), .B(
        n16706), .ZN(n16462) );
  AOI21_X1 U19689 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n16721), .A(n16462), .ZN(
        n16473) );
  INV_X1 U19690 ( .A(n16463), .ZN(n16464) );
  AOI211_X1 U19691 ( .C1(n17455), .C2(n16465), .A(n16464), .B(n18588), .ZN(
        n16468) );
  NOR3_X1 U19692 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16704), .A3(n16466), 
        .ZN(n16467) );
  AOI211_X1 U19693 ( .C1(n16725), .C2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16468), .B(n16467), .ZN(n16472) );
  OAI21_X1 U19694 ( .B1(n16469), .B2(n16704), .A(n16733), .ZN(n16479) );
  INV_X1 U19695 ( .A(n16479), .ZN(n16493) );
  INV_X1 U19696 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18645) );
  NAND3_X1 U19697 ( .A1(n18645), .A2(n16723), .A3(n16469), .ZN(n16476) );
  AOI21_X1 U19698 ( .B1(n16493), .B2(n16476), .A(n18646), .ZN(n16470) );
  INV_X1 U19699 ( .A(n16470), .ZN(n16471) );
  NAND3_X1 U19700 ( .A1(n16473), .A2(n16472), .A3(n16471), .ZN(P3_U2649) );
  AOI211_X1 U19701 ( .C1(n17461), .C2(n16475), .A(n16474), .B(n18588), .ZN(
        n16478) );
  OAI21_X1 U19702 ( .B1(n16693), .B2(n17458), .A(n16476), .ZN(n16477) );
  AOI211_X1 U19703 ( .C1(n16479), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16478), 
        .B(n16477), .ZN(n16482) );
  OAI211_X1 U19704 ( .C1(n16488), .C2(n16883), .A(n16731), .B(n16480), .ZN(
        n16481) );
  OAI211_X1 U19705 ( .C1(n16883), .C2(n16692), .A(n16482), .B(n16481), .ZN(
        P3_U2650) );
  AOI211_X1 U19706 ( .C1(n16485), .C2(n16484), .A(n16483), .B(n18588), .ZN(
        n16486) );
  AOI21_X1 U19707 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16721), .A(n16486), .ZN(
        n16492) );
  NOR3_X1 U19708 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16704), .A3(n16487), 
        .ZN(n16490) );
  AOI211_X1 U19709 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16501), .A(n16488), .B(
        n16706), .ZN(n16489) );
  AOI211_X1 U19710 ( .C1(n16725), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16490), .B(n16489), .ZN(n16491) );
  OAI211_X1 U19711 ( .C1(n20847), .C2(n16493), .A(n16492), .B(n16491), .ZN(
        P3_U2651) );
  AOI22_X1 U19712 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n16725), .B1(
        n16721), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n16505) );
  NOR2_X1 U19713 ( .A1(n16506), .A2(n16519), .ZN(n16495) );
  INV_X1 U19714 ( .A(n16494), .ZN(n17443) );
  OAI21_X1 U19715 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16495), .A(
        n17443), .ZN(n17490) );
  NOR2_X1 U19716 ( .A1(n16496), .A2(n16688), .ZN(n16497) );
  XNOR2_X1 U19717 ( .A(n17490), .B(n16497), .ZN(n16498) );
  AOI21_X1 U19718 ( .B1(n16498), .B2(n16713), .A(n18061), .ZN(n16504) );
  OAI21_X1 U19719 ( .B1(n16499), .B2(n16704), .A(n16733), .ZN(n16525) );
  INV_X1 U19720 ( .A(n16499), .ZN(n16516) );
  NOR2_X1 U19721 ( .A1(n16704), .A2(n16516), .ZN(n16512) );
  INV_X1 U19722 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18642) );
  INV_X1 U19723 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18639) );
  XOR2_X1 U19724 ( .A(n18642), .B(n18639), .Z(n16500) );
  AOI22_X1 U19725 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16525), .B1(n16512), 
        .B2(n16500), .ZN(n16503) );
  OAI211_X1 U19726 ( .C1(n16509), .C2(n20935), .A(n16731), .B(n16501), .ZN(
        n16502) );
  NAND4_X1 U19727 ( .A1(n16505), .A2(n16504), .A3(n16503), .A4(n16502), .ZN(
        P3_U2652) );
  AOI22_X1 U19728 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16725), .B1(
        n16721), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n16515) );
  AOI22_X1 U19729 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16519), .B1(
        n17486), .B2(n16506), .ZN(n17498) );
  NAND2_X1 U19730 ( .A1(n9710), .A2(n16507), .ZN(n16508) );
  XOR2_X1 U19731 ( .A(n17498), .B(n16508), .Z(n16511) );
  AOI211_X1 U19732 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16526), .A(n16509), .B(
        n16706), .ZN(n16510) );
  AOI211_X1 U19733 ( .C1(n16713), .C2(n16511), .A(n18061), .B(n16510), .ZN(
        n16514) );
  AOI22_X1 U19734 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16525), .B1(n16512), 
        .B2(n18639), .ZN(n16513) );
  NAND3_X1 U19735 ( .A1(n16515), .A2(n16514), .A3(n16513), .ZN(P3_U2653) );
  NAND2_X1 U19736 ( .A1(n16723), .A2(n16516), .ZN(n16522) );
  OR2_X1 U19737 ( .A1(n16517), .A2(n16688), .ZN(n16533) );
  INV_X1 U19738 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17526) );
  NOR2_X1 U19739 ( .A1(n17727), .A2(n17631), .ZN(n16602) );
  INV_X1 U19740 ( .A(n16602), .ZN(n16651) );
  NOR2_X1 U19741 ( .A1(n16518), .A2(n16651), .ZN(n16601) );
  NAND2_X1 U19742 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16601), .ZN(
        n16582) );
  OR2_X1 U19743 ( .A1(n17573), .A2(n16582), .ZN(n16571) );
  NOR2_X1 U19744 ( .A1(n17553), .A2(n16571), .ZN(n17528) );
  NAND2_X1 U19745 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17528), .ZN(
        n16542) );
  NOR2_X1 U19746 ( .A1(n17526), .A2(n16542), .ZN(n16531) );
  OAI21_X1 U19747 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16531), .A(
        n16519), .ZN(n17519) );
  XOR2_X1 U19748 ( .A(n16533), .B(n17519), .Z(n16520) );
  AOI22_X1 U19749 ( .A1(n16721), .A2(P3_EBX_REG_17__SCAN_IN), .B1(n16713), 
        .B2(n16520), .ZN(n16521) );
  OAI211_X1 U19750 ( .C1(n16523), .C2(n16522), .A(n16521), .B(n17892), .ZN(
        n16524) );
  AOI21_X1 U19751 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n16525), .A(n16524), 
        .ZN(n16529) );
  OAI211_X1 U19752 ( .C1(n16530), .C2(n16527), .A(n16731), .B(n16526), .ZN(
        n16528) );
  OAI211_X1 U19753 ( .C1(n16693), .C2(n17513), .A(n16529), .B(n16528), .ZN(
        P3_U2654) );
  AOI211_X1 U19754 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16549), .A(n16530), .B(
        n16706), .ZN(n16537) );
  INV_X1 U19755 ( .A(n17524), .ZN(n17527) );
  NOR2_X1 U19756 ( .A1(n17527), .A2(n16674), .ZN(n16544) );
  AOI21_X1 U19757 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n16544), .A(
        n16688), .ZN(n16543) );
  AOI21_X1 U19758 ( .B1(n17526), .B2(n16542), .A(n16531), .ZN(n17529) );
  INV_X1 U19759 ( .A(n17529), .ZN(n16532) );
  AOI221_X1 U19760 ( .B1(n16543), .B2(n17529), .C1(n16533), .C2(n16532), .A(
        n18588), .ZN(n16536) );
  INV_X1 U19761 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n21055) );
  INV_X1 U19762 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18635) );
  OAI21_X1 U19763 ( .B1(n16704), .B2(n16538), .A(n16733), .ZN(n16534) );
  INV_X1 U19764 ( .A(n16534), .ZN(n16553) );
  OAI22_X1 U19765 ( .A1(n16692), .A2(n21055), .B1(n18635), .B2(n16553), .ZN(
        n16535) );
  NOR4_X1 U19766 ( .A1(n18061), .A2(n16537), .A3(n16536), .A4(n16535), .ZN(
        n16540) );
  NAND3_X1 U19767 ( .A1(n16723), .A2(n16538), .A3(n18635), .ZN(n16539) );
  OAI211_X1 U19768 ( .C1(n16693), .C2(n17526), .A(n16540), .B(n16539), .ZN(
        P3_U2655) );
  OAI21_X1 U19769 ( .B1(n16704), .B2(n16558), .A(n18634), .ZN(n16541) );
  INV_X1 U19770 ( .A(n16541), .ZN(n16554) );
  OAI21_X1 U19771 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17528), .A(
        n16542), .ZN(n17538) );
  INV_X1 U19772 ( .A(n16543), .ZN(n16546) );
  NAND2_X1 U19773 ( .A1(n16688), .A2(n16713), .ZN(n16644) );
  OAI21_X1 U19774 ( .B1(n16544), .B2(n17538), .A(n16713), .ZN(n16545) );
  AOI22_X1 U19775 ( .A1(n17538), .A2(n16546), .B1(n16644), .B2(n16545), .ZN(
        n16548) );
  OAI21_X1 U19776 ( .B1(n16692), .B2(n16550), .A(n17892), .ZN(n16547) );
  AOI211_X1 U19777 ( .C1(n16725), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16548), .B(n16547), .ZN(n16552) );
  OAI211_X1 U19778 ( .C1(n16566), .C2(n16550), .A(n16731), .B(n16549), .ZN(
        n16551) );
  OAI211_X1 U19779 ( .C1(n16554), .C2(n16553), .A(n16552), .B(n16551), .ZN(
        P3_U2656) );
  AOI21_X1 U19780 ( .B1(n16576), .B2(P3_EBX_REG_14__SCAN_IN), .A(n16706), .ZN(
        n16555) );
  AOI21_X1 U19781 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n16721), .A(n16555), .ZN(
        n16565) );
  OAI21_X1 U19782 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16571), .A(
        n9710), .ZN(n16556) );
  AOI21_X1 U19783 ( .B1(n17553), .B2(n16571), .A(n17528), .ZN(n17555) );
  XOR2_X1 U19784 ( .A(n16556), .B(n17555), .Z(n16557) );
  OAI21_X1 U19785 ( .B1(n16557), .B2(n18588), .A(n18044), .ZN(n16563) );
  NAND3_X1 U19786 ( .A1(n16723), .A2(P3_REIP_REG_13__SCAN_IN), .A3(n16568), 
        .ZN(n16561) );
  INV_X1 U19787 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18632) );
  NOR2_X1 U19788 ( .A1(n16720), .A2(n16558), .ZN(n16559) );
  AOI211_X1 U19789 ( .C1(n16561), .C2(n18632), .A(n16560), .B(n16559), .ZN(
        n16562) );
  AOI211_X1 U19790 ( .C1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n16725), .A(
        n16563), .B(n16562), .ZN(n16564) );
  OAI21_X1 U19791 ( .B1(n16566), .B2(n16565), .A(n16564), .ZN(P3_U2657) );
  INV_X1 U19792 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16579) );
  INV_X1 U19793 ( .A(n16567), .ZN(n16586) );
  OAI21_X1 U19794 ( .B1(n16586), .B2(n16704), .A(n16733), .ZN(n16597) );
  NOR2_X1 U19795 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16704), .ZN(n16585) );
  NAND2_X1 U19796 ( .A1(n16723), .A2(n16568), .ZN(n16574) );
  AOI21_X1 U19797 ( .B1(n9710), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18588), .ZN(n16719) );
  INV_X1 U19798 ( .A(n16719), .ZN(n16653) );
  INV_X1 U19799 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17586) );
  NOR2_X1 U19800 ( .A1(n17586), .A2(n16582), .ZN(n16569) );
  OAI21_X1 U19801 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16569), .A(
        n16571), .ZN(n17576) );
  AOI211_X1 U19802 ( .C1(n9710), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16653), .B(n17576), .ZN(n16570) );
  AOI211_X1 U19803 ( .C1(n16721), .C2(P3_EBX_REG_13__SCAN_IN), .A(n18061), .B(
        n16570), .ZN(n16573) );
  OAI211_X1 U19804 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n16571), .A(
        n16724), .B(n17576), .ZN(n16572) );
  OAI211_X1 U19805 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16574), .A(n16573), 
        .B(n16572), .ZN(n16575) );
  AOI221_X1 U19806 ( .B1(n16597), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n16585), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n16575), .ZN(n16578) );
  OAI211_X1 U19807 ( .C1(n16580), .C2(n20869), .A(n16731), .B(n16576), .ZN(
        n16577) );
  OAI211_X1 U19808 ( .C1(n16693), .C2(n16579), .A(n16578), .B(n16577), .ZN(
        P3_U2658) );
  AOI211_X1 U19809 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16593), .A(n16580), .B(
        n16706), .ZN(n16581) );
  AOI21_X1 U19810 ( .B1(n16725), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16581), .ZN(n16589) );
  INV_X1 U19811 ( .A(n16582), .ZN(n17570) );
  AOI22_X1 U19812 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16582), .B1(
        n17570), .B2(n17586), .ZN(n17582) );
  INV_X1 U19813 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n20986) );
  NAND2_X1 U19814 ( .A1(n17592), .A2(n16714), .ZN(n16590) );
  OAI21_X1 U19815 ( .B1(n20986), .B2(n16590), .A(n9710), .ZN(n16583) );
  XOR2_X1 U19816 ( .A(n17582), .B(n16583), .Z(n16584) );
  AOI22_X1 U19817 ( .A1(n16721), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n16713), 
        .B2(n16584), .ZN(n16588) );
  AOI22_X1 U19818 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16597), .B1(n16586), 
        .B2(n16585), .ZN(n16587) );
  NAND4_X1 U19819 ( .A1(n16589), .A2(n16588), .A3(n16587), .A4(n17892), .ZN(
        P3_U2659) );
  NAND2_X1 U19820 ( .A1(n9710), .A2(n16590), .ZN(n16592) );
  INV_X1 U19821 ( .A(n16601), .ZN(n16591) );
  AOI21_X1 U19822 ( .B1(n20986), .B2(n16591), .A(n17570), .ZN(n17595) );
  XOR2_X1 U19823 ( .A(n16592), .B(n17595), .Z(n16595) );
  OAI211_X1 U19824 ( .C1(n16609), .C2(n20970), .A(n16731), .B(n16593), .ZN(
        n16594) );
  OAI21_X1 U19825 ( .B1(n16595), .B2(n18588), .A(n16594), .ZN(n16596) );
  AOI211_X1 U19826 ( .C1(n16721), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18061), .B(
        n16596), .ZN(n16600) );
  OAI221_X1 U19827 ( .B1(P3_REIP_REG_11__SCAN_IN), .B2(n16723), .C1(
        P3_REIP_REG_11__SCAN_IN), .C2(n16598), .A(n16597), .ZN(n16599) );
  OAI211_X1 U19828 ( .C1(n16693), .C2(n20986), .A(n16600), .B(n16599), .ZN(
        P3_U2660) );
  INV_X1 U19829 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n20951) );
  NAND2_X1 U19830 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16603) );
  NOR2_X1 U19831 ( .A1(n16603), .A2(n16651), .ZN(n16629) );
  NAND2_X1 U19832 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16629), .ZN(
        n16615) );
  AOI21_X1 U19833 ( .B1(n20951), .B2(n16615), .A(n16601), .ZN(n17607) );
  INV_X1 U19834 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16623) );
  INV_X1 U19835 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16689) );
  NAND2_X1 U19836 ( .A1(n16602), .A2(n16689), .ZN(n16652) );
  NOR3_X1 U19837 ( .A1(n16603), .A2(n16623), .A3(n16652), .ZN(n16618) );
  NOR2_X1 U19838 ( .A1(n16618), .A2(n16688), .ZN(n16604) );
  XOR2_X1 U19839 ( .A(n17607), .B(n16604), .Z(n16607) );
  NOR3_X1 U19840 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n16704), .A3(n16605), 
        .ZN(n16606) );
  AOI211_X1 U19841 ( .C1(n16713), .C2(n16607), .A(n18061), .B(n16606), .ZN(
        n16613) );
  INV_X1 U19842 ( .A(n16608), .ZN(n16627) );
  AOI21_X1 U19843 ( .B1(n16627), .B2(n16723), .A(n16720), .ZN(n16614) );
  INV_X1 U19844 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18623) );
  NAND2_X1 U19845 ( .A1(n16723), .A2(n18623), .ZN(n16626) );
  AOI21_X1 U19846 ( .B1(n16614), .B2(n16626), .A(n18624), .ZN(n16611) );
  AOI211_X1 U19847 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16620), .A(n16609), .B(
        n16706), .ZN(n16610) );
  AOI211_X1 U19848 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16721), .A(n16611), .B(
        n16610), .ZN(n16612) );
  OAI211_X1 U19849 ( .C1(n20951), .C2(n16693), .A(n16613), .B(n16612), .ZN(
        P3_U2661) );
  INV_X1 U19850 ( .A(n16614), .ZN(n16635) );
  OAI21_X1 U19851 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16629), .A(
        n16615), .ZN(n17622) );
  NOR2_X1 U19852 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18588), .ZN(
        n16616) );
  AOI22_X1 U19853 ( .A1(n16724), .A2(n17622), .B1(n16629), .B2(n16616), .ZN(
        n16617) );
  OAI22_X1 U19854 ( .A1(n16618), .A2(n16617), .B1(n17622), .B2(n16644), .ZN(
        n16619) );
  AOI211_X1 U19855 ( .C1(n16721), .C2(P3_EBX_REG_9__SCAN_IN), .A(n18061), .B(
        n16619), .ZN(n16622) );
  OAI211_X1 U19856 ( .C1(n16628), .C2(n20822), .A(n16731), .B(n16620), .ZN(
        n16621) );
  OAI211_X1 U19857 ( .C1(n16693), .C2(n16623), .A(n16622), .B(n16621), .ZN(
        n16624) );
  AOI21_X1 U19858 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n16635), .A(n16624), .ZN(
        n16625) );
  OAI21_X1 U19859 ( .B1(n16627), .B2(n16626), .A(n16625), .ZN(P3_U2662) );
  INV_X1 U19860 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17604) );
  AOI211_X1 U19861 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16642), .A(n16628), .B(
        n16706), .ZN(n16634) );
  INV_X1 U19862 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17649) );
  NOR2_X1 U19863 ( .A1(n17649), .A2(n16651), .ZN(n16643) );
  AOI21_X1 U19864 ( .B1(n16643), .B2(n16689), .A(n16688), .ZN(n16646) );
  INV_X1 U19865 ( .A(n16629), .ZN(n16630) );
  OAI21_X1 U19866 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16643), .A(
        n16630), .ZN(n17633) );
  XOR2_X1 U19867 ( .A(n16646), .B(n17633), .Z(n16631) );
  OAI22_X1 U19868 ( .A1(n16692), .A2(n16632), .B1(n18588), .B2(n16631), .ZN(
        n16633) );
  NOR3_X1 U19869 ( .A1(n18061), .A2(n16634), .A3(n16633), .ZN(n16637) );
  NAND3_X1 U19870 ( .A1(n16723), .A2(P3_REIP_REG_5__SCAN_IN), .A3(n16661), 
        .ZN(n16660) );
  NOR2_X1 U19871 ( .A1(n18617), .A2(n16660), .ZN(n16641) );
  OAI221_X1 U19872 ( .B1(P3_REIP_REG_8__SCAN_IN), .B2(P3_REIP_REG_7__SCAN_IN), 
        .C1(P3_REIP_REG_8__SCAN_IN), .C2(n16641), .A(n16635), .ZN(n16636) );
  OAI211_X1 U19873 ( .C1(n16693), .C2(n17604), .A(n16637), .B(n16636), .ZN(
        P3_U2663) );
  AOI21_X1 U19874 ( .B1(n16723), .B2(n16638), .A(n16720), .ZN(n16663) );
  OAI21_X1 U19875 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16660), .A(n16663), .ZN(
        n16640) );
  OAI22_X1 U19876 ( .A1(n17649), .A2(n16693), .B1(n16692), .B2(n17064), .ZN(
        n16639) );
  AOI221_X1 U19877 ( .B1(n16641), .B2(n18619), .C1(n16640), .C2(
        P3_REIP_REG_7__SCAN_IN), .A(n16639), .ZN(n16649) );
  OAI211_X1 U19878 ( .C1(n16650), .C2(n17064), .A(n16731), .B(n16642), .ZN(
        n16648) );
  AOI21_X1 U19879 ( .B1(n17649), .B2(n16651), .A(n16643), .ZN(n17654) );
  INV_X1 U19880 ( .A(n16644), .ZN(n16702) );
  AOI21_X1 U19881 ( .B1(n17654), .B2(n16652), .A(n18588), .ZN(n16645) );
  OAI22_X1 U19882 ( .A1(n17654), .A2(n16646), .B1(n16702), .B2(n16645), .ZN(
        n16647) );
  NAND4_X1 U19883 ( .A1(n16649), .A2(n17892), .A3(n16648), .A4(n16647), .ZN(
        P3_U2664) );
  AOI211_X1 U19884 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16665), .A(n16650), .B(
        n16706), .ZN(n16658) );
  INV_X1 U19885 ( .A(n17671), .ZN(n16687) );
  NOR3_X1 U19886 ( .A1(n17727), .A2(n16687), .A3(n17695), .ZN(n16672) );
  OAI221_X1 U19887 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n16672), .A(n16651), .ZN(n17663) );
  NAND3_X1 U19888 ( .A1(n17663), .A2(n16724), .A3(n16652), .ZN(n16656) );
  AOI211_X1 U19889 ( .C1(n9710), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16653), .B(n17663), .ZN(n16654) );
  AOI211_X1 U19890 ( .C1(n16721), .C2(P3_EBX_REG_6__SCAN_IN), .A(n18061), .B(
        n16654), .ZN(n16655) );
  NAND2_X1 U19891 ( .A1(n16656), .A2(n16655), .ZN(n16657) );
  AOI211_X1 U19892 ( .C1(n16725), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16658), .B(n16657), .ZN(n16659) );
  OAI221_X1 U19893 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16660), .C1(n18617), 
        .C2(n16663), .A(n16659), .ZN(P3_U2665) );
  AOI21_X1 U19894 ( .B1(n16723), .B2(n16661), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n16662) );
  OAI22_X1 U19895 ( .A1(n16663), .A2(n16662), .B1(n16692), .B2(n17067), .ZN(
        n16664) );
  AOI21_X1 U19896 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16725), .A(
        n16664), .ZN(n16670) );
  OAI211_X1 U19897 ( .C1(n16671), .C2(n17067), .A(n16731), .B(n16665), .ZN(
        n16669) );
  XOR2_X1 U19898 ( .A(n17672), .B(n16672), .Z(n17677) );
  INV_X1 U19899 ( .A(n17677), .ZN(n16667) );
  AOI21_X1 U19900 ( .B1(n16689), .B2(n16672), .A(n16688), .ZN(n16666) );
  INV_X1 U19901 ( .A(n16666), .ZN(n16675) );
  OAI221_X1 U19902 ( .B1(n16667), .B2(n16666), .C1(n17677), .C2(n16675), .A(
        n16713), .ZN(n16668) );
  NAND4_X1 U19903 ( .A1(n16670), .A2(n17892), .A3(n16669), .A4(n16668), .ZN(
        P3_U2666) );
  AOI211_X1 U19904 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16696), .A(n16671), .B(
        n16706), .ZN(n16682) );
  AOI21_X1 U19905 ( .B1(n16723), .B2(n16683), .A(n16720), .ZN(n16699) );
  NAND2_X1 U19906 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17671), .ZN(
        n16673) );
  AOI21_X1 U19907 ( .B1(n17695), .B2(n16673), .A(n16672), .ZN(n17692) );
  NAND2_X1 U19908 ( .A1(n17671), .A2(n17695), .ZN(n17686) );
  OAI22_X1 U19909 ( .A1(n17692), .A2(n16675), .B1(n16674), .B2(n17686), .ZN(
        n16676) );
  AOI22_X1 U19910 ( .A1(n16713), .A2(n16676), .B1(n17692), .B2(n16702), .ZN(
        n16680) );
  NOR2_X1 U19911 ( .A1(n16678), .A2(n16677), .ZN(n18747) );
  AOI221_X1 U19912 ( .B1(n17046), .B2(n18747), .C1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18747), .A(n18061), .ZN(
        n16679) );
  OAI211_X1 U19913 ( .C1(n18613), .C2(n16699), .A(n16680), .B(n16679), .ZN(
        n16681) );
  AOI211_X1 U19914 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16721), .A(n16682), .B(
        n16681), .ZN(n16685) );
  OR3_X1 U19915 ( .A1(n16704), .A2(n16683), .A3(P3_REIP_REG_4__SCAN_IN), .ZN(
        n16684) );
  OAI211_X1 U19916 ( .C1(n16693), .C2(n17695), .A(n16685), .B(n16684), .ZN(
        P3_U2667) );
  INV_X1 U19917 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18609) );
  NOR2_X1 U19918 ( .A1(n18711), .A2(n18609), .ZN(n16705) );
  AOI21_X1 U19919 ( .B1(n16723), .B2(n16705), .A(P3_REIP_REG_3__SCAN_IN), .ZN(
        n16700) );
  NOR2_X1 U19920 ( .A1(n18709), .A2(n18535), .ZN(n18532) );
  OAI21_X1 U19921 ( .B1(n18532), .B2(n18686), .A(n12553), .ZN(n18683) );
  NOR2_X1 U19922 ( .A1(n17727), .A2(n17718), .ZN(n16701) );
  OAI22_X1 U19923 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16701), .B1(
        n17727), .B2(n16687), .ZN(n17702) );
  AOI21_X1 U19924 ( .B1(n16689), .B2(n16701), .A(n16688), .ZN(n16712) );
  INV_X1 U19925 ( .A(n16712), .ZN(n16691) );
  OAI21_X1 U19926 ( .B1(n17702), .B2(n16691), .A(n16713), .ZN(n16690) );
  AOI21_X1 U19927 ( .B1(n17702), .B2(n16691), .A(n16690), .ZN(n16695) );
  OAI22_X1 U19928 ( .A1(n17704), .A2(n16693), .B1(n16692), .B2(n17075), .ZN(
        n16694) );
  AOI211_X1 U19929 ( .C1(n18747), .C2(n18683), .A(n16695), .B(n16694), .ZN(
        n16698) );
  OAI211_X1 U19930 ( .C1(n16707), .C2(n17075), .A(n16731), .B(n16696), .ZN(
        n16697) );
  OAI211_X1 U19931 ( .C1(n16700), .C2(n16699), .A(n16698), .B(n16697), .ZN(
        P3_U2668) );
  AOI22_X1 U19932 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n16725), .B1(
        n16721), .B2(P3_EBX_REG_2__SCAN_IN), .ZN(n16718) );
  NOR2_X1 U19933 ( .A1(n18709), .A2(n18703), .ZN(n18542) );
  OR2_X1 U19934 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18542), .ZN(
        n18531) );
  OAI21_X1 U19935 ( .B1(n18535), .B2(n18709), .A(n18531), .ZN(n18690) );
  INV_X1 U19936 ( .A(n18690), .ZN(n16703) );
  AOI21_X1 U19937 ( .B1(n17727), .B2(n17718), .A(n16701), .ZN(n16711) );
  AOI22_X1 U19938 ( .A1(n16703), .A2(n18747), .B1(n16711), .B2(n16702), .ZN(
        n16717) );
  AOI211_X1 U19939 ( .C1(n18711), .C2(n18609), .A(n16705), .B(n16704), .ZN(
        n16710) );
  NOR2_X1 U19940 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16722) );
  INV_X1 U19941 ( .A(n16722), .ZN(n16708) );
  AOI211_X1 U19942 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16708), .A(n16707), .B(
        n16706), .ZN(n16709) );
  AOI211_X1 U19943 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(n16720), .A(n16710), .B(
        n16709), .ZN(n16716) );
  INV_X1 U19944 ( .A(n16711), .ZN(n17714) );
  OAI211_X1 U19945 ( .C1(n16714), .C2(n17714), .A(n16713), .B(n16712), .ZN(
        n16715) );
  NAND4_X1 U19946 ( .A1(n16718), .A2(n16717), .A3(n16716), .A4(n16715), .ZN(
        P3_U2669) );
  OAI22_X1 U19947 ( .A1(n18709), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n18703), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18700) );
  AOI22_X1 U19948 ( .A1(n18747), .A2(n18700), .B1(n17727), .B2(n16719), .ZN(
        n16729) );
  AOI22_X1 U19949 ( .A1(n16721), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n16720), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n16728) );
  NOR2_X1 U19950 ( .A1(n16722), .A2(n17082), .ZN(n17086) );
  AOI22_X1 U19951 ( .A1(n16731), .A2(n17086), .B1(n16723), .B2(n18711), .ZN(
        n16727) );
  OAI221_X1 U19952 ( .B1(n16725), .B2(n16724), .C1(n16725), .C2(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16726) );
  NAND4_X1 U19953 ( .A1(n16729), .A2(n16728), .A3(n16727), .A4(n16726), .ZN(
        P3_U2670) );
  AOI22_X1 U19954 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16730), .B1(n18747), 
        .B2(n18709), .ZN(n16736) );
  OAI21_X1 U19955 ( .B1(n16732), .B2(n16731), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n16735) );
  INV_X1 U19956 ( .A(n18706), .ZN(n18692) );
  NAND3_X1 U19957 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18692), .A3(
        n16733), .ZN(n16734) );
  NAND3_X1 U19958 ( .A1(n16736), .A2(n16735), .A3(n16734), .ZN(P3_U2671) );
  NAND2_X1 U19959 ( .A1(n16738), .A2(n16737), .ZN(n16739) );
  NAND2_X1 U19960 ( .A1(n16739), .A2(n17079), .ZN(n16835) );
  AOI22_X1 U19961 ( .A1(n17033), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17044), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16744) );
  AOI22_X1 U19962 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16743) );
  AOI22_X1 U19963 ( .A1(n16755), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16742) );
  AOI22_X1 U19964 ( .A1(n9740), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16741) );
  NAND4_X1 U19965 ( .A1(n16744), .A2(n16743), .A3(n16742), .A4(n16741), .ZN(
        n16750) );
  AOI22_X1 U19966 ( .A1(n9715), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16748) );
  AOI22_X1 U19967 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16747) );
  AOI22_X1 U19968 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9711), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16746) );
  AOI22_X1 U19969 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16745) );
  NAND4_X1 U19970 ( .A1(n16748), .A2(n16747), .A3(n16746), .A4(n16745), .ZN(
        n16749) );
  NOR2_X1 U19971 ( .A1(n16750), .A2(n16749), .ZN(n16843) );
  AOI22_X1 U19972 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9716), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16754) );
  AOI22_X1 U19973 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12570), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16753) );
  AOI22_X1 U19974 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16752) );
  AOI22_X1 U19975 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16751) );
  NAND4_X1 U19976 ( .A1(n16754), .A2(n16753), .A3(n16752), .A4(n16751), .ZN(
        n16761) );
  AOI22_X1 U19977 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16759) );
  AOI22_X1 U19978 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17044), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16758) );
  AOI22_X1 U19979 ( .A1(n16740), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9711), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16757) );
  AOI22_X1 U19980 ( .A1(n16755), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16756) );
  NAND4_X1 U19981 ( .A1(n16759), .A2(n16758), .A3(n16757), .A4(n16756), .ZN(
        n16760) );
  NOR2_X1 U19982 ( .A1(n16761), .A2(n16760), .ZN(n16852) );
  AOI22_X1 U19983 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16765) );
  AOI22_X1 U19984 ( .A1(n17033), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16764) );
  AOI22_X1 U19985 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16763) );
  AOI22_X1 U19986 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9711), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16762) );
  NAND4_X1 U19987 ( .A1(n16765), .A2(n16764), .A3(n16763), .A4(n16762), .ZN(
        n16771) );
  AOI22_X1 U19988 ( .A1(n9716), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n16769) );
  AOI22_X1 U19989 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n16768) );
  AOI22_X1 U19990 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9740), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16767) );
  AOI22_X1 U19991 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16766) );
  NAND4_X1 U19992 ( .A1(n16769), .A2(n16768), .A3(n16767), .A4(n16766), .ZN(
        n16770) );
  NOR2_X1 U19993 ( .A1(n16771), .A2(n16770), .ZN(n16860) );
  AOI22_X1 U19994 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16781) );
  AOI22_X1 U19995 ( .A1(n12570), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16780) );
  AOI22_X1 U19996 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17033), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16772) );
  OAI21_X1 U19997 ( .B1(n9786), .B2(n18087), .A(n16772), .ZN(n16778) );
  AOI22_X1 U19998 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16776) );
  AOI22_X1 U19999 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9711), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16775) );
  AOI22_X1 U20000 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16774) );
  AOI22_X1 U20001 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16773) );
  NAND4_X1 U20002 ( .A1(n16776), .A2(n16775), .A3(n16774), .A4(n16773), .ZN(
        n16777) );
  AOI211_X1 U20003 ( .C1(n9716), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n16778), .B(n16777), .ZN(n16779) );
  NAND3_X1 U20004 ( .A1(n16781), .A2(n16780), .A3(n16779), .ZN(n16865) );
  AOI22_X1 U20005 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17017), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16791) );
  AOI22_X1 U20006 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n16740), .ZN(n16790) );
  INV_X1 U20007 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n20908) );
  AOI22_X1 U20008 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n12571), .ZN(n16782) );
  OAI21_X1 U20009 ( .B1(n20908), .B2(n9719), .A(n16782), .ZN(n16788) );
  AOI22_X1 U20010 ( .A1(n9715), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17044), .ZN(n16786) );
  AOI22_X1 U20011 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16785) );
  AOI22_X1 U20012 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n17033), .ZN(n16784) );
  AOI22_X1 U20013 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17048), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16783) );
  NAND4_X1 U20014 ( .A1(n16786), .A2(n16785), .A3(n16784), .A4(n16783), .ZN(
        n16787) );
  AOI211_X1 U20015 ( .C1(n17043), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n16788), .B(n16787), .ZN(n16789) );
  NAND3_X1 U20016 ( .A1(n16791), .A2(n16790), .A3(n16789), .ZN(n16866) );
  NAND2_X1 U20017 ( .A1(n16865), .A2(n16866), .ZN(n16864) );
  NOR2_X1 U20018 ( .A1(n16860), .A2(n16864), .ZN(n16857) );
  AOI22_X1 U20019 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16801) );
  AOI22_X1 U20020 ( .A1(n9740), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16800) );
  INV_X1 U20021 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n20924) );
  AOI22_X1 U20022 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16792) );
  OAI21_X1 U20023 ( .B1(n12519), .B2(n20924), .A(n16792), .ZN(n16798) );
  AOI22_X1 U20024 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16796) );
  AOI22_X1 U20025 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16795) );
  AOI22_X1 U20026 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16794) );
  AOI22_X1 U20027 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16793) );
  NAND4_X1 U20028 ( .A1(n16796), .A2(n16795), .A3(n16794), .A4(n16793), .ZN(
        n16797) );
  AOI211_X1 U20029 ( .C1(n9714), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n16798), .B(n16797), .ZN(n16799) );
  NAND3_X1 U20030 ( .A1(n16801), .A2(n16800), .A3(n16799), .ZN(n16856) );
  NAND2_X1 U20031 ( .A1(n16857), .A2(n16856), .ZN(n16855) );
  NOR2_X1 U20032 ( .A1(n16852), .A2(n16855), .ZN(n16848) );
  AOI22_X1 U20033 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16812) );
  AOI22_X1 U20034 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9709), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16811) );
  AOI22_X1 U20035 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17044), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16803) );
  OAI21_X1 U20036 ( .B1(n9786), .B2(n18107), .A(n16803), .ZN(n16809) );
  AOI22_X1 U20037 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16807) );
  AOI22_X1 U20038 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16806) );
  AOI22_X1 U20039 ( .A1(n9740), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16805) );
  AOI22_X1 U20040 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16804) );
  NAND4_X1 U20041 ( .A1(n16807), .A2(n16806), .A3(n16805), .A4(n16804), .ZN(
        n16808) );
  AOI211_X1 U20042 ( .C1(n17027), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n16809), .B(n16808), .ZN(n16810) );
  NAND3_X1 U20043 ( .A1(n16812), .A2(n16811), .A3(n16810), .ZN(n16847) );
  NAND2_X1 U20044 ( .A1(n16848), .A2(n16847), .ZN(n16846) );
  NOR2_X1 U20045 ( .A1(n16843), .A2(n16846), .ZN(n16842) );
  INV_X1 U20046 ( .A(n16842), .ZN(n16839) );
  AOI22_X1 U20047 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16816) );
  AOI22_X1 U20048 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16815) );
  AOI22_X1 U20049 ( .A1(n17033), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16814) );
  AOI22_X1 U20050 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16813) );
  NAND4_X1 U20051 ( .A1(n16816), .A2(n16815), .A3(n16814), .A4(n16813), .ZN(
        n16822) );
  AOI22_X1 U20052 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16820) );
  AOI22_X1 U20053 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17044), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16819) );
  AOI22_X1 U20054 ( .A1(n9716), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16818) );
  AOI22_X1 U20055 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16817) );
  NAND4_X1 U20056 ( .A1(n16820), .A2(n16819), .A3(n16818), .A4(n16817), .ZN(
        n16821) );
  NOR2_X1 U20057 ( .A1(n16822), .A2(n16821), .ZN(n16838) );
  NOR2_X1 U20058 ( .A1(n16839), .A2(n16838), .ZN(n16834) );
  AOI22_X1 U20059 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17044), .ZN(n16826) );
  AOI22_X1 U20060 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16825) );
  AOI22_X1 U20061 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n17043), .ZN(n16824) );
  AOI22_X1 U20062 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n16740), .ZN(n16823) );
  NAND4_X1 U20063 ( .A1(n16826), .A2(n16825), .A3(n16824), .A4(n16823), .ZN(
        n16832) );
  AOI22_X1 U20064 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17045), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16830) );
  AOI22_X1 U20065 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17048), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16829) );
  AOI22_X1 U20066 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17049), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16828) );
  AOI22_X1 U20067 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17046), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n12571), .ZN(n16827) );
  NAND4_X1 U20068 ( .A1(n16830), .A2(n16829), .A3(n16828), .A4(n16827), .ZN(
        n16831) );
  NOR2_X1 U20069 ( .A1(n16832), .A2(n16831), .ZN(n16833) );
  XOR2_X1 U20070 ( .A(n16834), .B(n16833), .Z(n17106) );
  OAI22_X1 U20071 ( .A1(n16836), .A2(n16835), .B1(n17106), .B2(n17079), .ZN(
        P3_U2673) );
  INV_X1 U20072 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n20981) );
  NAND2_X1 U20073 ( .A1(n17097), .A2(n16896), .ZN(n16882) );
  NAND3_X1 U20074 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n16854), .ZN(n16841) );
  XNOR2_X1 U20075 ( .A(n16839), .B(n16838), .ZN(n17110) );
  NAND3_X1 U20076 ( .A1(n16841), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n17079), 
        .ZN(n16840) );
  OAI221_X1 U20077 ( .B1(n16841), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n17079), 
        .C2(n17110), .A(n16840), .ZN(P3_U2674) );
  NAND2_X1 U20078 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16854), .ZN(n16849) );
  AND2_X1 U20079 ( .A1(n17079), .A2(n16841), .ZN(n16844) );
  AOI21_X1 U20080 ( .B1(n16843), .B2(n16846), .A(n16842), .ZN(n17111) );
  AOI22_X1 U20081 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16844), .B1(n17089), 
        .B2(n17111), .ZN(n16845) );
  OAI21_X1 U20082 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n16849), .A(n16845), .ZN(
        P3_U2675) );
  OAI21_X1 U20083 ( .B1(n16848), .B2(n16847), .A(n16846), .ZN(n17119) );
  OAI211_X1 U20084 ( .C1(n16854), .C2(P3_EBX_REG_27__SCAN_IN), .A(n17079), .B(
        n16849), .ZN(n16850) );
  OAI21_X1 U20085 ( .B1(n17119), .B2(n17079), .A(n16850), .ZN(P3_U2676) );
  INV_X1 U20086 ( .A(n16851), .ZN(n16859) );
  AOI21_X1 U20087 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17079), .A(n16859), .ZN(
        n16853) );
  XNOR2_X1 U20088 ( .A(n16852), .B(n16855), .ZN(n17124) );
  OAI22_X1 U20089 ( .A1(n16854), .A2(n16853), .B1(n17079), .B2(n17124), .ZN(
        P3_U2677) );
  AOI21_X1 U20090 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17079), .A(n16862), .ZN(
        n16858) );
  OAI21_X1 U20091 ( .B1(n16857), .B2(n16856), .A(n16855), .ZN(n17129) );
  OAI22_X1 U20092 ( .A1(n16859), .A2(n16858), .B1(n17079), .B2(n17129), .ZN(
        P3_U2678) );
  AOI21_X1 U20093 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17079), .A(n16868), .ZN(
        n16861) );
  XNOR2_X1 U20094 ( .A(n16860), .B(n16864), .ZN(n17134) );
  OAI22_X1 U20095 ( .A1(n16862), .A2(n16861), .B1(n17079), .B2(n17134), .ZN(
        P3_U2679) );
  AOI21_X1 U20096 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17079), .A(n16863), .ZN(
        n16867) );
  OAI21_X1 U20097 ( .B1(n16866), .B2(n16865), .A(n16864), .ZN(n17139) );
  OAI22_X1 U20098 ( .A1(n16868), .A2(n16867), .B1(n17079), .B2(n17139), .ZN(
        P3_U2680) );
  AOI22_X1 U20099 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16879) );
  AOI22_X1 U20100 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16878) );
  AOI22_X1 U20101 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16869) );
  OAI21_X1 U20102 ( .B1(n16870), .B2(n20853), .A(n16869), .ZN(n16876) );
  AOI22_X1 U20103 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16874) );
  AOI22_X1 U20104 ( .A1(n9740), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17033), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16873) );
  AOI22_X1 U20105 ( .A1(n16740), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16872) );
  AOI22_X1 U20106 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17044), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16871) );
  NAND4_X1 U20107 ( .A1(n16874), .A2(n16873), .A3(n16872), .A4(n16871), .ZN(
        n16875) );
  AOI211_X1 U20108 ( .C1(n17050), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n16876), .B(n16875), .ZN(n16877) );
  NAND3_X1 U20109 ( .A1(n16879), .A2(n16878), .A3(n16877), .ZN(n17140) );
  INV_X1 U20110 ( .A(n17140), .ZN(n16881) );
  NAND3_X1 U20111 ( .A1(n16882), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17079), 
        .ZN(n16880) );
  OAI221_X1 U20112 ( .B1(n16882), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17079), 
        .C2(n16881), .A(n16880), .ZN(P3_U2681) );
  AOI21_X1 U20113 ( .B1(n16883), .B2(n16907), .A(n17089), .ZN(n16884) );
  INV_X1 U20114 ( .A(n16884), .ZN(n16895) );
  AOI22_X1 U20115 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16888) );
  AOI22_X1 U20116 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16887) );
  AOI22_X1 U20117 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16886) );
  AOI22_X1 U20118 ( .A1(n17048), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16885) );
  NAND4_X1 U20119 ( .A1(n16888), .A2(n16887), .A3(n16886), .A4(n16885), .ZN(
        n16894) );
  AOI22_X1 U20120 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16892) );
  AOI22_X1 U20121 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16891) );
  AOI22_X1 U20122 ( .A1(n9716), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16890) );
  AOI22_X1 U20123 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17044), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16889) );
  NAND4_X1 U20124 ( .A1(n16892), .A2(n16891), .A3(n16890), .A4(n16889), .ZN(
        n16893) );
  NOR2_X1 U20125 ( .A1(n16894), .A2(n16893), .ZN(n17146) );
  OAI22_X1 U20126 ( .A1(n16896), .A2(n16895), .B1(n17146), .B2(n17079), .ZN(
        P3_U2682) );
  AOI22_X1 U20127 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16900) );
  AOI22_X1 U20128 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17033), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16899) );
  AOI22_X1 U20129 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16898) );
  AOI22_X1 U20130 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16897) );
  NAND4_X1 U20131 ( .A1(n16900), .A2(n16899), .A3(n16898), .A4(n16897), .ZN(
        n16906) );
  AOI22_X1 U20132 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9714), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16904) );
  AOI22_X1 U20133 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16903) );
  AOI22_X1 U20134 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16902) );
  AOI22_X1 U20135 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9709), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16901) );
  NAND4_X1 U20136 ( .A1(n16904), .A2(n16903), .A3(n16902), .A4(n16901), .ZN(
        n16905) );
  NOR2_X1 U20137 ( .A1(n16906), .A2(n16905), .ZN(n17153) );
  OAI21_X1 U20138 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16921), .A(n16907), .ZN(
        n16908) );
  AOI22_X1 U20139 ( .A1(n17089), .A2(n17153), .B1(n16908), .B2(n17079), .ZN(
        P3_U2683) );
  INV_X1 U20140 ( .A(n16909), .ZN(n16933) );
  OAI21_X1 U20141 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n16933), .A(n17079), .ZN(
        n16920) );
  AOI22_X1 U20142 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16913) );
  AOI22_X1 U20143 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16912) );
  AOI22_X1 U20144 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17044), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16911) );
  AOI22_X1 U20145 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16910) );
  NAND4_X1 U20146 ( .A1(n16913), .A2(n16912), .A3(n16911), .A4(n16910), .ZN(
        n16919) );
  AOI22_X1 U20147 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9709), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16917) );
  AOI22_X1 U20148 ( .A1(n17033), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16916) );
  AOI22_X1 U20149 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16755), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16915) );
  AOI22_X1 U20150 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16914) );
  NAND4_X1 U20151 ( .A1(n16917), .A2(n16916), .A3(n16915), .A4(n16914), .ZN(
        n16918) );
  NOR2_X1 U20152 ( .A1(n16919), .A2(n16918), .ZN(n17158) );
  OAI22_X1 U20153 ( .A1(n16921), .A2(n16920), .B1(n17158), .B2(n17079), .ZN(
        P3_U2684) );
  AOI22_X1 U20154 ( .A1(n17097), .A2(n16945), .B1(P3_EBX_REG_18__SCAN_IN), 
        .B2(n17079), .ZN(n16932) );
  AOI22_X1 U20155 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16925) );
  AOI22_X1 U20156 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16924) );
  AOI22_X1 U20157 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16923) );
  AOI22_X1 U20158 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9709), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16922) );
  NAND4_X1 U20159 ( .A1(n16925), .A2(n16924), .A3(n16923), .A4(n16922), .ZN(
        n16931) );
  AOI22_X1 U20160 ( .A1(n9714), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12535), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16929) );
  AOI22_X1 U20161 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16928) );
  AOI22_X1 U20162 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16927) );
  AOI22_X1 U20163 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16926) );
  NAND4_X1 U20164 ( .A1(n16929), .A2(n16928), .A3(n16927), .A4(n16926), .ZN(
        n16930) );
  NOR2_X1 U20165 ( .A1(n16931), .A2(n16930), .ZN(n17162) );
  OAI22_X1 U20166 ( .A1(n16933), .A2(n16932), .B1(n17162), .B2(n17079), .ZN(
        P3_U2685) );
  AOI22_X1 U20167 ( .A1(n17033), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17044), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16937) );
  AOI22_X1 U20168 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17051), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16936) );
  AOI22_X1 U20169 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9709), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16935) );
  AOI22_X1 U20170 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16934) );
  NAND4_X1 U20171 ( .A1(n16937), .A2(n16936), .A3(n16935), .A4(n16934), .ZN(
        n16943) );
  AOI22_X1 U20172 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16941) );
  AOI22_X1 U20173 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16940) );
  AOI22_X1 U20174 ( .A1(n9715), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16939) );
  AOI22_X1 U20175 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16938) );
  NAND4_X1 U20176 ( .A1(n16941), .A2(n16940), .A3(n16939), .A4(n16938), .ZN(
        n16942) );
  NOR2_X1 U20177 ( .A1(n16943), .A2(n16942), .ZN(n17168) );
  INV_X1 U20178 ( .A(n16944), .ZN(n16960) );
  INV_X1 U20179 ( .A(n16945), .ZN(n16946) );
  OAI21_X1 U20180 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n16960), .A(n16946), .ZN(
        n16947) );
  AOI22_X1 U20181 ( .A1(n17089), .A2(n17168), .B1(n16947), .B2(n17079), .ZN(
        P3_U2686) );
  AOI21_X1 U20182 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17079), .A(n16948), .ZN(
        n16959) );
  AOI22_X1 U20183 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16952) );
  AOI22_X1 U20184 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16951) );
  AOI22_X1 U20185 ( .A1(n12535), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16950) );
  AOI22_X1 U20186 ( .A1(n9716), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16949) );
  NAND4_X1 U20187 ( .A1(n16952), .A2(n16951), .A3(n16950), .A4(n16949), .ZN(
        n16958) );
  AOI22_X1 U20188 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16956) );
  AOI22_X1 U20189 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9717), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16955) );
  AOI22_X1 U20190 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16954) );
  AOI22_X1 U20191 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16953) );
  NAND4_X1 U20192 ( .A1(n16956), .A2(n16955), .A3(n16954), .A4(n16953), .ZN(
        n16957) );
  NOR2_X1 U20193 ( .A1(n16958), .A2(n16957), .ZN(n17175) );
  OAI22_X1 U20194 ( .A1(n16960), .A2(n16959), .B1(n17175), .B2(n17079), .ZN(
        P3_U2687) );
  NOR2_X1 U20195 ( .A1(n18119), .A2(n17085), .ZN(n17088) );
  INV_X1 U20196 ( .A(n17088), .ZN(n17073) );
  OAI22_X1 U20197 ( .A1(n17089), .A2(n16985), .B1(P3_EBX_REG_13__SCAN_IN), 
        .B2(n17073), .ZN(n16984) );
  AOI22_X1 U20198 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9716), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16970) );
  AOI22_X1 U20199 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16969) );
  INV_X1 U20200 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n20883) );
  AOI22_X1 U20201 ( .A1(n17048), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16961) );
  OAI21_X1 U20202 ( .B1(n9719), .B2(n20883), .A(n16961), .ZN(n16967) );
  AOI22_X1 U20203 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9717), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16965) );
  AOI22_X1 U20204 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16964) );
  AOI22_X1 U20205 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16963) );
  AOI22_X1 U20206 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16962) );
  NAND4_X1 U20207 ( .A1(n16965), .A2(n16964), .A3(n16963), .A4(n16962), .ZN(
        n16966) );
  AOI211_X1 U20208 ( .C1(n17027), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n16967), .B(n16966), .ZN(n16968) );
  NAND3_X1 U20209 ( .A1(n16970), .A2(n16969), .A3(n16968), .ZN(n17184) );
  AOI22_X1 U20210 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16984), .B1(n17089), 
        .B2(n17184), .ZN(n16973) );
  NAND4_X1 U20211 ( .A1(n17097), .A2(P3_EBX_REG_13__SCAN_IN), .A3(n16985), 
        .A4(n16971), .ZN(n16972) );
  NAND2_X1 U20212 ( .A1(n16973), .A2(n16972), .ZN(P3_U2689) );
  AOI22_X1 U20213 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16977) );
  AOI22_X1 U20214 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16976) );
  AOI22_X1 U20215 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16975) );
  AOI22_X1 U20216 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16974) );
  NAND4_X1 U20217 ( .A1(n16977), .A2(n16976), .A3(n16975), .A4(n16974), .ZN(
        n16983) );
  AOI22_X1 U20218 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9715), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16981) );
  AOI22_X1 U20219 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16980) );
  AOI22_X1 U20220 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16979) );
  AOI22_X1 U20221 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16978) );
  NAND4_X1 U20222 ( .A1(n16981), .A2(n16980), .A3(n16979), .A4(n16978), .ZN(
        n16982) );
  NOR2_X1 U20223 ( .A1(n16983), .A2(n16982), .ZN(n17188) );
  OAI21_X1 U20224 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n16985), .A(n16984), .ZN(
        n16986) );
  OAI21_X1 U20225 ( .B1(n17188), .B2(n17079), .A(n16986), .ZN(P3_U2690) );
  AOI22_X1 U20226 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16990) );
  AOI22_X1 U20227 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16989) );
  AOI22_X1 U20228 ( .A1(n9716), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17044), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16988) );
  AOI22_X1 U20229 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16987) );
  NAND4_X1 U20230 ( .A1(n16990), .A2(n16989), .A3(n16988), .A4(n16987), .ZN(
        n16996) );
  AOI22_X1 U20231 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16994) );
  AOI22_X1 U20232 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16993) );
  AOI22_X1 U20233 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17033), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16992) );
  AOI22_X1 U20234 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16991) );
  NAND4_X1 U20235 ( .A1(n16994), .A2(n16993), .A3(n16992), .A4(n16991), .ZN(
        n16995) );
  NOR2_X1 U20236 ( .A1(n16996), .A2(n16995), .ZN(n17192) );
  OAI211_X1 U20237 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16998), .A(n16997), .B(
        n17079), .ZN(n16999) );
  OAI21_X1 U20238 ( .B1(n17192), .B2(n17079), .A(n16999), .ZN(P3_U2691) );
  AOI22_X1 U20239 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20240 ( .A1(n9709), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17002) );
  AOI22_X1 U20241 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9718), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17001) );
  AOI22_X1 U20242 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17000) );
  NAND4_X1 U20243 ( .A1(n17003), .A2(n17002), .A3(n17001), .A4(n17000), .ZN(
        n17009) );
  AOI22_X1 U20244 ( .A1(n9716), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17017), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17007) );
  AOI22_X1 U20245 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17044), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17006) );
  AOI22_X1 U20246 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17005) );
  AOI22_X1 U20247 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17004) );
  NAND4_X1 U20248 ( .A1(n17007), .A2(n17006), .A3(n17005), .A4(n17004), .ZN(
        n17008) );
  NOR2_X1 U20249 ( .A1(n17009), .A2(n17008), .ZN(n17195) );
  OAI21_X1 U20250 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17025), .A(n17010), .ZN(
        n17011) );
  AOI22_X1 U20251 ( .A1(n17089), .A2(n17195), .B1(n17011), .B2(n17079), .ZN(
        P3_U2692) );
  OAI21_X1 U20252 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17012), .A(n17079), .ZN(
        n17024) );
  AOI22_X1 U20253 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17016) );
  AOI22_X1 U20254 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17015) );
  AOI22_X1 U20255 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17014) );
  AOI22_X1 U20256 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12544), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17013) );
  NAND4_X1 U20257 ( .A1(n17016), .A2(n17015), .A3(n17014), .A4(n17013), .ZN(
        n17023) );
  AOI22_X1 U20258 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17044), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17021) );
  AOI22_X1 U20259 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17020) );
  AOI22_X1 U20260 ( .A1(n17026), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17019) );
  AOI22_X1 U20261 ( .A1(n9716), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17017), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17018) );
  NAND4_X1 U20262 ( .A1(n17021), .A2(n17020), .A3(n17019), .A4(n17018), .ZN(
        n17022) );
  NOR2_X1 U20263 ( .A1(n17023), .A2(n17022), .ZN(n17202) );
  OAI22_X1 U20264 ( .A1(n17025), .A2(n17024), .B1(n17202), .B2(n17079), .ZN(
        P3_U2693) );
  AOI22_X1 U20265 ( .A1(n17026), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17031) );
  AOI22_X1 U20266 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17030) );
  AOI22_X1 U20267 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12571), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20268 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17028) );
  NAND4_X1 U20269 ( .A1(n17031), .A2(n17030), .A3(n17029), .A4(n17028), .ZN(
        n17039) );
  AOI22_X1 U20270 ( .A1(n17032), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17037) );
  AOI22_X1 U20271 ( .A1(n9716), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17036) );
  AOI22_X1 U20272 ( .A1(n17033), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17044), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17035) );
  AOI22_X1 U20273 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n9717), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17034) );
  NAND4_X1 U20274 ( .A1(n17037), .A2(n17036), .A3(n17035), .A4(n17034), .ZN(
        n17038) );
  NOR2_X1 U20275 ( .A1(n17039), .A2(n17038), .ZN(n17205) );
  OAI21_X1 U20276 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n9792), .A(n17040), .ZN(
        n17041) );
  AOI22_X1 U20277 ( .A1(n17089), .A2(n17205), .B1(n17041), .B2(n17079), .ZN(
        P3_U2694) );
  INV_X1 U20278 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17042) );
  NOR4_X1 U20279 ( .A1(n17042), .A2(n17067), .A3(n17074), .A4(n17073), .ZN(
        n17069) );
  AOI22_X1 U20280 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17079), .B1(
        P3_EBX_REG_7__SCAN_IN), .B2(n17069), .ZN(n17062) );
  AOI22_X1 U20281 ( .A1(n12590), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17060) );
  AOI22_X1 U20282 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16802), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17059) );
  AOI22_X1 U20283 ( .A1(n12585), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17047) );
  OAI21_X1 U20284 ( .B1(n9743), .B2(n18087), .A(n17047), .ZN(n17057) );
  AOI22_X1 U20285 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20286 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16740), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17054) );
  AOI22_X1 U20287 ( .A1(n17051), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U20288 ( .A1(n9718), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16755), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17052) );
  NAND4_X1 U20289 ( .A1(n17055), .A2(n17054), .A3(n17053), .A4(n17052), .ZN(
        n17056) );
  AOI211_X1 U20290 ( .C1(n9716), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n17057), .B(n17056), .ZN(n17058) );
  NAND3_X1 U20291 ( .A1(n17060), .A2(n17059), .A3(n17058), .ZN(n17209) );
  INV_X1 U20292 ( .A(n17209), .ZN(n17061) );
  OAI22_X1 U20293 ( .A1(n9792), .A2(n17062), .B1(n17061), .B2(n17079), .ZN(
        P3_U2695) );
  NAND3_X1 U20294 ( .A1(n17079), .A2(P3_EBX_REG_7__SCAN_IN), .A3(n17063), .ZN(
        n17066) );
  AOI22_X1 U20295 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17089), .B1(
        n17069), .B2(n17064), .ZN(n17065) );
  NAND2_X1 U20296 ( .A1(n17066), .A2(n17065), .ZN(P3_U2696) );
  NOR3_X1 U20297 ( .A1(n17067), .A2(n17074), .A3(n17073), .ZN(n17072) );
  AOI21_X1 U20298 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17079), .A(n17072), .ZN(
        n17068) );
  OAI22_X1 U20299 ( .A1(n17069), .A2(n17068), .B1(n20853), .B2(n17079), .ZN(
        P3_U2697) );
  OAI21_X1 U20300 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17070), .A(n17079), .ZN(
        n17071) );
  INV_X1 U20301 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18112) );
  OAI22_X1 U20302 ( .A1(n17072), .A2(n17071), .B1(n18112), .B2(n17079), .ZN(
        P3_U2698) );
  NOR2_X1 U20303 ( .A1(n17074), .A2(n17073), .ZN(n17077) );
  NAND3_X1 U20304 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17082), .A3(n17088), .ZN(
        n17078) );
  NOR2_X1 U20305 ( .A1(n17075), .A2(n17078), .ZN(n17081) );
  AOI21_X1 U20306 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17079), .A(n17081), .ZN(
        n17076) );
  OAI22_X1 U20307 ( .A1(n17077), .A2(n17076), .B1(n18107), .B2(n17079), .ZN(
        P3_U2699) );
  INV_X1 U20308 ( .A(n17078), .ZN(n17083) );
  AOI21_X1 U20309 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17079), .A(n17083), .ZN(
        n17080) );
  OAI22_X1 U20310 ( .A1(n17081), .A2(n17080), .B1(n18102), .B2(n17079), .ZN(
        P3_U2700) );
  INV_X1 U20311 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18097) );
  INV_X1 U20312 ( .A(n17085), .ZN(n17091) );
  AOI221_X1 U20313 ( .B1(n17082), .B2(n17091), .C1(n18119), .C2(n17091), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17084) );
  AOI211_X1 U20314 ( .C1(n17089), .C2(n18097), .A(n17084), .B(n17083), .ZN(
        P3_U2701) );
  AOI222_X1 U20315 ( .A1(n17086), .A2(n17088), .B1(P3_EBX_REG_1__SCAN_IN), 
        .B2(n17085), .C1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .C2(n17089), .ZN(
        n17087) );
  INV_X1 U20316 ( .A(n17087), .ZN(P3_U2702) );
  AOI22_X1 U20317 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17089), .B1(
        n17088), .B2(n20840), .ZN(n17090) );
  OAI21_X1 U20318 ( .B1(n17091), .B2(n20840), .A(n17090), .ZN(P3_U2703) );
  INV_X1 U20319 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17254) );
  INV_X1 U20320 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17258) );
  INV_X1 U20321 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17330) );
  INV_X1 U20322 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n20839) );
  INV_X1 U20323 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17337) );
  NAND4_X1 U20324 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17092) );
  NOR4_X1 U20325 ( .A1(n17330), .A2(n20839), .A3(n17337), .A4(n17092), .ZN(
        n17183) );
  NAND2_X1 U20326 ( .A1(n17242), .A2(n17183), .ZN(n17208) );
  NAND4_X1 U20327 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n17093)
         );
  NOR2_X1 U20328 ( .A1(n17208), .A2(n17093), .ZN(n17094) );
  NAND4_X1 U20329 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .A3(P3_EAX_REG_8__SCAN_IN), .A4(n17094), .ZN(n17176) );
  INV_X1 U20330 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17358) );
  INV_X1 U20331 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n20890) );
  INV_X1 U20332 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17265) );
  NAND4_X1 U20333 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17095)
         );
  NOR4_X2 U20334 ( .A1(n17171), .A2(n20890), .A3(n17265), .A4(n17095), .ZN(
        n17136) );
  NAND2_X1 U20335 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17136), .ZN(n17135) );
  NOR2_X2 U20336 ( .A1(n17254), .A2(n17116), .ZN(n17112) );
  NAND2_X1 U20337 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17112), .ZN(n17107) );
  NAND2_X1 U20338 ( .A1(n17103), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17102) );
  NAND2_X1 U20339 ( .A1(n17098), .A2(n17243), .ZN(n17145) );
  OAI22_X1 U20340 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17182), .B1(n17243), 
        .B2(n17103), .ZN(n17099) );
  AOI22_X1 U20341 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17169), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17099), .ZN(n17100) );
  OAI21_X1 U20342 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17102), .A(n17100), .ZN(
        P3_U2704) );
  AOI22_X1 U20343 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17170), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17169), .ZN(n17105) );
  OAI211_X1 U20344 ( .C1(n17103), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17234), .B(
        n17102), .ZN(n17104) );
  OAI211_X1 U20345 ( .C1(n17106), .C2(n17231), .A(n17105), .B(n17104), .ZN(
        P3_U2705) );
  AOI22_X1 U20346 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17170), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17169), .ZN(n17109) );
  OAI211_X1 U20347 ( .C1(n17112), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17234), .B(
        n17107), .ZN(n17108) );
  OAI211_X1 U20348 ( .C1(n17231), .C2(n17110), .A(n17109), .B(n17108), .ZN(
        P3_U2706) );
  INV_X1 U20349 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19105) );
  AOI22_X1 U20350 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17170), .B1(n17111), .B2(
        n17218), .ZN(n17115) );
  AOI211_X1 U20351 ( .C1(n17254), .C2(n17116), .A(n17112), .B(n17243), .ZN(
        n17113) );
  INV_X1 U20352 ( .A(n17113), .ZN(n17114) );
  OAI211_X1 U20353 ( .C1(n17145), .C2(n19105), .A(n17115), .B(n17114), .ZN(
        P3_U2707) );
  AOI22_X1 U20354 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17170), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17169), .ZN(n17118) );
  OAI211_X1 U20355 ( .C1(n17120), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17234), .B(
        n17116), .ZN(n17117) );
  OAI211_X1 U20356 ( .C1(n17119), .C2(n17231), .A(n17118), .B(n17117), .ZN(
        P3_U2708) );
  AOI22_X1 U20357 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17170), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17169), .ZN(n17123) );
  AOI211_X1 U20358 ( .C1(n17258), .C2(n17125), .A(n17120), .B(n17243), .ZN(
        n17121) );
  INV_X1 U20359 ( .A(n17121), .ZN(n17122) );
  OAI211_X1 U20360 ( .C1(n17124), .C2(n17231), .A(n17123), .B(n17122), .ZN(
        P3_U2709) );
  AOI22_X1 U20361 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17170), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17169), .ZN(n17128) );
  OAI211_X1 U20362 ( .C1(n17126), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17234), .B(
        n17125), .ZN(n17127) );
  OAI211_X1 U20363 ( .C1(n17129), .C2(n17231), .A(n17128), .B(n17127), .ZN(
        P3_U2710) );
  AOI22_X1 U20364 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17170), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17169), .ZN(n17133) );
  OAI211_X1 U20365 ( .C1(n17131), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17234), .B(
        n17130), .ZN(n17132) );
  OAI211_X1 U20366 ( .C1(n17134), .C2(n17231), .A(n17133), .B(n17132), .ZN(
        P3_U2711) );
  AOI22_X1 U20367 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17170), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17169), .ZN(n17138) );
  OAI211_X1 U20368 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17136), .A(n17234), .B(
        n17135), .ZN(n17137) );
  OAI211_X1 U20369 ( .C1(n17139), .C2(n17231), .A(n17138), .B(n17137), .ZN(
        P3_U2712) );
  INV_X1 U20370 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17269) );
  INV_X1 U20371 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17273) );
  NAND2_X1 U20372 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17163), .ZN(n17159) );
  NAND2_X1 U20373 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17154), .ZN(n17150) );
  NAND2_X1 U20374 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n20890), .ZN(n17144) );
  AOI22_X1 U20375 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17169), .B1(n17218), .B2(
        n17140), .ZN(n17143) );
  NAND2_X1 U20376 ( .A1(n17234), .A2(n17150), .ZN(n17149) );
  OAI21_X1 U20377 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17182), .A(n17149), .ZN(
        n17141) );
  AOI22_X1 U20378 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17170), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17141), .ZN(n17142) );
  OAI211_X1 U20379 ( .C1(n17150), .C2(n17144), .A(n17143), .B(n17142), .ZN(
        P3_U2713) );
  OAI22_X1 U20380 ( .A1(n17146), .A2(n17231), .B1(n14042), .B2(n17145), .ZN(
        n17147) );
  AOI21_X1 U20381 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17170), .A(n17147), .ZN(
        n17148) );
  OAI221_X1 U20382 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17150), .C1(n17265), 
        .C2(n17149), .A(n17148), .ZN(P3_U2714) );
  AOI22_X1 U20383 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17170), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17169), .ZN(n17152) );
  OAI211_X1 U20384 ( .C1(n17154), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17234), .B(
        n17150), .ZN(n17151) );
  OAI211_X1 U20385 ( .C1(n17153), .C2(n17231), .A(n17152), .B(n17151), .ZN(
        P3_U2715) );
  AOI22_X1 U20386 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17170), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17169), .ZN(n17157) );
  AOI211_X1 U20387 ( .C1(n17269), .C2(n17159), .A(n17154), .B(n17243), .ZN(
        n17155) );
  INV_X1 U20388 ( .A(n17155), .ZN(n17156) );
  OAI211_X1 U20389 ( .C1(n17158), .C2(n17231), .A(n17157), .B(n17156), .ZN(
        P3_U2716) );
  AOI22_X1 U20390 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17170), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17169), .ZN(n17161) );
  OAI211_X1 U20391 ( .C1(n17163), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17234), .B(
        n17159), .ZN(n17160) );
  OAI211_X1 U20392 ( .C1(n17162), .C2(n17231), .A(n17161), .B(n17160), .ZN(
        P3_U2717) );
  AOI22_X1 U20393 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17170), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17169), .ZN(n17167) );
  INV_X1 U20394 ( .A(n17171), .ZN(n17165) );
  INV_X1 U20395 ( .A(n17163), .ZN(n17164) );
  OAI211_X1 U20396 ( .C1(n17165), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17234), .B(
        n17164), .ZN(n17166) );
  OAI211_X1 U20397 ( .C1(n17168), .C2(n17231), .A(n17167), .B(n17166), .ZN(
        P3_U2718) );
  AOI22_X1 U20398 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17170), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17169), .ZN(n17174) );
  OAI211_X1 U20399 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17172), .A(n17234), .B(
        n17171), .ZN(n17173) );
  OAI211_X1 U20400 ( .C1(n17175), .C2(n17231), .A(n17174), .B(n17173), .ZN(
        P3_U2719) );
  NOR2_X1 U20401 ( .A1(n18119), .A2(n17176), .ZN(n17178) );
  NAND2_X1 U20402 ( .A1(n17234), .A2(n17176), .ZN(n17186) );
  INV_X1 U20403 ( .A(n17186), .ZN(n17177) );
  MUX2_X1 U20404 ( .A(n17178), .B(n17177), .S(P3_EAX_REG_15__SCAN_IN), .Z(
        n17179) );
  AOI21_X1 U20405 ( .B1(BUF2_REG_15__SCAN_IN), .B2(n17241), .A(n17179), .ZN(
        n17180) );
  OAI21_X1 U20406 ( .B1(n17181), .B2(n17231), .A(n17180), .ZN(P3_U2720) );
  INV_X1 U20407 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20848) );
  INV_X1 U20408 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17199) );
  INV_X1 U20409 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17339) );
  NAND2_X1 U20410 ( .A1(n17183), .A2(n17240), .ZN(n17213) );
  NOR2_X1 U20411 ( .A1(n17339), .A2(n17213), .ZN(n17204) );
  NAND2_X1 U20412 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17204), .ZN(n17203) );
  NAND2_X1 U20413 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17198), .ZN(n17191) );
  NOR2_X1 U20414 ( .A1(n20848), .A2(n17191), .ZN(n17194) );
  NAND2_X1 U20415 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17194), .ZN(n17187) );
  INV_X1 U20416 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U20417 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17241), .B1(n17218), .B2(
        n17184), .ZN(n17185) );
  OAI221_X1 U20418 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17187), .C1(n17353), 
        .C2(n17186), .A(n17185), .ZN(P3_U2721) );
  INV_X1 U20419 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17351) );
  INV_X1 U20420 ( .A(n17187), .ZN(n17190) );
  AOI21_X1 U20421 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17234), .A(n17194), .ZN(
        n17189) );
  OAI222_X1 U20422 ( .A1(n17239), .A2(n17351), .B1(n17190), .B2(n17189), .C1(
        n17231), .C2(n17188), .ZN(P3_U2722) );
  INV_X1 U20423 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17347) );
  INV_X1 U20424 ( .A(n17191), .ZN(n17197) );
  AOI21_X1 U20425 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17234), .A(n17197), .ZN(
        n17193) );
  OAI222_X1 U20426 ( .A1(n17239), .A2(n17347), .B1(n17194), .B2(n17193), .C1(
        n17231), .C2(n17192), .ZN(P3_U2723) );
  AOI21_X1 U20427 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17234), .A(n17198), .ZN(
        n17196) );
  OAI222_X1 U20428 ( .A1(n17239), .A2(n17345), .B1(n17197), .B2(n17196), .C1(
        n17231), .C2(n17195), .ZN(P3_U2724) );
  AOI211_X1 U20429 ( .C1(n17199), .C2(n17203), .A(n17243), .B(n17198), .ZN(
        n17200) );
  AOI21_X1 U20430 ( .B1(n17241), .B2(BUF2_REG_10__SCAN_IN), .A(n17200), .ZN(
        n17201) );
  OAI21_X1 U20431 ( .B1(n17202), .B2(n17231), .A(n17201), .ZN(P3_U2725) );
  INV_X1 U20432 ( .A(n17203), .ZN(n17207) );
  AOI21_X1 U20433 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17234), .A(n17204), .ZN(
        n17206) );
  OAI222_X1 U20434 ( .A1(n17239), .A2(n17341), .B1(n17207), .B2(n17206), .C1(
        n17231), .C2(n17205), .ZN(P3_U2726) );
  NAND2_X1 U20435 ( .A1(n17234), .A2(n17208), .ZN(n17211) );
  AOI22_X1 U20436 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17241), .B1(n17218), .B2(
        n17209), .ZN(n17210) );
  OAI221_X1 U20437 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n17213), .C1(n17339), 
        .C2(n17211), .A(n17210), .ZN(P3_U2727) );
  INV_X1 U20438 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17296) );
  NAND3_X1 U20439 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(n17240), .ZN(n17229) );
  NOR2_X1 U20440 ( .A1(n17296), .A2(n17229), .ZN(n17233) );
  NAND2_X1 U20441 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17228), .ZN(n17216) );
  INV_X1 U20442 ( .A(n17216), .ZN(n17224) );
  NAND2_X1 U20443 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17224), .ZN(n17220) );
  OAI21_X1 U20444 ( .B1(n17243), .B2(n17337), .A(n17220), .ZN(n17212) );
  AOI22_X1 U20445 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17241), .B1(n17213), .B2(
        n17212), .ZN(n17214) );
  OAI21_X1 U20446 ( .B1(n17215), .B2(n17231), .A(n17214), .ZN(P3_U2728) );
  INV_X1 U20447 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17291) );
  OAI21_X1 U20448 ( .B1(n17291), .B2(n17243), .A(n17216), .ZN(n17219) );
  AOI222_X1 U20449 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17241), .B1(n17220), .B2(
        n17219), .C1(n17218), .C2(n17217), .ZN(n17221) );
  INV_X1 U20450 ( .A(n17221), .ZN(P3_U2729) );
  INV_X1 U20451 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18108) );
  AOI21_X1 U20452 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17234), .A(n17228), .ZN(
        n17223) );
  OAI222_X1 U20453 ( .A1(n18108), .A2(n17239), .B1(n17224), .B2(n17223), .C1(
        n17231), .C2(n17222), .ZN(P3_U2730) );
  INV_X1 U20454 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18103) );
  AOI21_X1 U20455 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17234), .A(n17233), .ZN(
        n17227) );
  INV_X1 U20456 ( .A(n17225), .ZN(n17226) );
  OAI222_X1 U20457 ( .A1(n18103), .A2(n17239), .B1(n17228), .B2(n17227), .C1(
        n17231), .C2(n17226), .ZN(P3_U2731) );
  INV_X1 U20458 ( .A(n17229), .ZN(n17238) );
  AOI21_X1 U20459 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17234), .A(n17238), .ZN(
        n17232) );
  OAI222_X1 U20460 ( .A1(n18098), .A2(n17239), .B1(n17233), .B2(n17232), .C1(
        n17231), .C2(n17230), .ZN(P3_U2732) );
  AOI22_X1 U20461 ( .A1(n17240), .A2(P3_EAX_REG_1__SCAN_IN), .B1(
        P3_EAX_REG_2__SCAN_IN), .B2(n17234), .ZN(n17237) );
  INV_X1 U20462 ( .A(n17235), .ZN(n17236) );
  OAI222_X1 U20463 ( .A1(n18093), .A2(n17239), .B1(n17238), .B2(n17237), .C1(
        n17231), .C2(n17236), .ZN(P3_U2733) );
  AOI22_X1 U20464 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17241), .B1(n17240), .B2(
        n17330), .ZN(n17245) );
  OR3_X1 U20465 ( .A1(n17330), .A2(n17243), .A3(n17242), .ZN(n17244) );
  OAI211_X1 U20466 ( .C1(n17246), .C2(n17231), .A(n17245), .B(n17244), .ZN(
        P3_U2734) );
  INV_X1 U20467 ( .A(n18592), .ZN(n17444) );
  NAND2_X1 U20468 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17444), .ZN(n17287) );
  INV_X1 U20469 ( .A(n17307), .ZN(n17248) );
  NOR2_X1 U20470 ( .A1(n17272), .A2(n17249), .ZN(P3_U2736) );
  INV_X1 U20471 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17327) );
  NOR2_X1 U20472 ( .A1(n17303), .A2(n18084), .ZN(n17270) );
  INV_X1 U20473 ( .A(n17270), .ZN(n17275) );
  INV_X2 U20474 ( .A(n17287), .ZN(n17301) );
  AOI22_X1 U20475 ( .A1(n17301), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17250) );
  OAI21_X1 U20476 ( .B1(n17327), .B2(n17275), .A(n17250), .ZN(P3_U2737) );
  INV_X1 U20477 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17252) );
  AOI22_X1 U20478 ( .A1(n17301), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17251) );
  OAI21_X1 U20479 ( .B1(n17252), .B2(n17275), .A(n17251), .ZN(P3_U2738) );
  AOI22_X1 U20480 ( .A1(n17301), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17253) );
  OAI21_X1 U20481 ( .B1(n17254), .B2(n17275), .A(n17253), .ZN(P3_U2739) );
  INV_X1 U20482 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17256) );
  AOI22_X1 U20483 ( .A1(n17301), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17255) );
  OAI21_X1 U20484 ( .B1(n17256), .B2(n17275), .A(n17255), .ZN(P3_U2740) );
  AOI22_X1 U20485 ( .A1(n17301), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17257) );
  OAI21_X1 U20486 ( .B1(n17258), .B2(n17275), .A(n17257), .ZN(P3_U2741) );
  INV_X1 U20487 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17260) );
  AOI22_X1 U20488 ( .A1(P3_DATAO_REG_25__SCAN_IN), .A2(n17300), .B1(n17301), 
        .B2(P3_UWORD_REG_9__SCAN_IN), .ZN(n17259) );
  OAI21_X1 U20489 ( .B1(n17260), .B2(n17275), .A(n17259), .ZN(P3_U2742) );
  INV_X1 U20490 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17320) );
  AOI22_X1 U20491 ( .A1(n17301), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17261) );
  OAI21_X1 U20492 ( .B1(n17320), .B2(n17275), .A(n17261), .ZN(P3_U2743) );
  INV_X1 U20493 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17318) );
  AOI22_X1 U20494 ( .A1(n17301), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17262) );
  OAI21_X1 U20495 ( .B1(n17318), .B2(n17275), .A(n17262), .ZN(P3_U2744) );
  AOI22_X1 U20496 ( .A1(n17301), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17263) );
  OAI21_X1 U20497 ( .B1(n20890), .B2(n17275), .A(n17263), .ZN(P3_U2745) );
  AOI22_X1 U20498 ( .A1(n17301), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17264) );
  OAI21_X1 U20499 ( .B1(n17265), .B2(n17275), .A(n17264), .ZN(P3_U2746) );
  INV_X1 U20500 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17267) );
  AOI22_X1 U20501 ( .A1(n17301), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17266) );
  OAI21_X1 U20502 ( .B1(n17267), .B2(n17275), .A(n17266), .ZN(P3_U2747) );
  AOI22_X1 U20503 ( .A1(n17301), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17268) );
  OAI21_X1 U20504 ( .B1(n17269), .B2(n17275), .A(n17268), .ZN(P3_U2748) );
  INV_X1 U20505 ( .A(P3_UWORD_REG_2__SCAN_IN), .ZN(n20905) );
  AOI22_X1 U20506 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17270), .B1(n17300), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17271) );
  OAI21_X1 U20507 ( .B1(n20905), .B2(n17287), .A(n17271), .ZN(P3_U2749) );
  INV_X1 U20508 ( .A(P3_UWORD_REG_1__SCAN_IN), .ZN(n21046) );
  INV_X1 U20509 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n20954) );
  OAI222_X1 U20510 ( .A1(n17287), .A2(n21046), .B1(n17275), .B2(n17273), .C1(
        n20954), .C2(n17272), .ZN(P3_U2750) );
  INV_X1 U20511 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17276) );
  AOI22_X1 U20512 ( .A1(n17301), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17274) );
  OAI21_X1 U20513 ( .B1(n17276), .B2(n17275), .A(n17274), .ZN(P3_U2751) );
  AOI22_X1 U20514 ( .A1(n17301), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17277) );
  OAI21_X1 U20515 ( .B1(n17358), .B2(n17303), .A(n17277), .ZN(P3_U2752) );
  INV_X1 U20516 ( .A(P3_LWORD_REG_14__SCAN_IN), .ZN(n20972) );
  INV_X1 U20517 ( .A(n17303), .ZN(n17285) );
  AOI22_X1 U20518 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17285), .B1(n17300), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17278) );
  OAI21_X1 U20519 ( .B1(n20972), .B2(n17287), .A(n17278), .ZN(P3_U2753) );
  INV_X1 U20520 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17280) );
  AOI22_X1 U20521 ( .A1(n17301), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17279) );
  OAI21_X1 U20522 ( .B1(n17280), .B2(n17303), .A(n17279), .ZN(P3_U2754) );
  AOI22_X1 U20523 ( .A1(n17301), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17281) );
  OAI21_X1 U20524 ( .B1(n20848), .B2(n17303), .A(n17281), .ZN(P3_U2755) );
  INV_X1 U20525 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17283) );
  AOI22_X1 U20526 ( .A1(n17301), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17282) );
  OAI21_X1 U20527 ( .B1(n17283), .B2(n17303), .A(n17282), .ZN(P3_U2756) );
  INV_X1 U20528 ( .A(P3_LWORD_REG_10__SCAN_IN), .ZN(n20934) );
  AOI22_X1 U20529 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17285), .B1(n17300), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17284) );
  OAI21_X1 U20530 ( .B1(n20934), .B2(n17287), .A(n17284), .ZN(P3_U2757) );
  INV_X1 U20531 ( .A(P3_LWORD_REG_9__SCAN_IN), .ZN(n20836) );
  AOI22_X1 U20532 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17285), .B1(n17300), .B2(
        P3_DATAO_REG_9__SCAN_IN), .ZN(n17286) );
  OAI21_X1 U20533 ( .B1(n20836), .B2(n17287), .A(n17286), .ZN(P3_U2758) );
  AOI22_X1 U20534 ( .A1(n17301), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17288) );
  OAI21_X1 U20535 ( .B1(n17339), .B2(n17303), .A(n17288), .ZN(P3_U2759) );
  AOI22_X1 U20536 ( .A1(n17301), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17289) );
  OAI21_X1 U20537 ( .B1(n17337), .B2(n17303), .A(n17289), .ZN(P3_U2760) );
  AOI22_X1 U20538 ( .A1(n17301), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17290) );
  OAI21_X1 U20539 ( .B1(n17291), .B2(n17303), .A(n17290), .ZN(P3_U2761) );
  AOI22_X1 U20540 ( .A1(n17301), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17292) );
  OAI21_X1 U20541 ( .B1(n20839), .B2(n17303), .A(n17292), .ZN(P3_U2762) );
  INV_X1 U20542 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17294) );
  AOI22_X1 U20543 ( .A1(n17301), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17293) );
  OAI21_X1 U20544 ( .B1(n17294), .B2(n17303), .A(n17293), .ZN(P3_U2763) );
  AOI22_X1 U20545 ( .A1(n17301), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17295) );
  OAI21_X1 U20546 ( .B1(n17296), .B2(n17303), .A(n17295), .ZN(P3_U2764) );
  INV_X1 U20547 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17298) );
  AOI22_X1 U20548 ( .A1(n17301), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17297) );
  OAI21_X1 U20549 ( .B1(n17298), .B2(n17303), .A(n17297), .ZN(P3_U2765) );
  AOI22_X1 U20550 ( .A1(n17301), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17299) );
  OAI21_X1 U20551 ( .B1(n17330), .B2(n17303), .A(n17299), .ZN(P3_U2766) );
  AOI22_X1 U20552 ( .A1(n17301), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17300), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17302) );
  OAI21_X1 U20553 ( .B1(n17304), .B2(n17303), .A(n17302), .ZN(P3_U2767) );
  NAND2_X1 U20554 ( .A1(n17306), .A2(n17305), .ZN(n18572) );
  INV_X2 U20555 ( .A(n17311), .ZN(n17354) );
  NAND2_X1 U20556 ( .A1(n18090), .A2(n17311), .ZN(n17357) );
  AOI22_X1 U20557 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17348), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17354), .ZN(n17309) );
  OAI21_X1 U20558 ( .B1(n18081), .B2(n17350), .A(n17309), .ZN(P3_U2768) );
  AOI22_X1 U20559 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17355), .B1(
        P3_EAX_REG_17__SCAN_IN), .B2(n17348), .ZN(n17310) );
  OAI21_X1 U20560 ( .B1(n17311), .B2(n21046), .A(n17310), .ZN(P3_U2769) );
  AOI22_X1 U20561 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17348), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17354), .ZN(n17312) );
  OAI21_X1 U20562 ( .B1(n18093), .B2(n17350), .A(n17312), .ZN(P3_U2770) );
  AOI22_X1 U20563 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17348), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17354), .ZN(n17313) );
  OAI21_X1 U20564 ( .B1(n18098), .B2(n17350), .A(n17313), .ZN(P3_U2771) );
  AOI22_X1 U20565 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17348), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17354), .ZN(n17314) );
  OAI21_X1 U20566 ( .B1(n18103), .B2(n17350), .A(n17314), .ZN(P3_U2772) );
  AOI22_X1 U20567 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17348), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17354), .ZN(n17315) );
  OAI21_X1 U20568 ( .B1(n18108), .B2(n17350), .A(n17315), .ZN(P3_U2773) );
  AOI22_X1 U20569 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17348), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17354), .ZN(n17316) );
  OAI21_X1 U20570 ( .B1(n18113), .B2(n17350), .A(n17316), .ZN(P3_U2774) );
  AOI22_X1 U20571 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17355), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17354), .ZN(n17317) );
  OAI21_X1 U20572 ( .B1(n17318), .B2(n17357), .A(n17317), .ZN(P3_U2775) );
  AOI22_X1 U20573 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17355), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17354), .ZN(n17319) );
  OAI21_X1 U20574 ( .B1(n17320), .B2(n17357), .A(n17319), .ZN(P3_U2776) );
  AOI22_X1 U20575 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17348), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17354), .ZN(n17321) );
  OAI21_X1 U20576 ( .B1(n17341), .B2(n17350), .A(n17321), .ZN(P3_U2777) );
  INV_X1 U20577 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17343) );
  AOI22_X1 U20578 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17348), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17354), .ZN(n17322) );
  OAI21_X1 U20579 ( .B1(n17343), .B2(n17350), .A(n17322), .ZN(P3_U2778) );
  AOI22_X1 U20580 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17348), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17354), .ZN(n17323) );
  OAI21_X1 U20581 ( .B1(n17345), .B2(n17350), .A(n17323), .ZN(P3_U2779) );
  AOI22_X1 U20582 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17348), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17354), .ZN(n17324) );
  OAI21_X1 U20583 ( .B1(n17347), .B2(n17350), .A(n17324), .ZN(P3_U2780) );
  AOI22_X1 U20584 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17348), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17354), .ZN(n17325) );
  OAI21_X1 U20585 ( .B1(n17351), .B2(n17350), .A(n17325), .ZN(P3_U2781) );
  AOI22_X1 U20586 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17355), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17354), .ZN(n17326) );
  OAI21_X1 U20587 ( .B1(n17327), .B2(n17357), .A(n17326), .ZN(P3_U2782) );
  AOI22_X1 U20588 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17348), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17354), .ZN(n17328) );
  OAI21_X1 U20589 ( .B1(n18081), .B2(n17350), .A(n17328), .ZN(P3_U2783) );
  AOI22_X1 U20590 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17355), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17354), .ZN(n17329) );
  OAI21_X1 U20591 ( .B1(n17330), .B2(n17357), .A(n17329), .ZN(P3_U2784) );
  AOI22_X1 U20592 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17348), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17354), .ZN(n17331) );
  OAI21_X1 U20593 ( .B1(n18093), .B2(n17350), .A(n17331), .ZN(P3_U2785) );
  AOI22_X1 U20594 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17348), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17354), .ZN(n17332) );
  OAI21_X1 U20595 ( .B1(n18098), .B2(n17350), .A(n17332), .ZN(P3_U2786) );
  AOI22_X1 U20596 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17348), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17354), .ZN(n17333) );
  OAI21_X1 U20597 ( .B1(n18103), .B2(n17350), .A(n17333), .ZN(P3_U2787) );
  AOI22_X1 U20598 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17348), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17354), .ZN(n17334) );
  OAI21_X1 U20599 ( .B1(n18108), .B2(n17350), .A(n17334), .ZN(P3_U2788) );
  AOI22_X1 U20600 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17348), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17354), .ZN(n17335) );
  OAI21_X1 U20601 ( .B1(n18113), .B2(n17350), .A(n17335), .ZN(P3_U2789) );
  AOI22_X1 U20602 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17355), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17354), .ZN(n17336) );
  OAI21_X1 U20603 ( .B1(n17337), .B2(n17357), .A(n17336), .ZN(P3_U2790) );
  AOI22_X1 U20604 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17355), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17354), .ZN(n17338) );
  OAI21_X1 U20605 ( .B1(n17339), .B2(n17357), .A(n17338), .ZN(P3_U2791) );
  AOI22_X1 U20606 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17348), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17354), .ZN(n17340) );
  OAI21_X1 U20607 ( .B1(n17341), .B2(n17350), .A(n17340), .ZN(P3_U2792) );
  AOI22_X1 U20608 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17348), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17354), .ZN(n17342) );
  OAI21_X1 U20609 ( .B1(n17343), .B2(n17350), .A(n17342), .ZN(P3_U2793) );
  AOI22_X1 U20610 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17348), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17354), .ZN(n17344) );
  OAI21_X1 U20611 ( .B1(n17345), .B2(n17350), .A(n17344), .ZN(P3_U2794) );
  AOI22_X1 U20612 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17348), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17354), .ZN(n17346) );
  OAI21_X1 U20613 ( .B1(n17347), .B2(n17350), .A(n17346), .ZN(P3_U2795) );
  AOI22_X1 U20614 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17348), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17354), .ZN(n17349) );
  OAI21_X1 U20615 ( .B1(n17351), .B2(n17350), .A(n17349), .ZN(P3_U2796) );
  AOI22_X1 U20616 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17355), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17354), .ZN(n17352) );
  OAI21_X1 U20617 ( .B1(n17353), .B2(n17357), .A(n17352), .ZN(P3_U2797) );
  AOI22_X1 U20618 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17355), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17354), .ZN(n17356) );
  OAI21_X1 U20619 ( .B1(n17358), .B2(n17357), .A(n17356), .ZN(P3_U2798) );
  AOI21_X1 U20620 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17390), .A(
        n18592), .ZN(n17359) );
  AOI211_X1 U20621 ( .C1(n17705), .C2(n12349), .A(n17630), .B(n17359), .ZN(
        n17394) );
  OAI21_X1 U20622 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17508), .A(
        n17394), .ZN(n17384) );
  AOI22_X1 U20623 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17384), .B1(
        n17530), .B2(n17360), .ZN(n17374) );
  AOI21_X1 U20624 ( .B1(n17363), .B2(n17362), .A(n17361), .ZN(n17369) );
  NOR3_X1 U20625 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n9918), .A3(
        n17386), .ZN(n17368) );
  NOR3_X1 U20626 ( .A1(n17881), .A2(n17365), .A3(n17759), .ZN(n17742) );
  NOR3_X1 U20627 ( .A1(n17365), .A2(n17883), .A3(n17759), .ZN(n17741) );
  OAI22_X1 U20628 ( .A1(n17742), .A2(n17600), .B1(n17741), .B2(n17735), .ZN(
        n17396) );
  NOR2_X1 U20629 ( .A1(n9918), .A2(n17396), .ZN(n17387) );
  AOI211_X1 U20630 ( .C1(n17600), .C2(n17735), .A(n17387), .B(n17366), .ZN(
        n17367) );
  AOI211_X1 U20631 ( .C1(n17639), .C2(n17369), .A(n17368), .B(n17367), .ZN(
        n17373) );
  NOR2_X1 U20632 ( .A1(n17572), .A2(n12349), .ZN(n17376) );
  OAI211_X1 U20633 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17376), .B(n17370), .ZN(n17371) );
  NAND4_X1 U20634 ( .A1(n17374), .A2(n17373), .A3(n17372), .A4(n17371), .ZN(
        P3_U2802) );
  OAI22_X1 U20635 ( .A1(n17892), .A2(n18656), .B1(n17583), .B2(n17375), .ZN(
        n17383) );
  INV_X1 U20636 ( .A(n17376), .ZN(n17381) );
  INV_X1 U20637 ( .A(n17377), .ZN(n17379) );
  NAND2_X1 U20638 ( .A1(n17379), .A2(n17378), .ZN(n17380) );
  OAI22_X1 U20639 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17381), .B1(
        n17750), .B2(n17627), .ZN(n17382) );
  OAI221_X1 U20640 ( .B1(n17387), .B2(n9918), .C1(n17387), .C2(n17386), .A(
        n17385), .ZN(P3_U2803) );
  AOI21_X1 U20641 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17389), .A(
        n9724), .ZN(n17757) );
  AOI21_X1 U20642 ( .B1(n17390), .B2(n18460), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17393) );
  OAI21_X1 U20643 ( .B1(n17530), .B2(n17476), .A(n17391), .ZN(n17392) );
  NAND2_X1 U20644 ( .A1(n18061), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17755) );
  OAI211_X1 U20645 ( .C1(n17394), .C2(n17393), .A(n17392), .B(n17755), .ZN(
        n17395) );
  AOI221_X1 U20646 ( .B1(n17397), .B2(n17751), .C1(n17396), .C2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n17395), .ZN(n17398) );
  OAI21_X1 U20647 ( .B1(n17757), .B2(n17627), .A(n17398), .ZN(P3_U2804) );
  NOR3_X1 U20648 ( .A1(n17760), .A2(n17883), .A3(n17759), .ZN(n17399) );
  XOR2_X1 U20649 ( .A(n17763), .B(n17399), .Z(n17772) );
  AOI21_X1 U20650 ( .B1(n18460), .B2(n17401), .A(n17630), .ZN(n17423) );
  OAI21_X1 U20651 ( .B1(n17400), .B2(n18592), .A(n17423), .ZN(n17414) );
  NOR2_X1 U20652 ( .A1(n17572), .A2(n17401), .ZN(n17415) );
  OAI211_X1 U20653 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17415), .B(n17402), .ZN(n17404) );
  NOR2_X1 U20654 ( .A1(n18044), .A2(n18652), .ZN(n17767) );
  INV_X1 U20655 ( .A(n17767), .ZN(n17403) );
  OAI211_X1 U20656 ( .C1(n17583), .C2(n17405), .A(n17404), .B(n17403), .ZN(
        n17406) );
  AOI21_X1 U20657 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17414), .A(
        n17406), .ZN(n17412) );
  NOR3_X1 U20658 ( .A1(n17759), .A2(n17760), .A3(n17881), .ZN(n17407) );
  XOR2_X1 U20659 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17407), .Z(
        n17769) );
  AOI21_X1 U20660 ( .B1(n17409), .B2(n17636), .A(n17408), .ZN(n17410) );
  XOR2_X1 U20661 ( .A(n17410), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17768) );
  AOI22_X1 U20662 ( .A1(n17640), .A2(n17769), .B1(n17639), .B2(n17768), .ZN(
        n17411) );
  OAI211_X1 U20663 ( .C1(n17735), .C2(n17772), .A(n17412), .B(n17411), .ZN(
        P3_U2805) );
  NOR2_X1 U20664 ( .A1(n18044), .A2(n18650), .ZN(n17775) );
  AOI221_X1 U20665 ( .B1(n17415), .B2(n20851), .C1(n17414), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17775), .ZN(n17421) );
  INV_X1 U20666 ( .A(n17881), .ZN(n17800) );
  AOI21_X1 U20667 ( .B1(n17800), .B2(n17777), .A(n17600), .ZN(n17433) );
  NOR3_X1 U20668 ( .A1(n17782), .A2(n17883), .A3(n17759), .ZN(n17781) );
  NOR2_X1 U20669 ( .A1(n17781), .A2(n17735), .ZN(n17434) );
  AOI21_X1 U20670 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17417), .A(
        n17416), .ZN(n17774) );
  INV_X1 U20671 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17418) );
  NAND2_X1 U20672 ( .A1(n17777), .A2(n17418), .ZN(n17788) );
  OAI22_X1 U20673 ( .A1(n17774), .A2(n17627), .B1(n17536), .B2(n17788), .ZN(
        n17419) );
  AOI221_X1 U20674 ( .B1(n17433), .B2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), 
        .C1(n17434), .C2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A(n17419), .ZN(
        n17420) );
  OAI211_X1 U20675 ( .C1(n17583), .C2(n12365), .A(n17421), .B(n17420), .ZN(
        P3_U2806) );
  NAND2_X1 U20676 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17448) );
  INV_X1 U20677 ( .A(n17572), .ZN(n17523) );
  NAND2_X1 U20678 ( .A1(n17447), .A2(n17523), .ZN(n17459) );
  NOR3_X1 U20679 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17448), .A3(
        n17459), .ZN(n17426) );
  AOI221_X1 U20680 ( .B1(n17424), .B2(n17423), .C1(n18592), .C2(n17423), .A(
        n17422), .ZN(n17425) );
  AOI211_X1 U20681 ( .C1(n17530), .C2(n17427), .A(n17426), .B(n17425), .ZN(
        n17438) );
  AOI22_X1 U20682 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17636), .B1(
        n17429), .B2(n17441), .ZN(n17430) );
  NAND2_X1 U20683 ( .A1(n17428), .A2(n17430), .ZN(n17431) );
  XOR2_X1 U20684 ( .A(n17431), .B(n17782), .Z(n17789) );
  OAI21_X1 U20685 ( .B1(n17881), .B2(n17759), .A(n17782), .ZN(n17432) );
  AOI22_X1 U20686 ( .A1(n17639), .A2(n17789), .B1(n17433), .B2(n17432), .ZN(
        n17437) );
  NOR2_X1 U20687 ( .A1(n17883), .A2(n17759), .ZN(n17435) );
  OAI21_X1 U20688 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17435), .A(
        n17434), .ZN(n17436) );
  NAND2_X1 U20689 ( .A1(n18061), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17793) );
  NAND4_X1 U20690 ( .A1(n17438), .A2(n17437), .A3(n17436), .A4(n17793), .ZN(
        P3_U2807) );
  INV_X1 U20691 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17804) );
  NAND2_X1 U20692 ( .A1(n17439), .A2(n17471), .ZN(n17805) );
  INV_X1 U20693 ( .A(n17428), .ZN(n17440) );
  AOI221_X1 U20694 ( .B1(n17521), .B2(n17441), .C1(n17805), .C2(n17441), .A(
        n17440), .ZN(n17442) );
  XOR2_X1 U20695 ( .A(n17804), .B(n17442), .Z(n17811) );
  INV_X1 U20696 ( .A(n17705), .ZN(n17446) );
  AOI21_X1 U20697 ( .B1(n17444), .B2(n17443), .A(n17630), .ZN(n17445) );
  OAI21_X1 U20698 ( .B1(n17447), .B2(n17446), .A(n17445), .ZN(n17481) );
  AOI21_X1 U20699 ( .B1(n17476), .B2(n17474), .A(n17481), .ZN(n17457) );
  NAND2_X1 U20700 ( .A1(n18061), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17809) );
  INV_X1 U20701 ( .A(n17459), .ZN(n17449) );
  OAI211_X1 U20702 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17449), .B(n17448), .ZN(n17450) );
  OAI211_X1 U20703 ( .C1(n17457), .C2(n21049), .A(n17809), .B(n17450), .ZN(
        n17454) );
  NOR2_X1 U20704 ( .A1(n17536), .A2(n17805), .ZN(n17452) );
  NAND2_X1 U20705 ( .A1(n17600), .A2(n17735), .ZN(n17473) );
  AOI22_X1 U20706 ( .A1(n17881), .A2(n17640), .B1(n17883), .B2(n17537), .ZN(
        n17535) );
  INV_X1 U20707 ( .A(n17535), .ZN(n17472) );
  AOI21_X1 U20708 ( .B1(n17473), .B2(n17805), .A(n17472), .ZN(n17470) );
  INV_X1 U20709 ( .A(n17470), .ZN(n17451) );
  MUX2_X1 U20710 ( .A(n17452), .B(n17451), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17453) );
  AOI211_X1 U20711 ( .C1(n17530), .C2(n17455), .A(n17454), .B(n17453), .ZN(
        n17456) );
  OAI21_X1 U20712 ( .B1(n17627), .B2(n17811), .A(n17456), .ZN(P3_U2808) );
  NAND2_X1 U20713 ( .A1(n18061), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n17822) );
  OAI221_X1 U20714 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17459), .C1(
        n17458), .C2(n17457), .A(n17822), .ZN(n17460) );
  AOI21_X1 U20715 ( .B1(n17530), .B2(n17461), .A(n17460), .ZN(n17468) );
  NOR3_X1 U20716 ( .A1(n17636), .A2(n17850), .A3(n17462), .ZN(n17492) );
  INV_X1 U20717 ( .A(n17463), .ZN(n17504) );
  AOI22_X1 U20718 ( .A1(n17819), .A2(n17492), .B1(n17504), .B2(n17464), .ZN(
        n17465) );
  XOR2_X1 U20719 ( .A(n17469), .B(n17465), .Z(n17815) );
  NOR2_X1 U20720 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17466), .ZN(
        n17814) );
  NOR2_X1 U20721 ( .A1(n17813), .A2(n17536), .ZN(n17494) );
  AOI22_X1 U20722 ( .A1(n17639), .A2(n17815), .B1(n17814), .B2(n17494), .ZN(
        n17467) );
  OAI211_X1 U20723 ( .C1(n17470), .C2(n17469), .A(n17468), .B(n17467), .ZN(
        P3_U2809) );
  NAND2_X1 U20724 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17471), .ZN(
        n17825) );
  AOI21_X1 U20725 ( .B1(n17473), .B2(n17825), .A(n17472), .ZN(n17497) );
  OAI21_X1 U20726 ( .B1(n18190), .B2(n17475), .A(n17474), .ZN(n17480) );
  AOI21_X1 U20727 ( .B1(n17583), .B2(n17508), .A(n17477), .ZN(n17479) );
  NAND2_X1 U20728 ( .A1(n18061), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17831) );
  INV_X1 U20729 ( .A(n17831), .ZN(n17478) );
  AOI211_X1 U20730 ( .C1(n17481), .C2(n17480), .A(n17479), .B(n17478), .ZN(
        n17484) );
  OAI221_X1 U20731 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17503), 
        .C1(n17837), .C2(n17492), .A(n17428), .ZN(n17482) );
  XOR2_X1 U20732 ( .A(n17833), .B(n17482), .Z(n17830) );
  NOR2_X1 U20733 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17837), .ZN(
        n17829) );
  AOI22_X1 U20734 ( .A1(n17639), .A2(n17830), .B1(n17494), .B2(n17829), .ZN(
        n17483) );
  OAI211_X1 U20735 ( .C1(n17497), .C2(n17833), .A(n17484), .B(n17483), .ZN(
        P3_U2810) );
  AOI21_X1 U20736 ( .B1(n17705), .B2(n17485), .A(n17630), .ZN(n17511) );
  OAI21_X1 U20737 ( .B1(n17486), .B2(n18592), .A(n17511), .ZN(n17501) );
  NOR2_X1 U20738 ( .A1(n18044), .A2(n18642), .ZN(n17836) );
  NAND2_X1 U20739 ( .A1(n17487), .A2(n17523), .ZN(n17499) );
  OAI21_X1 U20740 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17488), .ZN(n17489) );
  OAI22_X1 U20741 ( .A1(n17583), .A2(n17490), .B1(n17499), .B2(n17489), .ZN(
        n17491) );
  AOI211_X1 U20742 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n17501), .A(
        n17836), .B(n17491), .ZN(n17496) );
  AOI21_X1 U20743 ( .B1(n17503), .B2(n17504), .A(n17492), .ZN(n17493) );
  XOR2_X1 U20744 ( .A(n17837), .B(n17493), .Z(n17835) );
  AOI22_X1 U20745 ( .A1(n17639), .A2(n17835), .B1(n17494), .B2(n17837), .ZN(
        n17495) );
  OAI211_X1 U20746 ( .C1(n17497), .C2(n17837), .A(n17496), .B(n17495), .ZN(
        P3_U2811) );
  NAND2_X1 U20747 ( .A1(n17502), .A2(n17850), .ZN(n17856) );
  NOR2_X1 U20748 ( .A1(n17892), .A2(n18639), .ZN(n17853) );
  OAI22_X1 U20749 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17499), .B1(
        n17498), .B2(n17583), .ZN(n17500) );
  AOI211_X1 U20750 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n17501), .A(
        n17853), .B(n17500), .ZN(n17507) );
  OAI21_X1 U20751 ( .B1(n17502), .B2(n17536), .A(n17535), .ZN(n17515) );
  AOI21_X1 U20752 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17638), .A(
        n17503), .ZN(n17505) );
  XOR2_X1 U20753 ( .A(n17505), .B(n17504), .Z(n17854) );
  AOI22_X1 U20754 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17515), .B1(
        n17639), .B2(n17854), .ZN(n17506) );
  OAI211_X1 U20755 ( .C1(n17536), .C2(n17856), .A(n17507), .B(n17506), .ZN(
        P3_U2812) );
  OAI21_X1 U20756 ( .B1(n17510), .B2(n17849), .A(n17509), .ZN(n17861) );
  NOR2_X1 U20757 ( .A1(n17892), .A2(n18637), .ZN(n17860) );
  AOI221_X1 U20758 ( .B1(n18190), .B2(n17513), .C1(n17512), .C2(n17513), .A(
        n17511), .ZN(n17514) );
  AOI211_X1 U20759 ( .C1(n17639), .C2(n17861), .A(n17860), .B(n17514), .ZN(
        n17518) );
  OAI221_X1 U20760 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17516), .A(n17515), .ZN(
        n17517) );
  OAI211_X1 U20761 ( .C1(n17715), .C2(n17519), .A(n17518), .B(n17517), .ZN(
        P3_U2813) );
  AOI21_X1 U20762 ( .B1(n17638), .B2(n17521), .A(n17520), .ZN(n17522) );
  XOR2_X1 U20763 ( .A(n17522), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Z(
        n17871) );
  NAND2_X1 U20764 ( .A1(n17524), .A2(n17523), .ZN(n17539) );
  INV_X1 U20765 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17525) );
  AOI22_X1 U20766 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17526), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17525), .ZN(n17532) );
  AOI21_X1 U20767 ( .B1(n17705), .B2(n17527), .A(n17630), .ZN(n17552) );
  OAI21_X1 U20768 ( .B1(n17528), .B2(n18592), .A(n17552), .ZN(n17542) );
  AOI22_X1 U20769 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17542), .B1(
        n17530), .B2(n17529), .ZN(n17531) );
  NAND2_X1 U20770 ( .A1(n18061), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n17873) );
  OAI211_X1 U20771 ( .C1(n17539), .C2(n17532), .A(n17531), .B(n17873), .ZN(
        n17533) );
  AOI21_X1 U20772 ( .B1(n17639), .B2(n17871), .A(n17533), .ZN(n17534) );
  OAI221_X1 U20773 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17536), 
        .C1(n17858), .C2(n17535), .A(n17534), .ZN(P3_U2814) );
  NOR2_X1 U20774 ( .A1(n17909), .A2(n17578), .ZN(n17912) );
  AOI21_X1 U20775 ( .B1(n17557), .B2(n17912), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17885) );
  NAND2_X1 U20776 ( .A1(n17537), .A2(n17883), .ZN(n17550) );
  NOR2_X1 U20777 ( .A1(n17892), .A2(n18634), .ZN(n17541) );
  OAI22_X1 U20778 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17539), .B1(
        n17538), .B2(n17583), .ZN(n17540) );
  AOI211_X1 U20779 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17542), .A(
        n17541), .B(n17540), .ZN(n17549) );
  INV_X1 U20780 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17922) );
  NAND2_X1 U20781 ( .A1(n17559), .A2(n17557), .ZN(n17543) );
  OAI21_X1 U20782 ( .B1(n17915), .B2(n17543), .A(n9818), .ZN(n17544) );
  OAI221_X1 U20783 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17898), 
        .C1(n17922), .C2(n17638), .A(n17544), .ZN(n17545) );
  XOR2_X1 U20784 ( .A(n17880), .B(n17545), .Z(n17876) );
  NOR2_X1 U20785 ( .A1(n17800), .A2(n17600), .ZN(n17547) );
  NOR2_X1 U20786 ( .A1(n17908), .A2(n17578), .ZN(n17913) );
  AOI21_X1 U20787 ( .B1(n17557), .B2(n17913), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17887) );
  INV_X1 U20788 ( .A(n17887), .ZN(n17546) );
  AOI22_X1 U20789 ( .A1(n17639), .A2(n17876), .B1(n17547), .B2(n17546), .ZN(
        n17548) );
  OAI211_X1 U20790 ( .C1(n17885), .C2(n17550), .A(n17549), .B(n17548), .ZN(
        P3_U2815) );
  NAND2_X1 U20791 ( .A1(n17557), .A2(n17912), .ZN(n17551) );
  OAI221_X1 U20792 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17912), .A(n17551), .ZN(
        n17905) );
  NAND3_X1 U20793 ( .A1(n18460), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        n17592), .ZN(n17594) );
  AOI221_X1 U20794 ( .B1(n17573), .B2(n17553), .C1(n17594), .C2(n17553), .A(
        n17552), .ZN(n17554) );
  NOR2_X1 U20795 ( .A1(n18044), .A2(n18632), .ZN(n17900) );
  AOI211_X1 U20796 ( .C1(n17555), .C2(n17723), .A(n17554), .B(n17900), .ZN(
        n17564) );
  AOI21_X1 U20797 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n17913), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17556) );
  AOI21_X1 U20798 ( .B1(n17913), .B2(n17557), .A(n17556), .ZN(n17902) );
  NOR2_X1 U20799 ( .A1(n17578), .A2(n17558), .ZN(n17561) );
  NAND2_X1 U20800 ( .A1(n17638), .A2(n17559), .ZN(n17617) );
  INV_X1 U20801 ( .A(n17617), .ZN(n17609) );
  AOI21_X1 U20802 ( .B1(n17561), .B2(n17609), .A(n17560), .ZN(n17562) );
  XOR2_X1 U20803 ( .A(n17898), .B(n17562), .Z(n17901) );
  AOI22_X1 U20804 ( .A1(n17640), .A2(n17902), .B1(n17639), .B2(n17901), .ZN(
        n17563) );
  OAI211_X1 U20805 ( .C1(n17735), .C2(n17905), .A(n17564), .B(n17563), .ZN(
        P3_U2816) );
  OAI22_X1 U20806 ( .A1(n17638), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n17578), .B2(n17566), .ZN(n17567) );
  OAI21_X1 U20807 ( .B1(n17638), .B2(n17565), .A(n17567), .ZN(n17568) );
  XOR2_X1 U20808 ( .A(n17568), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n17920) );
  AOI21_X1 U20809 ( .B1(n17705), .B2(n17571), .A(n17630), .ZN(n17569) );
  OAI21_X1 U20810 ( .B1(n17570), .B2(n18592), .A(n17569), .ZN(n17585) );
  NOR2_X1 U20811 ( .A1(n17572), .A2(n17571), .ZN(n17587) );
  OAI211_X1 U20812 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17587), .B(n17573), .ZN(n17575) );
  NAND2_X1 U20813 ( .A1(n18061), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17574) );
  OAI211_X1 U20814 ( .C1(n17583), .C2(n17576), .A(n17575), .B(n17574), .ZN(
        n17577) );
  AOI21_X1 U20815 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17585), .A(
        n17577), .ZN(n17580) );
  OAI22_X1 U20816 ( .A1(n17913), .A2(n17600), .B1(n17912), .B2(n17735), .ZN(
        n17589) );
  NOR2_X1 U20817 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17578), .ZN(
        n17911) );
  INV_X1 U20818 ( .A(n17598), .ZN(n17624) );
  AOI22_X1 U20819 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17589), .B1(
        n17911), .B2(n17624), .ZN(n17579) );
  OAI211_X1 U20820 ( .C1(n17627), .C2(n17920), .A(n17580), .B(n17579), .ZN(
        P3_U2817) );
  AOI21_X1 U20821 ( .B1(n17609), .B2(n17942), .A(n17565), .ZN(n17581) );
  XOR2_X1 U20822 ( .A(n17581), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n17929) );
  OAI22_X1 U20823 ( .A1(n17892), .A2(n18628), .B1(n17583), .B2(n17582), .ZN(
        n17584) );
  AOI221_X1 U20824 ( .B1(n17587), .B2(n17586), .C1(n17585), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17584), .ZN(n17591) );
  NOR2_X1 U20825 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17915), .ZN(
        n17588) );
  AOI22_X1 U20826 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17589), .B1(
        n17588), .B2(n17624), .ZN(n17590) );
  OAI211_X1 U20827 ( .C1(n17929), .C2(n17627), .A(n17591), .B(n17590), .ZN(
        P3_U2818) );
  NAND2_X1 U20828 ( .A1(n18460), .A2(n17592), .ZN(n17606) );
  OAI21_X1 U20829 ( .B1(n17728), .B2(n20986), .A(n17606), .ZN(n17593) );
  AOI22_X1 U20830 ( .A1(n17595), .A2(n17723), .B1(n17594), .B2(n17593), .ZN(
        n17603) );
  OAI21_X1 U20831 ( .B1(n17938), .B2(n17617), .A(n17596), .ZN(n17597) );
  XOR2_X1 U20832 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17597), .Z(
        n17931) );
  NOR2_X1 U20833 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17938), .ZN(
        n17930) );
  AOI22_X1 U20834 ( .A1(n17639), .A2(n17931), .B1(n17930), .B2(n17624), .ZN(
        n17602) );
  NOR2_X1 U20835 ( .A1(n17599), .A2(n17598), .ZN(n17611) );
  OAI22_X1 U20836 ( .A1(n17935), .A2(n17600), .B1(n17735), .B2(n17933), .ZN(
        n17625) );
  OAI21_X1 U20837 ( .B1(n17611), .B2(n17625), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17601) );
  NAND2_X1 U20838 ( .A1(n18061), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n17946) );
  NAND4_X1 U20839 ( .A1(n17603), .A2(n17602), .A3(n17601), .A4(n17946), .ZN(
        P3_U2819) );
  NOR2_X1 U20840 ( .A1(n18190), .A2(n17631), .ZN(n17650) );
  NAND2_X1 U20841 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17650), .ZN(
        n17632) );
  NOR2_X1 U20842 ( .A1(n17604), .A2(n17632), .ZN(n17620) );
  NAND2_X1 U20843 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17620), .ZN(
        n17619) );
  OAI21_X1 U20844 ( .B1(n17728), .B2(n20951), .A(n17619), .ZN(n17605) );
  AOI22_X1 U20845 ( .A1(n17607), .A2(n17723), .B1(n17606), .B2(n17605), .ZN(
        n17615) );
  AOI21_X1 U20846 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17609), .A(
        n17608), .ZN(n17610) );
  XOR2_X1 U20847 ( .A(n17953), .B(n17610), .Z(n17950) );
  AOI22_X1 U20848 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17625), .B1(
        n17639), .B2(n17950), .ZN(n17614) );
  NAND2_X1 U20849 ( .A1(n18061), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n17613) );
  OAI21_X1 U20850 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n17611), .ZN(n17612) );
  NAND4_X1 U20851 ( .A1(n17615), .A2(n17614), .A3(n17613), .A4(n17612), .ZN(
        P3_U2820) );
  NAND2_X1 U20852 ( .A1(n17617), .A2(n17616), .ZN(n17618) );
  INV_X1 U20853 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17959) );
  XOR2_X1 U20854 ( .A(n17618), .B(n17959), .Z(n17965) );
  INV_X1 U20855 ( .A(n17728), .ZN(n17683) );
  OAI211_X1 U20856 ( .C1(n17620), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17683), .B(n17619), .ZN(n17621) );
  NAND2_X1 U20857 ( .A1(n18061), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n17962) );
  OAI211_X1 U20858 ( .C1(n17715), .C2(n17622), .A(n17621), .B(n17962), .ZN(
        n17623) );
  AOI221_X1 U20859 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17625), .C1(
        n17959), .C2(n17624), .A(n17623), .ZN(n17626) );
  OAI21_X1 U20860 ( .B1(n17965), .B2(n17627), .A(n17626), .ZN(P3_U2821) );
  OAI21_X1 U20861 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17629), .A(
        n17628), .ZN(n17984) );
  AOI21_X1 U20862 ( .B1(n17705), .B2(n17631), .A(n17630), .ZN(n17647) );
  OAI21_X1 U20863 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18190), .A(
        n17647), .ZN(n17635) );
  NOR2_X1 U20864 ( .A1(n18044), .A2(n18621), .ZN(n17974) );
  OAI22_X1 U20865 ( .A1(n17715), .A2(n17633), .B1(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17632), .ZN(n17634) );
  AOI211_X1 U20866 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17635), .A(
        n17974), .B(n17634), .ZN(n17642) );
  INV_X1 U20867 ( .A(n17981), .ZN(n17637) );
  AOI22_X1 U20868 ( .A1(n17638), .A2(n17637), .B1(n17981), .B2(n17636), .ZN(
        n17978) );
  AOI22_X1 U20869 ( .A1(n17640), .A2(n17981), .B1(n17639), .B2(n17978), .ZN(
        n17641) );
  OAI211_X1 U20870 ( .C1(n17735), .C2(n17984), .A(n17642), .B(n17641), .ZN(
        P3_U2822) );
  OAI21_X1 U20871 ( .B1(n17645), .B2(n17644), .A(n17643), .ZN(n17646) );
  XOR2_X1 U20872 ( .A(n17646), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n17993) );
  INV_X1 U20873 ( .A(n17647), .ZN(n17648) );
  NOR2_X1 U20874 ( .A1(n18044), .A2(n18619), .ZN(n17985) );
  AOI221_X1 U20875 ( .B1(n17650), .B2(n17649), .C1(n17648), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n17985), .ZN(n17656) );
  AOI21_X1 U20876 ( .B1(n17988), .B2(n17653), .A(n17652), .ZN(n17989) );
  AOI22_X1 U20877 ( .A1(n9765), .A2(n17989), .B1(n17654), .B2(n17723), .ZN(
        n17655) );
  OAI211_X1 U20878 ( .C1(n17735), .C2(n17993), .A(n17656), .B(n17655), .ZN(
        P3_U2823) );
  NAND2_X1 U20879 ( .A1(n18460), .A2(n17660), .ZN(n17667) );
  AOI21_X1 U20880 ( .B1(n17659), .B2(n17658), .A(n17657), .ZN(n18000) );
  AOI22_X1 U20881 ( .A1(n9765), .A2(n18000), .B1(n18061), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n17666) );
  AOI21_X1 U20882 ( .B1(n17660), .B2(n18460), .A(n17728), .ZN(n17680) );
  OAI21_X1 U20883 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17662), .A(
        n17661), .ZN(n18002) );
  OAI22_X1 U20884 ( .A1(n17715), .A2(n17663), .B1(n17735), .B2(n18002), .ZN(
        n17664) );
  AOI21_X1 U20885 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17680), .A(
        n17664), .ZN(n17665) );
  OAI211_X1 U20886 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n17667), .A(
        n17666), .B(n17665), .ZN(P3_U2824) );
  OAI21_X1 U20887 ( .B1(n17670), .B2(n17669), .A(n17668), .ZN(n18003) );
  NAND2_X1 U20888 ( .A1(n17671), .A2(n17731), .ZN(n17682) );
  OAI21_X1 U20889 ( .B1(n17695), .B2(n17682), .A(n17672), .ZN(n17679) );
  INV_X1 U20890 ( .A(n9765), .ZN(n17734) );
  OAI21_X1 U20891 ( .B1(n17675), .B2(n17674), .A(n17673), .ZN(n17676) );
  XOR2_X1 U20892 ( .A(n17676), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18010) );
  OAI22_X1 U20893 ( .A1(n17715), .A2(n17677), .B1(n17734), .B2(n18010), .ZN(
        n17678) );
  AOI21_X1 U20894 ( .B1(n17680), .B2(n17679), .A(n17678), .ZN(n17681) );
  NAND2_X1 U20895 ( .A1(n18061), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18008) );
  OAI211_X1 U20896 ( .C1(n17735), .C2(n18003), .A(n17681), .B(n18008), .ZN(
        P3_U2825) );
  NAND2_X1 U20897 ( .A1(n17683), .A2(n17682), .ZN(n17701) );
  OAI21_X1 U20898 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n17685), .A(
        n17684), .ZN(n18018) );
  OAI22_X1 U20899 ( .A1(n17735), .A2(n18018), .B1(n18190), .B2(n17686), .ZN(
        n17687) );
  AOI21_X1 U20900 ( .B1(n18061), .B2(P3_REIP_REG_4__SCAN_IN), .A(n17687), .ZN(
        n17694) );
  NOR2_X1 U20901 ( .A1(n17688), .A2(n17699), .ZN(n17691) );
  NOR2_X1 U20902 ( .A1(n17691), .A2(n17690), .ZN(n17689) );
  AOI21_X1 U20903 ( .B1(n17691), .B2(n17690), .A(n17689), .ZN(n18011) );
  AOI22_X1 U20904 ( .A1(n9765), .A2(n18011), .B1(n17692), .B2(n17723), .ZN(
        n17693) );
  OAI211_X1 U20905 ( .C1(n17695), .C2(n17701), .A(n17694), .B(n17693), .ZN(
        P3_U2826) );
  OAI21_X1 U20906 ( .B1(n17698), .B2(n17697), .A(n17696), .ZN(n18027) );
  AOI21_X1 U20907 ( .B1(n18019), .B2(n17700), .A(n17699), .ZN(n18024) );
  INV_X1 U20908 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18611) );
  NOR2_X1 U20909 ( .A1(n17892), .A2(n18611), .ZN(n18023) );
  OAI22_X1 U20910 ( .A1(n17715), .A2(n17702), .B1(n17704), .B2(n17701), .ZN(
        n17703) );
  AOI211_X1 U20911 ( .C1(n9765), .C2(n18024), .A(n18023), .B(n17703), .ZN(
        n17707) );
  NAND4_X1 U20912 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17705), .A3(
        n17731), .A4(n17704), .ZN(n17706) );
  OAI211_X1 U20913 ( .C1(n17735), .C2(n18027), .A(n17707), .B(n17706), .ZN(
        P3_U2827) );
  AOI21_X1 U20914 ( .B1(n17710), .B2(n17709), .A(n17708), .ZN(n18040) );
  NOR2_X1 U20915 ( .A1(n18044), .A2(n18609), .ZN(n18039) );
  OAI21_X1 U20916 ( .B1(n17713), .B2(n17712), .A(n17711), .ZN(n18035) );
  OAI22_X1 U20917 ( .A1(n17715), .A2(n17714), .B1(n17735), .B2(n18035), .ZN(
        n17716) );
  AOI211_X1 U20918 ( .C1(n9765), .C2(n18040), .A(n18039), .B(n17716), .ZN(
        n17717) );
  OAI221_X1 U20919 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18190), .C1(
        n17718), .C2(n17731), .A(n17717), .ZN(P3_U2828) );
  NOR2_X1 U20920 ( .A1(n17730), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17719) );
  XOR2_X1 U20921 ( .A(n17719), .B(n17722), .Z(n18056) );
  OAI22_X1 U20922 ( .A1(n17735), .A2(n18056), .B1(n17892), .B2(n18711), .ZN(
        n17720) );
  INV_X1 U20923 ( .A(n17720), .ZN(n17726) );
  AOI21_X1 U20924 ( .B1(n17729), .B2(n17722), .A(n17721), .ZN(n18049) );
  AOI22_X1 U20925 ( .A1(n9765), .A2(n18049), .B1(n17727), .B2(n17723), .ZN(
        n17725) );
  OAI211_X1 U20926 ( .C1(n17728), .C2(n17727), .A(n17726), .B(n17725), .ZN(
        P3_U2829) );
  OAI21_X1 U20927 ( .B1(n17730), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17729), .ZN(n18064) );
  INV_X1 U20928 ( .A(n18064), .ZN(n17736) );
  NAND3_X1 U20929 ( .A1(n18689), .A2(n18592), .A3(n17731), .ZN(n17732) );
  AOI22_X1 U20930 ( .A1(n18061), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17732), .ZN(n17733) );
  OAI221_X1 U20931 ( .B1(n17736), .B2(n17735), .C1(n18064), .C2(n17734), .A(
        n17733), .ZN(P3_U2830) );
  NOR2_X1 U20932 ( .A1(n17806), .A2(n17759), .ZN(n17791) );
  NAND2_X1 U20933 ( .A1(n17737), .A2(n17791), .ZN(n17752) );
  AOI221_X1 U20934 ( .B1(n17751), .B2(n9918), .C1(n17752), .C2(n9918), .A(
        n18050), .ZN(n17747) );
  NOR2_X1 U20935 ( .A1(n17941), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17967) );
  INV_X1 U20936 ( .A(n17967), .ZN(n18029) );
  NAND2_X1 U20937 ( .A1(n18549), .A2(n17941), .ZN(n17969) );
  INV_X1 U20938 ( .A(n17969), .ZN(n18031) );
  AOI21_X1 U20939 ( .B1(n17738), .B2(n18029), .A(n18031), .ZN(n17778) );
  AOI22_X1 U20940 ( .A1(n18547), .A2(n17739), .B1(n17760), .B2(n17969), .ZN(
        n17740) );
  OAI21_X1 U20941 ( .B1(n18549), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17740), .ZN(n17744) );
  OAI22_X1 U20942 ( .A1(n17742), .A2(n17934), .B1(n17741), .B2(n18037), .ZN(
        n17743) );
  NOR4_X1 U20943 ( .A1(n17745), .A2(n17778), .A3(n17744), .A4(n17743), .ZN(
        n17753) );
  OAI211_X1 U20944 ( .C1(n18549), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17753), .ZN(n17746) );
  AOI22_X1 U20945 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18052), .B1(
        n17747), .B2(n17746), .ZN(n17749) );
  NAND2_X1 U20946 ( .A1(n18061), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17748) );
  OAI211_X1 U20947 ( .C1(n17750), .C2(n17964), .A(n17749), .B(n17748), .ZN(
        P3_U2835) );
  AOI221_X1 U20948 ( .B1(n17753), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), 
        .C1(n17752), .C2(n17751), .A(n18050), .ZN(n17754) );
  AOI21_X1 U20949 ( .B1(n18052), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17754), .ZN(n17756) );
  OAI211_X1 U20950 ( .C1(n17757), .C2(n17964), .A(n17756), .B(n17755), .ZN(
        P3_U2836) );
  AOI21_X1 U20951 ( .B1(n17758), .B2(n17848), .A(n17866), .ZN(n17783) );
  AOI211_X1 U20952 ( .C1(n17973), .C2(n17760), .A(n17783), .B(n17778), .ZN(
        n17765) );
  NOR2_X1 U20953 ( .A1(n17760), .A2(n17759), .ZN(n17762) );
  NAND2_X1 U20954 ( .A1(n17762), .A2(n17761), .ZN(n17764) );
  AOI221_X1 U20955 ( .B1(n17765), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n17764), .C2(n17763), .A(n18050), .ZN(n17766) );
  AOI211_X1 U20956 ( .C1(n18052), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17767), .B(n17766), .ZN(n17771) );
  AOI22_X1 U20957 ( .A1(n17980), .A2(n17769), .B1(n17979), .B2(n17768), .ZN(
        n17770) );
  OAI211_X1 U20958 ( .C1(n18055), .C2(n17772), .A(n17771), .B(n17770), .ZN(
        P3_U2837) );
  INV_X1 U20959 ( .A(n17773), .ZN(n17812) );
  INV_X1 U20960 ( .A(n17774), .ZN(n17776) );
  AOI21_X1 U20961 ( .B1(n17979), .B2(n17776), .A(n17775), .ZN(n17787) );
  NAND2_X1 U20962 ( .A1(n17800), .A2(n17777), .ZN(n17779) );
  AOI211_X1 U20963 ( .C1(n17882), .C2(n17779), .A(n17778), .B(n18052), .ZN(
        n17780) );
  OAI21_X1 U20964 ( .B1(n17781), .B2(n18037), .A(n17780), .ZN(n17785) );
  NOR3_X1 U20965 ( .A1(n17783), .A2(n17782), .A3(n17785), .ZN(n17784) );
  NOR2_X1 U20966 ( .A1(n18061), .A2(n17784), .ZN(n17790) );
  OAI211_X1 U20967 ( .C1(n17973), .C2(n17785), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17790), .ZN(n17786) );
  OAI211_X1 U20968 ( .C1(n17788), .C2(n17812), .A(n17787), .B(n17786), .ZN(
        P3_U2838) );
  INV_X1 U20969 ( .A(n17789), .ZN(n17794) );
  OAI221_X1 U20970 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17791), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n18042), .A(n17790), .ZN(
        n17792) );
  OAI211_X1 U20971 ( .C1(n17794), .C2(n17964), .A(n17793), .B(n17792), .ZN(
        P3_U2839) );
  NAND2_X1 U20972 ( .A1(n18037), .A2(n17934), .ZN(n17937) );
  OAI21_X1 U20973 ( .B1(n17795), .B2(n17813), .A(n18545), .ZN(n17796) );
  INV_X1 U20974 ( .A(n17796), .ZN(n17797) );
  AOI221_X1 U20975 ( .B1(n17844), .B2(n18534), .C1(n17825), .C2(n18534), .A(
        n17797), .ZN(n17827) );
  OAI21_X1 U20976 ( .B1(n18549), .B2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n17827), .ZN(n17798) );
  AOI21_X1 U20977 ( .B1(n17805), .B2(n17937), .A(n17798), .ZN(n17818) );
  OAI22_X1 U20978 ( .A1(n17800), .A2(n17934), .B1(n17799), .B2(n18037), .ZN(
        n17816) );
  INV_X1 U20979 ( .A(n17948), .ZN(n17943) );
  OAI22_X1 U20980 ( .A1(n17943), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n17819), .B2(n17866), .ZN(n17801) );
  NOR4_X1 U20981 ( .A1(n17804), .A2(n17802), .A3(n17816), .A4(n17801), .ZN(
        n17803) );
  AOI21_X1 U20982 ( .B1(n17818), .B2(n17803), .A(n18050), .ZN(n17808) );
  OAI21_X1 U20983 ( .B1(n17806), .B2(n17805), .A(n17804), .ZN(n17807) );
  AOI22_X1 U20984 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18052), .B1(
        n17808), .B2(n17807), .ZN(n17810) );
  OAI211_X1 U20985 ( .C1(n17811), .C2(n17964), .A(n17810), .B(n17809), .ZN(
        P3_U2840) );
  NOR2_X1 U20986 ( .A1(n17813), .A2(n17812), .ZN(n17838) );
  AOI22_X1 U20987 ( .A1(n17979), .A2(n17815), .B1(n17814), .B2(n17838), .ZN(
        n17823) );
  NOR2_X1 U20988 ( .A1(n18050), .A2(n17816), .ZN(n17870) );
  NAND2_X1 U20989 ( .A1(n17870), .A2(n17817), .ZN(n17824) );
  NOR2_X1 U20990 ( .A1(n18545), .A2(n18547), .ZN(n18051) );
  OAI21_X1 U20991 ( .B1(n17819), .B2(n18051), .A(n17818), .ZN(n17820) );
  OAI211_X1 U20992 ( .C1(n17824), .C2(n17820), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17892), .ZN(n17821) );
  NAND3_X1 U20993 ( .A1(n17823), .A2(n17822), .A3(n17821), .ZN(P3_U2841) );
  NOR3_X1 U20994 ( .A1(n18051), .A2(n18729), .A3(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17828) );
  AOI21_X1 U20995 ( .B1(n17825), .B2(n17937), .A(n17824), .ZN(n17826) );
  AOI21_X1 U20996 ( .B1(n17827), .B2(n17826), .A(n18061), .ZN(n17839) );
  NOR2_X1 U20997 ( .A1(n17828), .A2(n17839), .ZN(n17834) );
  AOI22_X1 U20998 ( .A1(n17979), .A2(n17830), .B1(n17838), .B2(n17829), .ZN(
        n17832) );
  OAI211_X1 U20999 ( .C1(n17834), .C2(n17833), .A(n17832), .B(n17831), .ZN(
        P3_U2842) );
  INV_X1 U21000 ( .A(n17835), .ZN(n17841) );
  AOI221_X1 U21001 ( .B1(n17839), .B2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), 
        .C1(n17838), .C2(n17837), .A(n17836), .ZN(n17840) );
  OAI21_X1 U21002 ( .B1(n17841), .B2(n17964), .A(n17840), .ZN(P3_U2843) );
  OAI22_X1 U21003 ( .A1(n17966), .A2(n17866), .B1(n18028), .B2(n17968), .ZN(
        n17906) );
  INV_X1 U21004 ( .A(n17906), .ZN(n18020) );
  NOR2_X1 U21005 ( .A1(n18020), .A2(n17910), .ZN(n17877) );
  OAI211_X1 U21006 ( .C1(n17843), .C2(n17877), .A(n17842), .B(n18057), .ZN(
        n17875) );
  OR3_X1 U21007 ( .A1(n17844), .A2(n17858), .A3(n17967), .ZN(n17845) );
  AOI22_X1 U21008 ( .A1(n17846), .A2(n17937), .B1(n17969), .B2(n17845), .ZN(
        n17847) );
  OAI211_X1 U21009 ( .C1(n17848), .C2(n17866), .A(n17870), .B(n17847), .ZN(
        n17857) );
  AOI21_X1 U21010 ( .B1(n17849), .B2(n17969), .A(n17857), .ZN(n17851) );
  NOR3_X1 U21011 ( .A1(n18061), .A2(n17851), .A3(n17850), .ZN(n17852) );
  AOI211_X1 U21012 ( .C1(n17854), .C2(n17979), .A(n17853), .B(n17852), .ZN(
        n17855) );
  OAI21_X1 U21013 ( .B1(n17856), .B2(n17875), .A(n17855), .ZN(P3_U2844) );
  NAND3_X1 U21014 ( .A1(n17892), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n17857), .ZN(n17863) );
  NOR3_X1 U21015 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17858), .A3(
        n17875), .ZN(n17859) );
  AOI211_X1 U21016 ( .C1(n17979), .C2(n17861), .A(n17860), .B(n17859), .ZN(
        n17862) );
  NAND2_X1 U21017 ( .A1(n17863), .A2(n17862), .ZN(P3_U2845) );
  OAI21_X1 U21018 ( .B1(n17880), .B2(n18547), .A(n17864), .ZN(n17865) );
  INV_X1 U21019 ( .A(n17865), .ZN(n17869) );
  OAI22_X1 U21020 ( .A1(n18549), .A2(n17868), .B1(n17867), .B2(n17866), .ZN(
        n17955) );
  AOI211_X1 U21021 ( .C1(n17948), .C2(n17895), .A(n17869), .B(n17955), .ZN(
        n17879) );
  AOI221_X1 U21022 ( .B1(n17971), .B2(n17870), .C1(n17879), .C2(n17870), .A(
        n18061), .ZN(n17872) );
  AOI22_X1 U21023 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17872), .B1(
        n17979), .B2(n17871), .ZN(n17874) );
  OAI211_X1 U21024 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n17875), .A(
        n17874), .B(n17873), .ZN(P3_U2846) );
  AOI22_X1 U21025 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18052), .B1(
        n17979), .B2(n17876), .ZN(n17891) );
  NAND3_X1 U21026 ( .A1(n17893), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n17877), .ZN(n17897) );
  AOI211_X1 U21027 ( .C1(n17880), .C2(n17897), .A(n17879), .B(n17878), .ZN(
        n17889) );
  NAND2_X1 U21028 ( .A1(n17882), .A2(n17881), .ZN(n17886) );
  NAND2_X1 U21029 ( .A1(n18515), .A2(n17883), .ZN(n17884) );
  OAI22_X1 U21030 ( .A1(n17887), .A2(n17886), .B1(n17885), .B2(n17884), .ZN(
        n17888) );
  OAI21_X1 U21031 ( .B1(n17889), .B2(n17888), .A(n18057), .ZN(n17890) );
  OAI211_X1 U21032 ( .C1(n18634), .C2(n17892), .A(n17891), .B(n17890), .ZN(
        P3_U2847) );
  INV_X1 U21033 ( .A(n17955), .ZN(n17940) );
  NAND2_X1 U21034 ( .A1(n17893), .A2(n17932), .ZN(n17921) );
  NAND2_X1 U21035 ( .A1(n18547), .A2(n17921), .ZN(n17916) );
  OAI211_X1 U21036 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18051), .A(
        n17940), .B(n17916), .ZN(n17894) );
  AOI211_X1 U21037 ( .C1(n17895), .C2(n17948), .A(n17894), .B(n17898), .ZN(
        n17896) );
  AOI211_X1 U21038 ( .C1(n17898), .C2(n17897), .A(n17896), .B(n18050), .ZN(
        n17899) );
  AOI211_X1 U21039 ( .C1(n18052), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17900), .B(n17899), .ZN(n17904) );
  AOI22_X1 U21040 ( .A1(n17980), .A2(n17902), .B1(n17979), .B2(n17901), .ZN(
        n17903) );
  OAI211_X1 U21041 ( .C1(n18055), .C2(n17905), .A(n17904), .B(n17903), .ZN(
        P3_U2848) );
  NAND2_X1 U21042 ( .A1(n18057), .A2(n17906), .ZN(n18012) );
  OAI222_X1 U21043 ( .A1(n18012), .A2(n17910), .B1(n18055), .B2(n17909), .C1(
        n17908), .C2(n17907), .ZN(n17960) );
  AOI22_X1 U21044 ( .A1(n18061), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n17911), 
        .B2(n17960), .ZN(n17919) );
  OAI22_X1 U21045 ( .A1(n17913), .A2(n17934), .B1(n17912), .B2(n18037), .ZN(
        n17914) );
  AOI211_X1 U21046 ( .C1(n17948), .C2(n17915), .A(n17955), .B(n17914), .ZN(
        n17925) );
  OAI211_X1 U21047 ( .C1(n17943), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17925), .B(n17916), .ZN(n17917) );
  OAI211_X1 U21048 ( .C1(n18050), .C2(n17917), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17892), .ZN(n17918) );
  OAI211_X1 U21049 ( .C1(n17920), .C2(n17964), .A(n17919), .B(n17918), .ZN(
        P3_U2849) );
  NOR2_X1 U21050 ( .A1(n18044), .A2(n18628), .ZN(n17927) );
  OAI21_X1 U21051 ( .B1(n17922), .B2(n18547), .A(n17921), .ZN(n17924) );
  AOI22_X1 U21052 ( .A1(n17942), .A2(n17960), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18057), .ZN(n17923) );
  AOI21_X1 U21053 ( .B1(n17925), .B2(n17924), .A(n17923), .ZN(n17926) );
  AOI211_X1 U21054 ( .C1(n18052), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17927), .B(n17926), .ZN(n17928) );
  OAI21_X1 U21055 ( .B1(n17929), .B2(n17964), .A(n17928), .ZN(P3_U2850) );
  AOI22_X1 U21056 ( .A1(n17979), .A2(n17931), .B1(n17930), .B2(n17960), .ZN(
        n17947) );
  AOI21_X1 U21057 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17932), .A(
        n17941), .ZN(n17936) );
  OAI22_X1 U21058 ( .A1(n17935), .A2(n17934), .B1(n18037), .B2(n17933), .ZN(
        n17956) );
  AOI211_X1 U21059 ( .C1(n17938), .C2(n17937), .A(n17936), .B(n17956), .ZN(
        n17939) );
  NAND3_X1 U21060 ( .A1(n18057), .A2(n17940), .A3(n17939), .ZN(n17949) );
  OAI22_X1 U21061 ( .A1(n17943), .A2(n17942), .B1(n17941), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17944) );
  OAI211_X1 U21062 ( .C1(n17949), .C2(n17944), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17892), .ZN(n17945) );
  NAND3_X1 U21063 ( .A1(n17947), .A2(n17946), .A3(n17945), .ZN(P3_U2851) );
  NAND2_X1 U21064 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17960), .ZN(
        n17954) );
  OAI221_X1 U21065 ( .B1(n17949), .B2(n17948), .C1(n17949), .C2(n17959), .A(
        n18044), .ZN(n17952) );
  AOI22_X1 U21066 ( .A1(n18061), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17979), 
        .B2(n17950), .ZN(n17951) );
  OAI221_X1 U21067 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17954), 
        .C1(n17953), .C2(n17952), .A(n17951), .ZN(P3_U2852) );
  AOI211_X1 U21068 ( .C1(n17957), .C2(n18547), .A(n17956), .B(n17955), .ZN(
        n17958) );
  AOI21_X1 U21069 ( .B1(n18057), .B2(n17958), .A(n18061), .ZN(n17961) );
  AOI22_X1 U21070 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17961), .B1(
        n17960), .B2(n17959), .ZN(n17963) );
  OAI211_X1 U21071 ( .C1(n17965), .C2(n17964), .A(n17963), .B(n17962), .ZN(
        P3_U2853) );
  NOR2_X1 U21072 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18012), .ZN(
        n17976) );
  AND2_X1 U21073 ( .A1(n18545), .A2(n17966), .ZN(n18032) );
  AOI211_X1 U21074 ( .C1(n17969), .C2(n17968), .A(n17967), .B(n18032), .ZN(
        n18021) );
  OAI21_X1 U21075 ( .B1(n17971), .B2(n17970), .A(n18021), .ZN(n17995) );
  AOI211_X1 U21076 ( .C1(n17973), .C2(n17972), .A(n17988), .B(n17995), .ZN(
        n17986) );
  AOI221_X1 U21077 ( .B1(n17986), .B2(n18042), .C1(n18045), .C2(n18042), .A(
        n9929), .ZN(n17975) );
  AOI211_X1 U21078 ( .C1(n17977), .C2(n17976), .A(n17975), .B(n17974), .ZN(
        n17983) );
  AOI22_X1 U21079 ( .A1(n17981), .A2(n17980), .B1(n17979), .B2(n17978), .ZN(
        n17982) );
  OAI211_X1 U21080 ( .C1(n18055), .C2(n17984), .A(n17983), .B(n17982), .ZN(
        P3_U2854) );
  AOI21_X1 U21081 ( .B1(n18052), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17985), .ZN(n17992) );
  AOI221_X1 U21082 ( .B1(n18020), .B2(n17988), .C1(n17987), .C2(n17988), .A(
        n17986), .ZN(n17990) );
  AOI22_X1 U21083 ( .A1(n18057), .A2(n17990), .B1(n18048), .B2(n17989), .ZN(
        n17991) );
  OAI211_X1 U21084 ( .C1(n18055), .C2(n17993), .A(n17992), .B(n17991), .ZN(
        P3_U2855) );
  NOR2_X1 U21085 ( .A1(n17892), .A2(n18617), .ZN(n17999) );
  NOR2_X1 U21086 ( .A1(n17994), .A2(n18012), .ZN(n17997) );
  AOI21_X1 U21087 ( .B1(n18057), .B2(n17995), .A(n18052), .ZN(n18005) );
  INV_X1 U21088 ( .A(n18005), .ZN(n17996) );
  MUX2_X1 U21089 ( .A(n17997), .B(n17996), .S(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n17998) );
  AOI211_X1 U21090 ( .C1(n18048), .C2(n18000), .A(n17999), .B(n17998), .ZN(
        n18001) );
  OAI21_X1 U21091 ( .B1(n18055), .B2(n18002), .A(n18001), .ZN(P3_U2856) );
  INV_X1 U21092 ( .A(n18048), .ZN(n18065) );
  NOR4_X1 U21093 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18019), .A3(
        n18013), .A4(n18012), .ZN(n18007) );
  INV_X1 U21094 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18004) );
  OAI22_X1 U21095 ( .A1(n18005), .A2(n18004), .B1(n18055), .B2(n18003), .ZN(
        n18006) );
  NOR2_X1 U21096 ( .A1(n18007), .A2(n18006), .ZN(n18009) );
  OAI211_X1 U21097 ( .C1(n18010), .C2(n18065), .A(n18009), .B(n18008), .ZN(
        P3_U2857) );
  AOI22_X1 U21098 ( .A1(n18061), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18048), 
        .B2(n18011), .ZN(n18017) );
  OAI221_X1 U21099 ( .B1(n18045), .B2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C1(
        n18045), .C2(n18021), .A(n18042), .ZN(n18015) );
  NOR2_X1 U21100 ( .A1(n18019), .A2(n18012), .ZN(n18014) );
  AOI22_X1 U21101 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18015), .B1(
        n18014), .B2(n18013), .ZN(n18016) );
  OAI211_X1 U21102 ( .C1(n18055), .C2(n18018), .A(n18017), .B(n18016), .ZN(
        P3_U2858) );
  AOI221_X1 U21103 ( .B1(n18021), .B2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C1(
        n18020), .C2(n18019), .A(n18050), .ZN(n18022) );
  AOI211_X1 U21104 ( .C1(n18048), .C2(n18024), .A(n18023), .B(n18022), .ZN(
        n18026) );
  NAND2_X1 U21105 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18052), .ZN(
        n18025) );
  OAI211_X1 U21106 ( .C1(n18027), .C2(n18055), .A(n18026), .B(n18025), .ZN(
        P3_U2859) );
  NOR2_X1 U21107 ( .A1(n18687), .A2(n18028), .ZN(n18034) );
  NAND3_X1 U21108 ( .A1(n18545), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18030) );
  OAI211_X1 U21109 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n18031), .A(
        n18030), .B(n18029), .ZN(n18033) );
  AOI221_X1 U21110 ( .B1(n18034), .B2(n18043), .C1(n18033), .C2(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n18032), .ZN(n18036) );
  AOI221_X1 U21111 ( .B1(n18037), .B2(n18036), .C1(n18035), .C2(n18036), .A(
        n18050), .ZN(n18038) );
  AOI211_X1 U21112 ( .C1(n18048), .C2(n18040), .A(n18039), .B(n18038), .ZN(
        n18041) );
  OAI21_X1 U21113 ( .B1(n18043), .B2(n18042), .A(n18041), .ZN(P3_U2860) );
  NOR2_X1 U21114 ( .A1(n18044), .A2(n18711), .ZN(n18047) );
  AOI211_X1 U21115 ( .C1(n18549), .C2(n21029), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18045), .ZN(n18046) );
  AOI211_X1 U21116 ( .C1(n18049), .C2(n18048), .A(n18047), .B(n18046), .ZN(
        n18054) );
  NOR3_X1 U21117 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18051), .A3(
        n18050), .ZN(n18059) );
  OAI21_X1 U21118 ( .B1(n18052), .B2(n18059), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18053) );
  OAI211_X1 U21119 ( .C1(n18056), .C2(n18055), .A(n18054), .B(n18053), .ZN(
        P3_U2861) );
  AOI211_X1 U21120 ( .C1(n18549), .C2(n18057), .A(n18061), .B(n21029), .ZN(
        n18058) );
  AOI211_X1 U21121 ( .C1(n18060), .C2(n18064), .A(n18059), .B(n18058), .ZN(
        n18063) );
  NAND2_X1 U21122 ( .A1(n18061), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18062) );
  OAI211_X1 U21123 ( .C1(n18065), .C2(n18064), .A(n18063), .B(n18062), .ZN(
        P3_U2862) );
  INV_X1 U21124 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18553) );
  AOI21_X1 U21125 ( .B1(n18068), .B2(n18067), .A(n18066), .ZN(n18574) );
  OAI21_X1 U21126 ( .B1(n18574), .B2(n18126), .A(n18078), .ZN(n18069) );
  OAI221_X1 U21127 ( .B1(n18553), .B2(n18725), .C1(n18553), .C2(n18078), .A(
        n18069), .ZN(P3_U2863) );
  NAND2_X1 U21128 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18235) );
  AOI221_X1 U21129 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18235), .C1(n18071), 
        .C2(n18235), .A(n18070), .ZN(n18077) );
  NOR2_X1 U21130 ( .A1(n18072), .A2(n18555), .ZN(n18074) );
  OAI21_X1 U21131 ( .B1(n18074), .B2(n18073), .A(n18078), .ZN(n18075) );
  AOI22_X1 U21132 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18077), .B1(
        n18075), .B2(n18560), .ZN(P3_U2865) );
  INV_X1 U21133 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18563) );
  NAND2_X1 U21134 ( .A1(n18560), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18325) );
  INV_X1 U21135 ( .A(n18325), .ZN(n18303) );
  NOR2_X1 U21136 ( .A1(n18560), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18258) );
  NOR2_X1 U21137 ( .A1(n18303), .A2(n18258), .ZN(n18076) );
  OAI22_X1 U21138 ( .A1(n18077), .A2(n18563), .B1(n18076), .B2(n18075), .ZN(
        P3_U2866) );
  NOR2_X1 U21139 ( .A1(n18564), .A2(n18078), .ZN(P3_U2867) );
  NAND2_X1 U21140 ( .A1(n18555), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18305) );
  NAND2_X1 U21141 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18395) );
  NOR2_X2 U21142 ( .A1(n18305), .A2(n18395), .ZN(n18507) );
  INV_X1 U21143 ( .A(n18507), .ZN(n18503) );
  NOR2_X1 U21144 ( .A1(n18563), .A2(n18235), .ZN(n18458) );
  NAND2_X1 U21145 ( .A1(n18553), .A2(n18458), .ZN(n18454) );
  NAND2_X1 U21146 ( .A1(n18503), .A2(n18454), .ZN(n18420) );
  NAND2_X1 U21147 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18458), .ZN(
        n18513) );
  INV_X1 U21148 ( .A(n18513), .ZN(n18499) );
  NOR2_X1 U21149 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18281) );
  INV_X1 U21150 ( .A(n18281), .ZN(n18556) );
  NAND2_X1 U21151 ( .A1(n18560), .A2(n18563), .ZN(n18147) );
  NOR2_X2 U21152 ( .A1(n18556), .A2(n18147), .ZN(n18185) );
  NOR2_X1 U21153 ( .A1(n18499), .A2(n18185), .ZN(n18148) );
  AOI211_X1 U21154 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18189), .B(n18148), .ZN(
        n18079) );
  AOI21_X1 U21155 ( .B1(n18420), .B2(n18460), .A(n18079), .ZN(n18123) );
  INV_X1 U21156 ( .A(n18123), .ZN(n18118) );
  NOR2_X1 U21157 ( .A1(n18080), .A2(n18190), .ZN(n18349) );
  NOR2_X2 U21158 ( .A1(n18189), .A2(n18081), .ZN(n18455) );
  NOR2_X1 U21159 ( .A1(n18421), .A2(n18148), .ZN(n18122) );
  AOI22_X1 U21160 ( .A1(n18349), .A2(n18507), .B1(n18455), .B2(n18122), .ZN(
        n18086) );
  NOR2_X1 U21161 ( .A1(n18083), .A2(n18082), .ZN(n18120) );
  INV_X1 U21162 ( .A(n18120), .ZN(n18114) );
  NOR2_X2 U21163 ( .A1(n18084), .A2(n18114), .ZN(n18461) );
  NAND2_X1 U21164 ( .A1(n18460), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18354) );
  INV_X1 U21165 ( .A(n18354), .ZN(n18456) );
  INV_X1 U21166 ( .A(n18454), .ZN(n18444) );
  AOI22_X1 U21167 ( .A1(n18461), .A2(n18185), .B1(n18456), .B2(n18444), .ZN(
        n18085) );
  OAI211_X1 U21168 ( .C1(n18087), .C2(n18118), .A(n18086), .B(n18085), .ZN(
        P3_U2868) );
  INV_X1 U21169 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20830) );
  INV_X1 U21170 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n18088) );
  NOR2_X2 U21171 ( .A1(n18190), .A2(n18088), .ZN(n18466) );
  NOR2_X2 U21172 ( .A1(n18189), .A2(n18089), .ZN(n18465) );
  AOI22_X1 U21173 ( .A1(n18466), .A2(n18444), .B1(n18465), .B2(n18122), .ZN(
        n18092) );
  NOR2_X1 U21174 ( .A1(n18114), .A2(n18090), .ZN(n18129) );
  AND2_X1 U21175 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18460), .ZN(n18467) );
  AOI22_X1 U21176 ( .A1(n18129), .A2(n18185), .B1(n18467), .B2(n18507), .ZN(
        n18091) );
  OAI211_X1 U21177 ( .C1(n20830), .C2(n18118), .A(n18092), .B(n18091), .ZN(
        P3_U2869) );
  NOR2_X2 U21178 ( .A1(n18190), .A2(n14000), .ZN(n18472) );
  NOR2_X2 U21179 ( .A1(n18189), .A2(n18093), .ZN(n18471) );
  AOI22_X1 U21180 ( .A1(n18472), .A2(n18444), .B1(n18471), .B2(n18122), .ZN(
        n18096) );
  NOR2_X1 U21181 ( .A1(n18114), .A2(n18094), .ZN(n18132) );
  AND2_X1 U21182 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18460), .ZN(n18473) );
  AOI22_X1 U21183 ( .A1(n18132), .A2(n18185), .B1(n18473), .B2(n18507), .ZN(
        n18095) );
  OAI211_X1 U21184 ( .C1(n18097), .C2(n18118), .A(n18096), .B(n18095), .ZN(
        P3_U2870) );
  INV_X1 U21185 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n21026) );
  NOR2_X1 U21186 ( .A1(n21026), .A2(n18190), .ZN(n18478) );
  NOR2_X2 U21187 ( .A1(n18189), .A2(n18098), .ZN(n18477) );
  AOI22_X1 U21188 ( .A1(n18478), .A2(n18507), .B1(n18477), .B2(n18122), .ZN(
        n18101) );
  NOR2_X2 U21189 ( .A1(n18099), .A2(n18114), .ZN(n18479) );
  NAND2_X1 U21190 ( .A1(n18460), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18482) );
  INV_X1 U21191 ( .A(n18482), .ZN(n18433) );
  AOI22_X1 U21192 ( .A1(n18479), .A2(n18185), .B1(n18433), .B2(n18444), .ZN(
        n18100) );
  OAI211_X1 U21193 ( .C1(n18102), .C2(n18118), .A(n18101), .B(n18100), .ZN(
        P3_U2871) );
  NOR2_X2 U21194 ( .A1(n18189), .A2(n18103), .ZN(n18484) );
  NAND2_X1 U21195 ( .A1(n18460), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18410) );
  INV_X1 U21196 ( .A(n18410), .ZN(n18483) );
  AOI22_X1 U21197 ( .A1(n18484), .A2(n18122), .B1(n18483), .B2(n18444), .ZN(
        n18106) );
  NOR2_X1 U21198 ( .A1(n19105), .A2(n18190), .ZN(n18407) );
  NOR2_X2 U21199 ( .A1(n18104), .A2(n18114), .ZN(n18485) );
  AOI22_X1 U21200 ( .A1(n18407), .A2(n18507), .B1(n18485), .B2(n18185), .ZN(
        n18105) );
  OAI211_X1 U21201 ( .C1(n18107), .C2(n18118), .A(n18106), .B(n18105), .ZN(
        P3_U2872) );
  NOR2_X1 U21202 ( .A1(n19110), .A2(n18190), .ZN(n18491) );
  NOR2_X2 U21203 ( .A1(n18189), .A2(n18108), .ZN(n18490) );
  AOI22_X1 U21204 ( .A1(n9703), .A2(n18507), .B1(n18490), .B2(n18122), .ZN(
        n18111) );
  NOR2_X2 U21205 ( .A1(n18109), .A2(n18114), .ZN(n18493) );
  NAND2_X1 U21206 ( .A1(n18460), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18496) );
  INV_X1 U21207 ( .A(n18496), .ZN(n18439) );
  AOI22_X1 U21208 ( .A1(n18493), .A2(n18185), .B1(n18439), .B2(n18444), .ZN(
        n18110) );
  OAI211_X1 U21209 ( .C1(n18112), .C2(n18118), .A(n18111), .B(n18110), .ZN(
        P3_U2873) );
  NOR2_X2 U21210 ( .A1(n18189), .A2(n18113), .ZN(n18497) );
  NAND2_X1 U21211 ( .A1(n18460), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18504) );
  INV_X1 U21212 ( .A(n18504), .ZN(n18443) );
  AOI22_X1 U21213 ( .A1(n18497), .A2(n18122), .B1(n18443), .B2(n18444), .ZN(
        n18117) );
  INV_X1 U21214 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n21048) );
  NOR2_X1 U21215 ( .A1(n21048), .A2(n18190), .ZN(n18498) );
  NOR2_X2 U21216 ( .A1(n18115), .A2(n18114), .ZN(n18500) );
  AOI22_X1 U21217 ( .A1(n18498), .A2(n18507), .B1(n18500), .B2(n18185), .ZN(
        n18116) );
  OAI211_X1 U21218 ( .C1(n20853), .C2(n18118), .A(n18117), .B(n18116), .ZN(
        P3_U2874) );
  NAND2_X1 U21219 ( .A1(n18120), .A2(n18119), .ZN(n18514) );
  INV_X1 U21220 ( .A(n18185), .ZN(n18183) );
  INV_X1 U21221 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n18121) );
  NOR2_X2 U21222 ( .A1(n18190), .A2(n18121), .ZN(n18508) );
  AND2_X1 U21223 ( .A1(n18426), .A2(BUF2_REG_7__SCAN_IN), .ZN(n18506) );
  AOI22_X1 U21224 ( .A1(n18508), .A2(n18444), .B1(n18506), .B2(n18122), .ZN(
        n18125) );
  NOR2_X2 U21225 ( .A1(n18190), .A2(n19122), .ZN(n18509) );
  AOI22_X1 U21226 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18123), .B1(
        n18509), .B2(n18507), .ZN(n18124) );
  OAI211_X1 U21227 ( .C1(n18514), .C2(n18183), .A(n18125), .B(n18124), .ZN(
        P3_U2875) );
  INV_X1 U21228 ( .A(n18349), .ZN(n18464) );
  NAND2_X1 U21229 ( .A1(n18555), .A2(n18582), .ZN(n18394) );
  NOR2_X1 U21230 ( .A1(n18147), .A2(n18394), .ZN(n18143) );
  AOI22_X1 U21231 ( .A1(n18456), .A2(n18499), .B1(n18455), .B2(n18143), .ZN(
        n18128) );
  INV_X1 U21232 ( .A(n18147), .ZN(n18168) );
  NOR2_X1 U21233 ( .A1(n18189), .A2(n18126), .ZN(n18457) );
  AND2_X1 U21234 ( .A1(n18555), .A2(n18457), .ZN(n18396) );
  AOI22_X1 U21235 ( .A1(n18460), .A2(n18458), .B1(n18168), .B2(n18396), .ZN(
        n18144) );
  NOR2_X2 U21236 ( .A1(n18305), .A2(n18147), .ZN(n18209) );
  AOI22_X1 U21237 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18144), .B1(
        n18461), .B2(n18209), .ZN(n18127) );
  OAI211_X1 U21238 ( .C1(n18464), .C2(n18454), .A(n18128), .B(n18127), .ZN(
        P3_U2876) );
  INV_X1 U21239 ( .A(n18209), .ZN(n18205) );
  AOI22_X1 U21240 ( .A1(n18467), .A2(n18444), .B1(n18465), .B2(n18143), .ZN(
        n18131) );
  AOI22_X1 U21241 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18144), .B1(
        n18466), .B2(n18499), .ZN(n18130) );
  OAI211_X1 U21242 ( .C1(n18470), .C2(n18205), .A(n18131), .B(n18130), .ZN(
        P3_U2877) );
  INV_X1 U21243 ( .A(n18132), .ZN(n18476) );
  AOI22_X1 U21244 ( .A1(n18472), .A2(n18499), .B1(n18471), .B2(n18143), .ZN(
        n18134) );
  AOI22_X1 U21245 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18144), .B1(
        n18473), .B2(n18444), .ZN(n18133) );
  OAI211_X1 U21246 ( .C1(n18476), .C2(n18205), .A(n18134), .B(n18133), .ZN(
        P3_U2878) );
  INV_X1 U21247 ( .A(n18478), .ZN(n18436) );
  AOI22_X1 U21248 ( .A1(n18477), .A2(n18143), .B1(n18433), .B2(n18499), .ZN(
        n18136) );
  AOI22_X1 U21249 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18144), .B1(
        n18479), .B2(n18209), .ZN(n18135) );
  OAI211_X1 U21250 ( .C1(n18436), .C2(n18454), .A(n18136), .B(n18135), .ZN(
        P3_U2879) );
  AOI22_X1 U21251 ( .A1(n18407), .A2(n18444), .B1(n18484), .B2(n18143), .ZN(
        n18138) );
  AOI22_X1 U21252 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18144), .B1(
        n18485), .B2(n18209), .ZN(n18137) );
  OAI211_X1 U21253 ( .C1(n18410), .C2(n18513), .A(n18138), .B(n18137), .ZN(
        P3_U2880) );
  AOI22_X1 U21254 ( .A1(n9703), .A2(n18444), .B1(n18490), .B2(n18143), .ZN(
        n18140) );
  AOI22_X1 U21255 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18144), .B1(
        n18493), .B2(n18209), .ZN(n18139) );
  OAI211_X1 U21256 ( .C1(n18496), .C2(n18513), .A(n18140), .B(n18139), .ZN(
        P3_U2881) );
  AOI22_X1 U21257 ( .A1(n18498), .A2(n18444), .B1(n18497), .B2(n18143), .ZN(
        n18142) );
  AOI22_X1 U21258 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18144), .B1(
        n18500), .B2(n18209), .ZN(n18141) );
  OAI211_X1 U21259 ( .C1(n18504), .C2(n18513), .A(n18142), .B(n18141), .ZN(
        P3_U2882) );
  AOI22_X1 U21260 ( .A1(n18508), .A2(n18499), .B1(n18506), .B2(n18143), .ZN(
        n18146) );
  AOI22_X1 U21261 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18144), .B1(
        n18509), .B2(n18444), .ZN(n18145) );
  OAI211_X1 U21262 ( .C1(n18514), .C2(n18205), .A(n18146), .B(n18145), .ZN(
        P3_U2883) );
  NOR2_X1 U21263 ( .A1(n18555), .A2(n18147), .ZN(n18213) );
  NAND2_X1 U21264 ( .A1(n18553), .A2(n18213), .ZN(n18225) );
  NOR2_X1 U21265 ( .A1(n18209), .A2(n18231), .ZN(n18191) );
  NOR2_X1 U21266 ( .A1(n18421), .A2(n18191), .ZN(n18164) );
  AOI22_X1 U21267 ( .A1(n18456), .A2(n18185), .B1(n18455), .B2(n18164), .ZN(
        n18151) );
  OAI21_X1 U21268 ( .B1(n18148), .B2(n18423), .A(n18191), .ZN(n18149) );
  OAI211_X1 U21269 ( .C1(n18231), .C2(n18678), .A(n18426), .B(n18149), .ZN(
        n18165) );
  AOI22_X1 U21270 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18165), .B1(
        n18461), .B2(n18231), .ZN(n18150) );
  OAI211_X1 U21271 ( .C1(n18464), .C2(n18513), .A(n18151), .B(n18150), .ZN(
        P3_U2884) );
  AOI22_X1 U21272 ( .A1(n18467), .A2(n18499), .B1(n18465), .B2(n18164), .ZN(
        n18153) );
  AOI22_X1 U21273 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18165), .B1(
        n18466), .B2(n18185), .ZN(n18152) );
  OAI211_X1 U21274 ( .C1(n18470), .C2(n18225), .A(n18153), .B(n18152), .ZN(
        P3_U2885) );
  AOI22_X1 U21275 ( .A1(n18471), .A2(n18164), .B1(n18473), .B2(n18499), .ZN(
        n18155) );
  AOI22_X1 U21276 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18165), .B1(
        n18472), .B2(n18185), .ZN(n18154) );
  OAI211_X1 U21277 ( .C1(n18476), .C2(n18225), .A(n18155), .B(n18154), .ZN(
        P3_U2886) );
  AOI22_X1 U21278 ( .A1(n18478), .A2(n18499), .B1(n18477), .B2(n18164), .ZN(
        n18157) );
  AOI22_X1 U21279 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18165), .B1(
        n18479), .B2(n18231), .ZN(n18156) );
  OAI211_X1 U21280 ( .C1(n18482), .C2(n18183), .A(n18157), .B(n18156), .ZN(
        P3_U2887) );
  AOI22_X1 U21281 ( .A1(n18407), .A2(n18499), .B1(n18484), .B2(n18164), .ZN(
        n18159) );
  AOI22_X1 U21282 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18165), .B1(
        n18485), .B2(n18231), .ZN(n18158) );
  OAI211_X1 U21283 ( .C1(n18410), .C2(n18183), .A(n18159), .B(n18158), .ZN(
        P3_U2888) );
  AOI22_X1 U21284 ( .A1(n9703), .A2(n18499), .B1(n18490), .B2(n18164), .ZN(
        n18161) );
  AOI22_X1 U21285 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18165), .B1(
        n18493), .B2(n18231), .ZN(n18160) );
  OAI211_X1 U21286 ( .C1(n18496), .C2(n18183), .A(n18161), .B(n18160), .ZN(
        P3_U2889) );
  AOI22_X1 U21287 ( .A1(n18498), .A2(n18499), .B1(n18497), .B2(n18164), .ZN(
        n18163) );
  AOI22_X1 U21288 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18165), .B1(
        n18500), .B2(n18231), .ZN(n18162) );
  OAI211_X1 U21289 ( .C1(n18504), .C2(n18183), .A(n18163), .B(n18162), .ZN(
        P3_U2890) );
  AOI22_X1 U21290 ( .A1(n18509), .A2(n18499), .B1(n18506), .B2(n18164), .ZN(
        n18167) );
  AOI22_X1 U21291 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18165), .B1(
        n18508), .B2(n18185), .ZN(n18166) );
  OAI211_X1 U21292 ( .C1(n18514), .C2(n18225), .A(n18167), .B(n18166), .ZN(
        P3_U2891) );
  AND2_X1 U21293 ( .A1(n18582), .A2(n18213), .ZN(n18184) );
  AOI22_X1 U21294 ( .A1(n18349), .A2(n18185), .B1(n18455), .B2(n18184), .ZN(
        n18170) );
  NAND2_X1 U21295 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18213), .ZN(
        n18252) );
  AOI21_X1 U21296 ( .B1(n18555), .B2(n18423), .A(n18189), .ZN(n18259) );
  OAI211_X1 U21297 ( .C1(n18254), .C2(n18678), .A(n18168), .B(n18259), .ZN(
        n18186) );
  AOI22_X1 U21298 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18186), .B1(
        n18461), .B2(n18254), .ZN(n18169) );
  OAI211_X1 U21299 ( .C1(n18354), .C2(n18205), .A(n18170), .B(n18169), .ZN(
        P3_U2892) );
  AOI22_X1 U21300 ( .A1(n18467), .A2(n18185), .B1(n18465), .B2(n18184), .ZN(
        n18172) );
  AOI22_X1 U21301 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18186), .B1(
        n18466), .B2(n18209), .ZN(n18171) );
  OAI211_X1 U21302 ( .C1(n18470), .C2(n18252), .A(n18172), .B(n18171), .ZN(
        P3_U2893) );
  AOI22_X1 U21303 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18186), .B1(
        n18471), .B2(n18184), .ZN(n18174) );
  AOI22_X1 U21304 ( .A1(n18472), .A2(n18209), .B1(n18473), .B2(n18185), .ZN(
        n18173) );
  OAI211_X1 U21305 ( .C1(n18476), .C2(n18252), .A(n18174), .B(n18173), .ZN(
        P3_U2894) );
  AOI22_X1 U21306 ( .A1(n18478), .A2(n18185), .B1(n18477), .B2(n18184), .ZN(
        n18176) );
  AOI22_X1 U21307 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18186), .B1(
        n18479), .B2(n18254), .ZN(n18175) );
  OAI211_X1 U21308 ( .C1(n18482), .C2(n18205), .A(n18176), .B(n18175), .ZN(
        P3_U2895) );
  AOI22_X1 U21309 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18186), .B1(
        n18484), .B2(n18184), .ZN(n18178) );
  AOI22_X1 U21310 ( .A1(n18407), .A2(n18185), .B1(n18485), .B2(n18254), .ZN(
        n18177) );
  OAI211_X1 U21311 ( .C1(n18410), .C2(n18205), .A(n18178), .B(n18177), .ZN(
        P3_U2896) );
  INV_X1 U21312 ( .A(n9703), .ZN(n18442) );
  AOI22_X1 U21313 ( .A1(n18439), .A2(n18209), .B1(n18490), .B2(n18184), .ZN(
        n18180) );
  AOI22_X1 U21314 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18186), .B1(
        n18493), .B2(n18254), .ZN(n18179) );
  OAI211_X1 U21315 ( .C1(n18442), .C2(n18183), .A(n18180), .B(n18179), .ZN(
        P3_U2897) );
  INV_X1 U21316 ( .A(n18498), .ZN(n18447) );
  AOI22_X1 U21317 ( .A1(n18497), .A2(n18184), .B1(n18443), .B2(n18209), .ZN(
        n18182) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18186), .B1(
        n18500), .B2(n18254), .ZN(n18181) );
  OAI211_X1 U21319 ( .C1(n18447), .C2(n18183), .A(n18182), .B(n18181), .ZN(
        P3_U2898) );
  AOI22_X1 U21320 ( .A1(n18509), .A2(n18185), .B1(n18506), .B2(n18184), .ZN(
        n18188) );
  AOI22_X1 U21321 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18186), .B1(
        n18508), .B2(n18209), .ZN(n18187) );
  OAI211_X1 U21322 ( .C1(n18514), .C2(n18252), .A(n18188), .B(n18187), .ZN(
        P3_U2899) );
  NAND2_X1 U21323 ( .A1(n18281), .A2(n18258), .ZN(n18270) );
  INV_X1 U21324 ( .A(n18270), .ZN(n18277) );
  NOR2_X1 U21325 ( .A1(n18254), .A2(n18277), .ZN(n18236) );
  NOR2_X1 U21326 ( .A1(n18421), .A2(n18236), .ZN(n18208) );
  AOI22_X1 U21327 ( .A1(n18456), .A2(n18231), .B1(n18455), .B2(n18208), .ZN(
        n18194) );
  OAI22_X1 U21328 ( .A1(n18191), .A2(n18190), .B1(n18236), .B2(n18189), .ZN(
        n18192) );
  OAI21_X1 U21329 ( .B1(n18277), .B2(n18678), .A(n18192), .ZN(n18210) );
  AOI22_X1 U21330 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18210), .B1(
        n18461), .B2(n18277), .ZN(n18193) );
  OAI211_X1 U21331 ( .C1(n18464), .C2(n18205), .A(n18194), .B(n18193), .ZN(
        P3_U2900) );
  AOI22_X1 U21332 ( .A1(n18466), .A2(n18231), .B1(n18465), .B2(n18208), .ZN(
        n18196) );
  AOI22_X1 U21333 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18210), .B1(
        n18467), .B2(n18209), .ZN(n18195) );
  OAI211_X1 U21334 ( .C1(n18470), .C2(n18270), .A(n18196), .B(n18195), .ZN(
        P3_U2901) );
  AOI22_X1 U21335 ( .A1(n18472), .A2(n18231), .B1(n18471), .B2(n18208), .ZN(
        n18198) );
  AOI22_X1 U21336 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18210), .B1(
        n18473), .B2(n18209), .ZN(n18197) );
  OAI211_X1 U21337 ( .C1(n18476), .C2(n18270), .A(n18198), .B(n18197), .ZN(
        P3_U2902) );
  AOI22_X1 U21338 ( .A1(n18478), .A2(n18209), .B1(n18477), .B2(n18208), .ZN(
        n18200) );
  AOI22_X1 U21339 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18210), .B1(
        n18479), .B2(n18277), .ZN(n18199) );
  OAI211_X1 U21340 ( .C1(n18482), .C2(n18225), .A(n18200), .B(n18199), .ZN(
        P3_U2903) );
  AOI22_X1 U21341 ( .A1(n18407), .A2(n18209), .B1(n18484), .B2(n18208), .ZN(
        n18202) );
  AOI22_X1 U21342 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18210), .B1(
        n18485), .B2(n18277), .ZN(n18201) );
  OAI211_X1 U21343 ( .C1(n18410), .C2(n18225), .A(n18202), .B(n18201), .ZN(
        P3_U2904) );
  AOI22_X1 U21344 ( .A1(n18439), .A2(n18231), .B1(n18490), .B2(n18208), .ZN(
        n18204) );
  AOI22_X1 U21345 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18210), .B1(
        n18493), .B2(n18277), .ZN(n18203) );
  OAI211_X1 U21346 ( .C1(n18442), .C2(n18205), .A(n18204), .B(n18203), .ZN(
        P3_U2905) );
  AOI22_X1 U21347 ( .A1(n18498), .A2(n18209), .B1(n18497), .B2(n18208), .ZN(
        n18207) );
  AOI22_X1 U21348 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18210), .B1(
        n18500), .B2(n18277), .ZN(n18206) );
  OAI211_X1 U21349 ( .C1(n18504), .C2(n18225), .A(n18207), .B(n18206), .ZN(
        P3_U2906) );
  AOI22_X1 U21350 ( .A1(n18509), .A2(n18209), .B1(n18506), .B2(n18208), .ZN(
        n18212) );
  AOI22_X1 U21351 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18210), .B1(
        n18508), .B2(n18231), .ZN(n18211) );
  OAI211_X1 U21352 ( .C1(n18514), .C2(n18270), .A(n18212), .B(n18211), .ZN(
        P3_U2907) );
  INV_X1 U21353 ( .A(n18258), .ZN(n18214) );
  NOR2_X1 U21354 ( .A1(n18394), .A2(n18214), .ZN(n18230) );
  AOI22_X1 U21355 ( .A1(n18349), .A2(n18231), .B1(n18455), .B2(n18230), .ZN(
        n18216) );
  AOI22_X1 U21356 ( .A1(n18460), .A2(n18213), .B1(n18396), .B2(n18258), .ZN(
        n18232) );
  NOR2_X2 U21357 ( .A1(n18305), .A2(n18214), .ZN(n18299) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18232), .B1(
        n18461), .B2(n18299), .ZN(n18215) );
  OAI211_X1 U21359 ( .C1(n18354), .C2(n18252), .A(n18216), .B(n18215), .ZN(
        P3_U2908) );
  INV_X1 U21360 ( .A(n18299), .ZN(n18275) );
  AOI22_X1 U21361 ( .A1(n18467), .A2(n18231), .B1(n18465), .B2(n18230), .ZN(
        n18218) );
  AOI22_X1 U21362 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18232), .B1(
        n18466), .B2(n18254), .ZN(n18217) );
  OAI211_X1 U21363 ( .C1(n18470), .C2(n18275), .A(n18218), .B(n18217), .ZN(
        P3_U2909) );
  AOI22_X1 U21364 ( .A1(n18472), .A2(n18254), .B1(n18471), .B2(n18230), .ZN(
        n18220) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18232), .B1(
        n18473), .B2(n18231), .ZN(n18219) );
  OAI211_X1 U21366 ( .C1(n18476), .C2(n18275), .A(n18220), .B(n18219), .ZN(
        P3_U2910) );
  AOI22_X1 U21367 ( .A1(n18478), .A2(n18231), .B1(n18477), .B2(n18230), .ZN(
        n18222) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18232), .B1(
        n18479), .B2(n18299), .ZN(n18221) );
  OAI211_X1 U21369 ( .C1(n18482), .C2(n18252), .A(n18222), .B(n18221), .ZN(
        P3_U2911) );
  INV_X1 U21370 ( .A(n18407), .ZN(n18488) );
  AOI22_X1 U21371 ( .A1(n18484), .A2(n18230), .B1(n18483), .B2(n18254), .ZN(
        n18224) );
  AOI22_X1 U21372 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18232), .B1(
        n18485), .B2(n18299), .ZN(n18223) );
  OAI211_X1 U21373 ( .C1(n18488), .C2(n18225), .A(n18224), .B(n18223), .ZN(
        P3_U2912) );
  AOI22_X1 U21374 ( .A1(n9703), .A2(n18231), .B1(n18490), .B2(n18230), .ZN(
        n18227) );
  AOI22_X1 U21375 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18232), .B1(
        n18493), .B2(n18299), .ZN(n18226) );
  OAI211_X1 U21376 ( .C1(n18496), .C2(n18252), .A(n18227), .B(n18226), .ZN(
        P3_U2913) );
  AOI22_X1 U21377 ( .A1(n18498), .A2(n18231), .B1(n18497), .B2(n18230), .ZN(
        n18229) );
  AOI22_X1 U21378 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18232), .B1(
        n18500), .B2(n18299), .ZN(n18228) );
  OAI211_X1 U21379 ( .C1(n18504), .C2(n18252), .A(n18229), .B(n18228), .ZN(
        P3_U2914) );
  AOI22_X1 U21380 ( .A1(n18509), .A2(n18231), .B1(n18506), .B2(n18230), .ZN(
        n18234) );
  AOI22_X1 U21381 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18232), .B1(
        n18508), .B2(n18254), .ZN(n18233) );
  OAI211_X1 U21382 ( .C1(n18514), .C2(n18275), .A(n18234), .B(n18233), .ZN(
        P3_U2915) );
  NOR2_X1 U21383 ( .A1(n18235), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18304) );
  NAND2_X1 U21384 ( .A1(n18553), .A2(n18304), .ZN(n18314) );
  INV_X1 U21385 ( .A(n18314), .ZN(n18321) );
  NOR2_X1 U21386 ( .A1(n18299), .A2(n18321), .ZN(n18282) );
  NOR2_X1 U21387 ( .A1(n18421), .A2(n18282), .ZN(n18253) );
  AOI22_X1 U21388 ( .A1(n18349), .A2(n18254), .B1(n18455), .B2(n18253), .ZN(
        n18239) );
  OAI21_X1 U21389 ( .B1(n18236), .B2(n18423), .A(n18282), .ZN(n18237) );
  OAI211_X1 U21390 ( .C1(n18321), .C2(n18678), .A(n18426), .B(n18237), .ZN(
        n18255) );
  AOI22_X1 U21391 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18255), .B1(
        n18461), .B2(n18321), .ZN(n18238) );
  OAI211_X1 U21392 ( .C1(n18354), .C2(n18270), .A(n18239), .B(n18238), .ZN(
        P3_U2916) );
  AOI22_X1 U21393 ( .A1(n18467), .A2(n18254), .B1(n18465), .B2(n18253), .ZN(
        n18241) );
  AOI22_X1 U21394 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18255), .B1(
        n18466), .B2(n18277), .ZN(n18240) );
  OAI211_X1 U21395 ( .C1(n18470), .C2(n18314), .A(n18241), .B(n18240), .ZN(
        P3_U2917) );
  AOI22_X1 U21396 ( .A1(n18472), .A2(n18277), .B1(n18471), .B2(n18253), .ZN(
        n18243) );
  AOI22_X1 U21397 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18255), .B1(
        n18473), .B2(n18254), .ZN(n18242) );
  OAI211_X1 U21398 ( .C1(n18476), .C2(n18314), .A(n18243), .B(n18242), .ZN(
        P3_U2918) );
  AOI22_X1 U21399 ( .A1(n18478), .A2(n18254), .B1(n18477), .B2(n18253), .ZN(
        n18245) );
  AOI22_X1 U21400 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18255), .B1(
        n18479), .B2(n18321), .ZN(n18244) );
  OAI211_X1 U21401 ( .C1(n18482), .C2(n18270), .A(n18245), .B(n18244), .ZN(
        P3_U2919) );
  AOI22_X1 U21402 ( .A1(n18407), .A2(n18254), .B1(n18484), .B2(n18253), .ZN(
        n18247) );
  AOI22_X1 U21403 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18255), .B1(
        n18485), .B2(n18321), .ZN(n18246) );
  OAI211_X1 U21404 ( .C1(n18410), .C2(n18270), .A(n18247), .B(n18246), .ZN(
        P3_U2920) );
  AOI22_X1 U21405 ( .A1(n9703), .A2(n18254), .B1(n18490), .B2(n18253), .ZN(
        n18249) );
  AOI22_X1 U21406 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18255), .B1(
        n18493), .B2(n18321), .ZN(n18248) );
  OAI211_X1 U21407 ( .C1(n18496), .C2(n18270), .A(n18249), .B(n18248), .ZN(
        P3_U2921) );
  AOI22_X1 U21408 ( .A1(n18497), .A2(n18253), .B1(n18443), .B2(n18277), .ZN(
        n18251) );
  AOI22_X1 U21409 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18255), .B1(
        n18500), .B2(n18321), .ZN(n18250) );
  OAI211_X1 U21410 ( .C1(n18447), .C2(n18252), .A(n18251), .B(n18250), .ZN(
        P3_U2922) );
  AOI22_X1 U21411 ( .A1(n18509), .A2(n18254), .B1(n18506), .B2(n18253), .ZN(
        n18257) );
  AOI22_X1 U21412 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18255), .B1(
        n18508), .B2(n18277), .ZN(n18256) );
  OAI211_X1 U21413 ( .C1(n18514), .C2(n18314), .A(n18257), .B(n18256), .ZN(
        P3_U2923) );
  NAND2_X1 U21414 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18304), .ZN(
        n18343) );
  INV_X1 U21415 ( .A(n18343), .ZN(n18345) );
  OAI211_X1 U21416 ( .C1(n18345), .C2(n18678), .A(n18259), .B(n18258), .ZN(
        n18278) );
  AND2_X1 U21417 ( .A1(n18582), .A2(n18304), .ZN(n18276) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18278), .B1(
        n18455), .B2(n18276), .ZN(n18261) );
  AOI22_X1 U21419 ( .A1(n18349), .A2(n18277), .B1(n18461), .B2(n18345), .ZN(
        n18260) );
  OAI211_X1 U21420 ( .C1(n18354), .C2(n18275), .A(n18261), .B(n18260), .ZN(
        P3_U2924) );
  AOI22_X1 U21421 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18278), .B1(
        n18465), .B2(n18276), .ZN(n18263) );
  AOI22_X1 U21422 ( .A1(n18466), .A2(n18299), .B1(n18467), .B2(n18277), .ZN(
        n18262) );
  OAI211_X1 U21423 ( .C1(n18470), .C2(n18343), .A(n18263), .B(n18262), .ZN(
        P3_U2925) );
  AOI22_X1 U21424 ( .A1(n18472), .A2(n18299), .B1(n18471), .B2(n18276), .ZN(
        n18265) );
  AOI22_X1 U21425 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18278), .B1(
        n18473), .B2(n18277), .ZN(n18264) );
  OAI211_X1 U21426 ( .C1(n18476), .C2(n18343), .A(n18265), .B(n18264), .ZN(
        P3_U2926) );
  AOI22_X1 U21427 ( .A1(n18477), .A2(n18276), .B1(n18433), .B2(n18299), .ZN(
        n18267) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18278), .B1(
        n18479), .B2(n18345), .ZN(n18266) );
  OAI211_X1 U21429 ( .C1(n18436), .C2(n18270), .A(n18267), .B(n18266), .ZN(
        P3_U2927) );
  AOI22_X1 U21430 ( .A1(n18484), .A2(n18276), .B1(n18483), .B2(n18299), .ZN(
        n18269) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18278), .B1(
        n18485), .B2(n18345), .ZN(n18268) );
  OAI211_X1 U21432 ( .C1(n18488), .C2(n18270), .A(n18269), .B(n18268), .ZN(
        P3_U2928) );
  AOI22_X1 U21433 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18278), .B1(
        n18490), .B2(n18276), .ZN(n18272) );
  AOI22_X1 U21434 ( .A1(n9703), .A2(n18277), .B1(n18493), .B2(n18345), .ZN(
        n18271) );
  OAI211_X1 U21435 ( .C1(n18496), .C2(n18275), .A(n18272), .B(n18271), .ZN(
        P3_U2929) );
  AOI22_X1 U21436 ( .A1(n18498), .A2(n18277), .B1(n18497), .B2(n18276), .ZN(
        n18274) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18278), .B1(
        n18500), .B2(n18345), .ZN(n18273) );
  OAI211_X1 U21438 ( .C1(n18504), .C2(n18275), .A(n18274), .B(n18273), .ZN(
        P3_U2930) );
  AOI22_X1 U21439 ( .A1(n18508), .A2(n18299), .B1(n18506), .B2(n18276), .ZN(
        n18280) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18278), .B1(
        n18509), .B2(n18277), .ZN(n18279) );
  OAI211_X1 U21441 ( .C1(n18514), .C2(n18343), .A(n18280), .B(n18279), .ZN(
        P3_U2931) );
  NAND2_X1 U21442 ( .A1(n18281), .A2(n18303), .ZN(n18336) );
  INV_X1 U21443 ( .A(n18336), .ZN(n18368) );
  NOR2_X1 U21444 ( .A1(n18345), .A2(n18368), .ZN(n18326) );
  NOR2_X1 U21445 ( .A1(n18421), .A2(n18326), .ZN(n18298) );
  AOI22_X1 U21446 ( .A1(n18349), .A2(n18299), .B1(n18455), .B2(n18298), .ZN(
        n18285) );
  OAI21_X1 U21447 ( .B1(n18282), .B2(n18423), .A(n18326), .ZN(n18283) );
  OAI211_X1 U21448 ( .C1(n18368), .C2(n18678), .A(n18426), .B(n18283), .ZN(
        n18300) );
  AOI22_X1 U21449 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18300), .B1(
        n18461), .B2(n18368), .ZN(n18284) );
  OAI211_X1 U21450 ( .C1(n18354), .C2(n18314), .A(n18285), .B(n18284), .ZN(
        P3_U2932) );
  AOI22_X1 U21451 ( .A1(n18466), .A2(n18321), .B1(n18465), .B2(n18298), .ZN(
        n18287) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18300), .B1(
        n18467), .B2(n18299), .ZN(n18286) );
  OAI211_X1 U21453 ( .C1(n18470), .C2(n18336), .A(n18287), .B(n18286), .ZN(
        P3_U2933) );
  AOI22_X1 U21454 ( .A1(n18472), .A2(n18321), .B1(n18471), .B2(n18298), .ZN(
        n18289) );
  AOI22_X1 U21455 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18300), .B1(
        n18473), .B2(n18299), .ZN(n18288) );
  OAI211_X1 U21456 ( .C1(n18476), .C2(n18336), .A(n18289), .B(n18288), .ZN(
        P3_U2934) );
  AOI22_X1 U21457 ( .A1(n18478), .A2(n18299), .B1(n18477), .B2(n18298), .ZN(
        n18291) );
  AOI22_X1 U21458 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18300), .B1(
        n18479), .B2(n18368), .ZN(n18290) );
  OAI211_X1 U21459 ( .C1(n18482), .C2(n18314), .A(n18291), .B(n18290), .ZN(
        P3_U2935) );
  AOI22_X1 U21460 ( .A1(n18407), .A2(n18299), .B1(n18484), .B2(n18298), .ZN(
        n18293) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18300), .B1(
        n18485), .B2(n18368), .ZN(n18292) );
  OAI211_X1 U21462 ( .C1(n18410), .C2(n18314), .A(n18293), .B(n18292), .ZN(
        P3_U2936) );
  AOI22_X1 U21463 ( .A1(n9703), .A2(n18299), .B1(n18490), .B2(n18298), .ZN(
        n18295) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18300), .B1(
        n18493), .B2(n18368), .ZN(n18294) );
  OAI211_X1 U21465 ( .C1(n18496), .C2(n18314), .A(n18295), .B(n18294), .ZN(
        P3_U2937) );
  AOI22_X1 U21466 ( .A1(n18498), .A2(n18299), .B1(n18497), .B2(n18298), .ZN(
        n18297) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18300), .B1(
        n18500), .B2(n18368), .ZN(n18296) );
  OAI211_X1 U21468 ( .C1(n18504), .C2(n18314), .A(n18297), .B(n18296), .ZN(
        P3_U2938) );
  AOI22_X1 U21469 ( .A1(n18509), .A2(n18299), .B1(n18506), .B2(n18298), .ZN(
        n18302) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18300), .B1(
        n18508), .B2(n18321), .ZN(n18301) );
  OAI211_X1 U21471 ( .C1(n18514), .C2(n18336), .A(n18302), .B(n18301), .ZN(
        P3_U2939) );
  NOR2_X1 U21472 ( .A1(n18325), .A2(n18394), .ZN(n18350) );
  AOI22_X1 U21473 ( .A1(n18456), .A2(n18345), .B1(n18455), .B2(n18350), .ZN(
        n18307) );
  AOI22_X1 U21474 ( .A1(n18460), .A2(n18304), .B1(n18303), .B2(n18396), .ZN(
        n18322) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18322), .B1(
        n18390), .B2(n18461), .ZN(n18306) );
  OAI211_X1 U21476 ( .C1(n18464), .C2(n18314), .A(n18307), .B(n18306), .ZN(
        P3_U2940) );
  INV_X1 U21477 ( .A(n18390), .ZN(n18388) );
  AOI22_X1 U21478 ( .A1(n18466), .A2(n18345), .B1(n18465), .B2(n18350), .ZN(
        n18309) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18322), .B1(
        n18467), .B2(n18321), .ZN(n18308) );
  OAI211_X1 U21480 ( .C1(n18388), .C2(n18470), .A(n18309), .B(n18308), .ZN(
        P3_U2941) );
  AOI22_X1 U21481 ( .A1(n18472), .A2(n18345), .B1(n18471), .B2(n18350), .ZN(
        n18311) );
  AOI22_X1 U21482 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18322), .B1(
        n18473), .B2(n18321), .ZN(n18310) );
  OAI211_X1 U21483 ( .C1(n18388), .C2(n18476), .A(n18311), .B(n18310), .ZN(
        P3_U2942) );
  AOI22_X1 U21484 ( .A1(n18477), .A2(n18350), .B1(n18433), .B2(n18345), .ZN(
        n18313) );
  AOI22_X1 U21485 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18322), .B1(
        n18390), .B2(n18479), .ZN(n18312) );
  OAI211_X1 U21486 ( .C1(n18436), .C2(n18314), .A(n18313), .B(n18312), .ZN(
        P3_U2943) );
  AOI22_X1 U21487 ( .A1(n18407), .A2(n18321), .B1(n18484), .B2(n18350), .ZN(
        n18316) );
  AOI22_X1 U21488 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18322), .B1(
        n18390), .B2(n18485), .ZN(n18315) );
  OAI211_X1 U21489 ( .C1(n18410), .C2(n18343), .A(n18316), .B(n18315), .ZN(
        P3_U2944) );
  AOI22_X1 U21490 ( .A1(n9703), .A2(n18321), .B1(n18490), .B2(n18350), .ZN(
        n18318) );
  AOI22_X1 U21491 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18322), .B1(
        n18390), .B2(n18493), .ZN(n18317) );
  OAI211_X1 U21492 ( .C1(n18496), .C2(n18343), .A(n18318), .B(n18317), .ZN(
        P3_U2945) );
  AOI22_X1 U21493 ( .A1(n18498), .A2(n18321), .B1(n18497), .B2(n18350), .ZN(
        n18320) );
  AOI22_X1 U21494 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18322), .B1(
        n18390), .B2(n18500), .ZN(n18319) );
  OAI211_X1 U21495 ( .C1(n18504), .C2(n18343), .A(n18320), .B(n18319), .ZN(
        P3_U2946) );
  AOI22_X1 U21496 ( .A1(n18509), .A2(n18321), .B1(n18506), .B2(n18350), .ZN(
        n18324) );
  AOI22_X1 U21497 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18322), .B1(
        n18508), .B2(n18345), .ZN(n18323) );
  OAI211_X1 U21498 ( .C1(n18388), .C2(n18514), .A(n18324), .B(n18323), .ZN(
        P3_U2947) );
  NOR2_X1 U21499 ( .A1(n18555), .A2(n18325), .ZN(n18398) );
  NAND2_X1 U21500 ( .A1(n18553), .A2(n18398), .ZN(n18415) );
  NOR2_X1 U21501 ( .A1(n18390), .A2(n18416), .ZN(n18372) );
  NOR2_X1 U21502 ( .A1(n18421), .A2(n18372), .ZN(n18344) );
  AOI22_X1 U21503 ( .A1(n18456), .A2(n18368), .B1(n18455), .B2(n18344), .ZN(
        n18329) );
  OAI21_X1 U21504 ( .B1(n18326), .B2(n18423), .A(n18372), .ZN(n18327) );
  OAI211_X1 U21505 ( .C1(n18416), .C2(n18678), .A(n18426), .B(n18327), .ZN(
        n18346) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18346), .B1(
        n18416), .B2(n18461), .ZN(n18328) );
  OAI211_X1 U21507 ( .C1(n18464), .C2(n18343), .A(n18329), .B(n18328), .ZN(
        P3_U2948) );
  AOI22_X1 U21508 ( .A1(n18466), .A2(n18368), .B1(n18465), .B2(n18344), .ZN(
        n18331) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18346), .B1(
        n18467), .B2(n18345), .ZN(n18330) );
  OAI211_X1 U21510 ( .C1(n18415), .C2(n18470), .A(n18331), .B(n18330), .ZN(
        P3_U2949) );
  AOI22_X1 U21511 ( .A1(n18471), .A2(n18344), .B1(n18473), .B2(n18345), .ZN(
        n18333) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18346), .B1(
        n18472), .B2(n18368), .ZN(n18332) );
  OAI211_X1 U21513 ( .C1(n18415), .C2(n18476), .A(n18333), .B(n18332), .ZN(
        P3_U2950) );
  AOI22_X1 U21514 ( .A1(n18478), .A2(n18345), .B1(n18477), .B2(n18344), .ZN(
        n18335) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18346), .B1(
        n18416), .B2(n18479), .ZN(n18334) );
  OAI211_X1 U21516 ( .C1(n18482), .C2(n18336), .A(n18335), .B(n18334), .ZN(
        P3_U2951) );
  AOI22_X1 U21517 ( .A1(n18484), .A2(n18344), .B1(n18483), .B2(n18368), .ZN(
        n18338) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18346), .B1(
        n18416), .B2(n18485), .ZN(n18337) );
  OAI211_X1 U21519 ( .C1(n18488), .C2(n18343), .A(n18338), .B(n18337), .ZN(
        P3_U2952) );
  AOI22_X1 U21520 ( .A1(n18439), .A2(n18368), .B1(n18490), .B2(n18344), .ZN(
        n18340) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18346), .B1(
        n18416), .B2(n18493), .ZN(n18339) );
  OAI211_X1 U21522 ( .C1(n18442), .C2(n18343), .A(n18340), .B(n18339), .ZN(
        P3_U2953) );
  AOI22_X1 U21523 ( .A1(n18497), .A2(n18344), .B1(n18443), .B2(n18368), .ZN(
        n18342) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18346), .B1(
        n18416), .B2(n18500), .ZN(n18341) );
  OAI211_X1 U21525 ( .C1(n18447), .C2(n18343), .A(n18342), .B(n18341), .ZN(
        P3_U2954) );
  AOI22_X1 U21526 ( .A1(n18509), .A2(n18345), .B1(n18506), .B2(n18344), .ZN(
        n18348) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18346), .B1(
        n18508), .B2(n18368), .ZN(n18347) );
  OAI211_X1 U21528 ( .C1(n18415), .C2(n18514), .A(n18348), .B(n18347), .ZN(
        P3_U2955) );
  INV_X1 U21529 ( .A(n18398), .ZN(n18351) );
  NOR2_X1 U21530 ( .A1(n18421), .A2(n18351), .ZN(n18367) );
  AOI22_X1 U21531 ( .A1(n18349), .A2(n18368), .B1(n18455), .B2(n18367), .ZN(
        n18353) );
  AOI22_X1 U21532 ( .A1(n18460), .A2(n18350), .B1(n18398), .B2(n18457), .ZN(
        n18369) );
  NOR2_X2 U21533 ( .A1(n18553), .A2(n18351), .ZN(n18450) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18369), .B1(
        n18450), .B2(n18461), .ZN(n18352) );
  OAI211_X1 U21535 ( .C1(n18388), .C2(n18354), .A(n18353), .B(n18352), .ZN(
        P3_U2956) );
  INV_X1 U21536 ( .A(n18450), .ZN(n18448) );
  AOI22_X1 U21537 ( .A1(n18390), .A2(n18466), .B1(n18465), .B2(n18367), .ZN(
        n18356) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18369), .B1(
        n18467), .B2(n18368), .ZN(n18355) );
  OAI211_X1 U21539 ( .C1(n18448), .C2(n18470), .A(n18356), .B(n18355), .ZN(
        P3_U2957) );
  AOI22_X1 U21540 ( .A1(n18471), .A2(n18367), .B1(n18473), .B2(n18368), .ZN(
        n18358) );
  AOI22_X1 U21541 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18369), .B1(
        n18390), .B2(n18472), .ZN(n18357) );
  OAI211_X1 U21542 ( .C1(n18448), .C2(n18476), .A(n18358), .B(n18357), .ZN(
        P3_U2958) );
  AOI22_X1 U21543 ( .A1(n18478), .A2(n18368), .B1(n18477), .B2(n18367), .ZN(
        n18360) );
  AOI22_X1 U21544 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18369), .B1(
        n18450), .B2(n18479), .ZN(n18359) );
  OAI211_X1 U21545 ( .C1(n18388), .C2(n18482), .A(n18360), .B(n18359), .ZN(
        P3_U2959) );
  AOI22_X1 U21546 ( .A1(n18407), .A2(n18368), .B1(n18484), .B2(n18367), .ZN(
        n18362) );
  AOI22_X1 U21547 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18369), .B1(
        n18450), .B2(n18485), .ZN(n18361) );
  OAI211_X1 U21548 ( .C1(n18388), .C2(n18410), .A(n18362), .B(n18361), .ZN(
        P3_U2960) );
  AOI22_X1 U21549 ( .A1(n9703), .A2(n18368), .B1(n18490), .B2(n18367), .ZN(
        n18364) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18369), .B1(
        n18450), .B2(n18493), .ZN(n18363) );
  OAI211_X1 U21551 ( .C1(n18388), .C2(n18496), .A(n18364), .B(n18363), .ZN(
        P3_U2961) );
  AOI22_X1 U21552 ( .A1(n18498), .A2(n18368), .B1(n18497), .B2(n18367), .ZN(
        n18366) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18369), .B1(
        n18450), .B2(n18500), .ZN(n18365) );
  OAI211_X1 U21554 ( .C1(n18388), .C2(n18504), .A(n18366), .B(n18365), .ZN(
        P3_U2962) );
  AOI22_X1 U21555 ( .A1(n18509), .A2(n18368), .B1(n18506), .B2(n18367), .ZN(
        n18371) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18369), .B1(
        n18390), .B2(n18508), .ZN(n18370) );
  OAI211_X1 U21557 ( .C1(n18448), .C2(n18514), .A(n18371), .B(n18370), .ZN(
        P3_U2963) );
  INV_X1 U21558 ( .A(n9702), .ZN(n18489) );
  AOI21_X1 U21559 ( .B1(n18489), .B2(n18448), .A(n18421), .ZN(n18389) );
  AOI22_X1 U21560 ( .A1(n18416), .A2(n18456), .B1(n18455), .B2(n18389), .ZN(
        n18375) );
  AOI221_X1 U21561 ( .B1(n18372), .B2(n18448), .C1(n18423), .C2(n18448), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18373) );
  OAI21_X1 U21562 ( .B1(n9702), .B2(n18373), .A(n18426), .ZN(n18391) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18391), .B1(
        n9702), .B2(n18461), .ZN(n18374) );
  OAI211_X1 U21564 ( .C1(n18464), .C2(n18388), .A(n18375), .B(n18374), .ZN(
        P3_U2964) );
  AOI22_X1 U21565 ( .A1(n18390), .A2(n18467), .B1(n18389), .B2(n18465), .ZN(
        n18377) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18391), .B1(
        n18416), .B2(n18466), .ZN(n18376) );
  OAI211_X1 U21567 ( .C1(n18489), .C2(n18470), .A(n18377), .B(n18376), .ZN(
        P3_U2965) );
  AOI22_X1 U21568 ( .A1(n18390), .A2(n18473), .B1(n18389), .B2(n18471), .ZN(
        n18379) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18391), .B1(
        n18416), .B2(n18472), .ZN(n18378) );
  OAI211_X1 U21570 ( .C1(n18489), .C2(n18476), .A(n18379), .B(n18378), .ZN(
        P3_U2966) );
  AOI22_X1 U21571 ( .A1(n18416), .A2(n18433), .B1(n18389), .B2(n18477), .ZN(
        n18381) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18391), .B1(
        n9702), .B2(n18479), .ZN(n18380) );
  OAI211_X1 U21573 ( .C1(n18388), .C2(n18436), .A(n18381), .B(n18380), .ZN(
        P3_U2967) );
  AOI22_X1 U21574 ( .A1(n18416), .A2(n18483), .B1(n18389), .B2(n18484), .ZN(
        n18383) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18391), .B1(
        n9702), .B2(n18485), .ZN(n18382) );
  OAI211_X1 U21576 ( .C1(n18388), .C2(n18488), .A(n18383), .B(n18382), .ZN(
        P3_U2968) );
  AOI22_X1 U21577 ( .A1(n18416), .A2(n18439), .B1(n18389), .B2(n18490), .ZN(
        n18385) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18391), .B1(
        n9702), .B2(n18493), .ZN(n18384) );
  OAI211_X1 U21579 ( .C1(n18388), .C2(n18442), .A(n18385), .B(n18384), .ZN(
        P3_U2969) );
  AOI22_X1 U21580 ( .A1(n18416), .A2(n18443), .B1(n18389), .B2(n18497), .ZN(
        n18387) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18391), .B1(
        n9702), .B2(n18500), .ZN(n18386) );
  OAI211_X1 U21582 ( .C1(n18388), .C2(n18447), .A(n18387), .B(n18386), .ZN(
        P3_U2970) );
  AOI22_X1 U21583 ( .A1(n18390), .A2(n18509), .B1(n18389), .B2(n18506), .ZN(
        n18393) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18391), .B1(
        n18416), .B2(n18508), .ZN(n18392) );
  OAI211_X1 U21585 ( .C1(n18489), .C2(n18514), .A(n18393), .B(n18392), .ZN(
        P3_U2971) );
  NOR2_X1 U21586 ( .A1(n18395), .A2(n18394), .ZN(n18459) );
  AOI22_X1 U21587 ( .A1(n18450), .A2(n18456), .B1(n18455), .B2(n18459), .ZN(
        n18400) );
  INV_X1 U21588 ( .A(n18395), .ZN(n18397) );
  AOI22_X1 U21589 ( .A1(n18460), .A2(n18398), .B1(n18397), .B2(n18396), .ZN(
        n18417) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18417), .B1(
        n18461), .B2(n18507), .ZN(n18399) );
  OAI211_X1 U21591 ( .C1(n18464), .C2(n18415), .A(n18400), .B(n18399), .ZN(
        P3_U2972) );
  AOI22_X1 U21592 ( .A1(n18416), .A2(n18467), .B1(n18465), .B2(n18459), .ZN(
        n18402) );
  AOI22_X1 U21593 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18417), .B1(
        n18450), .B2(n18466), .ZN(n18401) );
  OAI211_X1 U21594 ( .C1(n18470), .C2(n18503), .A(n18402), .B(n18401), .ZN(
        P3_U2973) );
  AOI22_X1 U21595 ( .A1(n18416), .A2(n18473), .B1(n18471), .B2(n18459), .ZN(
        n18404) );
  AOI22_X1 U21596 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18417), .B1(
        n18450), .B2(n18472), .ZN(n18403) );
  OAI211_X1 U21597 ( .C1(n18476), .C2(n18503), .A(n18404), .B(n18403), .ZN(
        P3_U2974) );
  AOI22_X1 U21598 ( .A1(n18450), .A2(n18433), .B1(n18477), .B2(n18459), .ZN(
        n18406) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18417), .B1(
        n18479), .B2(n18507), .ZN(n18405) );
  OAI211_X1 U21600 ( .C1(n18415), .C2(n18436), .A(n18406), .B(n18405), .ZN(
        P3_U2975) );
  AOI22_X1 U21601 ( .A1(n18416), .A2(n18407), .B1(n18484), .B2(n18459), .ZN(
        n18409) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18417), .B1(
        n18485), .B2(n18507), .ZN(n18408) );
  OAI211_X1 U21603 ( .C1(n18448), .C2(n18410), .A(n18409), .B(n18408), .ZN(
        P3_U2976) );
  AOI22_X1 U21604 ( .A1(n18416), .A2(n9703), .B1(n18490), .B2(n18459), .ZN(
        n18412) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18417), .B1(
        n18493), .B2(n18507), .ZN(n18411) );
  OAI211_X1 U21606 ( .C1(n18448), .C2(n18496), .A(n18412), .B(n18411), .ZN(
        P3_U2977) );
  AOI22_X1 U21607 ( .A1(n18450), .A2(n18443), .B1(n18497), .B2(n18459), .ZN(
        n18414) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18417), .B1(
        n18500), .B2(n18507), .ZN(n18413) );
  OAI211_X1 U21609 ( .C1(n18415), .C2(n18447), .A(n18414), .B(n18413), .ZN(
        P3_U2978) );
  AOI22_X1 U21610 ( .A1(n18450), .A2(n18508), .B1(n18506), .B2(n18459), .ZN(
        n18419) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18417), .B1(
        n18416), .B2(n18509), .ZN(n18418) );
  OAI211_X1 U21612 ( .C1(n18514), .C2(n18503), .A(n18419), .B(n18418), .ZN(
        P3_U2979) );
  INV_X1 U21613 ( .A(n18420), .ZN(n18422) );
  NOR2_X1 U21614 ( .A1(n18421), .A2(n18422), .ZN(n18449) );
  AOI22_X1 U21615 ( .A1(n9702), .A2(n18456), .B1(n18455), .B2(n18449), .ZN(
        n18428) );
  NOR2_X1 U21616 ( .A1(n9702), .A2(n18450), .ZN(n18424) );
  OAI21_X1 U21617 ( .B1(n18424), .B2(n18423), .A(n18422), .ZN(n18425) );
  OAI211_X1 U21618 ( .C1(n18444), .C2(n18678), .A(n18426), .B(n18425), .ZN(
        n18451) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18451), .B1(
        n18461), .B2(n18444), .ZN(n18427) );
  OAI211_X1 U21620 ( .C1(n18464), .C2(n18448), .A(n18428), .B(n18427), .ZN(
        P3_U2980) );
  AOI22_X1 U21621 ( .A1(n9702), .A2(n18466), .B1(n18465), .B2(n18449), .ZN(
        n18430) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18451), .B1(
        n18450), .B2(n18467), .ZN(n18429) );
  OAI211_X1 U21623 ( .C1(n18470), .C2(n18454), .A(n18430), .B(n18429), .ZN(
        P3_U2981) );
  AOI22_X1 U21624 ( .A1(n9702), .A2(n18472), .B1(n18471), .B2(n18449), .ZN(
        n18432) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18451), .B1(
        n18450), .B2(n18473), .ZN(n18431) );
  OAI211_X1 U21626 ( .C1(n18476), .C2(n18454), .A(n18432), .B(n18431), .ZN(
        P3_U2982) );
  AOI22_X1 U21627 ( .A1(n9702), .A2(n18433), .B1(n18477), .B2(n18449), .ZN(
        n18435) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18451), .B1(
        n18479), .B2(n18444), .ZN(n18434) );
  OAI211_X1 U21629 ( .C1(n18448), .C2(n18436), .A(n18435), .B(n18434), .ZN(
        P3_U2983) );
  AOI22_X1 U21630 ( .A1(n9702), .A2(n18483), .B1(n18484), .B2(n18449), .ZN(
        n18438) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18451), .B1(
        n18485), .B2(n18444), .ZN(n18437) );
  OAI211_X1 U21632 ( .C1(n18448), .C2(n18488), .A(n18438), .B(n18437), .ZN(
        P3_U2984) );
  AOI22_X1 U21633 ( .A1(n9702), .A2(n18439), .B1(n18490), .B2(n18449), .ZN(
        n18441) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18451), .B1(
        n18493), .B2(n18444), .ZN(n18440) );
  OAI211_X1 U21635 ( .C1(n18448), .C2(n18442), .A(n18441), .B(n18440), .ZN(
        P3_U2985) );
  AOI22_X1 U21636 ( .A1(n9702), .A2(n18443), .B1(n18497), .B2(n18449), .ZN(
        n18446) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18451), .B1(
        n18500), .B2(n18444), .ZN(n18445) );
  OAI211_X1 U21638 ( .C1(n18448), .C2(n18447), .A(n18446), .B(n18445), .ZN(
        P3_U2986) );
  AOI22_X1 U21639 ( .A1(n9702), .A2(n18508), .B1(n18506), .B2(n18449), .ZN(
        n18453) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18451), .B1(
        n18450), .B2(n18509), .ZN(n18452) );
  OAI211_X1 U21641 ( .C1(n18514), .C2(n18454), .A(n18453), .B(n18452), .ZN(
        P3_U2987) );
  AND2_X1 U21642 ( .A1(n18582), .A2(n18458), .ZN(n18505) );
  AOI22_X1 U21643 ( .A1(n18456), .A2(n18507), .B1(n18455), .B2(n18505), .ZN(
        n18463) );
  AOI22_X1 U21644 ( .A1(n18460), .A2(n18459), .B1(n18458), .B2(n18457), .ZN(
        n18510) );
  AOI22_X1 U21645 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18510), .B1(
        n18461), .B2(n18499), .ZN(n18462) );
  OAI211_X1 U21646 ( .C1(n18464), .C2(n18489), .A(n18463), .B(n18462), .ZN(
        P3_U2988) );
  AOI22_X1 U21647 ( .A1(n18466), .A2(n18507), .B1(n18465), .B2(n18505), .ZN(
        n18469) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18510), .B1(
        n9702), .B2(n18467), .ZN(n18468) );
  OAI211_X1 U21649 ( .C1(n18470), .C2(n18513), .A(n18469), .B(n18468), .ZN(
        P3_U2989) );
  AOI22_X1 U21650 ( .A1(n18472), .A2(n18507), .B1(n18471), .B2(n18505), .ZN(
        n18475) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18510), .B1(
        n9702), .B2(n18473), .ZN(n18474) );
  OAI211_X1 U21652 ( .C1(n18476), .C2(n18513), .A(n18475), .B(n18474), .ZN(
        P3_U2990) );
  AOI22_X1 U21653 ( .A1(n9702), .A2(n18478), .B1(n18477), .B2(n18505), .ZN(
        n18481) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18510), .B1(
        n18479), .B2(n18499), .ZN(n18480) );
  OAI211_X1 U21655 ( .C1(n18482), .C2(n18503), .A(n18481), .B(n18480), .ZN(
        P3_U2991) );
  AOI22_X1 U21656 ( .A1(n18484), .A2(n18505), .B1(n18483), .B2(n18507), .ZN(
        n18487) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18510), .B1(
        n18485), .B2(n18499), .ZN(n18486) );
  OAI211_X1 U21658 ( .C1(n18489), .C2(n18488), .A(n18487), .B(n18486), .ZN(
        P3_U2992) );
  AOI22_X1 U21659 ( .A1(n9703), .A2(n9702), .B1(n18490), .B2(n18505), .ZN(
        n18495) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18510), .B1(
        n18493), .B2(n18499), .ZN(n18494) );
  OAI211_X1 U21661 ( .C1(n18496), .C2(n18503), .A(n18495), .B(n18494), .ZN(
        P3_U2993) );
  AOI22_X1 U21662 ( .A1(n9702), .A2(n18498), .B1(n18497), .B2(n18505), .ZN(
        n18502) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18510), .B1(
        n18500), .B2(n18499), .ZN(n18501) );
  OAI211_X1 U21664 ( .C1(n18504), .C2(n18503), .A(n18502), .B(n18501), .ZN(
        P3_U2994) );
  AOI22_X1 U21665 ( .A1(n18508), .A2(n18507), .B1(n18506), .B2(n18505), .ZN(
        n18512) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18510), .B1(
        n9702), .B2(n18509), .ZN(n18511) );
  OAI211_X1 U21667 ( .C1(n18514), .C2(n18513), .A(n18512), .B(n18511), .ZN(
        P3_U2995) );
  NOR2_X1 U21668 ( .A1(n18545), .A2(n18515), .ZN(n18517) );
  OAI222_X1 U21669 ( .A1(n18521), .A2(n18520), .B1(n18519), .B2(n18518), .C1(
        n18517), .C2(n18516), .ZN(n18722) );
  OAI21_X1 U21670 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18522), .ZN(n18523) );
  OAI211_X1 U21671 ( .C1(n18525), .C2(n18546), .A(n18524), .B(n18523), .ZN(
        n18569) );
  AOI21_X1 U21672 ( .B1(n18547), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n18534), .ZN(n18550) );
  INV_X1 U21673 ( .A(n18550), .ZN(n18526) );
  AOI22_X1 U21674 ( .A1(n18527), .A2(n18526), .B1(n18545), .B2(n18531), .ZN(
        n18681) );
  NOR2_X1 U21675 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18681), .ZN(
        n18537) );
  AOI21_X1 U21676 ( .B1(n18530), .B2(n18529), .A(n18528), .ZN(n18541) );
  OAI21_X1 U21677 ( .B1(n18532), .B2(n18541), .A(n18531), .ZN(n18533) );
  AOI21_X1 U21678 ( .B1(n18535), .B2(n18534), .A(n18533), .ZN(n18679) );
  NAND2_X1 U21679 ( .A1(n18546), .A2(n18679), .ZN(n18536) );
  AOI22_X1 U21680 ( .A1(n18546), .A2(n18537), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18536), .ZN(n18567) );
  AOI21_X1 U21681 ( .B1(n18539), .B2(n18538), .A(n18550), .ZN(n18544) );
  NOR3_X1 U21682 ( .A1(n18542), .A2(n18541), .A3(n18540), .ZN(n18543) );
  AOI211_X1 U21683 ( .C1(n18545), .C2(n18690), .A(n18544), .B(n18543), .ZN(
        n18693) );
  AOI22_X1 U21684 ( .A1(n18558), .A2(n18697), .B1(n18693), .B2(n18546), .ZN(
        n18562) );
  NOR2_X1 U21685 ( .A1(n18548), .A2(n18547), .ZN(n18552) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18549), .B1(
        n18552), .B2(n18709), .ZN(n18705) );
  INV_X1 U21687 ( .A(n18700), .ZN(n18551) );
  OAI22_X1 U21688 ( .A1(n18552), .A2(n18551), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18550), .ZN(n18701) );
  OR3_X1 U21689 ( .A1(n18705), .A2(n18555), .A3(n18553), .ZN(n18554) );
  AOI22_X1 U21690 ( .A1(n18705), .A2(n18555), .B1(n18701), .B2(n18554), .ZN(
        n18557) );
  OAI21_X1 U21691 ( .B1(n18558), .B2(n18557), .A(n18556), .ZN(n18561) );
  AND2_X1 U21692 ( .A1(n18562), .A2(n18561), .ZN(n18559) );
  OAI221_X1 U21693 ( .B1(n18562), .B2(n18561), .C1(n18560), .C2(n18559), .A(
        n18564), .ZN(n18566) );
  AOI21_X1 U21694 ( .B1(n18564), .B2(n18563), .A(n18562), .ZN(n18565) );
  AOI222_X1 U21695 ( .A1(n18567), .A2(n18566), .B1(n18567), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18566), .C2(n18565), .ZN(
        n18568) );
  NOR4_X1 U21696 ( .A1(n18570), .A2(n18722), .A3(n18569), .A4(n18568), .ZN(
        n18580) );
  AOI22_X1 U21697 ( .A1(n18704), .A2(n18735), .B1(n18730), .B2(n17301), .ZN(
        n18571) );
  INV_X1 U21698 ( .A(n18571), .ZN(n18576) );
  OAI211_X1 U21699 ( .C1(n18573), .C2(n18572), .A(n18726), .B(n18580), .ZN(
        n18677) );
  OAI21_X1 U21700 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18723), .A(n18677), 
        .ZN(n18581) );
  NOR2_X1 U21701 ( .A1(n18574), .A2(n18581), .ZN(n18575) );
  MUX2_X1 U21702 ( .A(n18576), .B(n18575), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18578) );
  OAI211_X1 U21703 ( .C1(n18580), .C2(n18579), .A(n18578), .B(n18577), .ZN(
        P3_U2996) );
  NAND2_X1 U21704 ( .A1(n18730), .A2(n17301), .ZN(n18587) );
  NOR4_X1 U21705 ( .A1(n18732), .A2(n18689), .A3(n18723), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18590) );
  INV_X1 U21706 ( .A(n18590), .ZN(n18586) );
  INV_X1 U21707 ( .A(n18581), .ZN(n18583) );
  NAND3_X1 U21708 ( .A1(n18584), .A2(n18583), .A3(n18582), .ZN(n18585) );
  NAND4_X1 U21709 ( .A1(n18588), .A2(n18587), .A3(n18586), .A4(n18585), .ZN(
        P3_U2997) );
  OAI21_X1 U21710 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18589), .ZN(n18591) );
  AOI21_X1 U21711 ( .B1(n18592), .B2(n18591), .A(n18590), .ZN(P3_U2998) );
  INV_X1 U21712 ( .A(P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20997) );
  NOR2_X1 U21713 ( .A1(n20997), .A2(n18675), .ZN(P3_U2999) );
  AND2_X1 U21714 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18672), .ZN(
        P3_U3000) );
  AND2_X1 U21715 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18672), .ZN(
        P3_U3001) );
  AND2_X1 U21716 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18672), .ZN(
        P3_U3002) );
  AND2_X1 U21717 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18672), .ZN(
        P3_U3003) );
  AND2_X1 U21718 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18672), .ZN(
        P3_U3004) );
  AND2_X1 U21719 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18672), .ZN(
        P3_U3005) );
  AND2_X1 U21720 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18672), .ZN(
        P3_U3006) );
  INV_X1 U21721 ( .A(P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20940) );
  NOR2_X1 U21722 ( .A1(n20940), .A2(n18675), .ZN(P3_U3007) );
  AND2_X1 U21723 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18672), .ZN(
        P3_U3008) );
  INV_X1 U21724 ( .A(P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n20902) );
  NOR2_X1 U21725 ( .A1(n20902), .A2(n18675), .ZN(P3_U3009) );
  AND2_X1 U21726 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18672), .ZN(
        P3_U3010) );
  INV_X1 U21727 ( .A(P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20956) );
  NOR2_X1 U21728 ( .A1(n20956), .A2(n18675), .ZN(P3_U3011) );
  AND2_X1 U21729 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18672), .ZN(
        P3_U3012) );
  AND2_X1 U21730 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18672), .ZN(
        P3_U3013) );
  AND2_X1 U21731 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18672), .ZN(
        P3_U3014) );
  AND2_X1 U21732 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18672), .ZN(
        P3_U3015) );
  AND2_X1 U21733 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18672), .ZN(
        P3_U3016) );
  AND2_X1 U21734 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18672), .ZN(
        P3_U3017) );
  AND2_X1 U21735 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18672), .ZN(
        P3_U3018) );
  AND2_X1 U21736 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18672), .ZN(
        P3_U3019) );
  AND2_X1 U21737 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18672), .ZN(
        P3_U3020) );
  AND2_X1 U21738 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18672), .ZN(P3_U3021) );
  AND2_X1 U21739 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18672), .ZN(P3_U3022) );
  AND2_X1 U21740 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18672), .ZN(P3_U3023) );
  AND2_X1 U21741 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18672), .ZN(P3_U3024) );
  AND2_X1 U21742 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18672), .ZN(P3_U3025) );
  AND2_X1 U21743 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18672), .ZN(P3_U3026) );
  AND2_X1 U21744 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18672), .ZN(P3_U3027) );
  AND2_X1 U21745 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18672), .ZN(P3_U3028) );
  INV_X1 U21746 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18737) );
  AOI21_X1 U21747 ( .B1(HOLD), .B2(n18593), .A(n18737), .ZN(n18596) );
  AOI21_X1 U21748 ( .B1(n18730), .B2(P3_STATE_REG_1__SCAN_IN), .A(n18604), 
        .ZN(n18606) );
  INV_X1 U21749 ( .A(NA), .ZN(n20654) );
  OAI21_X1 U21750 ( .B1(n20654), .B2(n18594), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18605) );
  INV_X1 U21751 ( .A(n18605), .ZN(n18595) );
  OAI22_X1 U21752 ( .A1(n18719), .A2(n18596), .B1(n18606), .B2(n18595), .ZN(
        P3_U3029) );
  NOR2_X1 U21753 ( .A1(n18607), .A2(n20668), .ZN(n18602) );
  NOR3_X1 U21754 ( .A1(n18602), .A2(n18604), .A3(n18737), .ZN(n18597) );
  NOR2_X1 U21755 ( .A1(n18597), .A2(n18727), .ZN(n18598) );
  NAND2_X1 U21756 ( .A1(n18730), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18600) );
  OAI211_X1 U21757 ( .C1(n20668), .C2(n18599), .A(n18598), .B(n18600), .ZN(
        P3_U3030) );
  OAI22_X1 U21758 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18600), .ZN(n18601) );
  OAI22_X1 U21759 ( .A1(n18602), .A2(n18601), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18603) );
  OAI22_X1 U21760 ( .A1(n18606), .A2(n18605), .B1(n18604), .B2(n18603), .ZN(
        P3_U3031) );
  OAI222_X1 U21761 ( .A1(n18711), .A2(n18666), .B1(n18608), .B2(n18739), .C1(
        n18609), .C2(n18658), .ZN(P3_U3032) );
  OAI222_X1 U21762 ( .A1(n18658), .A2(n18611), .B1(n18610), .B2(n18719), .C1(
        n18609), .C2(n18666), .ZN(P3_U3033) );
  OAI222_X1 U21763 ( .A1(n18658), .A2(n18613), .B1(n18612), .B2(n18739), .C1(
        n18611), .C2(n18666), .ZN(P3_U3034) );
  INV_X1 U21764 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18615) );
  OAI222_X1 U21765 ( .A1(n18658), .A2(n18615), .B1(n18614), .B2(n18719), .C1(
        n18613), .C2(n18666), .ZN(P3_U3035) );
  OAI222_X1 U21766 ( .A1(n18658), .A2(n18617), .B1(n18616), .B2(n18739), .C1(
        n18615), .C2(n18666), .ZN(P3_U3036) );
  OAI222_X1 U21767 ( .A1(n18658), .A2(n18619), .B1(n18618), .B2(n18719), .C1(
        n18617), .C2(n18666), .ZN(P3_U3037) );
  OAI222_X1 U21768 ( .A1(n18658), .A2(n18621), .B1(n18620), .B2(n18739), .C1(
        n18619), .C2(n18666), .ZN(P3_U3038) );
  OAI222_X1 U21769 ( .A1(n18658), .A2(n18623), .B1(n18622), .B2(n18739), .C1(
        n18621), .C2(n18666), .ZN(P3_U3039) );
  OAI222_X1 U21770 ( .A1(n18658), .A2(n18624), .B1(n21056), .B2(n18739), .C1(
        n18623), .C2(n18666), .ZN(P3_U3040) );
  INV_X1 U21771 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18626) );
  OAI222_X1 U21772 ( .A1(n18658), .A2(n18626), .B1(n18625), .B2(n18739), .C1(
        n18624), .C2(n18666), .ZN(P3_U3041) );
  OAI222_X1 U21773 ( .A1(n18658), .A2(n18628), .B1(n18627), .B2(n18739), .C1(
        n18626), .C2(n18666), .ZN(P3_U3042) );
  INV_X1 U21774 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18630) );
  OAI222_X1 U21775 ( .A1(n18658), .A2(n18630), .B1(n18629), .B2(n18739), .C1(
        n18628), .C2(n18666), .ZN(P3_U3043) );
  OAI222_X1 U21776 ( .A1(n18658), .A2(n18632), .B1(n18631), .B2(n18739), .C1(
        n18630), .C2(n18666), .ZN(P3_U3044) );
  OAI222_X1 U21777 ( .A1(n18658), .A2(n18634), .B1(n18633), .B2(n18739), .C1(
        n18632), .C2(n18666), .ZN(P3_U3045) );
  OAI222_X1 U21778 ( .A1(n18658), .A2(n18635), .B1(n20870), .B2(n18739), .C1(
        n18634), .C2(n18666), .ZN(P3_U3046) );
  OAI222_X1 U21779 ( .A1(n18658), .A2(n18637), .B1(n18636), .B2(n18739), .C1(
        n18635), .C2(n18666), .ZN(P3_U3047) );
  OAI222_X1 U21780 ( .A1(n18658), .A2(n18639), .B1(n18638), .B2(n18739), .C1(
        n18637), .C2(n18666), .ZN(P3_U3048) );
  OAI222_X1 U21781 ( .A1(n18658), .A2(n18642), .B1(n18640), .B2(n18739), .C1(
        n18639), .C2(n18666), .ZN(P3_U3049) );
  OAI222_X1 U21782 ( .A1(n18642), .A2(n18666), .B1(n18641), .B2(n18739), .C1(
        n20847), .C2(n18658), .ZN(P3_U3050) );
  OAI222_X1 U21783 ( .A1(n18658), .A2(n18645), .B1(n18643), .B2(n18739), .C1(
        n20847), .C2(n18666), .ZN(P3_U3051) );
  OAI222_X1 U21784 ( .A1(n18645), .A2(n18666), .B1(n18644), .B2(n18739), .C1(
        n18646), .C2(n18658), .ZN(P3_U3052) );
  INV_X1 U21785 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18649) );
  OAI222_X1 U21786 ( .A1(n18658), .A2(n18649), .B1(n18647), .B2(n18719), .C1(
        n18646), .C2(n18666), .ZN(P3_U3053) );
  OAI222_X1 U21787 ( .A1(n18649), .A2(n18666), .B1(n18648), .B2(n18719), .C1(
        n18650), .C2(n18658), .ZN(P3_U3054) );
  OAI222_X1 U21788 ( .A1(n18658), .A2(n18652), .B1(n18651), .B2(n18719), .C1(
        n18650), .C2(n18666), .ZN(P3_U3055) );
  OAI222_X1 U21789 ( .A1(n18658), .A2(n18654), .B1(n18653), .B2(n18719), .C1(
        n18652), .C2(n18666), .ZN(P3_U3056) );
  OAI222_X1 U21790 ( .A1(n18658), .A2(n18656), .B1(n18655), .B2(n18719), .C1(
        n18654), .C2(n18666), .ZN(P3_U3057) );
  INV_X1 U21791 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18660) );
  OAI222_X1 U21792 ( .A1(n18658), .A2(n18660), .B1(n18657), .B2(n18719), .C1(
        n18656), .C2(n18666), .ZN(P3_U3058) );
  OAI222_X1 U21793 ( .A1(n18660), .A2(n18666), .B1(n18659), .B2(n18719), .C1(
        n18661), .C2(n18658), .ZN(P3_U3059) );
  OAI222_X1 U21794 ( .A1(n18658), .A2(n18665), .B1(n18662), .B2(n18719), .C1(
        n18661), .C2(n18666), .ZN(P3_U3060) );
  OAI222_X1 U21795 ( .A1(n18666), .A2(n18665), .B1(n18664), .B2(n18719), .C1(
        n18663), .C2(n18658), .ZN(P3_U3061) );
  OAI22_X1 U21796 ( .A1(n18740), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18739), .ZN(n18667) );
  INV_X1 U21797 ( .A(n18667), .ZN(P3_U3274) );
  OAI22_X1 U21798 ( .A1(n18740), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18739), .ZN(n18668) );
  INV_X1 U21799 ( .A(n18668), .ZN(P3_U3275) );
  OAI22_X1 U21800 ( .A1(n18740), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18739), .ZN(n18669) );
  INV_X1 U21801 ( .A(n18669), .ZN(P3_U3276) );
  OAI22_X1 U21802 ( .A1(n18740), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18739), .ZN(n18670) );
  INV_X1 U21803 ( .A(n18670), .ZN(P3_U3277) );
  INV_X1 U21804 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20900) );
  INV_X1 U21805 ( .A(n18673), .ZN(n18671) );
  AOI21_X1 U21806 ( .B1(n18672), .B2(n20900), .A(n18671), .ZN(P3_U3280) );
  OAI21_X1 U21807 ( .B1(n18675), .B2(n18674), .A(n18673), .ZN(P3_U3281) );
  OAI221_X1 U21808 ( .B1(n18678), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18678), 
        .C2(n18677), .A(n18676), .ZN(P3_U3282) );
  NOR2_X1 U21809 ( .A1(n18679), .A2(n18692), .ZN(n18680) );
  INV_X1 U21810 ( .A(n18707), .ZN(n18710) );
  NOR2_X1 U21811 ( .A1(n18680), .A2(n18710), .ZN(n18685) );
  NOR3_X1 U21812 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18681), .A3(
        n18692), .ZN(n18682) );
  AOI21_X1 U21813 ( .B1(n18704), .B2(n18683), .A(n18682), .ZN(n18684) );
  OAI22_X1 U21814 ( .A1(n18686), .A2(n18685), .B1(n18710), .B2(n18684), .ZN(
        P3_U3285) );
  OAI22_X1 U21815 ( .A1(n18688), .A2(n18687), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18699) );
  INV_X1 U21816 ( .A(n18699), .ZN(n18695) );
  NOR2_X1 U21817 ( .A1(n18689), .A2(n21029), .ZN(n18698) );
  OAI22_X1 U21818 ( .A1(n18693), .A2(n18692), .B1(n18691), .B2(n18690), .ZN(
        n18694) );
  AOI21_X1 U21819 ( .B1(n18695), .B2(n18698), .A(n18694), .ZN(n18696) );
  AOI22_X1 U21820 ( .A1(n18710), .A2(n18697), .B1(n18696), .B2(n18707), .ZN(
        P3_U3288) );
  AOI222_X1 U21821 ( .A1(n18701), .A2(n18706), .B1(n18704), .B2(n18700), .C1(
        n18699), .C2(n18698), .ZN(n18702) );
  AOI22_X1 U21822 ( .A1(n18710), .A2(n18703), .B1(n18702), .B2(n18707), .ZN(
        P3_U3289) );
  AOI222_X1 U21823 ( .A1(n21029), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18706), 
        .B2(n18705), .C1(n18709), .C2(n18704), .ZN(n18708) );
  AOI22_X1 U21824 ( .A1(n18710), .A2(n18709), .B1(n18708), .B2(n18707), .ZN(
        P3_U3290) );
  AOI21_X1 U21825 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18712) );
  AOI22_X1 U21826 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18712), .B2(n18711), .ZN(n18715) );
  INV_X1 U21827 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18714) );
  AOI22_X1 U21828 ( .A1(n18718), .A2(n18715), .B1(n18714), .B2(n18713), .ZN(
        P3_U3292) );
  INV_X1 U21829 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18717) );
  OAI21_X1 U21830 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18718), .ZN(n18716) );
  OAI21_X1 U21831 ( .B1(n18718), .B2(n18717), .A(n18716), .ZN(P3_U3293) );
  INV_X1 U21832 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18744) );
  OAI22_X1 U21833 ( .A1(n18740), .A2(n18744), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n18719), .ZN(n18720) );
  INV_X1 U21834 ( .A(n18720), .ZN(P3_U3294) );
  MUX2_X1 U21835 ( .A(P3_MORE_REG_SCAN_IN), .B(n18722), .S(n18721), .Z(
        P3_U3295) );
  AOI21_X1 U21836 ( .B1(n17301), .B2(n18723), .A(n18745), .ZN(n18724) );
  OAI21_X1 U21837 ( .B1(n18726), .B2(n18725), .A(n18724), .ZN(n18738) );
  OAI21_X1 U21838 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18728), .A(n18727), 
        .ZN(n18731) );
  AOI211_X1 U21839 ( .C1(n18746), .C2(n18731), .A(n18730), .B(n18729), .ZN(
        n18733) );
  NOR2_X1 U21840 ( .A1(n18733), .A2(n18732), .ZN(n18734) );
  OAI21_X1 U21841 ( .B1(n18735), .B2(n18734), .A(n18738), .ZN(n18736) );
  OAI21_X1 U21842 ( .B1(n18738), .B2(n18737), .A(n18736), .ZN(P3_U3296) );
  OAI22_X1 U21843 ( .A1(n18740), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18739), .ZN(n18741) );
  INV_X1 U21844 ( .A(n18741), .ZN(P3_U3297) );
  INV_X1 U21845 ( .A(n18742), .ZN(n18743) );
  NOR2_X1 U21846 ( .A1(n18743), .A2(n18745), .ZN(n18749) );
  AOI22_X1 U21847 ( .A1(n18746), .A2(n18745), .B1(n18749), .B2(n18744), .ZN(
        P3_U3298) );
  INV_X1 U21848 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18748) );
  AOI21_X1 U21849 ( .B1(n18749), .B2(n18748), .A(n18747), .ZN(P3_U3299) );
  INV_X1 U21850 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19621) );
  NAND2_X1 U21851 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19621), .ZN(n19612) );
  INV_X1 U21852 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19606) );
  AOI22_X1 U21853 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19612), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n19606), .ZN(n19679) );
  AOI21_X1 U21854 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19679), .ZN(n18750) );
  INV_X1 U21855 ( .A(n18750), .ZN(P2_U2815) );
  INV_X1 U21856 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18752) );
  OAI22_X1 U21857 ( .A1(n18753), .A2(n18752), .B1(n19727), .B2(n18751), .ZN(
        P2_U2816) );
  INV_X1 U21858 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20989) );
  OR2_X1 U21859 ( .A1(n20989), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n19748) );
  AOI22_X1 U21860 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(n19748), .B1(n19616), .B2(
        n19606), .ZN(n18754) );
  OAI21_X1 U21861 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n19748), .A(n18754), 
        .ZN(P2_U2817) );
  OAI21_X1 U21862 ( .B1(n19616), .B2(BS16), .A(n19679), .ZN(n19677) );
  OAI21_X1 U21863 ( .B1(n19679), .B2(n19738), .A(n19677), .ZN(P2_U2818) );
  NOR2_X1 U21864 ( .A1(n18756), .A2(n18755), .ZN(n19724) );
  OAI21_X1 U21865 ( .B1(n19724), .B2(n10577), .A(n18757), .ZN(P2_U2819) );
  NOR4_X1 U21866 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18767) );
  NOR4_X1 U21867 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18766) );
  AOI211_X1 U21868 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_4__SCAN_IN), .B(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n18758) );
  INV_X1 U21869 ( .A(P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n21064) );
  INV_X1 U21870 ( .A(P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n21018) );
  NAND3_X1 U21871 ( .A1(n18758), .A2(n21064), .A3(n21018), .ZN(n18764) );
  NOR4_X1 U21872 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18762) );
  NOR4_X1 U21873 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18761) );
  NOR4_X1 U21874 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18760) );
  NOR4_X1 U21875 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18759) );
  NAND4_X1 U21876 ( .A1(n18762), .A2(n18761), .A3(n18760), .A4(n18759), .ZN(
        n18763) );
  NOR4_X1 U21877 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(n18764), .A4(n18763), .ZN(n18765) );
  NAND3_X1 U21878 ( .A1(n18767), .A2(n18766), .A3(n18765), .ZN(n18774) );
  NOR2_X1 U21879 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18774), .ZN(n18769) );
  INV_X1 U21880 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20967) );
  AOI22_X1 U21881 ( .A1(n18769), .A2(n18928), .B1(n20967), .B2(n18774), .ZN(
        P2_U2820) );
  OR3_X1 U21882 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18773) );
  INV_X1 U21883 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18768) );
  AOI22_X1 U21884 ( .A1(n18769), .A2(n18773), .B1(n18774), .B2(n18768), .ZN(
        P2_U2821) );
  INV_X1 U21885 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19678) );
  NAND2_X1 U21886 ( .A1(n18769), .A2(n19678), .ZN(n18772) );
  INV_X1 U21887 ( .A(n18774), .ZN(n18776) );
  OAI21_X1 U21888 ( .B1(n18928), .B2(n19622), .A(n18776), .ZN(n18770) );
  OAI21_X1 U21889 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18776), .A(n18770), 
        .ZN(n18771) );
  OAI221_X1 U21890 ( .B1(n18772), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18772), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18771), .ZN(P2_U2822) );
  INV_X1 U21891 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18775) );
  OAI221_X1 U21892 ( .B1(n18776), .B2(n18775), .C1(n18774), .C2(n18773), .A(
        n18772), .ZN(P2_U2823) );
  INV_X1 U21893 ( .A(n18777), .ZN(n18783) );
  OAI22_X1 U21894 ( .A1(n18906), .A2(n10835), .B1(n18908), .B2(n18778), .ZN(
        n18779) );
  AOI21_X1 U21895 ( .B1(n18912), .B2(P2_REIP_REG_21__SCAN_IN), .A(n18779), 
        .ZN(n18780) );
  OAI21_X1 U21896 ( .B1(n18781), .B2(n18927), .A(n18780), .ZN(n18782) );
  AOI21_X1 U21897 ( .B1(n18783), .B2(n18933), .A(n18782), .ZN(n18790) );
  INV_X1 U21898 ( .A(n18784), .ZN(n18788) );
  NAND2_X1 U21899 ( .A1(n18785), .A2(n18870), .ZN(n18787) );
  AOI21_X1 U21900 ( .B1(n18788), .B2(n18787), .A(n19602), .ZN(n18786) );
  OAI21_X1 U21901 ( .B1(n18788), .B2(n18787), .A(n18786), .ZN(n18789) );
  OAI211_X1 U21902 ( .C1(n18921), .C2(n18791), .A(n18790), .B(n18789), .ZN(
        P2_U2834) );
  NAND2_X1 U21903 ( .A1(n18870), .A2(n18792), .ZN(n18793) );
  XOR2_X1 U21904 ( .A(n18794), .B(n18793), .Z(n18803) );
  OAI21_X1 U21905 ( .B1(n19648), .B2(n18929), .A(n11123), .ZN(n18798) );
  OAI22_X1 U21906 ( .A1(n18796), .A2(n18927), .B1(n18908), .B2(n18795), .ZN(
        n18797) );
  AOI211_X1 U21907 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n18922), .A(n18798), .B(
        n18797), .ZN(n18802) );
  AOI22_X1 U21908 ( .A1(n18800), .A2(n18923), .B1(n18799), .B2(n18933), .ZN(
        n18801) );
  OAI211_X1 U21909 ( .C1(n19602), .C2(n18803), .A(n18802), .B(n18801), .ZN(
        P2_U2836) );
  AOI22_X1 U21910 ( .A1(n18922), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18939), .ZN(n18804) );
  OAI21_X1 U21911 ( .B1(n18805), .B2(n18927), .A(n18804), .ZN(n18806) );
  AOI211_X1 U21912 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n18912), .A(n19044), 
        .B(n18806), .ZN(n18812) );
  NOR2_X1 U21913 ( .A1(n18896), .A2(n18807), .ZN(n18823) );
  XNOR2_X1 U21914 ( .A(n18823), .B(n18808), .ZN(n18810) );
  AOI22_X1 U21915 ( .A1(n18810), .A2(n18917), .B1(n18809), .B2(n18933), .ZN(
        n18811) );
  OAI211_X1 U21916 ( .C1(n18813), .C2(n18921), .A(n18812), .B(n18811), .ZN(
        P2_U2837) );
  AOI22_X1 U21917 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(n18922), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18939), .ZN(n18815) );
  OAI211_X1 U21918 ( .C1(n18824), .C2(n18816), .A(n18815), .B(n18814), .ZN(
        n18817) );
  AOI21_X1 U21919 ( .B1(n18912), .B2(P2_REIP_REG_17__SCAN_IN), .A(n18817), 
        .ZN(n18818) );
  OAI21_X1 U21920 ( .B1(n18819), .B2(n18927), .A(n18818), .ZN(n18820) );
  AOI21_X1 U21921 ( .B1(n18821), .B2(n18933), .A(n18820), .ZN(n18827) );
  INV_X1 U21922 ( .A(n18822), .ZN(n18825) );
  OAI211_X1 U21923 ( .C1(n18825), .C2(n18824), .A(n18917), .B(n18823), .ZN(
        n18826) );
  OAI211_X1 U21924 ( .C1(n18921), .C2(n18828), .A(n18827), .B(n18826), .ZN(
        P2_U2838) );
  AOI211_X1 U21925 ( .C1(n18838), .C2(n18831), .A(n18830), .B(n18829), .ZN(
        n18837) );
  AOI22_X1 U21926 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(n18922), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18939), .ZN(n18832) );
  NAND2_X1 U21927 ( .A1(n18814), .A2(n18832), .ZN(n18833) );
  AOI21_X1 U21928 ( .B1(n18912), .B2(P2_REIP_REG_15__SCAN_IN), .A(n18833), 
        .ZN(n18834) );
  OAI21_X1 U21929 ( .B1(n18835), .B2(n18927), .A(n18834), .ZN(n18836) );
  NOR2_X1 U21930 ( .A1(n18837), .A2(n18836), .ZN(n18841) );
  AOI22_X1 U21931 ( .A1(n18839), .A2(n18933), .B1(n18938), .B2(n18838), .ZN(
        n18840) );
  OAI211_X1 U21932 ( .C1(n18842), .C2(n18921), .A(n18841), .B(n18840), .ZN(
        P2_U2840) );
  NOR2_X1 U21933 ( .A1(n18896), .A2(n18843), .ZN(n18845) );
  XOR2_X1 U21934 ( .A(n18845), .B(n18844), .Z(n18852) );
  AOI22_X1 U21935 ( .A1(n18922), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n18939), .ZN(n18846) );
  OAI21_X1 U21936 ( .B1(n18847), .B2(n18927), .A(n18846), .ZN(n18848) );
  AOI211_X1 U21937 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n18912), .A(n19044), 
        .B(n18848), .ZN(n18851) );
  OAI22_X1 U21938 ( .A1(n18955), .A2(n18900), .B1(n18921), .B2(n18987), .ZN(
        n18849) );
  INV_X1 U21939 ( .A(n18849), .ZN(n18850) );
  OAI211_X1 U21940 ( .C1(n19602), .C2(n18852), .A(n18851), .B(n18850), .ZN(
        P2_U2841) );
  OAI21_X1 U21941 ( .B1(n19639), .B2(n18929), .A(n11123), .ZN(n18856) );
  OAI22_X1 U21942 ( .A1(n18854), .A2(n18927), .B1(n18908), .B2(n18853), .ZN(
        n18855) );
  AOI211_X1 U21943 ( .C1(P2_EBX_REG_13__SCAN_IN), .C2(n18922), .A(n18856), .B(
        n18855), .ZN(n18863) );
  NAND2_X1 U21944 ( .A1(n18870), .A2(n18857), .ZN(n18858) );
  XNOR2_X1 U21945 ( .A(n18859), .B(n18858), .ZN(n18861) );
  AOI22_X1 U21946 ( .A1(n18861), .A2(n18917), .B1(n18933), .B2(n18860), .ZN(
        n18862) );
  OAI211_X1 U21947 ( .C1(n18864), .C2(n18921), .A(n18863), .B(n18862), .ZN(
        P2_U2842) );
  OAI21_X1 U21948 ( .B1(n10963), .B2(n18929), .A(n11123), .ZN(n18868) );
  INV_X1 U21949 ( .A(n18865), .ZN(n18866) );
  OAI22_X1 U21950 ( .A1(n18866), .A2(n18927), .B1(n18908), .B2(n10781), .ZN(
        n18867) );
  AOI211_X1 U21951 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n18922), .A(n18868), .B(
        n18867), .ZN(n18876) );
  NAND2_X1 U21952 ( .A1(n18870), .A2(n18869), .ZN(n18871) );
  XNOR2_X1 U21953 ( .A(n18872), .B(n18871), .ZN(n18874) );
  AOI22_X1 U21954 ( .A1(n18874), .A2(n18917), .B1(n18933), .B2(n18873), .ZN(
        n18875) );
  OAI211_X1 U21955 ( .C1(n18877), .C2(n18921), .A(n18876), .B(n18875), .ZN(
        P2_U2846) );
  NAND2_X1 U21956 ( .A1(n18870), .A2(n18878), .ZN(n18880) );
  XOR2_X1 U21957 ( .A(n18880), .B(n18879), .Z(n18892) );
  NAND2_X1 U21958 ( .A1(n18881), .A2(n18933), .ZN(n18888) );
  NAND2_X1 U21959 ( .A1(n18922), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n18883) );
  AOI22_X1 U21960 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18939), .B1(
        P2_REIP_REG_7__SCAN_IN), .B2(n18912), .ZN(n18882) );
  NAND3_X1 U21961 ( .A1(n18883), .A2(n18882), .A3(n11123), .ZN(n18884) );
  AOI21_X1 U21962 ( .B1(n18886), .B2(n18885), .A(n18884), .ZN(n18887) );
  NAND2_X1 U21963 ( .A1(n18888), .A2(n18887), .ZN(n18889) );
  AOI21_X1 U21964 ( .B1(n18890), .B2(n18923), .A(n18889), .ZN(n18891) );
  OAI21_X1 U21965 ( .B1(n18892), .B2(n19602), .A(n18891), .ZN(P2_U2848) );
  OAI22_X1 U21966 ( .A1(n18893), .A2(n18927), .B1(n18908), .B2(n9871), .ZN(
        n18894) );
  AOI211_X1 U21967 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n18912), .A(n19044), .B(
        n18894), .ZN(n18905) );
  NOR2_X1 U21968 ( .A1(n18896), .A2(n18895), .ZN(n18897) );
  XNOR2_X1 U21969 ( .A(n18898), .B(n18897), .ZN(n18903) );
  OAI22_X1 U21970 ( .A1(n18901), .A2(n18921), .B1(n18900), .B2(n18899), .ZN(
        n18902) );
  AOI21_X1 U21971 ( .B1(n18903), .B2(n18917), .A(n18902), .ZN(n18904) );
  OAI211_X1 U21972 ( .C1(n10769), .C2(n18906), .A(n18905), .B(n18904), .ZN(
        P2_U2849) );
  OAI21_X1 U21973 ( .B1(n18907), .B2(n18906), .A(n11123), .ZN(n18911) );
  OAI22_X1 U21974 ( .A1(n18909), .A2(n18927), .B1(n18908), .B2(n10763), .ZN(
        n18910) );
  AOI211_X1 U21975 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18912), .A(n18911), .B(
        n18910), .ZN(n18920) );
  NAND2_X1 U21976 ( .A1(n18870), .A2(n18913), .ZN(n18914) );
  XNOR2_X1 U21977 ( .A(n18915), .B(n18914), .ZN(n18918) );
  AOI22_X1 U21978 ( .A1(n18918), .A2(n18917), .B1(n18933), .B2(n18916), .ZN(
        n18919) );
  OAI211_X1 U21979 ( .C1(n18921), .C2(n19003), .A(n18920), .B(n18919), .ZN(
        P2_U2850) );
  AOI22_X1 U21980 ( .A1(n18924), .A2(n18923), .B1(n18922), .B2(
        P2_EBX_REG_0__SCAN_IN), .ZN(n18925) );
  OAI21_X1 U21981 ( .B1(n18927), .B2(n18926), .A(n18925), .ZN(n18931) );
  NOR2_X1 U21982 ( .A1(n18929), .A2(n18928), .ZN(n18930) );
  AOI211_X1 U21983 ( .C1(n18933), .C2(n18932), .A(n18931), .B(n18930), .ZN(
        n18942) );
  AOI22_X1 U21984 ( .A1(n18937), .A2(n18936), .B1(n18935), .B2(n18934), .ZN(
        n18941) );
  OAI21_X1 U21985 ( .B1(n18939), .B2(n18938), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18940) );
  NAND3_X1 U21986 ( .A1(n18942), .A2(n18941), .A3(n18940), .ZN(P2_U2855) );
  NAND2_X1 U21987 ( .A1(n18944), .A2(n18943), .ZN(n18945) );
  NAND2_X1 U21988 ( .A1(n18946), .A2(n18945), .ZN(n18978) );
  OAI22_X1 U21989 ( .A1(n18978), .A2(n18951), .B1(n18965), .B2(n18947), .ZN(
        n18948) );
  INV_X1 U21990 ( .A(n18948), .ZN(n18949) );
  OAI21_X1 U21991 ( .B1(n13516), .B2(n18950), .A(n18949), .ZN(P2_U2871) );
  AOI211_X1 U21992 ( .C1(n18952), .C2(n13731), .A(n18951), .B(n9778), .ZN(
        n18953) );
  AOI21_X1 U21993 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n13516), .A(n18953), .ZN(
        n18954) );
  OAI21_X1 U21994 ( .B1(n18955), .B2(n13516), .A(n18954), .ZN(P2_U2873) );
  XNOR2_X1 U21995 ( .A(n13611), .B(n18956), .ZN(n18957) );
  AOI22_X1 U21996 ( .A1(n18957), .A2(n18966), .B1(P2_EBX_REG_12__SCAN_IN), 
        .B2(n13516), .ZN(n18958) );
  OAI21_X1 U21997 ( .B1(n18959), .B2(n13516), .A(n18958), .ZN(P2_U2875) );
  XNOR2_X1 U21998 ( .A(n13536), .B(n18960), .ZN(n18962) );
  AOI22_X1 U21999 ( .A1(n18962), .A2(n18966), .B1(n18965), .B2(n18961), .ZN(
        n18963) );
  OAI21_X1 U22000 ( .B1(n18965), .B2(n18964), .A(n18963), .ZN(P2_U2877) );
  INV_X1 U22001 ( .A(n18999), .ZN(n18967) );
  AOI22_X1 U22002 ( .A1(n18967), .A2(n18966), .B1(P2_EBX_REG_4__SCAN_IN), .B2(
        n13516), .ZN(n18968) );
  OAI21_X1 U22003 ( .B1(n13516), .B2(n18969), .A(n18968), .ZN(P2_U2883) );
  INV_X1 U22004 ( .A(n14467), .ZN(n18970) );
  AOI22_X1 U22005 ( .A1(n18980), .A2(n18970), .B1(n18976), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n18972) );
  AOI22_X1 U22006 ( .A1(n18977), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n18995), .ZN(n18971) );
  NAND2_X1 U22007 ( .A1(n18972), .A2(n18971), .ZN(P2_U2888) );
  INV_X1 U22008 ( .A(n18973), .ZN(n18975) );
  AOI22_X1 U22009 ( .A1(n18975), .A2(n18974), .B1(n18995), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n18984) );
  AOI22_X1 U22010 ( .A1(n18977), .A2(BUF1_REG_16__SCAN_IN), .B1(n18976), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n18983) );
  NOR2_X1 U22011 ( .A1(n18978), .A2(n18998), .ZN(n18979) );
  AOI21_X1 U22012 ( .B1(n18981), .B2(n18980), .A(n18979), .ZN(n18982) );
  NAND3_X1 U22013 ( .A1(n18984), .A2(n18983), .A3(n18982), .ZN(P2_U2903) );
  AOI22_X1 U22014 ( .A1(n18997), .A2(n18985), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n18995), .ZN(n18986) );
  OAI21_X1 U22015 ( .B1(n19004), .B2(n18987), .A(n18986), .ZN(P2_U2905) );
  AOI22_X1 U22016 ( .A1(n18997), .A2(n18988), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n18995), .ZN(n18989) );
  OAI21_X1 U22017 ( .B1(n19004), .B2(n18990), .A(n18989), .ZN(P2_U2907) );
  INV_X1 U22018 ( .A(n18991), .ZN(n18994) );
  AOI22_X1 U22019 ( .A1(n18997), .A2(n18992), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n18995), .ZN(n18993) );
  OAI21_X1 U22020 ( .B1(n19004), .B2(n18994), .A(n18993), .ZN(P2_U2909) );
  AOI22_X1 U22021 ( .A1(n18997), .A2(n18996), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n18995), .ZN(n19002) );
  OR3_X1 U22022 ( .A1(n19000), .A2(n18999), .A3(n18998), .ZN(n19001) );
  OAI211_X1 U22023 ( .C1(n19004), .C2(n19003), .A(n19002), .B(n19001), .ZN(
        P2_U2914) );
  NOR2_X1 U22024 ( .A1(n19016), .A2(n19005), .ZN(P2_U2920) );
  INV_X1 U22025 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n20856) );
  INV_X1 U22026 ( .A(n19006), .ZN(n19007) );
  AOI22_X1 U22027 ( .A1(n19040), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(n19007), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n19008) );
  OAI21_X1 U22028 ( .B1(n20856), .B2(n19031), .A(n19008), .ZN(P2_U2931) );
  AOI22_X1 U22029 ( .A1(n19041), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19009) );
  OAI21_X1 U22030 ( .B1(n13062), .B2(n19043), .A(n19009), .ZN(P2_U2936) );
  AOI22_X1 U22031 ( .A1(n19026), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19010) );
  OAI21_X1 U22032 ( .B1(n19011), .B2(n19043), .A(n19010), .ZN(P2_U2937) );
  AOI22_X1 U22033 ( .A1(n19026), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19012) );
  OAI21_X1 U22034 ( .B1(n20918), .B2(n19043), .A(n19012), .ZN(P2_U2938) );
  AOI22_X1 U22035 ( .A1(n19026), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19013) );
  OAI21_X1 U22036 ( .B1(n19014), .B2(n19043), .A(n19013), .ZN(P2_U2939) );
  INV_X1 U22037 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n20931) );
  OAI222_X1 U22038 ( .A1(n20931), .A2(n19031), .B1(n19043), .B2(n19017), .C1(
        n19016), .C2(n19015), .ZN(P2_U2940) );
  AOI22_X1 U22039 ( .A1(n19026), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19018) );
  OAI21_X1 U22040 ( .B1(n19019), .B2(n19043), .A(n19018), .ZN(P2_U2941) );
  AOI22_X1 U22041 ( .A1(n19026), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19020) );
  OAI21_X1 U22042 ( .B1(n19021), .B2(n19043), .A(n19020), .ZN(P2_U2942) );
  AOI22_X1 U22043 ( .A1(n19026), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19022) );
  OAI21_X1 U22044 ( .B1(n19023), .B2(n19043), .A(n19022), .ZN(P2_U2943) );
  AOI22_X1 U22045 ( .A1(n19026), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19024) );
  OAI21_X1 U22046 ( .B1(n19025), .B2(n19043), .A(n19024), .ZN(P2_U2944) );
  AOI22_X1 U22047 ( .A1(n19026), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19027) );
  OAI21_X1 U22048 ( .B1(n19028), .B2(n19043), .A(n19027), .ZN(P2_U2945) );
  INV_X1 U22049 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n20850) );
  AOI22_X1 U22050 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19029), .B1(n19040), .B2(
        P2_DATAO_REG_5__SCAN_IN), .ZN(n19030) );
  OAI21_X1 U22051 ( .B1(n20850), .B2(n19031), .A(n19030), .ZN(P2_U2946) );
  INV_X1 U22052 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19033) );
  AOI22_X1 U22053 ( .A1(n19041), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19032) );
  OAI21_X1 U22054 ( .B1(n19033), .B2(n19043), .A(n19032), .ZN(P2_U2947) );
  INV_X1 U22055 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19035) );
  AOI22_X1 U22056 ( .A1(n19041), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19034) );
  OAI21_X1 U22057 ( .B1(n19035), .B2(n19043), .A(n19034), .ZN(P2_U2948) );
  INV_X1 U22058 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19037) );
  AOI22_X1 U22059 ( .A1(n19041), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19036) );
  OAI21_X1 U22060 ( .B1(n19037), .B2(n19043), .A(n19036), .ZN(P2_U2949) );
  INV_X1 U22061 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19039) );
  AOI22_X1 U22062 ( .A1(n19041), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19038) );
  OAI21_X1 U22063 ( .B1(n19039), .B2(n19043), .A(n19038), .ZN(P2_U2950) );
  AOI22_X1 U22064 ( .A1(n19041), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19040), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19042) );
  OAI21_X1 U22065 ( .B1(n13063), .B2(n19043), .A(n19042), .ZN(P2_U2951) );
  AOI22_X1 U22066 ( .A1(n19055), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19044), .ZN(n19049) );
  AOI222_X1 U22067 ( .A1(n19047), .A2(n19056), .B1(n19063), .B2(n19046), .C1(
        n19045), .C2(n14248), .ZN(n19048) );
  OAI211_X1 U22068 ( .C1(n19061), .C2(n19050), .A(n19049), .B(n19048), .ZN(
        P2_U3010) );
  OAI21_X1 U22069 ( .B1(n19053), .B2(n19052), .A(n19051), .ZN(n19054) );
  XOR2_X1 U22070 ( .A(n19054), .B(n19059), .Z(n19068) );
  AOI22_X1 U22071 ( .A1(n19068), .A2(n19056), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19055), .ZN(n19066) );
  AOI21_X1 U22072 ( .B1(n19059), .B2(n19058), .A(n19057), .ZN(n19071) );
  NOR2_X1 U22073 ( .A1(n18814), .A2(n19622), .ZN(n19076) );
  AOI21_X1 U22074 ( .B1(n14248), .B2(n19071), .A(n19076), .ZN(n19060) );
  OAI21_X1 U22075 ( .B1(n19061), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n19060), .ZN(n19062) );
  AOI21_X1 U22076 ( .B1(n19064), .B2(n19063), .A(n19062), .ZN(n19065) );
  NAND2_X1 U22077 ( .A1(n19066), .A2(n19065), .ZN(P2_U3013) );
  AOI22_X1 U22078 ( .A1(n19069), .A2(n19068), .B1(n19067), .B2(n19706), .ZN(
        n19082) );
  INV_X1 U22079 ( .A(n19070), .ZN(n19077) );
  INV_X1 U22080 ( .A(n19071), .ZN(n19073) );
  OAI22_X1 U22081 ( .A1(n19074), .A2(n19073), .B1(n19072), .B2(n13206), .ZN(
        n19075) );
  AOI211_X1 U22082 ( .C1(n19077), .C2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n19076), .B(n19075), .ZN(n19081) );
  OAI211_X1 U22083 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n19079), .B(n19078), .ZN(n19080) );
  NAND3_X1 U22084 ( .A1(n19082), .A2(n19081), .A3(n19080), .ZN(P2_U3045) );
  INV_X1 U22085 ( .A(n19212), .ZN(n19083) );
  NOR2_X1 U22086 ( .A1(n19442), .A2(n19163), .ZN(n19126) );
  AOI22_X1 U22087 ( .A1(n19547), .A2(n19589), .B1(n19539), .B2(n19126), .ZN(
        n19094) );
  AOI21_X1 U22088 ( .B1(n19577), .B2(n19162), .A(n19738), .ZN(n19085) );
  NOR2_X1 U22089 ( .A1(n19085), .A2(n19685), .ZN(n19089) );
  INV_X1 U22090 ( .A(n19585), .ZN(n19087) );
  AOI21_X1 U22091 ( .B1(n19090), .B2(n19546), .A(n19697), .ZN(n19086) );
  AOI21_X1 U22092 ( .B1(n19089), .B2(n19087), .A(n19086), .ZN(n19088) );
  OAI21_X1 U22093 ( .B1(n19585), .B2(n19126), .A(n19089), .ZN(n19092) );
  OAI21_X1 U22094 ( .B1(n19090), .B2(n19126), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19091) );
  AOI22_X1 U22095 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19129), .B1(
        n19540), .B2(n19128), .ZN(n19093) );
  OAI211_X1 U22096 ( .C1(n19550), .C2(n19162), .A(n19094), .B(n19093), .ZN(
        P2_U3048) );
  AOI22_X1 U22097 ( .A1(n19512), .A2(n19589), .B1(n13769), .B2(n19126), .ZN(
        n19096) );
  AOI22_X1 U22098 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19129), .B1(
        n19551), .B2(n19128), .ZN(n19095) );
  OAI211_X1 U22099 ( .C1(n19488), .C2(n19162), .A(n19096), .B(n19095), .ZN(
        P2_U3049) );
  AOI22_X1 U22100 ( .A1(n19455), .A2(n19589), .B1(n19556), .B2(n19126), .ZN(
        n19098) );
  AOI22_X1 U22101 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19129), .B1(
        n19557), .B2(n19128), .ZN(n19097) );
  OAI211_X1 U22102 ( .C1(n19458), .C2(n19162), .A(n19098), .B(n19097), .ZN(
        P2_U3050) );
  AOI22_X1 U22103 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19120), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19119), .ZN(n19567) );
  OAI22_X2 U22104 ( .A1(n19099), .A2(n19123), .B1(n21026), .B2(n19121), .ZN(
        n19564) );
  AOI22_X1 U22105 ( .A1(n19564), .A2(n19589), .B1(n19562), .B2(n19126), .ZN(
        n19103) );
  NOR2_X2 U22106 ( .A1(n19101), .A2(n19447), .ZN(n19563) );
  AOI22_X1 U22107 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19129), .B1(
        n19563), .B2(n19128), .ZN(n19102) );
  OAI211_X1 U22108 ( .C1(n19567), .C2(n19162), .A(n19103), .B(n19102), .ZN(
        P2_U3051) );
  AOI22_X2 U22109 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19120), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19119), .ZN(n19573) );
  OAI22_X2 U22110 ( .A1(n19105), .A2(n19121), .B1(n19104), .B2(n19123), .ZN(
        n19570) );
  NOR2_X2 U22111 ( .A1(n19125), .A2(n10195), .ZN(n19568) );
  AOI22_X1 U22112 ( .A1(n19570), .A2(n19589), .B1(n19568), .B2(n19126), .ZN(
        n19108) );
  NOR2_X2 U22113 ( .A1(n19106), .A2(n19447), .ZN(n19569) );
  AOI22_X1 U22114 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19129), .B1(
        n19569), .B2(n19128), .ZN(n19107) );
  OAI211_X1 U22115 ( .C1(n19573), .C2(n19162), .A(n19108), .B(n19107), .ZN(
        P2_U3052) );
  AOI22_X2 U22116 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19120), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19119), .ZN(n21087) );
  OAI22_X2 U22117 ( .A1(n19110), .A2(n19121), .B1(n19109), .B2(n19123), .ZN(
        n21080) );
  NOR2_X2 U22118 ( .A1(n19125), .A2(n9757), .ZN(n21078) );
  AOI22_X1 U22119 ( .A1(n21080), .A2(n19589), .B1(n21078), .B2(n19126), .ZN(
        n19113) );
  NOR2_X2 U22120 ( .A1(n19111), .A2(n19447), .ZN(n21082) );
  AOI22_X1 U22121 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19129), .B1(
        n21082), .B2(n19128), .ZN(n19112) );
  OAI211_X1 U22122 ( .C1(n21087), .C2(n19162), .A(n19113), .B(n19112), .ZN(
        P2_U3053) );
  AOI22_X1 U22123 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19120), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19119), .ZN(n19467) );
  NOR2_X2 U22124 ( .A1(n19125), .A2(n19115), .ZN(n19578) );
  AOI22_X1 U22125 ( .A1(n19524), .A2(n19589), .B1(n19578), .B2(n19126), .ZN(
        n19118) );
  NOR2_X2 U22126 ( .A1(n19116), .A2(n19447), .ZN(n19579) );
  AOI22_X1 U22127 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19129), .B1(
        n19579), .B2(n19128), .ZN(n19117) );
  OAI211_X1 U22128 ( .C1(n19467), .C2(n19162), .A(n19118), .B(n19117), .ZN(
        P2_U3054) );
  AOI22_X1 U22129 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19120), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19119), .ZN(n19507) );
  NOR2_X2 U22130 ( .A1(n19125), .A2(n10558), .ZN(n19584) );
  AOI22_X1 U22131 ( .A1(n19502), .A2(n19589), .B1(n19584), .B2(n19126), .ZN(
        n19131) );
  NOR2_X2 U22132 ( .A1(n19127), .A2(n19447), .ZN(n19586) );
  AOI22_X1 U22133 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19129), .B1(
        n19586), .B2(n19128), .ZN(n19130) );
  OAI211_X1 U22134 ( .C1(n19507), .C2(n19162), .A(n19131), .B(n19130), .ZN(
        P2_U3055) );
  NOR2_X2 U22135 ( .A1(n19132), .A2(n19250), .ZN(n19189) );
  INV_X1 U22136 ( .A(n19189), .ZN(n19156) );
  NOR2_X1 U22137 ( .A1(n19163), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19135) );
  INV_X1 U22138 ( .A(n19135), .ZN(n19134) );
  NAND2_X1 U22139 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19135), .ZN(
        n19137) );
  NAND2_X1 U22140 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19137), .ZN(n19133) );
  NOR2_X1 U22141 ( .A1(n10431), .A2(n19133), .ZN(n19139) );
  AOI211_X2 U22142 ( .C1(n19134), .C2(n19732), .A(n19477), .B(n19139), .ZN(
        n19158) );
  INV_X1 U22143 ( .A(n19137), .ZN(n19157) );
  AOI22_X1 U22144 ( .A1(n19158), .A2(n19540), .B1(n19539), .B2(n19157), .ZN(
        n19142) );
  AOI21_X1 U22145 ( .B1(n19136), .B2(n19479), .A(n19135), .ZN(n19140) );
  AND2_X1 U22146 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19137), .ZN(n19138) );
  OR4_X1 U22147 ( .A1(n19140), .A2(n19447), .A3(n19139), .A4(n19138), .ZN(
        n19159) );
  AOI22_X1 U22148 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19159), .B1(
        n19153), .B2(n19547), .ZN(n19141) );
  OAI211_X1 U22149 ( .C1(n19550), .C2(n19156), .A(n19142), .B(n19141), .ZN(
        P2_U3056) );
  AOI22_X1 U22150 ( .A1(n19158), .A2(n19551), .B1(n13769), .B2(n19157), .ZN(
        n19144) );
  AOI22_X1 U22151 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19159), .B1(
        n19189), .B2(n19552), .ZN(n19143) );
  OAI211_X1 U22152 ( .C1(n19555), .C2(n19162), .A(n19144), .B(n19143), .ZN(
        P2_U3057) );
  AOI22_X1 U22153 ( .A1(n19158), .A2(n19557), .B1(n19556), .B2(n19157), .ZN(
        n19146) );
  AOI22_X1 U22154 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19159), .B1(
        n19153), .B2(n19455), .ZN(n19145) );
  OAI211_X1 U22155 ( .C1(n19458), .C2(n19156), .A(n19146), .B(n19145), .ZN(
        P2_U3058) );
  AOI22_X1 U22156 ( .A1(n19158), .A2(n19563), .B1(n19562), .B2(n19157), .ZN(
        n19148) );
  INV_X1 U22157 ( .A(n19567), .ZN(n19515) );
  AOI22_X1 U22158 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19159), .B1(
        n19189), .B2(n19515), .ZN(n19147) );
  OAI211_X1 U22159 ( .C1(n19424), .C2(n19162), .A(n19148), .B(n19147), .ZN(
        P2_U3059) );
  AOI22_X1 U22160 ( .A1(n19158), .A2(n19569), .B1(n19568), .B2(n19157), .ZN(
        n19150) );
  AOI22_X1 U22161 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19159), .B1(
        n19153), .B2(n19570), .ZN(n19149) );
  OAI211_X1 U22162 ( .C1(n19573), .C2(n19156), .A(n19150), .B(n19149), .ZN(
        P2_U3060) );
  AOI22_X1 U22163 ( .A1(n19158), .A2(n21082), .B1(n21078), .B2(n19157), .ZN(
        n19152) );
  AOI22_X1 U22164 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19159), .B1(
        n19153), .B2(n21080), .ZN(n19151) );
  OAI211_X1 U22165 ( .C1(n21087), .C2(n19156), .A(n19152), .B(n19151), .ZN(
        P2_U3061) );
  AOI22_X1 U22166 ( .A1(n19158), .A2(n19579), .B1(n19578), .B2(n19157), .ZN(
        n19155) );
  AOI22_X1 U22167 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19159), .B1(
        n19153), .B2(n19524), .ZN(n19154) );
  OAI211_X1 U22168 ( .C1(n19467), .C2(n19156), .A(n19155), .B(n19154), .ZN(
        P2_U3062) );
  AOI22_X1 U22169 ( .A1(n19158), .A2(n19586), .B1(n19584), .B2(n19157), .ZN(
        n19161) );
  INV_X1 U22170 ( .A(n19507), .ZN(n19588) );
  AOI22_X1 U22171 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19159), .B1(
        n19189), .B2(n19588), .ZN(n19160) );
  OAI211_X1 U22172 ( .C1(n19594), .C2(n19162), .A(n19161), .B(n19160), .ZN(
        P2_U3063) );
  NOR3_X2 U22173 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19708), .A3(
        n19163), .ZN(n19187) );
  OAI21_X1 U22174 ( .B1(n10425), .B2(n19187), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19165) );
  NAND2_X1 U22175 ( .A1(n19376), .A2(n19164), .ZN(n19168) );
  NAND2_X1 U22176 ( .A1(n19165), .A2(n19168), .ZN(n19188) );
  AOI22_X1 U22177 ( .A1(n19188), .A2(n19540), .B1(n19539), .B2(n19187), .ZN(
        n19174) );
  INV_X1 U22178 ( .A(n19187), .ZN(n19166) );
  OAI21_X1 U22179 ( .B1(n19167), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19166), 
        .ZN(n19171) );
  OAI21_X1 U22180 ( .B1(n19201), .B2(n19189), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19169) );
  NAND2_X1 U22181 ( .A1(n19169), .A2(n19168), .ZN(n19170) );
  MUX2_X1 U22182 ( .A(n19171), .B(n19170), .S(n19697), .Z(n19172) );
  NAND2_X1 U22183 ( .A1(n19172), .A2(n19545), .ZN(n19190) );
  AOI22_X1 U22184 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19190), .B1(
        n19189), .B2(n19547), .ZN(n19173) );
  OAI211_X1 U22185 ( .C1(n19550), .C2(n19211), .A(n19174), .B(n19173), .ZN(
        P2_U3064) );
  AOI22_X1 U22186 ( .A1(n19188), .A2(n19551), .B1(n13769), .B2(n19187), .ZN(
        n19176) );
  AOI22_X1 U22187 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19190), .B1(
        n19189), .B2(n19512), .ZN(n19175) );
  OAI211_X1 U22188 ( .C1(n19488), .C2(n19211), .A(n19176), .B(n19175), .ZN(
        P2_U3065) );
  AOI22_X1 U22189 ( .A1(n19188), .A2(n19557), .B1(n19556), .B2(n19187), .ZN(
        n19178) );
  AOI22_X1 U22190 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19190), .B1(
        n19189), .B2(n19455), .ZN(n19177) );
  OAI211_X1 U22191 ( .C1(n19458), .C2(n19211), .A(n19178), .B(n19177), .ZN(
        P2_U3066) );
  AOI22_X1 U22192 ( .A1(n19188), .A2(n19563), .B1(n19562), .B2(n19187), .ZN(
        n19180) );
  AOI22_X1 U22193 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19190), .B1(
        n19189), .B2(n19564), .ZN(n19179) );
  OAI211_X1 U22194 ( .C1(n19567), .C2(n19211), .A(n19180), .B(n19179), .ZN(
        P2_U3067) );
  AOI22_X1 U22195 ( .A1(n19188), .A2(n19569), .B1(n19568), .B2(n19187), .ZN(
        n19182) );
  AOI22_X1 U22196 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19190), .B1(
        n19189), .B2(n19570), .ZN(n19181) );
  OAI211_X1 U22197 ( .C1(n19573), .C2(n19211), .A(n19182), .B(n19181), .ZN(
        P2_U3068) );
  AOI22_X1 U22198 ( .A1(n19188), .A2(n21082), .B1(n21078), .B2(n19187), .ZN(
        n19184) );
  AOI22_X1 U22199 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19190), .B1(
        n19189), .B2(n21080), .ZN(n19183) );
  OAI211_X1 U22200 ( .C1(n21087), .C2(n19211), .A(n19184), .B(n19183), .ZN(
        P2_U3069) );
  AOI22_X1 U22201 ( .A1(n19188), .A2(n19579), .B1(n19578), .B2(n19187), .ZN(
        n19186) );
  AOI22_X1 U22202 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19190), .B1(
        n19189), .B2(n19524), .ZN(n19185) );
  OAI211_X1 U22203 ( .C1(n19467), .C2(n19211), .A(n19186), .B(n19185), .ZN(
        P2_U3070) );
  AOI22_X1 U22204 ( .A1(n19188), .A2(n19586), .B1(n19584), .B2(n19187), .ZN(
        n19192) );
  AOI22_X1 U22205 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19190), .B1(
        n19189), .B2(n19502), .ZN(n19191) );
  OAI211_X1 U22206 ( .C1(n19507), .C2(n19211), .A(n19192), .B(n19191), .ZN(
        P2_U3071) );
  AOI22_X1 U22207 ( .A1(n19512), .A2(n19201), .B1(n19206), .B2(n13769), .ZN(
        n19194) );
  AOI22_X1 U22208 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19208), .B1(
        n19551), .B2(n19207), .ZN(n19193) );
  OAI211_X1 U22209 ( .C1(n19488), .C2(n19243), .A(n19194), .B(n19193), .ZN(
        P2_U3073) );
  AOI22_X1 U22210 ( .A1(n19455), .A2(n19201), .B1(n19556), .B2(n19206), .ZN(
        n19196) );
  AOI22_X1 U22211 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19208), .B1(
        n19557), .B2(n19207), .ZN(n19195) );
  OAI211_X1 U22212 ( .C1(n19458), .C2(n19243), .A(n19196), .B(n19195), .ZN(
        P2_U3074) );
  AOI22_X1 U22213 ( .A1(n19515), .A2(n19245), .B1(n19206), .B2(n19562), .ZN(
        n19198) );
  AOI22_X1 U22214 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19208), .B1(
        n19563), .B2(n19207), .ZN(n19197) );
  OAI211_X1 U22215 ( .C1(n19424), .C2(n19211), .A(n19198), .B(n19197), .ZN(
        P2_U3075) );
  AOI22_X1 U22216 ( .A1(n19570), .A2(n19201), .B1(n19206), .B2(n19568), .ZN(
        n19200) );
  AOI22_X1 U22217 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19208), .B1(
        n19569), .B2(n19207), .ZN(n19199) );
  OAI211_X1 U22218 ( .C1(n19573), .C2(n19243), .A(n19200), .B(n19199), .ZN(
        P2_U3076) );
  AOI22_X1 U22219 ( .A1(n21080), .A2(n19201), .B1(n19206), .B2(n21078), .ZN(
        n19203) );
  AOI22_X1 U22220 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19208), .B1(
        n21082), .B2(n19207), .ZN(n19202) );
  OAI211_X1 U22221 ( .C1(n21087), .C2(n19243), .A(n19203), .B(n19202), .ZN(
        P2_U3077) );
  AOI22_X1 U22222 ( .A1(n19580), .A2(n19245), .B1(n19206), .B2(n19578), .ZN(
        n19205) );
  AOI22_X1 U22223 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19208), .B1(
        n19579), .B2(n19207), .ZN(n19204) );
  OAI211_X1 U22224 ( .C1(n19583), .C2(n19211), .A(n19205), .B(n19204), .ZN(
        P2_U3078) );
  AOI22_X1 U22225 ( .A1(n19588), .A2(n19245), .B1(n19206), .B2(n19584), .ZN(
        n19210) );
  AOI22_X1 U22226 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19208), .B1(
        n19586), .B2(n19207), .ZN(n19209) );
  OAI211_X1 U22227 ( .C1(n19594), .C2(n19211), .A(n19210), .B(n19209), .ZN(
        P2_U3079) );
  INV_X1 U22228 ( .A(n19439), .ZN(n19252) );
  OAI21_X1 U22229 ( .B1(n19245), .B2(n21079), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19213) );
  NAND2_X1 U22230 ( .A1(n19213), .A2(n19697), .ZN(n19224) );
  INV_X1 U22231 ( .A(n19284), .ZN(n19214) );
  AND2_X1 U22232 ( .A1(n19215), .A2(n19214), .ZN(n19445) );
  AND2_X1 U22233 ( .A1(n19445), .A2(n19689), .ZN(n19220) );
  OR2_X1 U22234 ( .A1(n19224), .A2(n19220), .ZN(n19219) );
  NAND2_X1 U22235 ( .A1(n19221), .A2(n19546), .ZN(n19217) );
  NOR2_X1 U22236 ( .A1(n19442), .A2(n19251), .ZN(n19244) );
  NOR2_X1 U22237 ( .A1(n19697), .A2(n19244), .ZN(n19216) );
  AOI21_X1 U22238 ( .B1(n19217), .B2(n19216), .A(n19447), .ZN(n19218) );
  AOI22_X1 U22239 ( .A1(n19508), .A2(n21079), .B1(n19539), .B2(n19244), .ZN(
        n19226) );
  INV_X1 U22240 ( .A(n19220), .ZN(n19223) );
  OAI21_X1 U22241 ( .B1(n19221), .B2(n19244), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19222) );
  AOI22_X1 U22242 ( .A1(n19540), .A2(n19246), .B1(n19245), .B2(n19547), .ZN(
        n19225) );
  OAI211_X1 U22243 ( .C1(n19236), .C2(n19227), .A(n19226), .B(n19225), .ZN(
        P2_U3080) );
  AOI22_X1 U22244 ( .A1(n19552), .A2(n21079), .B1(n13769), .B2(n19244), .ZN(
        n19229) );
  AOI22_X1 U22245 ( .A1(n19551), .A2(n19246), .B1(n19245), .B2(n19512), .ZN(
        n19228) );
  OAI211_X1 U22246 ( .C1(n19236), .C2(n10342), .A(n19229), .B(n19228), .ZN(
        P2_U3081) );
  INV_X1 U22247 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n19232) );
  AOI22_X1 U22248 ( .A1(n19455), .A2(n19245), .B1(n19556), .B2(n19244), .ZN(
        n19231) );
  AOI22_X1 U22249 ( .A1(n19557), .A2(n19246), .B1(n21079), .B2(n19558), .ZN(
        n19230) );
  OAI211_X1 U22250 ( .C1(n19236), .C2(n19232), .A(n19231), .B(n19230), .ZN(
        P2_U3082) );
  INV_X1 U22251 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n19235) );
  AOI22_X1 U22252 ( .A1(n19564), .A2(n19245), .B1(n19562), .B2(n19244), .ZN(
        n19234) );
  AOI22_X1 U22253 ( .A1(n19563), .A2(n19246), .B1(n21079), .B2(n19515), .ZN(
        n19233) );
  OAI211_X1 U22254 ( .C1(n19236), .C2(n19235), .A(n19234), .B(n19233), .ZN(
        P2_U3083) );
  AOI22_X1 U22255 ( .A1(n19570), .A2(n19245), .B1(n19568), .B2(n19244), .ZN(
        n19238) );
  AOI22_X1 U22256 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19247), .B1(
        n19569), .B2(n19246), .ZN(n19237) );
  OAI211_X1 U22257 ( .C1(n19573), .C2(n19273), .A(n19238), .B(n19237), .ZN(
        P2_U3084) );
  AOI22_X1 U22258 ( .A1(n21080), .A2(n19245), .B1(n21078), .B2(n19244), .ZN(
        n19240) );
  AOI22_X1 U22259 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19247), .B1(
        n21082), .B2(n19246), .ZN(n19239) );
  OAI211_X1 U22260 ( .C1(n21087), .C2(n19273), .A(n19240), .B(n19239), .ZN(
        P2_U3085) );
  AOI22_X1 U22261 ( .A1(n19580), .A2(n21079), .B1(n19578), .B2(n19244), .ZN(
        n19242) );
  AOI22_X1 U22262 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19247), .B1(
        n19579), .B2(n19246), .ZN(n19241) );
  OAI211_X1 U22263 ( .C1(n19583), .C2(n19243), .A(n19242), .B(n19241), .ZN(
        P2_U3086) );
  AOI22_X1 U22264 ( .A1(n19502), .A2(n19245), .B1(n19584), .B2(n19244), .ZN(
        n19249) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19247), .B1(
        n19586), .B2(n19246), .ZN(n19248) );
  OAI211_X1 U22266 ( .C1(n19507), .C2(n19273), .A(n19249), .B(n19248), .ZN(
        P2_U3087) );
  NOR2_X1 U22267 ( .A1(n19251), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19256) );
  INV_X1 U22268 ( .A(n19256), .ZN(n19259) );
  NOR2_X1 U22269 ( .A1(n19715), .A2(n19259), .ZN(n21077) );
  AOI22_X1 U22270 ( .A1(n19547), .A2(n21079), .B1(n19539), .B2(n21077), .ZN(
        n19262) );
  NAND2_X1 U22271 ( .A1(n19252), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19480) );
  OAI21_X1 U22272 ( .B1(n19480), .B2(n19681), .A(n19697), .ZN(n19260) );
  INV_X1 U22273 ( .A(n21077), .ZN(n19253) );
  OAI211_X1 U22274 ( .C1(n19254), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19685), 
        .B(n19253), .ZN(n19255) );
  OAI211_X1 U22275 ( .C1(n19260), .C2(n19256), .A(n19545), .B(n19255), .ZN(
        n21083) );
  OAI21_X1 U22276 ( .B1(n19257), .B2(n21077), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19258) );
  OAI21_X1 U22277 ( .B1(n19260), .B2(n19259), .A(n19258), .ZN(n21081) );
  AOI22_X1 U22278 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n21083), .B1(
        n19540), .B2(n21081), .ZN(n19261) );
  OAI211_X1 U22279 ( .C1(n19550), .C2(n21086), .A(n19262), .B(n19261), .ZN(
        P2_U3088) );
  AOI22_X1 U22280 ( .A1(n19512), .A2(n21079), .B1(n13769), .B2(n21077), .ZN(
        n19264) );
  AOI22_X1 U22281 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n21083), .B1(
        n19551), .B2(n21081), .ZN(n19263) );
  OAI211_X1 U22282 ( .C1(n19488), .C2(n21086), .A(n19264), .B(n19263), .ZN(
        P2_U3089) );
  AOI22_X1 U22283 ( .A1(n19558), .A2(n19305), .B1(n19556), .B2(n21077), .ZN(
        n19266) );
  AOI22_X1 U22284 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n21083), .B1(
        n19557), .B2(n21081), .ZN(n19265) );
  OAI211_X1 U22285 ( .C1(n19561), .C2(n19273), .A(n19266), .B(n19265), .ZN(
        P2_U3090) );
  AOI22_X1 U22286 ( .A1(n19515), .A2(n19305), .B1(n19562), .B2(n21077), .ZN(
        n19268) );
  AOI22_X1 U22287 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n21083), .B1(
        n19563), .B2(n21081), .ZN(n19267) );
  OAI211_X1 U22288 ( .C1(n19424), .C2(n19273), .A(n19268), .B(n19267), .ZN(
        P2_U3091) );
  AOI22_X1 U22289 ( .A1(n19570), .A2(n21079), .B1(n19568), .B2(n21077), .ZN(
        n19270) );
  AOI22_X1 U22290 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n21083), .B1(
        n19569), .B2(n21081), .ZN(n19269) );
  OAI211_X1 U22291 ( .C1(n19573), .C2(n21086), .A(n19270), .B(n19269), .ZN(
        P2_U3092) );
  AOI22_X1 U22292 ( .A1(n19580), .A2(n19305), .B1(n19578), .B2(n21077), .ZN(
        n19272) );
  AOI22_X1 U22293 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n21083), .B1(
        n19579), .B2(n21081), .ZN(n19271) );
  OAI211_X1 U22294 ( .C1(n19583), .C2(n19273), .A(n19272), .B(n19271), .ZN(
        P2_U3094) );
  AOI22_X1 U22295 ( .A1(n19502), .A2(n21079), .B1(n19584), .B2(n21077), .ZN(
        n19275) );
  AOI22_X1 U22296 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n21083), .B1(
        n19586), .B2(n21081), .ZN(n19274) );
  OAI211_X1 U22297 ( .C1(n19507), .C2(n21086), .A(n19275), .B(n19274), .ZN(
        P2_U3095) );
  NOR2_X1 U22298 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19276), .ZN(
        n19303) );
  NAND2_X1 U22299 ( .A1(n19284), .A2(n19283), .ZN(n19278) );
  OAI21_X1 U22300 ( .B1(n19305), .B2(n19318), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19277) );
  NAND2_X1 U22301 ( .A1(n19278), .A2(n19277), .ZN(n19279) );
  OAI21_X1 U22302 ( .B1(n19303), .B2(n19546), .A(n19279), .ZN(n19280) );
  NOR2_X1 U22303 ( .A1(n19447), .A2(n19280), .ZN(n19282) );
  INV_X1 U22304 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n20921) );
  NAND3_X1 U22305 ( .A1(n19284), .A2(n19283), .A3(n19546), .ZN(n19287) );
  INV_X1 U22306 ( .A(n19285), .ZN(n19286) );
  AOI22_X1 U22307 ( .A1(n19304), .A2(n19540), .B1(n19539), .B2(n19303), .ZN(
        n19289) );
  AOI22_X1 U22308 ( .A1(n19305), .A2(n19547), .B1(n19318), .B2(n19508), .ZN(
        n19288) );
  OAI211_X1 U22309 ( .C1(n19290), .C2(n20921), .A(n19289), .B(n19288), .ZN(
        P2_U3096) );
  AOI22_X1 U22310 ( .A1(n19304), .A2(n19551), .B1(n13769), .B2(n19303), .ZN(
        n19292) );
  AOI22_X1 U22311 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19306), .B1(
        n19318), .B2(n19552), .ZN(n19291) );
  OAI211_X1 U22312 ( .C1(n19555), .C2(n21086), .A(n19292), .B(n19291), .ZN(
        P2_U3097) );
  AOI22_X1 U22313 ( .A1(n19304), .A2(n19557), .B1(n19556), .B2(n19303), .ZN(
        n19294) );
  AOI22_X1 U22314 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19306), .B1(
        n19318), .B2(n19558), .ZN(n19293) );
  OAI211_X1 U22315 ( .C1(n19561), .C2(n21086), .A(n19294), .B(n19293), .ZN(
        P2_U3098) );
  AOI22_X1 U22316 ( .A1(n19304), .A2(n19563), .B1(n19562), .B2(n19303), .ZN(
        n19296) );
  AOI22_X1 U22317 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19306), .B1(
        n19318), .B2(n19515), .ZN(n19295) );
  OAI211_X1 U22318 ( .C1(n19424), .C2(n21086), .A(n19296), .B(n19295), .ZN(
        P2_U3099) );
  AOI22_X1 U22319 ( .A1(n19304), .A2(n19569), .B1(n19568), .B2(n19303), .ZN(
        n19298) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19306), .B1(
        n19305), .B2(n19570), .ZN(n19297) );
  OAI211_X1 U22321 ( .C1(n19573), .C2(n19327), .A(n19298), .B(n19297), .ZN(
        P2_U3100) );
  AOI22_X1 U22322 ( .A1(n19304), .A2(n21082), .B1(n21078), .B2(n19303), .ZN(
        n19300) );
  AOI22_X1 U22323 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19306), .B1(
        n19305), .B2(n21080), .ZN(n19299) );
  OAI211_X1 U22324 ( .C1(n21087), .C2(n19327), .A(n19300), .B(n19299), .ZN(
        P2_U3101) );
  AOI22_X1 U22325 ( .A1(n19304), .A2(n19579), .B1(n19578), .B2(n19303), .ZN(
        n19302) );
  AOI22_X1 U22326 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19306), .B1(
        n19318), .B2(n19580), .ZN(n19301) );
  OAI211_X1 U22327 ( .C1(n19583), .C2(n21086), .A(n19302), .B(n19301), .ZN(
        P2_U3102) );
  AOI22_X1 U22328 ( .A1(n19304), .A2(n19586), .B1(n19584), .B2(n19303), .ZN(
        n19308) );
  AOI22_X1 U22329 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19306), .B1(
        n19305), .B2(n19502), .ZN(n19307) );
  OAI211_X1 U22330 ( .C1(n19507), .C2(n19327), .A(n19308), .B(n19307), .ZN(
        P2_U3103) );
  INV_X1 U22331 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n20903) );
  AOI22_X1 U22332 ( .A1(n19323), .A2(n19540), .B1(n19539), .B2(n19333), .ZN(
        n19310) );
  AOI22_X1 U22333 ( .A1(n19347), .A2(n19508), .B1(n19318), .B2(n19547), .ZN(
        n19309) );
  OAI211_X1 U22334 ( .C1(n19313), .C2(n20903), .A(n19310), .B(n19309), .ZN(
        P2_U3104) );
  AOI22_X1 U22335 ( .A1(n19323), .A2(n19551), .B1(n13769), .B2(n19333), .ZN(
        n19312) );
  AOI22_X1 U22336 ( .A1(n19347), .A2(n19552), .B1(n19318), .B2(n19512), .ZN(
        n19311) );
  OAI211_X1 U22337 ( .C1(n19313), .C2(n10318), .A(n19312), .B(n19311), .ZN(
        P2_U3105) );
  AOI22_X1 U22338 ( .A1(n19323), .A2(n19563), .B1(n19562), .B2(n19333), .ZN(
        n19315) );
  AOI22_X1 U22339 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19324), .B1(
        n19318), .B2(n19564), .ZN(n19314) );
  OAI211_X1 U22340 ( .C1(n19567), .C2(n19357), .A(n19315), .B(n19314), .ZN(
        P2_U3107) );
  AOI22_X1 U22341 ( .A1(n19323), .A2(n19569), .B1(n19568), .B2(n19333), .ZN(
        n19317) );
  AOI22_X1 U22342 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19324), .B1(
        n19318), .B2(n19570), .ZN(n19316) );
  OAI211_X1 U22343 ( .C1(n19573), .C2(n19357), .A(n19317), .B(n19316), .ZN(
        P2_U3108) );
  AOI22_X1 U22344 ( .A1(n19323), .A2(n21082), .B1(n21078), .B2(n19333), .ZN(
        n19320) );
  AOI22_X1 U22345 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19324), .B1(
        n19318), .B2(n21080), .ZN(n19319) );
  OAI211_X1 U22346 ( .C1(n21087), .C2(n19357), .A(n19320), .B(n19319), .ZN(
        P2_U3109) );
  AOI22_X1 U22347 ( .A1(n19323), .A2(n19579), .B1(n19578), .B2(n19333), .ZN(
        n19322) );
  AOI22_X1 U22348 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19324), .B1(
        n19347), .B2(n19580), .ZN(n19321) );
  OAI211_X1 U22349 ( .C1(n19583), .C2(n19327), .A(n19322), .B(n19321), .ZN(
        P2_U3110) );
  AOI22_X1 U22350 ( .A1(n19323), .A2(n19586), .B1(n19584), .B2(n19333), .ZN(
        n19326) );
  AOI22_X1 U22351 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19324), .B1(
        n19347), .B2(n19588), .ZN(n19325) );
  OAI211_X1 U22352 ( .C1(n19594), .C2(n19327), .A(n19326), .B(n19325), .ZN(
        P2_U3111) );
  NOR2_X1 U22353 ( .A1(n19442), .A2(n19409), .ZN(n19352) );
  AOI22_X1 U22354 ( .A1(n19547), .A2(n19347), .B1(n19539), .B2(n19352), .ZN(
        n19338) );
  AOI21_X1 U22355 ( .B1(n19369), .B2(n19357), .A(n19738), .ZN(n19328) );
  NOR2_X1 U22356 ( .A1(n19328), .A2(n19685), .ZN(n19332) );
  OAI21_X1 U22357 ( .B1(n19334), .B2(n19732), .A(n19546), .ZN(n19329) );
  AOI21_X1 U22358 ( .B1(n19332), .B2(n19330), .A(n19329), .ZN(n19331) );
  OAI21_X1 U22359 ( .B1(n19333), .B2(n19352), .A(n19332), .ZN(n19336) );
  OAI21_X1 U22360 ( .B1(n19334), .B2(n19352), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19335) );
  AOI22_X1 U22361 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19354), .B1(
        n19540), .B2(n19353), .ZN(n19337) );
  OAI211_X1 U22362 ( .C1(n19550), .C2(n19369), .A(n19338), .B(n19337), .ZN(
        P2_U3112) );
  AOI22_X1 U22363 ( .A1(n19552), .A2(n19370), .B1(n13769), .B2(n19352), .ZN(
        n19340) );
  AOI22_X1 U22364 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19354), .B1(
        n19353), .B2(n19551), .ZN(n19339) );
  OAI211_X1 U22365 ( .C1(n19555), .C2(n19357), .A(n19340), .B(n19339), .ZN(
        P2_U3113) );
  AOI22_X1 U22366 ( .A1(n19558), .A2(n19370), .B1(n19556), .B2(n19352), .ZN(
        n19342) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19354), .B1(
        n19353), .B2(n19557), .ZN(n19341) );
  OAI211_X1 U22368 ( .C1(n19561), .C2(n19357), .A(n19342), .B(n19341), .ZN(
        P2_U3114) );
  AOI22_X1 U22369 ( .A1(n19515), .A2(n19370), .B1(n19352), .B2(n19562), .ZN(
        n19344) );
  AOI22_X1 U22370 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19354), .B1(
        n19353), .B2(n19563), .ZN(n19343) );
  OAI211_X1 U22371 ( .C1(n19424), .C2(n19357), .A(n19344), .B(n19343), .ZN(
        P2_U3115) );
  AOI22_X1 U22372 ( .A1(n19570), .A2(n19347), .B1(n19352), .B2(n19568), .ZN(
        n19346) );
  AOI22_X1 U22373 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19354), .B1(
        n19353), .B2(n19569), .ZN(n19345) );
  OAI211_X1 U22374 ( .C1(n19573), .C2(n19369), .A(n19346), .B(n19345), .ZN(
        P2_U3116) );
  AOI22_X1 U22375 ( .A1(n21080), .A2(n19347), .B1(n19352), .B2(n21078), .ZN(
        n19349) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19354), .B1(
        n19353), .B2(n21082), .ZN(n19348) );
  OAI211_X1 U22377 ( .C1(n21087), .C2(n19369), .A(n19349), .B(n19348), .ZN(
        P2_U3117) );
  AOI22_X1 U22378 ( .A1(n19580), .A2(n19370), .B1(n19352), .B2(n19578), .ZN(
        n19351) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19354), .B1(
        n19353), .B2(n19579), .ZN(n19350) );
  OAI211_X1 U22380 ( .C1(n19583), .C2(n19357), .A(n19351), .B(n19350), .ZN(
        P2_U3118) );
  AOI22_X1 U22381 ( .A1(n19588), .A2(n19370), .B1(n19352), .B2(n19584), .ZN(
        n19356) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19354), .B1(
        n19353), .B2(n19586), .ZN(n19355) );
  OAI211_X1 U22383 ( .C1(n19594), .C2(n19357), .A(n19356), .B(n19355), .ZN(
        P2_U3119) );
  INV_X1 U22384 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n19360) );
  AOI22_X1 U22385 ( .A1(n19564), .A2(n19370), .B1(n19379), .B2(n19562), .ZN(
        n19359) );
  AOI22_X1 U22386 ( .A1(n19563), .A2(n19371), .B1(n19400), .B2(n19515), .ZN(
        n19358) );
  OAI211_X1 U22387 ( .C1(n19364), .C2(n19360), .A(n19359), .B(n19358), .ZN(
        P2_U3123) );
  INV_X1 U22388 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n19363) );
  AOI22_X1 U22389 ( .A1(n19570), .A2(n19370), .B1(n19379), .B2(n19568), .ZN(
        n19362) );
  INV_X1 U22390 ( .A(n19573), .ZN(n19519) );
  AOI22_X1 U22391 ( .A1(n19569), .A2(n19371), .B1(n19400), .B2(n19519), .ZN(
        n19361) );
  OAI211_X1 U22392 ( .C1(n19364), .C2(n19363), .A(n19362), .B(n19361), .ZN(
        P2_U3124) );
  AOI22_X1 U22393 ( .A1(n21080), .A2(n19370), .B1(n19379), .B2(n21078), .ZN(
        n19366) );
  AOI22_X1 U22394 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19372), .B1(
        n21082), .B2(n19371), .ZN(n19365) );
  OAI211_X1 U22395 ( .C1(n21087), .C2(n19375), .A(n19366), .B(n19365), .ZN(
        P2_U3125) );
  AOI22_X1 U22396 ( .A1(n19580), .A2(n19400), .B1(n19379), .B2(n19578), .ZN(
        n19368) );
  AOI22_X1 U22397 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19372), .B1(
        n19579), .B2(n19371), .ZN(n19367) );
  OAI211_X1 U22398 ( .C1(n19583), .C2(n19369), .A(n19368), .B(n19367), .ZN(
        P2_U3126) );
  AOI22_X1 U22399 ( .A1(n19502), .A2(n19370), .B1(n19379), .B2(n19584), .ZN(
        n19374) );
  AOI22_X1 U22400 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19372), .B1(
        n19586), .B2(n19371), .ZN(n19373) );
  OAI211_X1 U22401 ( .C1(n19507), .C2(n19375), .A(n19374), .B(n19373), .ZN(
        P2_U3127) );
  INV_X1 U22402 ( .A(n19376), .ZN(n19378) );
  NOR3_X2 U22403 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19708), .A3(
        n19409), .ZN(n19398) );
  OAI21_X1 U22404 ( .B1(n10424), .B2(n19398), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19377) );
  OAI21_X1 U22405 ( .B1(n19409), .B2(n19378), .A(n19377), .ZN(n19399) );
  AOI22_X1 U22406 ( .A1(n19399), .A2(n19540), .B1(n19539), .B2(n19398), .ZN(
        n19385) );
  AOI221_X1 U22407 ( .B1(n19400), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19427), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19379), .ZN(n19381) );
  MUX2_X1 U22408 ( .A(n19381), .B(n19380), .S(P2_STATE2_REG_2__SCAN_IN), .Z(
        n19382) );
  NOR2_X1 U22409 ( .A1(n19382), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19383) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19401), .B1(
        n19400), .B2(n19547), .ZN(n19384) );
  OAI211_X1 U22411 ( .C1(n19550), .C2(n19438), .A(n19385), .B(n19384), .ZN(
        P2_U3128) );
  AOI22_X1 U22412 ( .A1(n19399), .A2(n19551), .B1(n13769), .B2(n19398), .ZN(
        n19387) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19401), .B1(
        n19400), .B2(n19512), .ZN(n19386) );
  OAI211_X1 U22414 ( .C1(n19488), .C2(n19438), .A(n19387), .B(n19386), .ZN(
        P2_U3129) );
  AOI22_X1 U22415 ( .A1(n19399), .A2(n19557), .B1(n19556), .B2(n19398), .ZN(
        n19389) );
  AOI22_X1 U22416 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19401), .B1(
        n19400), .B2(n19455), .ZN(n19388) );
  OAI211_X1 U22417 ( .C1(n19458), .C2(n19438), .A(n19389), .B(n19388), .ZN(
        P2_U3130) );
  AOI22_X1 U22418 ( .A1(n19399), .A2(n19563), .B1(n19562), .B2(n19398), .ZN(
        n19391) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19401), .B1(
        n19400), .B2(n19564), .ZN(n19390) );
  OAI211_X1 U22420 ( .C1(n19567), .C2(n19438), .A(n19391), .B(n19390), .ZN(
        P2_U3131) );
  AOI22_X1 U22421 ( .A1(n19399), .A2(n19569), .B1(n19568), .B2(n19398), .ZN(
        n19393) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19401), .B1(
        n19400), .B2(n19570), .ZN(n19392) );
  OAI211_X1 U22423 ( .C1(n19573), .C2(n19438), .A(n19393), .B(n19392), .ZN(
        P2_U3132) );
  AOI22_X1 U22424 ( .A1(n19399), .A2(n21082), .B1(n21078), .B2(n19398), .ZN(
        n19395) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19401), .B1(
        n19400), .B2(n21080), .ZN(n19394) );
  OAI211_X1 U22426 ( .C1(n21087), .C2(n19438), .A(n19395), .B(n19394), .ZN(
        P2_U3133) );
  AOI22_X1 U22427 ( .A1(n19399), .A2(n19579), .B1(n19578), .B2(n19398), .ZN(
        n19397) );
  AOI22_X1 U22428 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19401), .B1(
        n19400), .B2(n19524), .ZN(n19396) );
  OAI211_X1 U22429 ( .C1(n19467), .C2(n19438), .A(n19397), .B(n19396), .ZN(
        P2_U3134) );
  AOI22_X1 U22430 ( .A1(n19399), .A2(n19586), .B1(n19584), .B2(n19398), .ZN(
        n19403) );
  AOI22_X1 U22431 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19401), .B1(
        n19400), .B2(n19502), .ZN(n19402) );
  OAI211_X1 U22432 ( .C1(n19507), .C2(n19438), .A(n19403), .B(n19402), .ZN(
        P2_U3135) );
  NOR2_X2 U22433 ( .A1(n19405), .A2(n19404), .ZN(n19470) );
  INV_X1 U22434 ( .A(n19470), .ZN(n19430) );
  NAND2_X1 U22435 ( .A1(n19407), .A2(n19406), .ZN(n19412) );
  NAND2_X1 U22436 ( .A1(n19412), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19408) );
  OR2_X1 U22437 ( .A1(n19708), .A2(n19409), .ZN(n19411) );
  OAI21_X1 U22438 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19411), .A(n19732), 
        .ZN(n19410) );
  INV_X1 U22439 ( .A(n19412), .ZN(n19433) );
  AOI22_X1 U22440 ( .A1(n19434), .A2(n19540), .B1(n19539), .B2(n19433), .ZN(
        n19417) );
  OAI21_X1 U22441 ( .B1(n19680), .B2(n19479), .A(n19411), .ZN(n19415) );
  NAND2_X1 U22442 ( .A1(n19412), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19413) );
  NAND4_X1 U22443 ( .A1(n19415), .A2(n19545), .A3(n19414), .A4(n19413), .ZN(
        n19435) );
  AOI22_X1 U22444 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19435), .B1(
        n19427), .B2(n19547), .ZN(n19416) );
  OAI211_X1 U22445 ( .C1(n19550), .C2(n19430), .A(n19417), .B(n19416), .ZN(
        P2_U3136) );
  AOI22_X1 U22446 ( .A1(n19434), .A2(n19551), .B1(n13769), .B2(n19433), .ZN(
        n19419) );
  AOI22_X1 U22447 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19435), .B1(
        n19470), .B2(n19552), .ZN(n19418) );
  OAI211_X1 U22448 ( .C1(n19555), .C2(n19438), .A(n19419), .B(n19418), .ZN(
        P2_U3137) );
  AOI22_X1 U22449 ( .A1(n19434), .A2(n19557), .B1(n19556), .B2(n19433), .ZN(
        n19421) );
  AOI22_X1 U22450 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19435), .B1(
        n19427), .B2(n19455), .ZN(n19420) );
  OAI211_X1 U22451 ( .C1(n19458), .C2(n19430), .A(n19421), .B(n19420), .ZN(
        P2_U3138) );
  AOI22_X1 U22452 ( .A1(n19434), .A2(n19563), .B1(n19562), .B2(n19433), .ZN(
        n19423) );
  AOI22_X1 U22453 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19435), .B1(
        n19470), .B2(n19515), .ZN(n19422) );
  OAI211_X1 U22454 ( .C1(n19424), .C2(n19438), .A(n19423), .B(n19422), .ZN(
        P2_U3139) );
  AOI22_X1 U22455 ( .A1(n19434), .A2(n19569), .B1(n19568), .B2(n19433), .ZN(
        n19426) );
  AOI22_X1 U22456 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19435), .B1(
        n19427), .B2(n19570), .ZN(n19425) );
  OAI211_X1 U22457 ( .C1(n19573), .C2(n19430), .A(n19426), .B(n19425), .ZN(
        P2_U3140) );
  AOI22_X1 U22458 ( .A1(n19434), .A2(n21082), .B1(n21078), .B2(n19433), .ZN(
        n19429) );
  AOI22_X1 U22459 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19435), .B1(
        n19427), .B2(n21080), .ZN(n19428) );
  OAI211_X1 U22460 ( .C1(n21087), .C2(n19430), .A(n19429), .B(n19428), .ZN(
        P2_U3141) );
  AOI22_X1 U22461 ( .A1(n19434), .A2(n19579), .B1(n19578), .B2(n19433), .ZN(
        n19432) );
  AOI22_X1 U22462 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19435), .B1(
        n19470), .B2(n19580), .ZN(n19431) );
  OAI211_X1 U22463 ( .C1(n19583), .C2(n19438), .A(n19432), .B(n19431), .ZN(
        P2_U3142) );
  AOI22_X1 U22464 ( .A1(n19434), .A2(n19586), .B1(n19584), .B2(n19433), .ZN(
        n19437) );
  AOI22_X1 U22465 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19435), .B1(
        n19470), .B2(n19588), .ZN(n19436) );
  OAI211_X1 U22466 ( .C1(n19594), .C2(n19438), .A(n19437), .B(n19436), .ZN(
        P2_U3143) );
  NAND3_X1 U22467 ( .A1(n19445), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        n19546), .ZN(n19444) );
  NOR2_X1 U22468 ( .A1(n19442), .A2(n19441), .ZN(n19468) );
  NOR3_X1 U22469 ( .A1(n19443), .A2(n19468), .A3(n19732), .ZN(n19446) );
  AOI21_X1 U22470 ( .B1(n19732), .B2(n19444), .A(n19446), .ZN(n19469) );
  AOI22_X1 U22471 ( .A1(n19469), .A2(n19540), .B1(n19539), .B2(n19468), .ZN(
        n19452) );
  OAI21_X1 U22472 ( .B1(n19503), .B2(n19470), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19449) );
  NAND2_X1 U22473 ( .A1(n19445), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19448) );
  AOI211_X1 U22474 ( .C1(n19449), .C2(n19448), .A(n19447), .B(n19446), .ZN(
        n19450) );
  AOI22_X1 U22475 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19471), .B1(
        n19470), .B2(n19547), .ZN(n19451) );
  OAI211_X1 U22476 ( .C1(n19550), .C2(n19499), .A(n19452), .B(n19451), .ZN(
        P2_U3144) );
  AOI22_X1 U22477 ( .A1(n19469), .A2(n19551), .B1(n13769), .B2(n19468), .ZN(
        n19454) );
  AOI22_X1 U22478 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19471), .B1(
        n19470), .B2(n19512), .ZN(n19453) );
  OAI211_X1 U22479 ( .C1(n19488), .C2(n19499), .A(n19454), .B(n19453), .ZN(
        P2_U3145) );
  AOI22_X1 U22480 ( .A1(n19469), .A2(n19557), .B1(n19556), .B2(n19468), .ZN(
        n19457) );
  AOI22_X1 U22481 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19471), .B1(
        n19470), .B2(n19455), .ZN(n19456) );
  OAI211_X1 U22482 ( .C1(n19458), .C2(n19499), .A(n19457), .B(n19456), .ZN(
        P2_U3146) );
  AOI22_X1 U22483 ( .A1(n19469), .A2(n19563), .B1(n19562), .B2(n19468), .ZN(
        n19460) );
  AOI22_X1 U22484 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19471), .B1(
        n19470), .B2(n19564), .ZN(n19459) );
  OAI211_X1 U22485 ( .C1(n19567), .C2(n19499), .A(n19460), .B(n19459), .ZN(
        P2_U3147) );
  AOI22_X1 U22486 ( .A1(n19469), .A2(n19569), .B1(n19568), .B2(n19468), .ZN(
        n19462) );
  AOI22_X1 U22487 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19471), .B1(
        n19470), .B2(n19570), .ZN(n19461) );
  OAI211_X1 U22488 ( .C1(n19573), .C2(n19499), .A(n19462), .B(n19461), .ZN(
        P2_U3148) );
  AOI22_X1 U22489 ( .A1(n19469), .A2(n21082), .B1(n21078), .B2(n19468), .ZN(
        n19464) );
  AOI22_X1 U22490 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19471), .B1(
        n19470), .B2(n21080), .ZN(n19463) );
  OAI211_X1 U22491 ( .C1(n21087), .C2(n19499), .A(n19464), .B(n19463), .ZN(
        P2_U3149) );
  AOI22_X1 U22492 ( .A1(n19469), .A2(n19579), .B1(n19578), .B2(n19468), .ZN(
        n19466) );
  AOI22_X1 U22493 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19471), .B1(
        n19470), .B2(n19524), .ZN(n19465) );
  OAI211_X1 U22494 ( .C1(n19467), .C2(n19499), .A(n19466), .B(n19465), .ZN(
        P2_U3150) );
  AOI22_X1 U22495 ( .A1(n19469), .A2(n19586), .B1(n19584), .B2(n19468), .ZN(
        n19473) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19471), .B1(
        n19470), .B2(n19502), .ZN(n19472) );
  OAI211_X1 U22497 ( .C1(n19507), .C2(n19499), .A(n19473), .B(n19472), .ZN(
        P2_U3151) );
  NAND2_X1 U22498 ( .A1(n19474), .A2(n19708), .ZN(n19478) );
  NOR2_X1 U22499 ( .A1(n19715), .A2(n19478), .ZN(n19500) );
  INV_X1 U22500 ( .A(n19481), .ZN(n19476) );
  AOI211_X2 U22501 ( .C1(n19478), .C2(n19732), .A(n19477), .B(n19476), .ZN(
        n19501) );
  AOI22_X1 U22502 ( .A1(n19501), .A2(n19540), .B1(n19539), .B2(n19500), .ZN(
        n19485) );
  OAI21_X1 U22503 ( .B1(n19480), .B2(n19479), .A(n19478), .ZN(n19482) );
  AND2_X1 U22504 ( .A1(n19482), .A2(n19481), .ZN(n19483) );
  OAI211_X1 U22505 ( .C1(n19500), .C2(n19546), .A(n19545), .B(n19483), .ZN(
        n19504) );
  AOI22_X1 U22506 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19504), .B1(
        n19503), .B2(n19547), .ZN(n19484) );
  OAI211_X1 U22507 ( .C1(n19550), .C2(n19535), .A(n19485), .B(n19484), .ZN(
        P2_U3152) );
  AOI22_X1 U22508 ( .A1(n19501), .A2(n19551), .B1(n13769), .B2(n19500), .ZN(
        n19487) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19504), .B1(
        n19503), .B2(n19512), .ZN(n19486) );
  OAI211_X1 U22510 ( .C1(n19488), .C2(n19535), .A(n19487), .B(n19486), .ZN(
        P2_U3153) );
  AOI22_X1 U22511 ( .A1(n19501), .A2(n19557), .B1(n19556), .B2(n19500), .ZN(
        n19490) );
  AOI22_X1 U22512 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19504), .B1(
        n19525), .B2(n19558), .ZN(n19489) );
  OAI211_X1 U22513 ( .C1(n19561), .C2(n19499), .A(n19490), .B(n19489), .ZN(
        P2_U3154) );
  AOI22_X1 U22514 ( .A1(n19501), .A2(n19563), .B1(n19562), .B2(n19500), .ZN(
        n19492) );
  AOI22_X1 U22515 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19504), .B1(
        n19503), .B2(n19564), .ZN(n19491) );
  OAI211_X1 U22516 ( .C1(n19567), .C2(n19535), .A(n19492), .B(n19491), .ZN(
        P2_U3155) );
  AOI22_X1 U22517 ( .A1(n19501), .A2(n19569), .B1(n19568), .B2(n19500), .ZN(
        n19494) );
  AOI22_X1 U22518 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19504), .B1(
        n19503), .B2(n19570), .ZN(n19493) );
  OAI211_X1 U22519 ( .C1(n19573), .C2(n19535), .A(n19494), .B(n19493), .ZN(
        P2_U3156) );
  AOI22_X1 U22520 ( .A1(n19501), .A2(n21082), .B1(n21078), .B2(n19500), .ZN(
        n19496) );
  AOI22_X1 U22521 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19504), .B1(
        n19503), .B2(n21080), .ZN(n19495) );
  OAI211_X1 U22522 ( .C1(n21087), .C2(n19535), .A(n19496), .B(n19495), .ZN(
        P2_U3157) );
  AOI22_X1 U22523 ( .A1(n19501), .A2(n19579), .B1(n19578), .B2(n19500), .ZN(
        n19498) );
  AOI22_X1 U22524 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19504), .B1(
        n19525), .B2(n19580), .ZN(n19497) );
  OAI211_X1 U22525 ( .C1(n19583), .C2(n19499), .A(n19498), .B(n19497), .ZN(
        P2_U3158) );
  AOI22_X1 U22526 ( .A1(n19501), .A2(n19586), .B1(n19584), .B2(n19500), .ZN(
        n19506) );
  AOI22_X1 U22527 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19504), .B1(
        n19503), .B2(n19502), .ZN(n19505) );
  OAI211_X1 U22528 ( .C1(n19507), .C2(n19535), .A(n19506), .B(n19505), .ZN(
        P2_U3159) );
  AOI22_X1 U22529 ( .A1(n19547), .A2(n19525), .B1(n19530), .B2(n19539), .ZN(
        n19510) );
  AOI22_X1 U22530 ( .A1(n19540), .A2(n19531), .B1(n19574), .B2(n19508), .ZN(
        n19509) );
  OAI211_X1 U22531 ( .C1(n19529), .C2(n19511), .A(n19510), .B(n19509), .ZN(
        P2_U3160) );
  AOI22_X1 U22532 ( .A1(n19552), .A2(n19574), .B1(n19530), .B2(n13769), .ZN(
        n19514) );
  AOI22_X1 U22533 ( .A1(n19551), .A2(n19531), .B1(n19525), .B2(n19512), .ZN(
        n19513) );
  OAI211_X1 U22534 ( .C1(n19529), .C2(n10325), .A(n19514), .B(n19513), .ZN(
        P2_U3161) );
  INV_X1 U22535 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n19518) );
  AOI22_X1 U22536 ( .A1(n19564), .A2(n19525), .B1(n19530), .B2(n19562), .ZN(
        n19517) );
  AOI22_X1 U22537 ( .A1(n19563), .A2(n19531), .B1(n19574), .B2(n19515), .ZN(
        n19516) );
  OAI211_X1 U22538 ( .C1(n19529), .C2(n19518), .A(n19517), .B(n19516), .ZN(
        P2_U3163) );
  AOI22_X1 U22539 ( .A1(n19519), .A2(n19574), .B1(n19530), .B2(n19568), .ZN(
        n19521) );
  AOI22_X1 U22540 ( .A1(n19569), .A2(n19531), .B1(n19525), .B2(n19570), .ZN(
        n19520) );
  OAI211_X1 U22541 ( .C1(n19529), .C2(n20817), .A(n19521), .B(n19520), .ZN(
        P2_U3164) );
  AOI22_X1 U22542 ( .A1(n21080), .A2(n19525), .B1(n19530), .B2(n21078), .ZN(
        n19523) );
  AOI22_X1 U22543 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19532), .B1(
        n21082), .B2(n19531), .ZN(n19522) );
  OAI211_X1 U22544 ( .C1(n21087), .C2(n19593), .A(n19523), .B(n19522), .ZN(
        P2_U3165) );
  INV_X1 U22545 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n19528) );
  AOI22_X1 U22546 ( .A1(n19580), .A2(n19574), .B1(n19530), .B2(n19578), .ZN(
        n19527) );
  AOI22_X1 U22547 ( .A1(n19579), .A2(n19531), .B1(n19525), .B2(n19524), .ZN(
        n19526) );
  OAI211_X1 U22548 ( .C1(n19529), .C2(n19528), .A(n19527), .B(n19526), .ZN(
        P2_U3166) );
  AOI22_X1 U22549 ( .A1(n19588), .A2(n19574), .B1(n19530), .B2(n19584), .ZN(
        n19534) );
  AOI22_X1 U22550 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19532), .B1(
        n19586), .B2(n19531), .ZN(n19533) );
  OAI211_X1 U22551 ( .C1(n19594), .C2(n19535), .A(n19534), .B(n19533), .ZN(
        P2_U3167) );
  INV_X1 U22552 ( .A(n19542), .ZN(n19537) );
  AOI21_X1 U22553 ( .B1(n19546), .B2(n19537), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19538) );
  AOI22_X1 U22554 ( .A1(n19587), .A2(n19540), .B1(n19585), .B2(n19539), .ZN(
        n19549) );
  NAND2_X1 U22555 ( .A1(n19681), .A2(n19541), .ZN(n19543) );
  AOI21_X1 U22556 ( .B1(n19543), .B2(n19542), .A(n9823), .ZN(n19544) );
  OAI211_X1 U22557 ( .C1(n19585), .C2(n19546), .A(n19545), .B(n19544), .ZN(
        n19590) );
  AOI22_X1 U22558 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19590), .B1(
        n19574), .B2(n19547), .ZN(n19548) );
  OAI211_X1 U22559 ( .C1(n19550), .C2(n19577), .A(n19549), .B(n19548), .ZN(
        P2_U3168) );
  AOI22_X1 U22560 ( .A1(n19587), .A2(n19551), .B1(n19585), .B2(n13769), .ZN(
        n19554) );
  AOI22_X1 U22561 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19590), .B1(
        n19589), .B2(n19552), .ZN(n19553) );
  OAI211_X1 U22562 ( .C1(n19555), .C2(n19593), .A(n19554), .B(n19553), .ZN(
        P2_U3169) );
  AOI22_X1 U22563 ( .A1(n19587), .A2(n19557), .B1(n19585), .B2(n19556), .ZN(
        n19560) );
  AOI22_X1 U22564 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19590), .B1(
        n19589), .B2(n19558), .ZN(n19559) );
  OAI211_X1 U22565 ( .C1(n19561), .C2(n19593), .A(n19560), .B(n19559), .ZN(
        P2_U3170) );
  AOI22_X1 U22566 ( .A1(n19587), .A2(n19563), .B1(n19585), .B2(n19562), .ZN(
        n19566) );
  AOI22_X1 U22567 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19590), .B1(
        n19574), .B2(n19564), .ZN(n19565) );
  OAI211_X1 U22568 ( .C1(n19567), .C2(n19577), .A(n19566), .B(n19565), .ZN(
        P2_U3171) );
  AOI22_X1 U22569 ( .A1(n19587), .A2(n19569), .B1(n19585), .B2(n19568), .ZN(
        n19572) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19590), .B1(
        n19574), .B2(n19570), .ZN(n19571) );
  OAI211_X1 U22571 ( .C1(n19573), .C2(n19577), .A(n19572), .B(n19571), .ZN(
        P2_U3172) );
  AOI22_X1 U22572 ( .A1(n19587), .A2(n21082), .B1(n19585), .B2(n21078), .ZN(
        n19576) );
  AOI22_X1 U22573 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19590), .B1(
        n19574), .B2(n21080), .ZN(n19575) );
  OAI211_X1 U22574 ( .C1(n21087), .C2(n19577), .A(n19576), .B(n19575), .ZN(
        P2_U3173) );
  AOI22_X1 U22575 ( .A1(n19587), .A2(n19579), .B1(n19585), .B2(n19578), .ZN(
        n19582) );
  AOI22_X1 U22576 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19590), .B1(
        n19589), .B2(n19580), .ZN(n19581) );
  OAI211_X1 U22577 ( .C1(n19583), .C2(n19593), .A(n19582), .B(n19581), .ZN(
        P2_U3174) );
  AOI22_X1 U22578 ( .A1(n19587), .A2(n19586), .B1(n19585), .B2(n19584), .ZN(
        n19592) );
  AOI22_X1 U22579 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19590), .B1(
        n19589), .B2(n19588), .ZN(n19591) );
  OAI211_X1 U22580 ( .C1(n19594), .C2(n19593), .A(n19592), .B(n19591), .ZN(
        P2_U3175) );
  AOI21_X1 U22581 ( .B1(n19596), .B2(n19595), .A(n19731), .ZN(n19604) );
  AOI211_X1 U22582 ( .C1(n19599), .C2(n19598), .A(n19726), .B(n19597), .ZN(
        n19600) );
  INV_X1 U22583 ( .A(n19600), .ZN(n19601) );
  OAI211_X1 U22584 ( .C1(n19604), .C2(n19603), .A(n19602), .B(n19601), .ZN(
        P2_U3177) );
  INV_X1 U22585 ( .A(n19679), .ZN(n19605) );
  AND2_X1 U22586 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19605), .ZN(
        P2_U3179) );
  AND2_X1 U22587 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19605), .ZN(
        P2_U3180) );
  AND2_X1 U22588 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19605), .ZN(
        P2_U3181) );
  AND2_X1 U22589 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19605), .ZN(
        P2_U3182) );
  AND2_X1 U22590 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19605), .ZN(
        P2_U3183) );
  AND2_X1 U22591 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19605), .ZN(
        P2_U3184) );
  AND2_X1 U22592 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19605), .ZN(
        P2_U3185) );
  AND2_X1 U22593 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19605), .ZN(
        P2_U3186) );
  AND2_X1 U22594 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19605), .ZN(
        P2_U3187) );
  AND2_X1 U22595 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19605), .ZN(
        P2_U3188) );
  AND2_X1 U22596 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19605), .ZN(
        P2_U3189) );
  AND2_X1 U22597 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19605), .ZN(
        P2_U3190) );
  AND2_X1 U22598 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19605), .ZN(
        P2_U3191) );
  AND2_X1 U22599 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19605), .ZN(
        P2_U3192) );
  AND2_X1 U22600 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19605), .ZN(
        P2_U3193) );
  AND2_X1 U22601 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19605), .ZN(
        P2_U3194) );
  AND2_X1 U22602 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19605), .ZN(
        P2_U3195) );
  AND2_X1 U22603 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19605), .ZN(
        P2_U3196) );
  AND2_X1 U22604 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19605), .ZN(
        P2_U3197) );
  AND2_X1 U22605 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19605), .ZN(
        P2_U3198) );
  INV_X1 U22606 ( .A(P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20887) );
  NOR2_X1 U22607 ( .A1(n20887), .A2(n19679), .ZN(P2_U3199) );
  AND2_X1 U22608 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19605), .ZN(
        P2_U3200) );
  NOR2_X1 U22609 ( .A1(n21064), .A2(n19679), .ZN(P2_U3201) );
  AND2_X1 U22610 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19605), .ZN(P2_U3202) );
  AND2_X1 U22611 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19605), .ZN(P2_U3203) );
  AND2_X1 U22612 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19605), .ZN(P2_U3204) );
  AND2_X1 U22613 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19605), .ZN(P2_U3205) );
  AND2_X1 U22614 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19605), .ZN(P2_U3206) );
  AND2_X1 U22615 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19605), .ZN(P2_U3207) );
  NOR2_X1 U22616 ( .A1(n21018), .A2(n19679), .ZN(P2_U3208) );
  NOR2_X1 U22617 ( .A1(n20989), .A2(n19726), .ZN(n19615) );
  INV_X1 U22618 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19746) );
  OR3_X1 U22619 ( .A1(n19615), .A2(n19746), .A3(n19606), .ZN(n19608) );
  INV_X2 U22620 ( .A(n19748), .ZN(n19665) );
  AOI211_X1 U22621 ( .C1(n20668), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n19616), .B(n19665), .ZN(n19607) );
  NOR3_X1 U22622 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n20654), .ZN(n19620) );
  AOI211_X1 U22623 ( .C1(n19621), .C2(n19608), .A(n19607), .B(n19620), .ZN(
        n19609) );
  INV_X1 U22624 ( .A(n19609), .ZN(P2_U3209) );
  AOI21_X1 U22625 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20668), .A(n19621), 
        .ZN(n19613) );
  NOR3_X1 U22626 ( .A1(n19613), .A2(n19746), .A3(n19606), .ZN(n19610) );
  NOR2_X1 U22627 ( .A1(n19610), .A2(n19615), .ZN(n19611) );
  OAI211_X1 U22628 ( .C1(n20668), .C2(n19612), .A(n19611), .B(n19739), .ZN(
        P2_U3210) );
  NOR2_X1 U22629 ( .A1(n20989), .A2(n19621), .ZN(n19614) );
  AOI21_X1 U22630 ( .B1(n19733), .B2(n19614), .A(n19613), .ZN(n19619) );
  AOI22_X1 U22631 ( .A1(n19616), .A2(n19746), .B1(n19615), .B2(n20654), .ZN(
        n19618) );
  OAI21_X1 U22632 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n19617) );
  OAI22_X1 U22633 ( .A1(n19620), .A2(n19619), .B1(n19618), .B2(n19617), .ZN(
        P2_U3211) );
  OAI222_X1 U22634 ( .A1(n19672), .A2(n19624), .B1(n19623), .B2(n19665), .C1(
        n19622), .C2(n19669), .ZN(P2_U3212) );
  OAI222_X1 U22635 ( .A1(n19672), .A2(n10914), .B1(n19625), .B2(n19665), .C1(
        n19624), .C2(n19669), .ZN(P2_U3213) );
  OAI222_X1 U22636 ( .A1(n19672), .A2(n10920), .B1(n19626), .B2(n19665), .C1(
        n10914), .C2(n19669), .ZN(P2_U3214) );
  INV_X1 U22637 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19628) );
  OAI222_X1 U22638 ( .A1(n19672), .A2(n19628), .B1(n19627), .B2(n19665), .C1(
        n10920), .C2(n19669), .ZN(P2_U3215) );
  OAI222_X1 U22639 ( .A1(n19672), .A2(n19630), .B1(n19629), .B2(n19665), .C1(
        n19628), .C2(n19669), .ZN(P2_U3216) );
  OAI222_X1 U22640 ( .A1(n19672), .A2(n19632), .B1(n19631), .B2(n19665), .C1(
        n19630), .C2(n19669), .ZN(P2_U3217) );
  OAI222_X1 U22641 ( .A1(n19672), .A2(n10939), .B1(n19633), .B2(n19665), .C1(
        n19632), .C2(n19669), .ZN(P2_U3218) );
  OAI222_X1 U22642 ( .A1(n19672), .A2(n10963), .B1(n19634), .B2(n19665), .C1(
        n10939), .C2(n19669), .ZN(P2_U3219) );
  OAI222_X1 U22643 ( .A1(n19672), .A2(n10966), .B1(n19635), .B2(n19665), .C1(
        n10963), .C2(n19669), .ZN(P2_U3220) );
  OAI222_X1 U22644 ( .A1(n19672), .A2(n10990), .B1(n19636), .B2(n19665), .C1(
        n10966), .C2(n19669), .ZN(P2_U3221) );
  OAI222_X1 U22645 ( .A1(n19672), .A2(n10994), .B1(n19637), .B2(n19665), .C1(
        n10990), .C2(n19669), .ZN(P2_U3222) );
  OAI222_X1 U22646 ( .A1(n19672), .A2(n19639), .B1(n19638), .B2(n19665), .C1(
        n10994), .C2(n19669), .ZN(P2_U3223) );
  OAI222_X1 U22647 ( .A1(n19672), .A2(n11020), .B1(n19640), .B2(n19665), .C1(
        n19639), .C2(n19669), .ZN(P2_U3224) );
  OAI222_X1 U22648 ( .A1(n19672), .A2(n19642), .B1(n19641), .B2(n19665), .C1(
        n11020), .C2(n19669), .ZN(P2_U3225) );
  OAI222_X1 U22649 ( .A1(n19672), .A2(n15346), .B1(n19643), .B2(n19665), .C1(
        n19642), .C2(n19669), .ZN(P2_U3226) );
  OAI222_X1 U22650 ( .A1(n19672), .A2(n19644), .B1(n21063), .B2(n19665), .C1(
        n15346), .C2(n19669), .ZN(P2_U3227) );
  OAI222_X1 U22651 ( .A1(n19672), .A2(n19646), .B1(n19645), .B2(n19665), .C1(
        n19644), .C2(n19669), .ZN(P2_U3228) );
  OAI222_X1 U22652 ( .A1(n19672), .A2(n19648), .B1(n19647), .B2(n19665), .C1(
        n19646), .C2(n19669), .ZN(P2_U3229) );
  INV_X1 U22653 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19650) );
  OAI222_X1 U22654 ( .A1(n19672), .A2(n19650), .B1(n19649), .B2(n19665), .C1(
        n19648), .C2(n19669), .ZN(P2_U3230) );
  OAI222_X1 U22655 ( .A1(n19672), .A2(n19652), .B1(n19651), .B2(n19665), .C1(
        n19650), .C2(n19669), .ZN(P2_U3231) );
  OAI222_X1 U22656 ( .A1(n19672), .A2(n11059), .B1(n19653), .B2(n19665), .C1(
        n19652), .C2(n19669), .ZN(P2_U3232) );
  OAI222_X1 U22657 ( .A1(n19672), .A2(n19655), .B1(n19654), .B2(n19665), .C1(
        n11059), .C2(n19669), .ZN(P2_U3233) );
  OAI222_X1 U22658 ( .A1(n19672), .A2(n19657), .B1(n19656), .B2(n19665), .C1(
        n19655), .C2(n19669), .ZN(P2_U3234) );
  INV_X1 U22659 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19659) );
  OAI222_X1 U22660 ( .A1(n19672), .A2(n19659), .B1(n19658), .B2(n19665), .C1(
        n19657), .C2(n19669), .ZN(P2_U3235) );
  OAI222_X1 U22661 ( .A1(n19672), .A2(n19661), .B1(n19660), .B2(n19665), .C1(
        n19659), .C2(n19669), .ZN(P2_U3236) );
  OAI222_X1 U22662 ( .A1(n19672), .A2(n19664), .B1(n19662), .B2(n19665), .C1(
        n19661), .C2(n19669), .ZN(P2_U3237) );
  OAI222_X1 U22663 ( .A1(n19669), .A2(n19664), .B1(n19663), .B2(n19665), .C1(
        n15192), .C2(n19672), .ZN(P2_U3238) );
  OAI222_X1 U22664 ( .A1(n19672), .A2(n19667), .B1(n19666), .B2(n19665), .C1(
        n15192), .C2(n19669), .ZN(P2_U3239) );
  OAI222_X1 U22665 ( .A1(n19672), .A2(n12927), .B1(n19668), .B2(n19665), .C1(
        n19667), .C2(n19669), .ZN(P2_U3240) );
  INV_X1 U22666 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19671) );
  OAI222_X1 U22667 ( .A1(n19672), .A2(n19671), .B1(n19670), .B2(n19665), .C1(
        n12927), .C2(n19669), .ZN(P2_U3241) );
  OAI22_X1 U22668 ( .A1(n19748), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19665), .ZN(n19673) );
  INV_X1 U22669 ( .A(n19673), .ZN(P2_U3585) );
  MUX2_X1 U22670 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19748), .Z(P2_U3586) );
  OAI22_X1 U22671 ( .A1(n19748), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19665), .ZN(n19674) );
  INV_X1 U22672 ( .A(n19674), .ZN(P2_U3587) );
  OAI22_X1 U22673 ( .A1(n19748), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19665), .ZN(n19675) );
  INV_X1 U22674 ( .A(n19675), .ZN(P2_U3588) );
  OAI21_X1 U22675 ( .B1(n19679), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19677), 
        .ZN(n19676) );
  INV_X1 U22676 ( .A(n19676), .ZN(P2_U3591) );
  OAI21_X1 U22677 ( .B1(n19679), .B2(n19678), .A(n19677), .ZN(P2_U3592) );
  NOR2_X1 U22678 ( .A1(n19680), .A2(n19685), .ZN(n19693) );
  INV_X1 U22679 ( .A(n19701), .ZN(n19730) );
  AOI21_X1 U22680 ( .B1(n19702), .B2(n19699), .A(n19730), .ZN(n19691) );
  OAI21_X1 U22681 ( .B1(n19693), .B2(n19691), .A(n19681), .ZN(n19684) );
  NAND2_X1 U22682 ( .A1(n19682), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19683) );
  OAI211_X1 U22683 ( .C1(n19686), .C2(n19685), .A(n19684), .B(n19683), .ZN(
        n19687) );
  INV_X1 U22684 ( .A(n19687), .ZN(n19688) );
  AOI22_X1 U22685 ( .A1(n19713), .A2(n19689), .B1(n19688), .B2(n19714), .ZN(
        P2_U3602) );
  AOI22_X1 U22686 ( .A1(n19692), .A2(n19691), .B1(n19690), .B2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19695) );
  NOR2_X1 U22687 ( .A1(n19713), .A2(n19693), .ZN(n19694) );
  AOI22_X1 U22688 ( .A1(n19696), .A2(n19713), .B1(n19695), .B2(n19694), .ZN(
        P2_U3603) );
  NAND3_X1 U22689 ( .A1(n19698), .A2(n19697), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19704) );
  INV_X1 U22690 ( .A(n19699), .ZN(n19700) );
  NAND3_X1 U22691 ( .A1(n19702), .A2(n19701), .A3(n19700), .ZN(n19703) );
  NAND2_X1 U22692 ( .A1(n19704), .A2(n19703), .ZN(n19705) );
  AOI21_X1 U22693 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19706), .A(n19705), 
        .ZN(n19707) );
  AOI22_X1 U22694 ( .A1(n19713), .A2(n19708), .B1(n19707), .B2(n19714), .ZN(
        P2_U3604) );
  OAI22_X1 U22695 ( .A1(n19710), .A2(n19730), .B1(n19732), .B2(n19709), .ZN(
        n19711) );
  AOI21_X1 U22696 ( .B1(n19715), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19711), 
        .ZN(n19712) );
  OAI22_X1 U22697 ( .A1(n19715), .A2(n19714), .B1(n19713), .B2(n19712), .ZN(
        P2_U3605) );
  INV_X1 U22698 ( .A(P2_READREQUEST_REG_SCAN_IN), .ZN(n20915) );
  OAI22_X1 U22699 ( .A1(n19748), .A2(n20915), .B1(P2_W_R_N_REG_SCAN_IN), .B2(
        n19665), .ZN(n19716) );
  INV_X1 U22700 ( .A(n19716), .ZN(P2_U3608) );
  INV_X1 U22701 ( .A(n19717), .ZN(n19721) );
  AOI22_X1 U22702 ( .A1(n19721), .A2(n19720), .B1(n19719), .B2(n19718), .ZN(
        n19722) );
  NAND2_X1 U22703 ( .A1(n19723), .A2(n19722), .ZN(n19725) );
  MUX2_X1 U22704 ( .A(P2_MORE_REG_SCAN_IN), .B(n19725), .S(n19724), .Z(
        P2_U3609) );
  NAND4_X1 U22705 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .A3(n19727), .A4(n19726), .ZN(n19728) );
  OAI211_X1 U22706 ( .C1(n19731), .C2(n19730), .A(n19729), .B(n19728), .ZN(
        n19747) );
  NOR2_X1 U22707 ( .A1(n19733), .A2(n19732), .ZN(n19743) );
  INV_X1 U22708 ( .A(n19734), .ZN(n19736) );
  NAND2_X1 U22709 ( .A1(n19736), .A2(n19735), .ZN(n19741) );
  OAI211_X1 U22710 ( .C1(n19739), .C2(n19738), .A(n9776), .B(n19737), .ZN(
        n19740) );
  OAI211_X1 U22711 ( .C1(n19743), .C2(n19742), .A(n19741), .B(n19740), .ZN(
        n19744) );
  NAND2_X1 U22712 ( .A1(n19747), .A2(n19744), .ZN(n19745) );
  OAI21_X1 U22713 ( .B1(n19747), .B2(n19746), .A(n19745), .ZN(P2_U3610) );
  OAI22_X1 U22714 ( .A1(n19748), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19665), .ZN(n19749) );
  INV_X1 U22715 ( .A(n19749), .ZN(P2_U3611) );
  INV_X1 U22716 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20663) );
  AOI21_X1 U22717 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20959), .A(n20663), 
        .ZN(n20666) );
  INV_X1 U22718 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19750) );
  AND2_X1 U22719 ( .A1(n20663), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20769) );
  AOI21_X1 U22720 ( .B1(n20666), .B2(n19750), .A(n20769), .ZN(P1_U2802) );
  OAI21_X1 U22721 ( .B1(n19752), .B2(n19751), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19753) );
  OAI21_X1 U22722 ( .B1(n19754), .B2(n15945), .A(n19753), .ZN(P1_U2803) );
  INV_X2 U22723 ( .A(n20769), .ZN(n20770) );
  NAND2_X1 U22724 ( .A1(n20959), .A2(n20663), .ZN(n20657) );
  INV_X1 U22725 ( .A(n20657), .ZN(n19756) );
  OAI21_X1 U22726 ( .B1(n19756), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20770), .ZN(
        n19755) );
  OAI21_X1 U22727 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20770), .A(n19755), 
        .ZN(P1_U2804) );
  NOR2_X1 U22728 ( .A1(n20666), .A2(n20769), .ZN(n20724) );
  OAI21_X1 U22729 ( .B1(BS16), .B2(n19756), .A(n20724), .ZN(n20722) );
  OAI21_X1 U22730 ( .B1(n20724), .B2(n20516), .A(n20722), .ZN(P1_U2805) );
  OAI21_X1 U22731 ( .B1(n19759), .B2(n19758), .A(n19757), .ZN(P1_U2806) );
  NOR4_X1 U22732 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19763) );
  NOR4_X1 U22733 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19762) );
  NOR4_X1 U22734 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19761) );
  NOR4_X1 U22735 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19760) );
  NAND4_X1 U22736 ( .A1(n19763), .A2(n19762), .A3(n19761), .A4(n19760), .ZN(
        n19769) );
  NOR4_X1 U22737 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n19767) );
  AOI211_X1 U22738 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_12__SCAN_IN), .B(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19766) );
  NOR4_X1 U22739 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19765) );
  NOR4_X1 U22740 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19764) );
  NAND4_X1 U22741 ( .A1(n19767), .A2(n19766), .A3(n19765), .A4(n19764), .ZN(
        n19768) );
  NOR2_X1 U22742 ( .A1(n19769), .A2(n19768), .ZN(n20752) );
  INV_X1 U22743 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21025) );
  NOR3_X1 U22744 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19771) );
  OAI21_X1 U22745 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19771), .A(n20752), .ZN(
        n19770) );
  OAI21_X1 U22746 ( .B1(n20752), .B2(n21025), .A(n19770), .ZN(P1_U2807) );
  INV_X1 U22747 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20723) );
  AOI21_X1 U22748 ( .B1(n20748), .B2(n20723), .A(n19771), .ZN(n19772) );
  INV_X1 U22749 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21035) );
  INV_X1 U22750 ( .A(n20752), .ZN(n20755) );
  AOI22_X1 U22751 ( .A1(n20752), .A2(n19772), .B1(n21035), .B2(n20755), .ZN(
        P1_U2808) );
  OAI21_X1 U22752 ( .B1(n19774), .B2(n19845), .A(n19773), .ZN(n19847) );
  AOI21_X1 U22753 ( .B1(n19816), .B2(n19775), .A(n19847), .ZN(n19798) );
  NOR2_X1 U22754 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19775), .ZN(n19781) );
  AOI22_X1 U22755 ( .A1(n19776), .A2(n19863), .B1(n19837), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n19778) );
  OAI211_X1 U22756 ( .C1(n19840), .C2(n19779), .A(n19778), .B(n19777), .ZN(
        n19780) );
  AOI21_X1 U22757 ( .B1(n19781), .B2(n19826), .A(n19780), .ZN(n19786) );
  INV_X1 U22758 ( .A(n19782), .ZN(n19784) );
  AOI22_X1 U22759 ( .A1(n19784), .A2(n19821), .B1(n19865), .B2(n19783), .ZN(
        n19785) );
  OAI211_X1 U22760 ( .C1(n19798), .C2(n14008), .A(n19786), .B(n19785), .ZN(
        P1_U2831) );
  NAND3_X1 U22761 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n19787) );
  NOR2_X1 U22762 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n19787), .ZN(n19788) );
  AOI22_X1 U22763 ( .A1(n19826), .A2(n19788), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n19837), .ZN(n19789) );
  OAI21_X1 U22764 ( .B1(n19791), .B2(n19790), .A(n19789), .ZN(n19792) );
  AOI211_X1 U22765 ( .C1(n19858), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n19836), .B(n19792), .ZN(n19797) );
  INV_X1 U22766 ( .A(n19793), .ZN(n19794) );
  AOI22_X1 U22767 ( .A1(n19795), .A2(n19821), .B1(n19865), .B2(n19794), .ZN(
        n19796) );
  OAI211_X1 U22768 ( .C1(n19798), .C2(n20681), .A(n19797), .B(n19796), .ZN(
        P1_U2832) );
  INV_X1 U22769 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20679) );
  INV_X1 U22770 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20677) );
  NOR2_X1 U22771 ( .A1(n20679), .A2(n20677), .ZN(n19805) );
  INV_X1 U22772 ( .A(n19805), .ZN(n19799) );
  NOR2_X1 U22773 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19799), .ZN(n19800) );
  AOI22_X1 U22774 ( .A1(n19863), .A2(n19801), .B1(n19826), .B2(n19800), .ZN(
        n19811) );
  INV_X1 U22775 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20923) );
  AOI21_X1 U22776 ( .B1(n19837), .B2(P1_EBX_REG_7__SCAN_IN), .A(n19836), .ZN(
        n19807) );
  NOR2_X1 U22777 ( .A1(n19803), .A2(n19802), .ZN(n19804) );
  NAND2_X1 U22778 ( .A1(n19805), .A2(n19804), .ZN(n19815) );
  NAND3_X1 U22779 ( .A1(n19816), .A2(P1_REIP_REG_7__SCAN_IN), .A3(n19815), 
        .ZN(n19806) );
  OAI211_X1 U22780 ( .C1(n19840), .C2(n20923), .A(n19807), .B(n19806), .ZN(
        n19808) );
  AOI21_X1 U22781 ( .B1(n19809), .B2(n19821), .A(n19808), .ZN(n19810) );
  OAI211_X1 U22782 ( .C1(n19812), .C2(n19851), .A(n19811), .B(n19810), .ZN(
        P1_U2833) );
  NOR2_X1 U22783 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20677), .ZN(n19813) );
  AOI22_X1 U22784 ( .A1(n19863), .A2(n19814), .B1(n19826), .B2(n19813), .ZN(
        n19824) );
  AOI21_X1 U22785 ( .B1(n19837), .B2(P1_EBX_REG_6__SCAN_IN), .A(n19836), .ZN(
        n19818) );
  NAND3_X1 U22786 ( .A1(n19816), .A2(P1_REIP_REG_6__SCAN_IN), .A3(n19815), 
        .ZN(n19817) );
  OAI211_X1 U22787 ( .C1(n19840), .C2(n19819), .A(n19818), .B(n19817), .ZN(
        n19820) );
  AOI21_X1 U22788 ( .B1(n19822), .B2(n19821), .A(n19820), .ZN(n19823) );
  OAI211_X1 U22789 ( .C1(n19825), .C2(n19851), .A(n19824), .B(n19823), .ZN(
        P1_U2834) );
  AOI22_X1 U22790 ( .A1(n19863), .A2(n19827), .B1(n19826), .B2(n20677), .ZN(
        n19834) );
  AOI21_X1 U22791 ( .B1(n19837), .B2(P1_EBX_REG_5__SCAN_IN), .A(n19836), .ZN(
        n19829) );
  NAND2_X1 U22792 ( .A1(n19847), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n19828) );
  OAI211_X1 U22793 ( .C1(n19840), .C2(n19830), .A(n19829), .B(n19828), .ZN(
        n19831) );
  AOI21_X1 U22794 ( .B1(n19832), .B2(n19867), .A(n19831), .ZN(n19833) );
  OAI211_X1 U22795 ( .C1(n19835), .C2(n19851), .A(n19834), .B(n19833), .ZN(
        P1_U2835) );
  AOI21_X1 U22796 ( .B1(n19837), .B2(P1_EBX_REG_4__SCAN_IN), .A(n19836), .ZN(
        n19838) );
  OAI21_X1 U22797 ( .B1(n19840), .B2(n19839), .A(n19838), .ZN(n19843) );
  NOR2_X1 U22798 ( .A1(n19841), .A2(n19860), .ZN(n19842) );
  AOI211_X1 U22799 ( .C1(n19863), .C2(n19946), .A(n19843), .B(n19842), .ZN(
        n19850) );
  OAI21_X1 U22800 ( .B1(n19845), .B2(n19844), .A(n20673), .ZN(n19846) );
  AOI22_X1 U22801 ( .A1(n19848), .A2(n19867), .B1(n19847), .B2(n19846), .ZN(
        n19849) );
  OAI211_X1 U22802 ( .C1(n19852), .C2(n19851), .A(n19850), .B(n19849), .ZN(
        P1_U2836) );
  INV_X1 U22803 ( .A(n20736), .ZN(n19861) );
  NAND4_X1 U22804 ( .A1(n19853), .A2(n13486), .A3(P1_REIP_REG_2__SCAN_IN), 
        .A4(P1_REIP_REG_1__SCAN_IN), .ZN(n19854) );
  OAI21_X1 U22805 ( .B1(n19856), .B2(n19855), .A(n19854), .ZN(n19857) );
  AOI21_X1 U22806 ( .B1(n19858), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n19857), .ZN(n19859) );
  OAI21_X1 U22807 ( .B1(n19861), .B2(n19860), .A(n19859), .ZN(n19862) );
  AOI21_X1 U22808 ( .B1(n19863), .B2(n19954), .A(n19862), .ZN(n19870) );
  INV_X1 U22809 ( .A(n19864), .ZN(n19868) );
  AOI22_X1 U22810 ( .A1(n19868), .A2(n19867), .B1(n19866), .B2(n19865), .ZN(
        n19869) );
  OAI211_X1 U22811 ( .C1(n13486), .C2(n19871), .A(n19870), .B(n19869), .ZN(
        P1_U2837) );
  INV_X1 U22812 ( .A(n19872), .ZN(n19876) );
  AOI22_X1 U22813 ( .A1(n19876), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n13187), .ZN(n19873) );
  OAI21_X1 U22814 ( .B1(n20987), .B2(n19888), .A(n19873), .ZN(P1_U2907) );
  INV_X1 U22815 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n20892) );
  AOI22_X1 U22816 ( .A1(n19876), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n13187), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n19874) );
  OAI21_X1 U22817 ( .B1(n20892), .B2(n19888), .A(n19874), .ZN(P1_U2911) );
  INV_X1 U22818 ( .A(P1_UWORD_REG_6__SCAN_IN), .ZN(n20873) );
  AOI22_X1 U22819 ( .A1(n19896), .A2(P1_DATAO_REG_22__SCAN_IN), .B1(n19876), 
        .B2(P1_EAX_REG_22__SCAN_IN), .ZN(n19875) );
  OAI21_X1 U22820 ( .B1(n20873), .B2(n19889), .A(n19875), .ZN(P1_U2914) );
  INV_X1 U22821 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n21015) );
  AOI22_X1 U22822 ( .A1(n19876), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n13187), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n19877) );
  OAI21_X1 U22823 ( .B1(n21015), .B2(n19888), .A(n19877), .ZN(P1_U2915) );
  AOI22_X1 U22824 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19878) );
  OAI21_X1 U22825 ( .B1(n13261), .B2(n19895), .A(n19878), .ZN(P1_U2921) );
  INV_X1 U22826 ( .A(P1_LWORD_REG_14__SCAN_IN), .ZN(n20886) );
  AOI22_X1 U22827 ( .A1(P1_EAX_REG_14__SCAN_IN), .A2(n19897), .B1(n19896), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19879) );
  OAI21_X1 U22828 ( .B1(n20886), .B2(n19889), .A(n19879), .ZN(P1_U2922) );
  AOI222_X1 U22829 ( .A1(n13187), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n19897), 
        .B2(P1_EAX_REG_13__SCAN_IN), .C1(P1_DATAO_REG_13__SCAN_IN), .C2(n19896), .ZN(n19880) );
  INV_X1 U22830 ( .A(n19880), .ZN(P1_U2923) );
  AOI22_X1 U22831 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19881) );
  OAI21_X1 U22832 ( .B1(n12045), .B2(n19895), .A(n19881), .ZN(P1_U2924) );
  AOI22_X1 U22833 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19882) );
  OAI21_X1 U22834 ( .B1(n14019), .B2(n19895), .A(n19882), .ZN(P1_U2925) );
  AOI22_X1 U22835 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19883) );
  OAI21_X1 U22836 ( .B1(n13974), .B2(n19895), .A(n19883), .ZN(P1_U2926) );
  AOI22_X1 U22837 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19884) );
  OAI21_X1 U22838 ( .B1(n13867), .B2(n19895), .A(n19884), .ZN(P1_U2927) );
  AOI22_X1 U22839 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19885) );
  OAI21_X1 U22840 ( .B1(n13842), .B2(n19895), .A(n19885), .ZN(P1_U2928) );
  AOI222_X1 U22841 ( .A1(n13187), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n19897), 
        .B2(P1_EAX_REG_7__SCAN_IN), .C1(P1_DATAO_REG_7__SCAN_IN), .C2(n19896), 
        .ZN(n19886) );
  INV_X1 U22842 ( .A(n19886), .ZN(P1_U2929) );
  AOI22_X1 U22843 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19887) );
  OAI21_X1 U22844 ( .B1(n11962), .B2(n19895), .A(n19887), .ZN(P1_U2930) );
  INV_X1 U22845 ( .A(P1_LWORD_REG_5__SCAN_IN), .ZN(n20854) );
  OAI222_X1 U22846 ( .A1(n19889), .A2(n20854), .B1(n19895), .B2(n13583), .C1(
        n20979), .C2(n19888), .ZN(P1_U2931) );
  AOI22_X1 U22847 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19890) );
  OAI21_X1 U22848 ( .B1(n19891), .B2(n19895), .A(n19890), .ZN(P1_U2932) );
  AOI22_X1 U22849 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19892) );
  OAI21_X1 U22850 ( .B1(n13440), .B2(n19895), .A(n19892), .ZN(P1_U2933) );
  AOI22_X1 U22851 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19893) );
  OAI21_X1 U22852 ( .B1(n11917), .B2(n19895), .A(n19893), .ZN(P1_U2934) );
  AOI22_X1 U22853 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n13187), .B1(n19896), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19894) );
  OAI21_X1 U22854 ( .B1(n11923), .B2(n19895), .A(n19894), .ZN(P1_U2935) );
  AOI222_X1 U22855 ( .A1(n13187), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n19897), 
        .B2(P1_EAX_REG_0__SCAN_IN), .C1(P1_DATAO_REG_0__SCAN_IN), .C2(n19896), 
        .ZN(n19898) );
  INV_X1 U22856 ( .A(n19898), .ZN(P1_U2936) );
  AOI22_X1 U22857 ( .A1(n19923), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n13470), .ZN(n19901) );
  INV_X1 U22858 ( .A(n19899), .ZN(n19900) );
  NAND2_X1 U22859 ( .A1(n19915), .A2(n19900), .ZN(n19917) );
  NAND2_X1 U22860 ( .A1(n19901), .A2(n19917), .ZN(P1_U2945) );
  AOI22_X1 U22861 ( .A1(n19923), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n13470), .ZN(n19904) );
  INV_X1 U22862 ( .A(n19902), .ZN(n19903) );
  NAND2_X1 U22863 ( .A1(n19915), .A2(n19903), .ZN(n19919) );
  NAND2_X1 U22864 ( .A1(n19904), .A2(n19919), .ZN(P1_U2946) );
  AOI22_X1 U22865 ( .A1(n19923), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n13470), .ZN(n19907) );
  INV_X1 U22866 ( .A(n19905), .ZN(n19906) );
  NAND2_X1 U22867 ( .A1(n19915), .A2(n19906), .ZN(n19921) );
  NAND2_X1 U22868 ( .A1(n19907), .A2(n19921), .ZN(P1_U2947) );
  AOI22_X1 U22869 ( .A1(n19923), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n13470), .ZN(n19910) );
  INV_X1 U22870 ( .A(n19908), .ZN(n19909) );
  NAND2_X1 U22871 ( .A1(n19915), .A2(n19909), .ZN(n19924) );
  NAND2_X1 U22872 ( .A1(n19910), .A2(n19924), .ZN(P1_U2948) );
  AOI22_X1 U22873 ( .A1(n19923), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n19928), .ZN(n19912) );
  NAND2_X1 U22874 ( .A1(n19915), .A2(n19911), .ZN(n19926) );
  NAND2_X1 U22875 ( .A1(n19912), .A2(n19926), .ZN(P1_U2949) );
  AOI22_X1 U22876 ( .A1(n19923), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n19928), .ZN(n19916) );
  INV_X1 U22877 ( .A(n19913), .ZN(n19914) );
  NAND2_X1 U22878 ( .A1(n19915), .A2(n19914), .ZN(n19929) );
  NAND2_X1 U22879 ( .A1(n19916), .A2(n19929), .ZN(P1_U2951) );
  AOI22_X1 U22880 ( .A1(n19923), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n19928), .ZN(n19918) );
  NAND2_X1 U22881 ( .A1(n19918), .A2(n19917), .ZN(P1_U2960) );
  AOI22_X1 U22882 ( .A1(n19923), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n19928), .ZN(n19920) );
  NAND2_X1 U22883 ( .A1(n19920), .A2(n19919), .ZN(P1_U2961) );
  AOI22_X1 U22884 ( .A1(n19923), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n19928), .ZN(n19922) );
  NAND2_X1 U22885 ( .A1(n19922), .A2(n19921), .ZN(P1_U2962) );
  AOI22_X1 U22886 ( .A1(n19923), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n19928), .ZN(n19925) );
  NAND2_X1 U22887 ( .A1(n19925), .A2(n19924), .ZN(P1_U2963) );
  AOI22_X1 U22888 ( .A1(n19923), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n19928), .ZN(n19927) );
  NAND2_X1 U22889 ( .A1(n19927), .A2(n19926), .ZN(P1_U2964) );
  AOI22_X1 U22890 ( .A1(n19923), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n19928), .ZN(n19930) );
  NAND2_X1 U22891 ( .A1(n19930), .A2(n19929), .ZN(P1_U2966) );
  INV_X1 U22892 ( .A(n19931), .ZN(n19934) );
  AOI21_X1 U22893 ( .B1(n19934), .B2(n19933), .A(n11361), .ZN(n19966) );
  OR2_X1 U22894 ( .A1(n19936), .A2(n19935), .ZN(n19937) );
  AOI22_X1 U22895 ( .A1(n19966), .A2(n19938), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19937), .ZN(n19940) );
  NAND2_X1 U22896 ( .A1(n19939), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n19971) );
  OAI211_X1 U22897 ( .C1(n19941), .C2(n19975), .A(n19940), .B(n19971), .ZN(
        P1_U2999) );
  OAI21_X1 U22898 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n19942), .ZN(n19952) );
  AOI21_X1 U22899 ( .B1(n19945), .B2(n19944), .A(n19943), .ZN(n19962) );
  NAND2_X1 U22900 ( .A1(n19946), .A2(n19964), .ZN(n19948) );
  OAI211_X1 U22901 ( .C1(n19962), .C2(n11472), .A(n19948), .B(n19947), .ZN(
        n19949) );
  AOI21_X1 U22902 ( .B1(n19950), .B2(n19965), .A(n19949), .ZN(n19951) );
  OAI21_X1 U22903 ( .B1(n19958), .B2(n19952), .A(n19951), .ZN(P1_U3027) );
  AOI22_X1 U22904 ( .A1(n19964), .A2(n19954), .B1(n19953), .B2(
        P1_REIP_REG_3__SCAN_IN), .ZN(n19957) );
  NAND2_X1 U22905 ( .A1(n19955), .A2(n19965), .ZN(n19956) );
  OAI211_X1 U22906 ( .C1(n19958), .C2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n19957), .B(n19956), .ZN(n19959) );
  INV_X1 U22907 ( .A(n19959), .ZN(n19960) );
  OAI21_X1 U22908 ( .B1(n19962), .B2(n19961), .A(n19960), .ZN(P1_U3028) );
  AOI22_X1 U22909 ( .A1(n19966), .A2(n19965), .B1(n19964), .B2(n19963), .ZN(
        n19972) );
  OAI22_X1 U22910 ( .A1(n19969), .A2(n19968), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19967), .ZN(n19970) );
  NAND3_X1 U22911 ( .A1(n19972), .A2(n19971), .A3(n19970), .ZN(P1_U3031) );
  NOR2_X1 U22912 ( .A1(n19973), .A2(n20747), .ZN(P1_U3032) );
  NOR2_X2 U22913 ( .A1(n19975), .A2(n19974), .ZN(n20015) );
  NOR2_X2 U22914 ( .A1(n19976), .A2(n19975), .ZN(n20016) );
  AOI22_X1 U22915 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20015), .B1(DATAI_16_), 
        .B2(n20016), .ZN(n20528) );
  NAND2_X1 U22916 ( .A1(n20735), .A2(n14974), .ZN(n20092) );
  NAND2_X1 U22917 ( .A1(n20014), .A2(n19978), .ZN(n20585) );
  INV_X1 U22918 ( .A(n20585), .ZN(n20515) );
  NAND2_X1 U22919 ( .A1(n20746), .A2(n20284), .ZN(n20050) );
  AOI22_X1 U22920 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20015), .B1(DATAI_24_), 
        .B2(n20016), .ZN(n20595) );
  INV_X1 U22921 ( .A(n20595), .ZN(n20525) );
  AOI22_X1 U22922 ( .A1(n20515), .A2(n10066), .B1(n20644), .B2(n20525), .ZN(
        n19991) );
  OR2_X1 U22923 ( .A1(n19987), .A2(n20244), .ZN(n20447) );
  INV_X1 U22924 ( .A(n20447), .ZN(n20511) );
  INV_X1 U22925 ( .A(n20644), .ZN(n19980) );
  NAND3_X1 U22926 ( .A1(n20048), .A2(n20128), .A3(n19980), .ZN(n19981) );
  NAND2_X1 U22927 ( .A1(n20580), .A2(n20516), .ZN(n20441) );
  NAND2_X1 U22928 ( .A1(n19981), .A2(n20441), .ZN(n19986) );
  NAND2_X1 U22929 ( .A1(n9822), .A2(n20508), .ZN(n19988) );
  INV_X1 U22930 ( .A(n20285), .ZN(n19983) );
  NAND2_X1 U22931 ( .A1(n19983), .A2(n20362), .ZN(n20129) );
  AOI22_X1 U22932 ( .A1(n19986), .A2(n19988), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20129), .ZN(n19984) );
  INV_X1 U22933 ( .A(n19986), .ZN(n19989) );
  AND2_X1 U22934 ( .A1(n19987), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20136) );
  INV_X1 U22935 ( .A(n20136), .ZN(n20366) );
  AOI22_X1 U22936 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20019), .B1(
        n20514), .B2(n20018), .ZN(n19990) );
  OAI211_X1 U22937 ( .C1(n20528), .C2(n20048), .A(n19991), .B(n19990), .ZN(
        P1_U3033) );
  NAND2_X1 U22938 ( .A1(n20014), .A2(n19992), .ZN(n20597) );
  INV_X1 U22939 ( .A(n20597), .ZN(n20530) );
  AOI22_X1 U22940 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20015), .B1(DATAI_25_), 
        .B2(n20016), .ZN(n20602) );
  INV_X1 U22941 ( .A(n20602), .ZN(n20531) );
  AOI22_X1 U22942 ( .A1(n20530), .A2(n10066), .B1(n20644), .B2(n20531), .ZN(
        n19995) );
  AOI22_X1 U22943 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20019), .B1(
        n20529), .B2(n20018), .ZN(n19994) );
  OAI211_X1 U22944 ( .C1(n20534), .C2(n20048), .A(n19995), .B(n19994), .ZN(
        P1_U3034) );
  NAND2_X1 U22945 ( .A1(n20014), .A2(n19996), .ZN(n20604) );
  INV_X1 U22946 ( .A(n20604), .ZN(n20536) );
  AOI22_X1 U22947 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20015), .B1(DATAI_26_), 
        .B2(n20016), .ZN(n20609) );
  INV_X1 U22948 ( .A(n20609), .ZN(n20537) );
  AOI22_X1 U22949 ( .A1(n20536), .A2(n10066), .B1(n20644), .B2(n20537), .ZN(
        n19999) );
  AOI22_X1 U22950 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20019), .B1(
        n20535), .B2(n20018), .ZN(n19998) );
  OAI211_X1 U22951 ( .C1(n20540), .C2(n20048), .A(n19999), .B(n19998), .ZN(
        P1_U3035) );
  AOI22_X1 U22952 ( .A1(DATAI_19_), .A2(n20016), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20015), .ZN(n20546) );
  NAND2_X1 U22953 ( .A1(n20014), .A2(n11272), .ZN(n20611) );
  INV_X1 U22954 ( .A(n20611), .ZN(n20542) );
  AOI22_X1 U22955 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20015), .B1(DATAI_27_), 
        .B2(n20016), .ZN(n20616) );
  INV_X1 U22956 ( .A(n20616), .ZN(n20543) );
  AOI22_X1 U22957 ( .A1(n20542), .A2(n10066), .B1(n20644), .B2(n20543), .ZN(
        n20002) );
  AOI22_X1 U22958 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20019), .B1(
        n20541), .B2(n20018), .ZN(n20001) );
  OAI211_X1 U22959 ( .C1(n20546), .C2(n20048), .A(n20002), .B(n20001), .ZN(
        P1_U3036) );
  AOI22_X1 U22960 ( .A1(DATAI_20_), .A2(n20016), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20015), .ZN(n20552) );
  NAND2_X1 U22961 ( .A1(n20014), .A2(n11277), .ZN(n20618) );
  INV_X1 U22962 ( .A(n20618), .ZN(n20548) );
  AOI22_X1 U22963 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20015), .B1(DATAI_28_), 
        .B2(n20016), .ZN(n20623) );
  INV_X1 U22964 ( .A(n20623), .ZN(n20549) );
  AOI22_X1 U22965 ( .A1(n20548), .A2(n10066), .B1(n20644), .B2(n20549), .ZN(
        n20005) );
  AOI22_X1 U22966 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20019), .B1(
        n20547), .B2(n20018), .ZN(n20004) );
  OAI211_X1 U22967 ( .C1(n20552), .C2(n20048), .A(n20005), .B(n20004), .ZN(
        P1_U3037) );
  AOI22_X1 U22968 ( .A1(DATAI_21_), .A2(n20016), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20015), .ZN(n20558) );
  NAND2_X1 U22969 ( .A1(n20014), .A2(n20006), .ZN(n20625) );
  INV_X1 U22970 ( .A(n20625), .ZN(n20554) );
  INV_X1 U22971 ( .A(n20630), .ZN(n20555) );
  AOI22_X1 U22972 ( .A1(n20554), .A2(n10066), .B1(n20644), .B2(n20555), .ZN(
        n20009) );
  AOI22_X1 U22973 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20019), .B1(
        n20553), .B2(n20018), .ZN(n20008) );
  OAI211_X1 U22974 ( .C1(n20558), .C2(n20048), .A(n20009), .B(n20008), .ZN(
        P1_U3038) );
  NAND2_X1 U22975 ( .A1(n20014), .A2(n11262), .ZN(n20632) );
  INV_X1 U22976 ( .A(n20632), .ZN(n20560) );
  AOI22_X1 U22977 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20015), .B1(DATAI_30_), 
        .B2(n20016), .ZN(n20637) );
  INV_X1 U22978 ( .A(n20637), .ZN(n20561) );
  AOI22_X1 U22979 ( .A1(n20560), .A2(n10066), .B1(n20644), .B2(n20561), .ZN(
        n20012) );
  AOI22_X1 U22980 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20019), .B1(
        n20559), .B2(n20018), .ZN(n20011) );
  OAI211_X1 U22981 ( .C1(n20564), .C2(n20048), .A(n20012), .B(n20011), .ZN(
        P1_U3039) );
  AOI22_X1 U22982 ( .A1(DATAI_23_), .A2(n20016), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n20015), .ZN(n20574) );
  NAND2_X1 U22983 ( .A1(n20014), .A2(n20013), .ZN(n20641) );
  INV_X1 U22984 ( .A(n20641), .ZN(n20568) );
  AOI22_X1 U22985 ( .A1(DATAI_31_), .A2(n20016), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20015), .ZN(n20649) );
  INV_X1 U22986 ( .A(n20649), .ZN(n20569) );
  AOI22_X1 U22987 ( .A1(n20568), .A2(n10066), .B1(n20644), .B2(n20569), .ZN(
        n20021) );
  AOI22_X1 U22988 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20019), .B1(
        n20566), .B2(n20018), .ZN(n20020) );
  OAI211_X1 U22989 ( .C1(n20574), .C2(n20048), .A(n20021), .B(n20020), .ZN(
        P1_U3040) );
  NOR2_X1 U22990 ( .A1(n20050), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20027) );
  INV_X1 U22991 ( .A(n20027), .ZN(n20024) );
  NOR2_X1 U22992 ( .A1(n20471), .A2(n20024), .ZN(n20044) );
  INV_X1 U22993 ( .A(n20023), .ZN(n20322) );
  AOI21_X1 U22994 ( .B1(n9822), .B2(n20322), .A(n20044), .ZN(n20025) );
  OAI22_X1 U22995 ( .A1(n20025), .A2(n20743), .B1(n20024), .B2(n20244), .ZN(
        n20043) );
  AOI22_X1 U22996 ( .A1(n20515), .A2(n20044), .B1(n20514), .B2(n20043), .ZN(
        n20029) );
  OAI21_X1 U22997 ( .B1(n20092), .B2(n20516), .A(n20025), .ZN(n20026) );
  OAI221_X1 U22998 ( .B1(n20580), .B2(n20027), .C1(n20743), .C2(n20026), .A(
        n20589), .ZN(n20045) );
  INV_X1 U22999 ( .A(n20048), .ZN(n20034) );
  AOI22_X1 U23000 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20045), .B1(
        n20034), .B2(n20525), .ZN(n20028) );
  OAI211_X1 U23001 ( .C1(n20528), .C2(n20086), .A(n20029), .B(n20028), .ZN(
        P1_U3041) );
  AOI22_X1 U23002 ( .A1(n20530), .A2(n20044), .B1(n20529), .B2(n20043), .ZN(
        n20031) );
  AOI22_X1 U23003 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20045), .B1(
        n20034), .B2(n20531), .ZN(n20030) );
  OAI211_X1 U23004 ( .C1(n20534), .C2(n20086), .A(n20031), .B(n20030), .ZN(
        P1_U3042) );
  AOI22_X1 U23005 ( .A1(n20536), .A2(n20044), .B1(n20535), .B2(n20043), .ZN(
        n20033) );
  AOI22_X1 U23006 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20045), .B1(
        n20034), .B2(n20537), .ZN(n20032) );
  OAI211_X1 U23007 ( .C1(n20540), .C2(n20086), .A(n20033), .B(n20032), .ZN(
        P1_U3043) );
  AOI22_X1 U23008 ( .A1(n20542), .A2(n20044), .B1(n20541), .B2(n20043), .ZN(
        n20036) );
  AOI22_X1 U23009 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20045), .B1(
        n20034), .B2(n20543), .ZN(n20035) );
  OAI211_X1 U23010 ( .C1(n20546), .C2(n20086), .A(n20036), .B(n20035), .ZN(
        P1_U3044) );
  AOI22_X1 U23011 ( .A1(n20548), .A2(n20044), .B1(n20547), .B2(n20043), .ZN(
        n20038) );
  INV_X1 U23012 ( .A(n20552), .ZN(n20620) );
  AOI22_X1 U23013 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20045), .B1(
        n20053), .B2(n20620), .ZN(n20037) );
  OAI211_X1 U23014 ( .C1(n20623), .C2(n20048), .A(n20038), .B(n20037), .ZN(
        P1_U3045) );
  AOI22_X1 U23015 ( .A1(n20554), .A2(n20044), .B1(n20553), .B2(n20043), .ZN(
        n20040) );
  INV_X1 U23016 ( .A(n20558), .ZN(n20627) );
  AOI22_X1 U23017 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20045), .B1(
        n20053), .B2(n20627), .ZN(n20039) );
  OAI211_X1 U23018 ( .C1(n20630), .C2(n20048), .A(n20040), .B(n20039), .ZN(
        P1_U3046) );
  AOI22_X1 U23019 ( .A1(n20560), .A2(n20044), .B1(n20559), .B2(n20043), .ZN(
        n20042) );
  INV_X1 U23020 ( .A(n20564), .ZN(n20634) );
  AOI22_X1 U23021 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20045), .B1(
        n20053), .B2(n20634), .ZN(n20041) );
  OAI211_X1 U23022 ( .C1(n20637), .C2(n20048), .A(n20042), .B(n20041), .ZN(
        P1_U3047) );
  AOI22_X1 U23023 ( .A1(n20568), .A2(n20044), .B1(n20566), .B2(n20043), .ZN(
        n20047) );
  INV_X1 U23024 ( .A(n20574), .ZN(n20643) );
  AOI22_X1 U23025 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20045), .B1(
        n20053), .B2(n20643), .ZN(n20046) );
  OAI211_X1 U23026 ( .C1(n20649), .C2(n20048), .A(n20047), .B(n20046), .ZN(
        P1_U3048) );
  INV_X1 U23027 ( .A(n20506), .ZN(n20049) );
  INV_X1 U23028 ( .A(n20050), .ZN(n20087) );
  NAND2_X1 U23029 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20087), .ZN(
        n20096) );
  OR2_X1 U23030 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20096), .ZN(
        n20080) );
  OAI22_X1 U23031 ( .A1(n20086), .A2(n20595), .B1(n20585), .B2(n20080), .ZN(
        n20051) );
  INV_X1 U23032 ( .A(n20051), .ZN(n20061) );
  INV_X1 U23033 ( .A(n20120), .ZN(n20052) );
  OAI21_X1 U23034 ( .B1(n20053), .B2(n20052), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20054) );
  NAND2_X1 U23035 ( .A1(n20054), .A2(n20580), .ZN(n20059) );
  INV_X1 U23036 ( .A(n20059), .ZN(n20055) );
  INV_X1 U23037 ( .A(n20508), .ZN(n20518) );
  NAND2_X1 U23038 ( .A1(n9822), .A2(n20518), .ZN(n20058) );
  AOI22_X1 U23039 ( .A1(n20055), .A2(n20058), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20080), .ZN(n20056) );
  OAI21_X1 U23040 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20362), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20209) );
  NAND3_X1 U23041 ( .A1(n20364), .A2(n20056), .A3(n20209), .ZN(n20083) );
  NAND2_X1 U23042 ( .A1(n20057), .A2(n20746), .ZN(n20212) );
  AOI22_X1 U23043 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20083), .B1(
        n20514), .B2(n20082), .ZN(n20060) );
  OAI211_X1 U23044 ( .C1(n20528), .C2(n20120), .A(n20061), .B(n20060), .ZN(
        P1_U3049) );
  OAI22_X1 U23045 ( .A1(n20086), .A2(n20602), .B1(n20080), .B2(n20597), .ZN(
        n20062) );
  INV_X1 U23046 ( .A(n20062), .ZN(n20064) );
  AOI22_X1 U23047 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20083), .B1(
        n20529), .B2(n20082), .ZN(n20063) );
  OAI211_X1 U23048 ( .C1(n20534), .C2(n20120), .A(n20064), .B(n20063), .ZN(
        P1_U3050) );
  OAI22_X1 U23049 ( .A1(n20086), .A2(n20609), .B1(n20080), .B2(n20604), .ZN(
        n20065) );
  INV_X1 U23050 ( .A(n20065), .ZN(n20067) );
  AOI22_X1 U23051 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20083), .B1(
        n20535), .B2(n20082), .ZN(n20066) );
  OAI211_X1 U23052 ( .C1(n20540), .C2(n20120), .A(n20067), .B(n20066), .ZN(
        P1_U3051) );
  OAI22_X1 U23053 ( .A1(n20546), .A2(n20120), .B1(n20611), .B2(n20080), .ZN(
        n20068) );
  INV_X1 U23054 ( .A(n20068), .ZN(n20070) );
  AOI22_X1 U23055 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20083), .B1(
        n20541), .B2(n20082), .ZN(n20069) );
  OAI211_X1 U23056 ( .C1(n20616), .C2(n20086), .A(n20070), .B(n20069), .ZN(
        P1_U3052) );
  OAI22_X1 U23057 ( .A1(n20086), .A2(n20623), .B1(n20080), .B2(n20618), .ZN(
        n20071) );
  INV_X1 U23058 ( .A(n20071), .ZN(n20073) );
  AOI22_X1 U23059 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20083), .B1(
        n20547), .B2(n20082), .ZN(n20072) );
  OAI211_X1 U23060 ( .C1(n20552), .C2(n20120), .A(n20073), .B(n20072), .ZN(
        P1_U3053) );
  OAI22_X1 U23061 ( .A1(n20086), .A2(n20630), .B1(n20080), .B2(n20625), .ZN(
        n20074) );
  INV_X1 U23062 ( .A(n20074), .ZN(n20076) );
  AOI22_X1 U23063 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20083), .B1(
        n20553), .B2(n20082), .ZN(n20075) );
  OAI211_X1 U23064 ( .C1(n20558), .C2(n20120), .A(n20076), .B(n20075), .ZN(
        P1_U3054) );
  OAI22_X1 U23065 ( .A1(n20086), .A2(n20637), .B1(n20080), .B2(n20632), .ZN(
        n20077) );
  INV_X1 U23066 ( .A(n20077), .ZN(n20079) );
  AOI22_X1 U23067 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20083), .B1(
        n20559), .B2(n20082), .ZN(n20078) );
  OAI211_X1 U23068 ( .C1(n20564), .C2(n20120), .A(n20079), .B(n20078), .ZN(
        P1_U3055) );
  OAI22_X1 U23069 ( .A1(n20574), .A2(n20120), .B1(n20641), .B2(n20080), .ZN(
        n20081) );
  INV_X1 U23070 ( .A(n20081), .ZN(n20085) );
  AOI22_X1 U23071 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20083), .B1(
        n20566), .B2(n20082), .ZN(n20084) );
  OAI211_X1 U23072 ( .C1(n20649), .C2(n20086), .A(n20085), .B(n20084), .ZN(
        P1_U3056) );
  NAND2_X1 U23073 ( .A1(n20398), .A2(n20087), .ZN(n20119) );
  OAI22_X1 U23074 ( .A1(n20528), .A2(n20166), .B1(n20585), .B2(n20119), .ZN(
        n20088) );
  INV_X1 U23075 ( .A(n20088), .ZN(n20100) );
  AND2_X1 U23076 ( .A1(n20090), .A2(n20089), .ZN(n20575) );
  INV_X1 U23077 ( .A(n20119), .ZN(n20091) );
  AOI21_X1 U23078 ( .B1(n9822), .B2(n20575), .A(n20091), .ZN(n20097) );
  OR2_X1 U23079 ( .A1(n20092), .A2(n20587), .ZN(n20093) );
  AND2_X1 U23080 ( .A1(n20093), .A2(n20580), .ZN(n20095) );
  AOI22_X1 U23081 ( .A1(n20097), .A2(n20095), .B1(n20743), .B2(n20096), .ZN(
        n20094) );
  NAND2_X1 U23082 ( .A1(n20589), .A2(n20094), .ZN(n20123) );
  INV_X1 U23083 ( .A(n20095), .ZN(n20098) );
  OAI22_X1 U23084 ( .A1(n20098), .A2(n20097), .B1(n20244), .B2(n20096), .ZN(
        n20122) );
  AOI22_X1 U23085 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20123), .B1(
        n20514), .B2(n20122), .ZN(n20099) );
  OAI211_X1 U23086 ( .C1(n20595), .C2(n20120), .A(n20100), .B(n20099), .ZN(
        P1_U3057) );
  OAI22_X1 U23087 ( .A1(n20602), .A2(n20120), .B1(n20597), .B2(n20119), .ZN(
        n20101) );
  INV_X1 U23088 ( .A(n20101), .ZN(n20103) );
  AOI22_X1 U23089 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20123), .B1(
        n20529), .B2(n20122), .ZN(n20102) );
  OAI211_X1 U23090 ( .C1(n20534), .C2(n20166), .A(n20103), .B(n20102), .ZN(
        P1_U3058) );
  OAI22_X1 U23091 ( .A1(n20609), .A2(n20120), .B1(n20604), .B2(n20119), .ZN(
        n20104) );
  INV_X1 U23092 ( .A(n20104), .ZN(n20106) );
  AOI22_X1 U23093 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20123), .B1(
        n20535), .B2(n20122), .ZN(n20105) );
  OAI211_X1 U23094 ( .C1(n20540), .C2(n20166), .A(n20106), .B(n20105), .ZN(
        P1_U3059) );
  OAI22_X1 U23095 ( .A1(n20546), .A2(n20166), .B1(n20611), .B2(n20119), .ZN(
        n20107) );
  INV_X1 U23096 ( .A(n20107), .ZN(n20109) );
  AOI22_X1 U23097 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20123), .B1(
        n20541), .B2(n20122), .ZN(n20108) );
  OAI211_X1 U23098 ( .C1(n20616), .C2(n20120), .A(n20109), .B(n20108), .ZN(
        P1_U3060) );
  OAI22_X1 U23099 ( .A1(n20623), .A2(n20120), .B1(n20618), .B2(n20119), .ZN(
        n20110) );
  INV_X1 U23100 ( .A(n20110), .ZN(n20112) );
  AOI22_X1 U23101 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20123), .B1(
        n20547), .B2(n20122), .ZN(n20111) );
  OAI211_X1 U23102 ( .C1(n20552), .C2(n20166), .A(n20112), .B(n20111), .ZN(
        P1_U3061) );
  OAI22_X1 U23103 ( .A1(n20630), .A2(n20120), .B1(n20625), .B2(n20119), .ZN(
        n20113) );
  INV_X1 U23104 ( .A(n20113), .ZN(n20115) );
  AOI22_X1 U23105 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20123), .B1(
        n20553), .B2(n20122), .ZN(n20114) );
  OAI211_X1 U23106 ( .C1(n20558), .C2(n20166), .A(n20115), .B(n20114), .ZN(
        P1_U3062) );
  OAI22_X1 U23107 ( .A1(n20637), .A2(n20120), .B1(n20632), .B2(n20119), .ZN(
        n20116) );
  INV_X1 U23108 ( .A(n20116), .ZN(n20118) );
  AOI22_X1 U23109 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20123), .B1(
        n20559), .B2(n20122), .ZN(n20117) );
  OAI211_X1 U23110 ( .C1(n20564), .C2(n20166), .A(n20118), .B(n20117), .ZN(
        P1_U3063) );
  OAI22_X1 U23111 ( .A1(n20649), .A2(n20120), .B1(n20641), .B2(n20119), .ZN(
        n20121) );
  INV_X1 U23112 ( .A(n20121), .ZN(n20125) );
  AOI22_X1 U23113 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20123), .B1(
        n20566), .B2(n20122), .ZN(n20124) );
  OAI211_X1 U23114 ( .C1(n20574), .C2(n20166), .A(n20125), .B(n20124), .ZN(
        P1_U3064) );
  OR2_X1 U23115 ( .A1(n14974), .A2(n20126), .ZN(n20249) );
  OR2_X1 U23116 ( .A1(n20439), .A2(n20206), .ZN(n20161) );
  NOR2_X1 U23117 ( .A1(n13262), .A2(n20127), .ZN(n20242) );
  NAND3_X1 U23118 ( .A1(n20242), .A2(n20128), .A3(n20508), .ZN(n20131) );
  OR2_X1 U23119 ( .A1(n20447), .A2(n20129), .ZN(n20130) );
  OAI22_X1 U23120 ( .A1(n20585), .A2(n20161), .B1(n20160), .B2(n20584), .ZN(
        n20132) );
  INV_X1 U23121 ( .A(n20132), .ZN(n20140) );
  INV_X1 U23122 ( .A(n20161), .ZN(n20138) );
  AOI21_X1 U23123 ( .B1(n20198), .B2(n20166), .A(n20516), .ZN(n20133) );
  AOI21_X1 U23124 ( .B1(n20242), .B2(n20508), .A(n20133), .ZN(n20134) );
  NOR2_X1 U23125 ( .A1(n20134), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20137) );
  AOI22_X1 U23126 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20163), .B1(
        n20157), .B2(n20525), .ZN(n20139) );
  OAI211_X1 U23127 ( .C1(n20528), .C2(n20198), .A(n20140), .B(n20139), .ZN(
        P1_U3065) );
  OAI22_X1 U23128 ( .A1(n20597), .A2(n20161), .B1(n20160), .B2(n20596), .ZN(
        n20141) );
  INV_X1 U23129 ( .A(n20141), .ZN(n20143) );
  AOI22_X1 U23130 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20163), .B1(
        n20157), .B2(n20531), .ZN(n20142) );
  OAI211_X1 U23131 ( .C1(n20534), .C2(n20198), .A(n20143), .B(n20142), .ZN(
        P1_U3066) );
  OAI22_X1 U23132 ( .A1(n20604), .A2(n20161), .B1(n20160), .B2(n20603), .ZN(
        n20144) );
  INV_X1 U23133 ( .A(n20144), .ZN(n20146) );
  AOI22_X1 U23134 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20163), .B1(
        n20157), .B2(n20537), .ZN(n20145) );
  OAI211_X1 U23135 ( .C1(n20540), .C2(n20198), .A(n20146), .B(n20145), .ZN(
        P1_U3067) );
  OAI22_X1 U23136 ( .A1(n20611), .A2(n20161), .B1(n20160), .B2(n20610), .ZN(
        n20147) );
  INV_X1 U23137 ( .A(n20147), .ZN(n20149) );
  INV_X1 U23138 ( .A(n20198), .ZN(n20202) );
  INV_X1 U23139 ( .A(n20546), .ZN(n20613) );
  AOI22_X1 U23140 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20163), .B1(
        n20202), .B2(n20613), .ZN(n20148) );
  OAI211_X1 U23141 ( .C1(n20616), .C2(n20166), .A(n20149), .B(n20148), .ZN(
        P1_U3068) );
  OAI22_X1 U23142 ( .A1(n20618), .A2(n20161), .B1(n20160), .B2(n20617), .ZN(
        n20150) );
  INV_X1 U23143 ( .A(n20150), .ZN(n20152) );
  AOI22_X1 U23144 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20163), .B1(
        n20157), .B2(n20549), .ZN(n20151) );
  OAI211_X1 U23145 ( .C1(n20552), .C2(n20198), .A(n20152), .B(n20151), .ZN(
        P1_U3069) );
  OAI22_X1 U23146 ( .A1(n20625), .A2(n20161), .B1(n20160), .B2(n20624), .ZN(
        n20153) );
  INV_X1 U23147 ( .A(n20153), .ZN(n20155) );
  AOI22_X1 U23148 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20163), .B1(
        n20157), .B2(n20555), .ZN(n20154) );
  OAI211_X1 U23149 ( .C1(n20558), .C2(n20198), .A(n20155), .B(n20154), .ZN(
        P1_U3070) );
  OAI22_X1 U23150 ( .A1(n20632), .A2(n20161), .B1(n20160), .B2(n20631), .ZN(
        n20156) );
  INV_X1 U23151 ( .A(n20156), .ZN(n20159) );
  AOI22_X1 U23152 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20163), .B1(
        n20157), .B2(n20561), .ZN(n20158) );
  OAI211_X1 U23153 ( .C1(n20564), .C2(n20198), .A(n20159), .B(n20158), .ZN(
        P1_U3071) );
  OAI22_X1 U23154 ( .A1(n20641), .A2(n20161), .B1(n20160), .B2(n20638), .ZN(
        n20162) );
  INV_X1 U23155 ( .A(n20162), .ZN(n20165) );
  AOI22_X1 U23156 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20163), .B1(
        n20202), .B2(n20643), .ZN(n20164) );
  OAI211_X1 U23157 ( .C1(n20649), .C2(n20166), .A(n20165), .B(n20164), .ZN(
        P1_U3072) );
  NOR2_X1 U23158 ( .A1(n20206), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20175) );
  INV_X1 U23159 ( .A(n20175), .ZN(n20167) );
  OR2_X1 U23160 ( .A1(n20471), .A2(n20167), .ZN(n20200) );
  NAND2_X1 U23161 ( .A1(n20242), .A2(n20322), .ZN(n20168) );
  NAND2_X1 U23162 ( .A1(n20168), .A2(n20200), .ZN(n20172) );
  NAND2_X1 U23163 ( .A1(n20172), .A2(n20128), .ZN(n20170) );
  NAND2_X1 U23164 ( .A1(n20175), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20169) );
  OAI22_X1 U23165 ( .A1(n20585), .A2(n20200), .B1(n20199), .B2(n20584), .ZN(
        n20171) );
  INV_X1 U23166 ( .A(n20171), .ZN(n20178) );
  INV_X1 U23167 ( .A(n20172), .ZN(n20173) );
  OAI21_X1 U23168 ( .B1(n20249), .B2(n20516), .A(n20173), .ZN(n20174) );
  OAI221_X1 U23169 ( .B1(n20128), .B2(n20175), .C1(n20743), .C2(n20174), .A(
        n20589), .ZN(n20203) );
  INV_X1 U23170 ( .A(n20528), .ZN(n20592) );
  AOI22_X1 U23171 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20203), .B1(
        n20195), .B2(n20592), .ZN(n20177) );
  OAI211_X1 U23172 ( .C1(n20595), .C2(n20198), .A(n20178), .B(n20177), .ZN(
        P1_U3073) );
  OAI22_X1 U23173 ( .A1(n20597), .A2(n20200), .B1(n20199), .B2(n20596), .ZN(
        n20179) );
  INV_X1 U23174 ( .A(n20179), .ZN(n20181) );
  AOI22_X1 U23175 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20531), .ZN(n20180) );
  OAI211_X1 U23176 ( .C1(n20534), .C2(n20236), .A(n20181), .B(n20180), .ZN(
        P1_U3074) );
  OAI22_X1 U23177 ( .A1(n20604), .A2(n20200), .B1(n20199), .B2(n20603), .ZN(
        n20182) );
  INV_X1 U23178 ( .A(n20182), .ZN(n20184) );
  INV_X1 U23179 ( .A(n20540), .ZN(n20606) );
  AOI22_X1 U23180 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20203), .B1(
        n20195), .B2(n20606), .ZN(n20183) );
  OAI211_X1 U23181 ( .C1(n20609), .C2(n20198), .A(n20184), .B(n20183), .ZN(
        P1_U3075) );
  OAI22_X1 U23182 ( .A1(n20611), .A2(n20200), .B1(n20199), .B2(n20610), .ZN(
        n20185) );
  INV_X1 U23183 ( .A(n20185), .ZN(n20187) );
  AOI22_X1 U23184 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20203), .B1(
        n20195), .B2(n20613), .ZN(n20186) );
  OAI211_X1 U23185 ( .C1(n20616), .C2(n20198), .A(n20187), .B(n20186), .ZN(
        P1_U3076) );
  OAI22_X1 U23186 ( .A1(n20618), .A2(n20200), .B1(n20199), .B2(n20617), .ZN(
        n20188) );
  INV_X1 U23187 ( .A(n20188), .ZN(n20190) );
  AOI22_X1 U23188 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20203), .B1(
        n20195), .B2(n20620), .ZN(n20189) );
  OAI211_X1 U23189 ( .C1(n20623), .C2(n20198), .A(n20190), .B(n20189), .ZN(
        P1_U3077) );
  OAI22_X1 U23190 ( .A1(n20625), .A2(n20200), .B1(n20199), .B2(n20624), .ZN(
        n20191) );
  INV_X1 U23191 ( .A(n20191), .ZN(n20193) );
  AOI22_X1 U23192 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20203), .B1(
        n20195), .B2(n20627), .ZN(n20192) );
  OAI211_X1 U23193 ( .C1(n20630), .C2(n20198), .A(n20193), .B(n20192), .ZN(
        P1_U3078) );
  OAI22_X1 U23194 ( .A1(n20632), .A2(n20200), .B1(n20199), .B2(n20631), .ZN(
        n20194) );
  INV_X1 U23195 ( .A(n20194), .ZN(n20197) );
  AOI22_X1 U23196 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20203), .B1(
        n20195), .B2(n20634), .ZN(n20196) );
  OAI211_X1 U23197 ( .C1(n20637), .C2(n20198), .A(n20197), .B(n20196), .ZN(
        P1_U3079) );
  OAI22_X1 U23198 ( .A1(n20641), .A2(n20200), .B1(n20199), .B2(n20638), .ZN(
        n20201) );
  INV_X1 U23199 ( .A(n20201), .ZN(n20205) );
  AOI22_X1 U23200 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20569), .ZN(n20204) );
  OAI211_X1 U23201 ( .C1(n20574), .C2(n20236), .A(n20205), .B(n20204), .ZN(
        P1_U3080) );
  NOR2_X1 U23202 ( .A1(n20579), .A2(n20206), .ZN(n20252) );
  NAND2_X1 U23203 ( .A1(n20471), .A2(n20252), .ZN(n20235) );
  INV_X1 U23204 ( .A(n20249), .ZN(n20254) );
  OAI22_X1 U23205 ( .A1(n20585), .A2(n20235), .B1(n20283), .B2(n20528), .ZN(
        n20207) );
  INV_X1 U23206 ( .A(n20207), .ZN(n20216) );
  NAND2_X1 U23207 ( .A1(n20236), .A2(n20283), .ZN(n20208) );
  AOI21_X1 U23208 ( .B1(n20208), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20743), 
        .ZN(n20211) );
  NAND2_X1 U23209 ( .A1(n20242), .A2(n20518), .ZN(n20213) );
  AOI22_X1 U23210 ( .A1(n20211), .A2(n20213), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20235), .ZN(n20210) );
  NAND3_X1 U23211 ( .A1(n20522), .A2(n20210), .A3(n20209), .ZN(n20239) );
  INV_X1 U23212 ( .A(n20211), .ZN(n20214) );
  AOI22_X1 U23213 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20239), .B1(
        n20514), .B2(n20238), .ZN(n20215) );
  OAI211_X1 U23214 ( .C1(n20595), .C2(n20236), .A(n20216), .B(n20215), .ZN(
        P1_U3081) );
  OAI22_X1 U23215 ( .A1(n20597), .A2(n20235), .B1(n20283), .B2(n20534), .ZN(
        n20217) );
  INV_X1 U23216 ( .A(n20217), .ZN(n20219) );
  AOI22_X1 U23217 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20239), .B1(
        n20529), .B2(n20238), .ZN(n20218) );
  OAI211_X1 U23218 ( .C1(n20602), .C2(n20236), .A(n20219), .B(n20218), .ZN(
        P1_U3082) );
  OAI22_X1 U23219 ( .A1(n20236), .A2(n20609), .B1(n20604), .B2(n20235), .ZN(
        n20220) );
  INV_X1 U23220 ( .A(n20220), .ZN(n20222) );
  AOI22_X1 U23221 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20239), .B1(
        n20535), .B2(n20238), .ZN(n20221) );
  OAI211_X1 U23222 ( .C1(n20540), .C2(n20283), .A(n20222), .B(n20221), .ZN(
        P1_U3083) );
  OAI22_X1 U23223 ( .A1(n20611), .A2(n20235), .B1(n20283), .B2(n20546), .ZN(
        n20223) );
  INV_X1 U23224 ( .A(n20223), .ZN(n20225) );
  AOI22_X1 U23225 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20239), .B1(
        n20541), .B2(n20238), .ZN(n20224) );
  OAI211_X1 U23226 ( .C1(n20616), .C2(n20236), .A(n20225), .B(n20224), .ZN(
        P1_U3084) );
  OAI22_X1 U23227 ( .A1(n20618), .A2(n20235), .B1(n20283), .B2(n20552), .ZN(
        n20226) );
  INV_X1 U23228 ( .A(n20226), .ZN(n20228) );
  AOI22_X1 U23229 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20239), .B1(
        n20547), .B2(n20238), .ZN(n20227) );
  OAI211_X1 U23230 ( .C1(n20623), .C2(n20236), .A(n20228), .B(n20227), .ZN(
        P1_U3085) );
  OAI22_X1 U23231 ( .A1(n20236), .A2(n20630), .B1(n20625), .B2(n20235), .ZN(
        n20229) );
  INV_X1 U23232 ( .A(n20229), .ZN(n20231) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20239), .B1(
        n20553), .B2(n20238), .ZN(n20230) );
  OAI211_X1 U23234 ( .C1(n20558), .C2(n20283), .A(n20231), .B(n20230), .ZN(
        P1_U3086) );
  OAI22_X1 U23235 ( .A1(n20632), .A2(n20235), .B1(n20283), .B2(n20564), .ZN(
        n20232) );
  INV_X1 U23236 ( .A(n20232), .ZN(n20234) );
  AOI22_X1 U23237 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20239), .B1(
        n20559), .B2(n20238), .ZN(n20233) );
  OAI211_X1 U23238 ( .C1(n20637), .C2(n20236), .A(n20234), .B(n20233), .ZN(
        P1_U3087) );
  OAI22_X1 U23239 ( .A1(n20236), .A2(n20649), .B1(n20641), .B2(n20235), .ZN(
        n20237) );
  INV_X1 U23240 ( .A(n20237), .ZN(n20241) );
  AOI22_X1 U23241 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20239), .B1(
        n20566), .B2(n20238), .ZN(n20240) );
  OAI211_X1 U23242 ( .C1(n20574), .C2(n20283), .A(n20241), .B(n20240), .ZN(
        P1_U3088) );
  NAND2_X1 U23243 ( .A1(n20242), .A2(n20575), .ZN(n20243) );
  NAND2_X1 U23244 ( .A1(n20243), .A2(n20278), .ZN(n20247) );
  INV_X1 U23245 ( .A(n20252), .ZN(n20245) );
  NOR2_X1 U23246 ( .A1(n20245), .A2(n20244), .ZN(n20246) );
  AOI21_X1 U23247 ( .B1(n20247), .B2(n20580), .A(n20246), .ZN(n20277) );
  OAI22_X1 U23248 ( .A1(n20585), .A2(n20278), .B1(n20277), .B2(n20584), .ZN(
        n20248) );
  INV_X1 U23249 ( .A(n20248), .ZN(n20256) );
  NOR2_X1 U23250 ( .A1(n20249), .A2(n20743), .ZN(n20251) );
  INV_X1 U23251 ( .A(n20587), .ZN(n20250) );
  AND2_X1 U23252 ( .A1(n20251), .A2(n20250), .ZN(n20733) );
  OAI21_X1 U23253 ( .B1(n20252), .B2(n20733), .A(n20589), .ZN(n20280) );
  NAND2_X1 U23254 ( .A1(n20254), .A2(n20408), .ZN(n20276) );
  AOI22_X1 U23255 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20280), .B1(
        n20317), .B2(n20592), .ZN(n20255) );
  OAI211_X1 U23256 ( .C1(n20595), .C2(n20283), .A(n20256), .B(n20255), .ZN(
        P1_U3089) );
  OAI22_X1 U23257 ( .A1(n20597), .A2(n20278), .B1(n20277), .B2(n20596), .ZN(
        n20257) );
  INV_X1 U23258 ( .A(n20257), .ZN(n20259) );
  INV_X1 U23259 ( .A(n20534), .ZN(n20599) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20280), .B1(
        n20317), .B2(n20599), .ZN(n20258) );
  OAI211_X1 U23261 ( .C1(n20602), .C2(n20283), .A(n20259), .B(n20258), .ZN(
        P1_U3090) );
  OAI22_X1 U23262 ( .A1(n20604), .A2(n20278), .B1(n20277), .B2(n20603), .ZN(
        n20260) );
  INV_X1 U23263 ( .A(n20260), .ZN(n20262) );
  INV_X1 U23264 ( .A(n20283), .ZN(n20273) );
  AOI22_X1 U23265 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20280), .B1(
        n20273), .B2(n20537), .ZN(n20261) );
  OAI211_X1 U23266 ( .C1(n20540), .C2(n20276), .A(n20262), .B(n20261), .ZN(
        P1_U3091) );
  OAI22_X1 U23267 ( .A1(n20611), .A2(n20278), .B1(n20277), .B2(n20610), .ZN(
        n20263) );
  INV_X1 U23268 ( .A(n20263), .ZN(n20265) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20280), .B1(
        n20317), .B2(n20613), .ZN(n20264) );
  OAI211_X1 U23270 ( .C1(n20616), .C2(n20283), .A(n20265), .B(n20264), .ZN(
        P1_U3092) );
  OAI22_X1 U23271 ( .A1(n20618), .A2(n20278), .B1(n20277), .B2(n20617), .ZN(
        n20266) );
  INV_X1 U23272 ( .A(n20266), .ZN(n20268) );
  AOI22_X1 U23273 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20280), .B1(
        n20317), .B2(n20620), .ZN(n20267) );
  OAI211_X1 U23274 ( .C1(n20623), .C2(n20283), .A(n20268), .B(n20267), .ZN(
        P1_U3093) );
  OAI22_X1 U23275 ( .A1(n20625), .A2(n20278), .B1(n20277), .B2(n20624), .ZN(
        n20269) );
  INV_X1 U23276 ( .A(n20269), .ZN(n20271) );
  AOI22_X1 U23277 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20280), .B1(
        n20317), .B2(n20627), .ZN(n20270) );
  OAI211_X1 U23278 ( .C1(n20630), .C2(n20283), .A(n20271), .B(n20270), .ZN(
        P1_U3094) );
  OAI22_X1 U23279 ( .A1(n20632), .A2(n20278), .B1(n20277), .B2(n20631), .ZN(
        n20272) );
  INV_X1 U23280 ( .A(n20272), .ZN(n20275) );
  AOI22_X1 U23281 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20280), .B1(
        n20273), .B2(n20561), .ZN(n20274) );
  OAI211_X1 U23282 ( .C1(n20564), .C2(n20276), .A(n20275), .B(n20274), .ZN(
        P1_U3095) );
  OAI22_X1 U23283 ( .A1(n20641), .A2(n20278), .B1(n20277), .B2(n20638), .ZN(
        n20279) );
  INV_X1 U23284 ( .A(n20279), .ZN(n20282) );
  AOI22_X1 U23285 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20280), .B1(
        n20317), .B2(n20643), .ZN(n20281) );
  OAI211_X1 U23286 ( .C1(n20649), .C2(n20283), .A(n20282), .B(n20281), .ZN(
        P1_U3096) );
  NAND2_X1 U23287 ( .A1(n20284), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20396) );
  OR2_X1 U23288 ( .A1(n20439), .A2(n20396), .ZN(n20315) );
  AND2_X1 U23289 ( .A1(n20736), .A2(n13262), .ZN(n20399) );
  INV_X1 U23290 ( .A(n20315), .ZN(n20293) );
  AOI21_X1 U23291 ( .B1(n20399), .B2(n20508), .A(n20293), .ZN(n20290) );
  OR2_X1 U23292 ( .A1(n20290), .A2(n20743), .ZN(n20287) );
  NAND2_X1 U23293 ( .A1(n20285), .A2(n20362), .ZN(n20448) );
  OR2_X1 U23294 ( .A1(n20448), .A2(n20366), .ZN(n20286) );
  OAI22_X1 U23295 ( .A1(n20585), .A2(n20315), .B1(n20314), .B2(n20584), .ZN(
        n20288) );
  INV_X1 U23296 ( .A(n20288), .ZN(n20295) );
  INV_X1 U23297 ( .A(n20359), .ZN(n20289) );
  OAI21_X1 U23298 ( .B1(n20289), .B2(n20317), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20291) );
  NAND2_X1 U23299 ( .A1(n20291), .A2(n20290), .ZN(n20292) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20318), .B1(
        n20317), .B2(n20525), .ZN(n20294) );
  OAI211_X1 U23301 ( .C1(n20528), .C2(n20359), .A(n20295), .B(n20294), .ZN(
        P1_U3097) );
  OAI22_X1 U23302 ( .A1(n20597), .A2(n20315), .B1(n20314), .B2(n20596), .ZN(
        n20296) );
  INV_X1 U23303 ( .A(n20296), .ZN(n20298) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20318), .B1(
        n20317), .B2(n20531), .ZN(n20297) );
  OAI211_X1 U23305 ( .C1(n20534), .C2(n20359), .A(n20298), .B(n20297), .ZN(
        P1_U3098) );
  OAI22_X1 U23306 ( .A1(n20604), .A2(n20315), .B1(n20314), .B2(n20603), .ZN(
        n20299) );
  INV_X1 U23307 ( .A(n20299), .ZN(n20301) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20318), .B1(
        n20317), .B2(n20537), .ZN(n20300) );
  OAI211_X1 U23309 ( .C1(n20540), .C2(n20359), .A(n20301), .B(n20300), .ZN(
        P1_U3099) );
  OAI22_X1 U23310 ( .A1(n20611), .A2(n20315), .B1(n20314), .B2(n20610), .ZN(
        n20302) );
  INV_X1 U23311 ( .A(n20302), .ZN(n20304) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20318), .B1(
        n20317), .B2(n20543), .ZN(n20303) );
  OAI211_X1 U23313 ( .C1(n20546), .C2(n20359), .A(n20304), .B(n20303), .ZN(
        P1_U3100) );
  OAI22_X1 U23314 ( .A1(n20618), .A2(n20315), .B1(n20314), .B2(n20617), .ZN(
        n20305) );
  INV_X1 U23315 ( .A(n20305), .ZN(n20307) );
  AOI22_X1 U23316 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20318), .B1(
        n20317), .B2(n20549), .ZN(n20306) );
  OAI211_X1 U23317 ( .C1(n20552), .C2(n20359), .A(n20307), .B(n20306), .ZN(
        P1_U3101) );
  OAI22_X1 U23318 ( .A1(n20625), .A2(n20315), .B1(n20314), .B2(n20624), .ZN(
        n20308) );
  INV_X1 U23319 ( .A(n20308), .ZN(n20310) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20318), .B1(
        n20317), .B2(n20555), .ZN(n20309) );
  OAI211_X1 U23321 ( .C1(n20558), .C2(n20359), .A(n20310), .B(n20309), .ZN(
        P1_U3102) );
  OAI22_X1 U23322 ( .A1(n20632), .A2(n20315), .B1(n20314), .B2(n20631), .ZN(
        n20311) );
  INV_X1 U23323 ( .A(n20311), .ZN(n20313) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20318), .B1(
        n20317), .B2(n20561), .ZN(n20312) );
  OAI211_X1 U23325 ( .C1(n20564), .C2(n20359), .A(n20313), .B(n20312), .ZN(
        P1_U3103) );
  OAI22_X1 U23326 ( .A1(n20641), .A2(n20315), .B1(n20314), .B2(n20638), .ZN(
        n20316) );
  INV_X1 U23327 ( .A(n20316), .ZN(n20320) );
  AOI22_X1 U23328 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20318), .B1(
        n20317), .B2(n20569), .ZN(n20319) );
  OAI211_X1 U23329 ( .C1(n20574), .C2(n20359), .A(n20320), .B(n20319), .ZN(
        P1_U3104) );
  NOR2_X1 U23330 ( .A1(n20396), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20330) );
  INV_X1 U23331 ( .A(n20330), .ZN(n20321) );
  OR2_X1 U23332 ( .A1(n20471), .A2(n20321), .ZN(n20353) );
  NAND2_X1 U23333 ( .A1(n20399), .A2(n20322), .ZN(n20323) );
  NAND2_X1 U23334 ( .A1(n20323), .A2(n20353), .ZN(n20327) );
  NAND2_X1 U23335 ( .A1(n20327), .A2(n20128), .ZN(n20325) );
  NAND2_X1 U23336 ( .A1(n20330), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20324) );
  AND2_X1 U23337 ( .A1(n20325), .A2(n20324), .ZN(n20352) );
  OAI22_X1 U23338 ( .A1(n20585), .A2(n20353), .B1(n20352), .B2(n20584), .ZN(
        n20326) );
  INV_X1 U23339 ( .A(n20326), .ZN(n20333) );
  INV_X1 U23340 ( .A(n20327), .ZN(n20328) );
  OAI21_X1 U23341 ( .B1(n20742), .B2(n20516), .A(n20328), .ZN(n20329) );
  OAI221_X1 U23342 ( .B1(n20128), .B2(n20330), .C1(n20743), .C2(n20329), .A(
        n20589), .ZN(n20356) );
  AOI22_X1 U23343 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20356), .B1(
        n20355), .B2(n20592), .ZN(n20332) );
  OAI211_X1 U23344 ( .C1(n20595), .C2(n20359), .A(n20333), .B(n20332), .ZN(
        P1_U3105) );
  OAI22_X1 U23345 ( .A1(n20597), .A2(n20353), .B1(n20352), .B2(n20596), .ZN(
        n20334) );
  INV_X1 U23346 ( .A(n20334), .ZN(n20336) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20356), .B1(
        n20355), .B2(n20599), .ZN(n20335) );
  OAI211_X1 U23348 ( .C1(n20602), .C2(n20359), .A(n20336), .B(n20335), .ZN(
        P1_U3106) );
  OAI22_X1 U23349 ( .A1(n20604), .A2(n20353), .B1(n20352), .B2(n20603), .ZN(
        n20337) );
  INV_X1 U23350 ( .A(n20337), .ZN(n20339) );
  AOI22_X1 U23351 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20356), .B1(
        n20355), .B2(n20606), .ZN(n20338) );
  OAI211_X1 U23352 ( .C1(n20609), .C2(n20359), .A(n20339), .B(n20338), .ZN(
        P1_U3107) );
  OAI22_X1 U23353 ( .A1(n20611), .A2(n20353), .B1(n20352), .B2(n20610), .ZN(
        n20340) );
  INV_X1 U23354 ( .A(n20340), .ZN(n20342) );
  AOI22_X1 U23355 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20356), .B1(
        n20355), .B2(n20613), .ZN(n20341) );
  OAI211_X1 U23356 ( .C1(n20616), .C2(n20359), .A(n20342), .B(n20341), .ZN(
        P1_U3108) );
  OAI22_X1 U23357 ( .A1(n20618), .A2(n20353), .B1(n20352), .B2(n20617), .ZN(
        n20343) );
  INV_X1 U23358 ( .A(n20343), .ZN(n20345) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20356), .B1(
        n20355), .B2(n20620), .ZN(n20344) );
  OAI211_X1 U23360 ( .C1(n20623), .C2(n20359), .A(n20345), .B(n20344), .ZN(
        P1_U3109) );
  OAI22_X1 U23361 ( .A1(n20625), .A2(n20353), .B1(n20352), .B2(n20624), .ZN(
        n20346) );
  INV_X1 U23362 ( .A(n20346), .ZN(n20348) );
  AOI22_X1 U23363 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20356), .B1(
        n20355), .B2(n20627), .ZN(n20347) );
  OAI211_X1 U23364 ( .C1(n20630), .C2(n20359), .A(n20348), .B(n20347), .ZN(
        P1_U3110) );
  OAI22_X1 U23365 ( .A1(n20632), .A2(n20353), .B1(n20352), .B2(n20631), .ZN(
        n20349) );
  INV_X1 U23366 ( .A(n20349), .ZN(n20351) );
  AOI22_X1 U23367 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20356), .B1(
        n20355), .B2(n20634), .ZN(n20350) );
  OAI211_X1 U23368 ( .C1(n20637), .C2(n20359), .A(n20351), .B(n20350), .ZN(
        P1_U3111) );
  OAI22_X1 U23369 ( .A1(n20641), .A2(n20353), .B1(n20352), .B2(n20638), .ZN(
        n20354) );
  INV_X1 U23370 ( .A(n20354), .ZN(n20358) );
  AOI22_X1 U23371 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20356), .B1(
        n20355), .B2(n20643), .ZN(n20357) );
  OAI211_X1 U23372 ( .C1(n20649), .C2(n20359), .A(n20358), .B(n20357), .ZN(
        P1_U3112) );
  NOR2_X1 U23373 ( .A1(n20579), .A2(n20396), .ZN(n20407) );
  NAND2_X1 U23374 ( .A1(n20471), .A2(n20407), .ZN(n20389) );
  OAI22_X1 U23375 ( .A1(n20395), .A2(n20595), .B1(n20585), .B2(n20389), .ZN(
        n20360) );
  INV_X1 U23376 ( .A(n20360), .ZN(n20370) );
  NAND2_X1 U23377 ( .A1(n20395), .A2(n20427), .ZN(n20361) );
  AOI21_X1 U23378 ( .B1(n20361), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20743), 
        .ZN(n20365) );
  NAND2_X1 U23379 ( .A1(n20399), .A2(n20518), .ZN(n20367) );
  AOI22_X1 U23380 ( .A1(n20365), .A2(n20367), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20389), .ZN(n20363) );
  OR2_X1 U23381 ( .A1(n20362), .A2(n20746), .ZN(n20509) );
  NAND2_X1 U23382 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20509), .ZN(n20521) );
  NAND3_X1 U23383 ( .A1(n20364), .A2(n20363), .A3(n20521), .ZN(n20392) );
  INV_X1 U23384 ( .A(n20365), .ZN(n20368) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20392), .B1(
        n20514), .B2(n20391), .ZN(n20369) );
  OAI211_X1 U23386 ( .C1(n20528), .C2(n20427), .A(n20370), .B(n20369), .ZN(
        P1_U3113) );
  OAI22_X1 U23387 ( .A1(n20395), .A2(n20602), .B1(n20597), .B2(n20389), .ZN(
        n20371) );
  INV_X1 U23388 ( .A(n20371), .ZN(n20373) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20392), .B1(
        n20529), .B2(n20391), .ZN(n20372) );
  OAI211_X1 U23390 ( .C1(n20534), .C2(n20427), .A(n20373), .B(n20372), .ZN(
        P1_U3114) );
  OAI22_X1 U23391 ( .A1(n20427), .A2(n20540), .B1(n20604), .B2(n20389), .ZN(
        n20374) );
  INV_X1 U23392 ( .A(n20374), .ZN(n20376) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20392), .B1(
        n20535), .B2(n20391), .ZN(n20375) );
  OAI211_X1 U23394 ( .C1(n20609), .C2(n20395), .A(n20376), .B(n20375), .ZN(
        P1_U3115) );
  OAI22_X1 U23395 ( .A1(n20395), .A2(n20616), .B1(n20389), .B2(n20611), .ZN(
        n20377) );
  INV_X1 U23396 ( .A(n20377), .ZN(n20379) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20392), .B1(
        n20541), .B2(n20391), .ZN(n20378) );
  OAI211_X1 U23398 ( .C1(n20546), .C2(n20427), .A(n20379), .B(n20378), .ZN(
        P1_U3116) );
  OAI22_X1 U23399 ( .A1(n20395), .A2(n20623), .B1(n20618), .B2(n20389), .ZN(
        n20380) );
  INV_X1 U23400 ( .A(n20380), .ZN(n20382) );
  AOI22_X1 U23401 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20392), .B1(
        n20547), .B2(n20391), .ZN(n20381) );
  OAI211_X1 U23402 ( .C1(n20552), .C2(n20427), .A(n20382), .B(n20381), .ZN(
        P1_U3117) );
  OAI22_X1 U23403 ( .A1(n20427), .A2(n20558), .B1(n20625), .B2(n20389), .ZN(
        n20383) );
  INV_X1 U23404 ( .A(n20383), .ZN(n20385) );
  AOI22_X1 U23405 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20392), .B1(
        n20553), .B2(n20391), .ZN(n20384) );
  OAI211_X1 U23406 ( .C1(n20630), .C2(n20395), .A(n20385), .B(n20384), .ZN(
        P1_U3118) );
  OAI22_X1 U23407 ( .A1(n20395), .A2(n20637), .B1(n20632), .B2(n20389), .ZN(
        n20386) );
  INV_X1 U23408 ( .A(n20386), .ZN(n20388) );
  AOI22_X1 U23409 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20392), .B1(
        n20559), .B2(n20391), .ZN(n20387) );
  OAI211_X1 U23410 ( .C1(n20564), .C2(n20427), .A(n20388), .B(n20387), .ZN(
        P1_U3119) );
  OAI22_X1 U23411 ( .A1(n20427), .A2(n20574), .B1(n20389), .B2(n20641), .ZN(
        n20390) );
  INV_X1 U23412 ( .A(n20390), .ZN(n20394) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20392), .B1(
        n20566), .B2(n20391), .ZN(n20393) );
  OAI211_X1 U23414 ( .C1(n20649), .C2(n20395), .A(n20394), .B(n20393), .ZN(
        P1_U3120) );
  INV_X1 U23415 ( .A(n20396), .ZN(n20397) );
  NAND2_X1 U23416 ( .A1(n20398), .A2(n20397), .ZN(n20432) );
  NAND2_X1 U23417 ( .A1(n20399), .A2(n20575), .ZN(n20400) );
  NAND2_X1 U23418 ( .A1(n20400), .A2(n20432), .ZN(n20404) );
  INV_X1 U23419 ( .A(n20407), .ZN(n20401) );
  NOR2_X1 U23420 ( .A1(n20401), .A2(n20244), .ZN(n20402) );
  AOI21_X1 U23421 ( .B1(n20404), .B2(n20580), .A(n20402), .ZN(n20431) );
  OAI22_X1 U23422 ( .A1(n20585), .A2(n20432), .B1(n20431), .B2(n20584), .ZN(
        n20403) );
  INV_X1 U23423 ( .A(n20403), .ZN(n20411) );
  INV_X1 U23424 ( .A(n20404), .ZN(n20405) );
  OAI21_X1 U23425 ( .B1(n20742), .B2(n20587), .A(n20405), .ZN(n20406) );
  OAI221_X1 U23426 ( .B1(n20128), .B2(n20407), .C1(n20743), .C2(n20406), .A(
        n20589), .ZN(n20435) );
  AOI22_X1 U23427 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20435), .B1(
        n20440), .B2(n20592), .ZN(n20410) );
  OAI211_X1 U23428 ( .C1(n20595), .C2(n20427), .A(n20411), .B(n20410), .ZN(
        P1_U3121) );
  OAI22_X1 U23429 ( .A1(n20597), .A2(n20432), .B1(n20431), .B2(n20596), .ZN(
        n20412) );
  INV_X1 U23430 ( .A(n20412), .ZN(n20414) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20435), .B1(
        n20440), .B2(n20599), .ZN(n20413) );
  OAI211_X1 U23432 ( .C1(n20602), .C2(n20427), .A(n20414), .B(n20413), .ZN(
        P1_U3122) );
  OAI22_X1 U23433 ( .A1(n20604), .A2(n20432), .B1(n20431), .B2(n20603), .ZN(
        n20415) );
  INV_X1 U23434 ( .A(n20415), .ZN(n20417) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20435), .B1(
        n20440), .B2(n20606), .ZN(n20416) );
  OAI211_X1 U23436 ( .C1(n20609), .C2(n20427), .A(n20417), .B(n20416), .ZN(
        P1_U3123) );
  OAI22_X1 U23437 ( .A1(n20611), .A2(n20432), .B1(n20431), .B2(n20610), .ZN(
        n20418) );
  INV_X1 U23438 ( .A(n20418), .ZN(n20420) );
  INV_X1 U23439 ( .A(n20427), .ZN(n20434) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20435), .B1(
        n20434), .B2(n20543), .ZN(n20419) );
  OAI211_X1 U23441 ( .C1(n20546), .C2(n20469), .A(n20420), .B(n20419), .ZN(
        P1_U3124) );
  OAI22_X1 U23442 ( .A1(n20618), .A2(n20432), .B1(n20431), .B2(n20617), .ZN(
        n20421) );
  INV_X1 U23443 ( .A(n20421), .ZN(n20423) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20435), .B1(
        n20434), .B2(n20549), .ZN(n20422) );
  OAI211_X1 U23445 ( .C1(n20552), .C2(n20469), .A(n20423), .B(n20422), .ZN(
        P1_U3125) );
  OAI22_X1 U23446 ( .A1(n20625), .A2(n20432), .B1(n20431), .B2(n20624), .ZN(
        n20424) );
  INV_X1 U23447 ( .A(n20424), .ZN(n20426) );
  AOI22_X1 U23448 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20435), .B1(
        n20440), .B2(n20627), .ZN(n20425) );
  OAI211_X1 U23449 ( .C1(n20630), .C2(n20427), .A(n20426), .B(n20425), .ZN(
        P1_U3126) );
  OAI22_X1 U23450 ( .A1(n20632), .A2(n20432), .B1(n20431), .B2(n20631), .ZN(
        n20428) );
  INV_X1 U23451 ( .A(n20428), .ZN(n20430) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20435), .B1(
        n20434), .B2(n20561), .ZN(n20429) );
  OAI211_X1 U23453 ( .C1(n20564), .C2(n20469), .A(n20430), .B(n20429), .ZN(
        P1_U3127) );
  OAI22_X1 U23454 ( .A1(n20641), .A2(n20432), .B1(n20431), .B2(n20638), .ZN(
        n20433) );
  INV_X1 U23455 ( .A(n20433), .ZN(n20437) );
  AOI22_X1 U23456 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20435), .B1(
        n20434), .B2(n20569), .ZN(n20436) );
  OAI211_X1 U23457 ( .C1(n20574), .C2(n20469), .A(n20437), .B(n20436), .ZN(
        P1_U3128) );
  AOI22_X1 U23458 ( .A1(n20502), .A2(n20592), .B1(n20515), .B2(n10081), .ZN(
        n20452) );
  NOR3_X1 U23459 ( .A1(n20440), .A2(n20502), .A3(n20743), .ZN(n20442) );
  INV_X1 U23460 ( .A(n20441), .ZN(n20738) );
  NOR2_X1 U23461 ( .A1(n20442), .A2(n20738), .ZN(n20450) );
  INV_X1 U23462 ( .A(n20450), .ZN(n20444) );
  NOR2_X1 U23463 ( .A1(n13262), .A2(n20443), .ZN(n20519) );
  NAND2_X1 U23464 ( .A1(n20519), .A2(n20508), .ZN(n20449) );
  AOI22_X1 U23465 ( .A1(n20444), .A2(n20449), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20448), .ZN(n20445) );
  AOI22_X1 U23466 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20466), .B1(
        n20514), .B2(n20465), .ZN(n20451) );
  OAI211_X1 U23467 ( .C1(n20595), .C2(n20469), .A(n20452), .B(n20451), .ZN(
        P1_U3129) );
  AOI22_X1 U23468 ( .A1(n20502), .A2(n20599), .B1(n20530), .B2(n10081), .ZN(
        n20454) );
  AOI22_X1 U23469 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20466), .B1(
        n20529), .B2(n20465), .ZN(n20453) );
  OAI211_X1 U23470 ( .C1(n20602), .C2(n20469), .A(n20454), .B(n20453), .ZN(
        P1_U3130) );
  AOI22_X1 U23471 ( .A1(n20502), .A2(n20606), .B1(n20536), .B2(n10081), .ZN(
        n20456) );
  AOI22_X1 U23472 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20466), .B1(
        n20535), .B2(n20465), .ZN(n20455) );
  OAI211_X1 U23473 ( .C1(n20609), .C2(n20469), .A(n20456), .B(n20455), .ZN(
        P1_U3131) );
  AOI22_X1 U23474 ( .A1(n20502), .A2(n20613), .B1(n20542), .B2(n10081), .ZN(
        n20458) );
  AOI22_X1 U23475 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20466), .B1(
        n20541), .B2(n20465), .ZN(n20457) );
  OAI211_X1 U23476 ( .C1(n20616), .C2(n20469), .A(n20458), .B(n20457), .ZN(
        P1_U3132) );
  AOI22_X1 U23477 ( .A1(n20502), .A2(n20620), .B1(n20548), .B2(n10081), .ZN(
        n20460) );
  AOI22_X1 U23478 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20466), .B1(
        n20547), .B2(n20465), .ZN(n20459) );
  OAI211_X1 U23479 ( .C1(n20623), .C2(n20469), .A(n20460), .B(n20459), .ZN(
        P1_U3133) );
  AOI22_X1 U23480 ( .A1(n20502), .A2(n20627), .B1(n20554), .B2(n10081), .ZN(
        n20462) );
  AOI22_X1 U23481 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20466), .B1(
        n20553), .B2(n20465), .ZN(n20461) );
  OAI211_X1 U23482 ( .C1(n20630), .C2(n20469), .A(n20462), .B(n20461), .ZN(
        P1_U3134) );
  AOI22_X1 U23483 ( .A1(n20502), .A2(n20634), .B1(n20560), .B2(n10081), .ZN(
        n20464) );
  AOI22_X1 U23484 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20466), .B1(
        n20559), .B2(n20465), .ZN(n20463) );
  OAI211_X1 U23485 ( .C1(n20637), .C2(n20469), .A(n20464), .B(n20463), .ZN(
        P1_U3135) );
  AOI22_X1 U23486 ( .A1(n20502), .A2(n20643), .B1(n20568), .B2(n10081), .ZN(
        n20468) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20466), .B1(
        n20566), .B2(n20465), .ZN(n20467) );
  OAI211_X1 U23488 ( .C1(n20649), .C2(n20469), .A(n20468), .B(n20467), .ZN(
        P1_U3136) );
  NOR3_X1 U23489 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20471), .A3(
        n20578), .ZN(n20472) );
  INV_X1 U23490 ( .A(n20472), .ZN(n20500) );
  NAND2_X1 U23491 ( .A1(n20519), .A2(n20128), .ZN(n20577) );
  OR2_X1 U23492 ( .A1(n20577), .A2(n20023), .ZN(n20474) );
  NOR2_X1 U23493 ( .A1(n20578), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20478) );
  AOI22_X1 U23494 ( .A1(n20580), .A2(n20472), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20478), .ZN(n20473) );
  OAI22_X1 U23495 ( .A1(n20585), .A2(n20500), .B1(n20499), .B2(n20584), .ZN(
        n20475) );
  INV_X1 U23496 ( .A(n20475), .ZN(n20480) );
  INV_X1 U23497 ( .A(n20476), .ZN(n20477) );
  NOR3_X1 U23498 ( .A1(n20477), .A2(n20743), .A3(n20516), .ZN(n20734) );
  OAI21_X1 U23499 ( .B1(n20734), .B2(n20478), .A(n20589), .ZN(n20503) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20525), .ZN(n20479) );
  OAI211_X1 U23501 ( .C1(n20528), .C2(n20524), .A(n20480), .B(n20479), .ZN(
        P1_U3137) );
  OAI22_X1 U23502 ( .A1(n20597), .A2(n20500), .B1(n20499), .B2(n20596), .ZN(
        n20481) );
  INV_X1 U23503 ( .A(n20481), .ZN(n20483) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20531), .ZN(n20482) );
  OAI211_X1 U23505 ( .C1(n20534), .C2(n20524), .A(n20483), .B(n20482), .ZN(
        P1_U3138) );
  OAI22_X1 U23506 ( .A1(n20604), .A2(n20500), .B1(n20499), .B2(n20603), .ZN(
        n20484) );
  INV_X1 U23507 ( .A(n20484), .ZN(n20486) );
  AOI22_X1 U23508 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20537), .ZN(n20485) );
  OAI211_X1 U23509 ( .C1(n20540), .C2(n20524), .A(n20486), .B(n20485), .ZN(
        P1_U3139) );
  OAI22_X1 U23510 ( .A1(n20611), .A2(n20500), .B1(n20499), .B2(n20610), .ZN(
        n20487) );
  INV_X1 U23511 ( .A(n20487), .ZN(n20489) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20543), .ZN(n20488) );
  OAI211_X1 U23513 ( .C1(n20546), .C2(n20524), .A(n20489), .B(n20488), .ZN(
        P1_U3140) );
  OAI22_X1 U23514 ( .A1(n20618), .A2(n20500), .B1(n20499), .B2(n20617), .ZN(
        n20490) );
  INV_X1 U23515 ( .A(n20490), .ZN(n20492) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20549), .ZN(n20491) );
  OAI211_X1 U23517 ( .C1(n20552), .C2(n20524), .A(n20492), .B(n20491), .ZN(
        P1_U3141) );
  OAI22_X1 U23518 ( .A1(n20625), .A2(n20500), .B1(n20499), .B2(n20624), .ZN(
        n20493) );
  INV_X1 U23519 ( .A(n20493), .ZN(n20495) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20555), .ZN(n20494) );
  OAI211_X1 U23521 ( .C1(n20558), .C2(n20524), .A(n20495), .B(n20494), .ZN(
        P1_U3142) );
  OAI22_X1 U23522 ( .A1(n20632), .A2(n20500), .B1(n20499), .B2(n20631), .ZN(
        n20496) );
  INV_X1 U23523 ( .A(n20496), .ZN(n20498) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20561), .ZN(n20497) );
  OAI211_X1 U23525 ( .C1(n20564), .C2(n20524), .A(n20498), .B(n20497), .ZN(
        P1_U3143) );
  OAI22_X1 U23526 ( .A1(n20641), .A2(n20500), .B1(n20499), .B2(n20638), .ZN(
        n20501) );
  INV_X1 U23527 ( .A(n20501), .ZN(n20505) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20569), .ZN(n20504) );
  OAI211_X1 U23529 ( .C1(n20574), .C2(n20524), .A(n20505), .B(n20504), .ZN(
        P1_U3144) );
  INV_X1 U23530 ( .A(n20588), .ZN(n20507) );
  NOR3_X2 U23531 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20579), .A3(
        n20578), .ZN(n20567) );
  OR2_X1 U23532 ( .A1(n20577), .A2(n20508), .ZN(n20513) );
  INV_X1 U23533 ( .A(n20509), .ZN(n20510) );
  NAND2_X1 U23534 ( .A1(n20511), .A2(n20510), .ZN(n20512) );
  NAND2_X1 U23535 ( .A1(n20513), .A2(n20512), .ZN(n20565) );
  AOI22_X1 U23536 ( .A1(n20515), .A2(n20567), .B1(n20514), .B2(n20565), .ZN(
        n20527) );
  AOI21_X1 U23537 ( .B1(n20524), .B2(n20648), .A(n20516), .ZN(n20517) );
  AOI21_X1 U23538 ( .B1(n20519), .B2(n20518), .A(n20517), .ZN(n20520) );
  NOR2_X1 U23539 ( .A1(n20520), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20523) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20525), .ZN(n20526) );
  OAI211_X1 U23541 ( .C1(n20528), .C2(n20648), .A(n20527), .B(n20526), .ZN(
        P1_U3145) );
  AOI22_X1 U23542 ( .A1(n20530), .A2(n20567), .B1(n20529), .B2(n20565), .ZN(
        n20533) );
  AOI22_X1 U23543 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20531), .ZN(n20532) );
  OAI211_X1 U23544 ( .C1(n20534), .C2(n20648), .A(n20533), .B(n20532), .ZN(
        P1_U3146) );
  AOI22_X1 U23545 ( .A1(n20536), .A2(n20567), .B1(n20535), .B2(n20565), .ZN(
        n20539) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20537), .ZN(n20538) );
  OAI211_X1 U23547 ( .C1(n20540), .C2(n20648), .A(n20539), .B(n20538), .ZN(
        P1_U3147) );
  AOI22_X1 U23548 ( .A1(n20542), .A2(n20567), .B1(n20541), .B2(n20565), .ZN(
        n20545) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20543), .ZN(n20544) );
  OAI211_X1 U23550 ( .C1(n20546), .C2(n20648), .A(n20545), .B(n20544), .ZN(
        P1_U3148) );
  AOI22_X1 U23551 ( .A1(n20548), .A2(n20567), .B1(n20547), .B2(n20565), .ZN(
        n20551) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20549), .ZN(n20550) );
  OAI211_X1 U23553 ( .C1(n20552), .C2(n20648), .A(n20551), .B(n20550), .ZN(
        P1_U3149) );
  AOI22_X1 U23554 ( .A1(n20554), .A2(n20567), .B1(n20553), .B2(n20565), .ZN(
        n20557) );
  AOI22_X1 U23555 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20555), .ZN(n20556) );
  OAI211_X1 U23556 ( .C1(n20558), .C2(n20648), .A(n20557), .B(n20556), .ZN(
        P1_U3150) );
  AOI22_X1 U23557 ( .A1(n20560), .A2(n20567), .B1(n20559), .B2(n20565), .ZN(
        n20563) );
  AOI22_X1 U23558 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20561), .ZN(n20562) );
  OAI211_X1 U23559 ( .C1(n20564), .C2(n20648), .A(n20563), .B(n20562), .ZN(
        P1_U3151) );
  AOI22_X1 U23560 ( .A1(n20568), .A2(n20567), .B1(n20566), .B2(n20565), .ZN(
        n20573) );
  AOI22_X1 U23561 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20569), .ZN(n20572) );
  OAI211_X1 U23562 ( .C1(n20574), .C2(n20648), .A(n20573), .B(n20572), .ZN(
        P1_U3152) );
  INV_X1 U23563 ( .A(n20575), .ZN(n20576) );
  OR2_X1 U23564 ( .A1(n20577), .A2(n20576), .ZN(n20583) );
  INV_X1 U23565 ( .A(n20640), .ZN(n20581) );
  NOR2_X1 U23566 ( .A1(n20579), .A2(n20578), .ZN(n20590) );
  AOI22_X1 U23567 ( .A1(n20581), .A2(n20580), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20590), .ZN(n20582) );
  AND2_X1 U23568 ( .A1(n20583), .A2(n20582), .ZN(n20639) );
  OAI22_X1 U23569 ( .A1(n20585), .A2(n20640), .B1(n20639), .B2(n20584), .ZN(
        n20586) );
  INV_X1 U23570 ( .A(n20586), .ZN(n20594) );
  NOR3_X1 U23571 ( .A1(n20588), .A2(n20743), .A3(n20587), .ZN(n20591) );
  OAI21_X1 U23572 ( .B1(n20591), .B2(n20590), .A(n20589), .ZN(n20645) );
  AOI22_X1 U23573 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20592), .ZN(n20593) );
  OAI211_X1 U23574 ( .C1(n20595), .C2(n20648), .A(n20594), .B(n20593), .ZN(
        P1_U3153) );
  OAI22_X1 U23575 ( .A1(n20597), .A2(n20640), .B1(n20639), .B2(n20596), .ZN(
        n20598) );
  INV_X1 U23576 ( .A(n20598), .ZN(n20601) );
  AOI22_X1 U23577 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20599), .ZN(n20600) );
  OAI211_X1 U23578 ( .C1(n20602), .C2(n20648), .A(n20601), .B(n20600), .ZN(
        P1_U3154) );
  OAI22_X1 U23579 ( .A1(n20604), .A2(n20640), .B1(n20639), .B2(n20603), .ZN(
        n20605) );
  INV_X1 U23580 ( .A(n20605), .ZN(n20608) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20606), .ZN(n20607) );
  OAI211_X1 U23582 ( .C1(n20609), .C2(n20648), .A(n20608), .B(n20607), .ZN(
        P1_U3155) );
  OAI22_X1 U23583 ( .A1(n20611), .A2(n20640), .B1(n20639), .B2(n20610), .ZN(
        n20612) );
  INV_X1 U23584 ( .A(n20612), .ZN(n20615) );
  AOI22_X1 U23585 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20613), .ZN(n20614) );
  OAI211_X1 U23586 ( .C1(n20616), .C2(n20648), .A(n20615), .B(n20614), .ZN(
        P1_U3156) );
  OAI22_X1 U23587 ( .A1(n20618), .A2(n20640), .B1(n20639), .B2(n20617), .ZN(
        n20619) );
  INV_X1 U23588 ( .A(n20619), .ZN(n20622) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20620), .ZN(n20621) );
  OAI211_X1 U23590 ( .C1(n20623), .C2(n20648), .A(n20622), .B(n20621), .ZN(
        P1_U3157) );
  OAI22_X1 U23591 ( .A1(n20625), .A2(n20640), .B1(n20639), .B2(n20624), .ZN(
        n20626) );
  INV_X1 U23592 ( .A(n20626), .ZN(n20629) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20627), .ZN(n20628) );
  OAI211_X1 U23594 ( .C1(n20630), .C2(n20648), .A(n20629), .B(n20628), .ZN(
        P1_U3158) );
  OAI22_X1 U23595 ( .A1(n20632), .A2(n20640), .B1(n20639), .B2(n20631), .ZN(
        n20633) );
  INV_X1 U23596 ( .A(n20633), .ZN(n20636) );
  AOI22_X1 U23597 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20634), .ZN(n20635) );
  OAI211_X1 U23598 ( .C1(n20637), .C2(n20648), .A(n20636), .B(n20635), .ZN(
        P1_U3159) );
  OAI22_X1 U23599 ( .A1(n20641), .A2(n20640), .B1(n20639), .B2(n20638), .ZN(
        n20642) );
  INV_X1 U23600 ( .A(n20642), .ZN(n20647) );
  AOI22_X1 U23601 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20645), .B1(
        n20644), .B2(n20643), .ZN(n20646) );
  OAI211_X1 U23602 ( .C1(n20649), .C2(n20648), .A(n20647), .B(n20646), .ZN(
        P1_U3160) );
  NOR2_X1 U23603 ( .A1(n15945), .A2(n20957), .ZN(n20652) );
  INV_X1 U23604 ( .A(n20650), .ZN(n20651) );
  OAI21_X1 U23605 ( .B1(n20652), .B2(n20244), .A(n20651), .ZN(P1_U3163) );
  AND2_X1 U23606 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20720), .ZN(
        P1_U3164) );
  AND2_X1 U23607 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20720), .ZN(
        P1_U3165) );
  AND2_X1 U23608 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20720), .ZN(
        P1_U3166) );
  AND2_X1 U23609 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20720), .ZN(
        P1_U3167) );
  AND2_X1 U23610 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20720), .ZN(
        P1_U3168) );
  AND2_X1 U23611 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20720), .ZN(
        P1_U3169) );
  AND2_X1 U23612 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20720), .ZN(
        P1_U3170) );
  AND2_X1 U23613 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20720), .ZN(
        P1_U3171) );
  AND2_X1 U23614 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20720), .ZN(
        P1_U3172) );
  AND2_X1 U23615 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20720), .ZN(
        P1_U3173) );
  AND2_X1 U23616 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20720), .ZN(
        P1_U3174) );
  AND2_X1 U23617 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20720), .ZN(
        P1_U3175) );
  AND2_X1 U23618 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20720), .ZN(
        P1_U3176) );
  AND2_X1 U23619 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20720), .ZN(
        P1_U3177) );
  AND2_X1 U23620 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20720), .ZN(
        P1_U3178) );
  AND2_X1 U23621 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20720), .ZN(
        P1_U3179) );
  AND2_X1 U23622 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20720), .ZN(
        P1_U3180) );
  AND2_X1 U23623 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20720), .ZN(
        P1_U3181) );
  AND2_X1 U23624 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20720), .ZN(
        P1_U3182) );
  INV_X1 U23625 ( .A(P1_DATAWIDTH_REG_12__SCAN_IN), .ZN(n21034) );
  NOR2_X1 U23626 ( .A1(n20724), .A2(n21034), .ZN(P1_U3183) );
  AND2_X1 U23627 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20720), .ZN(
        P1_U3184) );
  AND2_X1 U23628 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20720), .ZN(
        P1_U3185) );
  AND2_X1 U23629 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20720), .ZN(P1_U3186) );
  AND2_X1 U23630 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20720), .ZN(P1_U3187) );
  INV_X1 U23631 ( .A(P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20824) );
  NOR2_X1 U23632 ( .A1(n20724), .A2(n20824), .ZN(P1_U3188) );
  AND2_X1 U23633 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20720), .ZN(P1_U3189) );
  AND2_X1 U23634 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20720), .ZN(P1_U3190) );
  AND2_X1 U23635 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20720), .ZN(P1_U3191) );
  AND2_X1 U23636 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20720), .ZN(P1_U3192) );
  AND2_X1 U23637 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20720), .ZN(P1_U3193) );
  NAND2_X1 U23638 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20959), .ZN(n20658) );
  INV_X1 U23639 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20664) );
  NOR2_X1 U23640 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_1__SCAN_IN), 
        .ZN(n20653) );
  OAI22_X1 U23641 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20654), .B1(n20653), 
        .B2(n20668), .ZN(n20655) );
  OAI21_X1 U23642 ( .B1(n20664), .B2(n20655), .A(n20770), .ZN(n20656) );
  OAI211_X1 U23643 ( .C1(n20658), .C2(n20760), .A(n20657), .B(n20656), .ZN(
        P1_U3194) );
  NOR2_X1 U23644 ( .A1(NA), .A2(n20663), .ZN(n20659) );
  AOI21_X1 U23645 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20659), .A(
        P1_STATE_REG_2__SCAN_IN), .ZN(n20670) );
  AOI21_X1 U23646 ( .B1(NA), .B2(n20660), .A(P1_STATE_REG_0__SCAN_IN), .ZN(
        n20661) );
  AOI21_X1 U23647 ( .B1(n20662), .B2(P1_STATE_REG_1__SCAN_IN), .A(n20661), 
        .ZN(n20669) );
  NOR3_X1 U23648 ( .A1(NA), .A2(n20663), .A3(n20760), .ZN(n20665) );
  OAI22_X1 U23649 ( .A1(n20666), .A2(n20665), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20664), .ZN(n20667) );
  OAI22_X1 U23650 ( .A1(n20670), .A2(n20669), .B1(n20668), .B2(n20667), .ZN(
        P1_U3196) );
  OR2_X1 U23651 ( .A1(n20770), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20706) );
  INV_X1 U23652 ( .A(n20706), .ZN(n20712) );
  AOI222_X1 U23653 ( .A1(n20712), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20713), .ZN(n20671) );
  INV_X1 U23654 ( .A(n20671), .ZN(P1_U3197) );
  AOI222_X1 U23655 ( .A1(n20713), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20712), .ZN(n20672) );
  INV_X1 U23656 ( .A(n20672), .ZN(P1_U3198) );
  INV_X1 U23657 ( .A(n20713), .ZN(n20709) );
  OAI222_X1 U23658 ( .A1(n20709), .A2(n13486), .B1(n20674), .B2(n20769), .C1(
        n20673), .C2(n20706), .ZN(P1_U3199) );
  AOI222_X1 U23659 ( .A1(n20712), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20713), .ZN(n20675) );
  INV_X1 U23660 ( .A(n20675), .ZN(P1_U3200) );
  AOI22_X1 U23661 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20712), .ZN(n20676) );
  OAI21_X1 U23662 ( .B1(n20677), .B2(n20709), .A(n20676), .ZN(P1_U3201) );
  AOI22_X1 U23663 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20712), .ZN(n20678) );
  OAI21_X1 U23664 ( .B1(n20679), .B2(n20709), .A(n20678), .ZN(P1_U3202) );
  AOI22_X1 U23665 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20713), .ZN(n20680) );
  OAI21_X1 U23666 ( .B1(n20681), .B2(n20706), .A(n20680), .ZN(P1_U3203) );
  AOI222_X1 U23667 ( .A1(n20713), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n20712), .ZN(n20682) );
  INV_X1 U23668 ( .A(n20682), .ZN(P1_U3204) );
  AOI222_X1 U23669 ( .A1(n20713), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20712), .ZN(n20683) );
  INV_X1 U23670 ( .A(n20683), .ZN(P1_U3205) );
  AOI222_X1 U23671 ( .A1(n20712), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20713), .ZN(n20684) );
  INV_X1 U23672 ( .A(n20684), .ZN(P1_U3206) );
  AOI22_X1 U23673 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20712), .ZN(n20685) );
  OAI21_X1 U23674 ( .B1(n20686), .B2(n20709), .A(n20685), .ZN(P1_U3207) );
  AOI22_X1 U23675 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20713), .ZN(n20687) );
  OAI21_X1 U23676 ( .B1(n14167), .B2(n20706), .A(n20687), .ZN(P1_U3208) );
  AOI222_X1 U23677 ( .A1(n20713), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20712), .ZN(n20688) );
  INV_X1 U23678 ( .A(n20688), .ZN(P1_U3209) );
  AOI222_X1 U23679 ( .A1(n20712), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20713), .ZN(n20689) );
  INV_X1 U23680 ( .A(n20689), .ZN(P1_U3210) );
  AOI222_X1 U23681 ( .A1(n20713), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20712), .ZN(n20690) );
  INV_X1 U23682 ( .A(n20690), .ZN(P1_U3211) );
  AOI22_X1 U23683 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20712), .ZN(n20691) );
  OAI21_X1 U23684 ( .B1(n20692), .B2(n20709), .A(n20691), .ZN(P1_U3212) );
  AOI22_X1 U23685 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20713), .ZN(n20693) );
  OAI21_X1 U23686 ( .B1(n20694), .B2(n20706), .A(n20693), .ZN(P1_U3213) );
  AOI222_X1 U23687 ( .A1(n20713), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20712), .ZN(n20695) );
  INV_X1 U23688 ( .A(n20695), .ZN(P1_U3214) );
  AOI222_X1 U23689 ( .A1(n20713), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20712), .ZN(n20696) );
  INV_X1 U23690 ( .A(n20696), .ZN(P1_U3215) );
  AOI22_X1 U23691 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(n20712), .ZN(n20697) );
  OAI21_X1 U23692 ( .B1(n20698), .B2(n20709), .A(n20697), .ZN(P1_U3216) );
  AOI22_X1 U23693 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(n20713), .ZN(n20699) );
  OAI21_X1 U23694 ( .B1(n14939), .B2(n20706), .A(n20699), .ZN(P1_U3217) );
  AOI22_X1 U23695 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20712), .ZN(n20700) );
  OAI21_X1 U23696 ( .B1(n14939), .B2(n20709), .A(n20700), .ZN(P1_U3218) );
  AOI22_X1 U23697 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20713), .ZN(n20701) );
  OAI21_X1 U23698 ( .B1(n20702), .B2(n20706), .A(n20701), .ZN(P1_U3219) );
  AOI222_X1 U23699 ( .A1(n20713), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20712), .ZN(n20703) );
  INV_X1 U23700 ( .A(n20703), .ZN(P1_U3220) );
  AOI222_X1 U23701 ( .A1(n20713), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20712), .ZN(n20704) );
  INV_X1 U23702 ( .A(n20704), .ZN(P1_U3221) );
  AOI222_X1 U23703 ( .A1(n20713), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20712), .ZN(n20705) );
  INV_X1 U23704 ( .A(n20705), .ZN(P1_U3222) );
  INV_X1 U23705 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20998) );
  OAI222_X1 U23706 ( .A1(n20709), .A2(n20708), .B1(n20998), .B2(n20769), .C1(
        n20707), .C2(n20706), .ZN(P1_U3223) );
  AOI222_X1 U23707 ( .A1(n20713), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20712), .ZN(n20710) );
  INV_X1 U23708 ( .A(n20710), .ZN(P1_U3224) );
  AOI222_X1 U23709 ( .A1(n20712), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20713), .ZN(n20711) );
  INV_X1 U23710 ( .A(n20711), .ZN(P1_U3225) );
  AOI222_X1 U23711 ( .A1(n20713), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20712), .ZN(n20714) );
  INV_X1 U23712 ( .A(n20714), .ZN(P1_U3226) );
  OAI22_X1 U23713 ( .A1(n20770), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20769), .ZN(n20715) );
  INV_X1 U23714 ( .A(n20715), .ZN(P1_U3458) );
  OAI22_X1 U23715 ( .A1(n20770), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20769), .ZN(n20716) );
  INV_X1 U23716 ( .A(n20716), .ZN(P1_U3459) );
  OAI22_X1 U23717 ( .A1(n20770), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20769), .ZN(n20717) );
  INV_X1 U23718 ( .A(n20717), .ZN(P1_U3460) );
  OAI22_X1 U23719 ( .A1(n20770), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20769), .ZN(n20718) );
  INV_X1 U23720 ( .A(n20718), .ZN(P1_U3461) );
  INV_X1 U23721 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20721) );
  INV_X1 U23722 ( .A(n20722), .ZN(n20719) );
  AOI21_X1 U23723 ( .B1(n20721), .B2(n20720), .A(n20719), .ZN(P1_U3464) );
  OAI21_X1 U23724 ( .B1(n20724), .B2(n20723), .A(n20722), .ZN(P1_U3465) );
  INV_X1 U23725 ( .A(n20725), .ZN(n20729) );
  OAI22_X1 U23726 ( .A1(n20729), .A2(n20728), .B1(n20727), .B2(n20726), .ZN(
        n20731) );
  MUX2_X1 U23727 ( .A(n20732), .B(n20731), .S(n20730), .Z(P1_U3469) );
  NOR2_X1 U23728 ( .A1(n20734), .A2(n20733), .ZN(n20741) );
  INV_X1 U23729 ( .A(n20735), .ZN(n20739) );
  AOI22_X1 U23730 ( .A1(n20739), .A2(n20738), .B1(n20737), .B2(n20736), .ZN(
        n20740) );
  OAI211_X1 U23731 ( .C1(n20743), .C2(n20742), .A(n20741), .B(n20740), .ZN(
        n20744) );
  NAND2_X1 U23732 ( .A1(n20747), .A2(n20744), .ZN(n20745) );
  OAI21_X1 U23733 ( .B1(n20747), .B2(n20746), .A(n20745), .ZN(P1_U3475) );
  AOI21_X1 U23734 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20749) );
  AOI22_X1 U23735 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20749), .B2(n20748), .ZN(n20751) );
  INV_X1 U23736 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20750) );
  AOI22_X1 U23737 ( .A1(n20752), .A2(n20751), .B1(n20750), .B2(n20755), .ZN(
        P1_U3481) );
  INV_X1 U23738 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20756) );
  NOR2_X1 U23739 ( .A1(n20755), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20753) );
  AOI22_X1 U23740 ( .A1(n20756), .A2(n20755), .B1(n20754), .B2(n20753), .ZN(
        P1_U3482) );
  INV_X1 U23741 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20757) );
  AOI22_X1 U23742 ( .A1(n20769), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20757), 
        .B2(n20770), .ZN(P1_U3483) );
  AOI211_X1 U23743 ( .C1(n13187), .C2(n20760), .A(n20759), .B(n20758), .ZN(
        n20768) );
  OAI211_X1 U23744 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20763), .A(n20762), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20765) );
  AOI21_X1 U23745 ( .B1(n20765), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20764), 
        .ZN(n20767) );
  NAND2_X1 U23746 ( .A1(n20768), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20766) );
  OAI21_X1 U23747 ( .B1(n20768), .B2(n20767), .A(n20766), .ZN(P1_U3485) );
  OAI22_X1 U23748 ( .A1(n20770), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n20769), .ZN(n20771) );
  INV_X1 U23749 ( .A(n20771), .ZN(P1_U3486) );
  NOR4_X1 U23750 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_0__4__SCAN_IN), .A3(P1_INSTQUEUE_REG_3__3__SCAN_IN), 
        .A4(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n20772) );
  NAND3_X1 U23751 ( .A1(n20772), .A2(n20923), .A3(n12062), .ZN(n20781) );
  NAND4_X1 U23752 ( .A1(DATAI_4_), .A2(P1_DATAO_REG_21__SCAN_IN), .A3(
        P1_DATAO_REG_29__SCAN_IN), .A4(P1_DATAO_REG_5__SCAN_IN), .ZN(n20773)
         );
  NOR3_X1 U23753 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20966), .A3(
        n20773), .ZN(n20779) );
  NAND4_X1 U23754 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n20777) );
  NAND4_X1 U23755 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(
        P3_DATAO_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_M_IO_N_REG_SCAN_IN), .ZN(n20776) );
  NAND4_X1 U23756 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(P2_LWORD_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(
        n20775) );
  NAND4_X1 U23757 ( .A1(P2_EAX_REG_13__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .A3(P1_EBX_REG_28__SCAN_IN), .A4(P1_UWORD_REG_6__SCAN_IN), .ZN(n20774)
         );
  NOR4_X1 U23758 ( .A1(n20777), .A2(n20776), .A3(n20775), .A4(n20774), .ZN(
        n20778) );
  NAND4_X1 U23759 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_BYTEENABLE_REG_3__SCAN_IN), .A3(n20779), .A4(n20778), .ZN(n20780)
         );
  NOR4_X1 U23760 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n20781), .A4(n20780), .ZN(
        n20814) );
  NAND4_X1 U23761 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(BUF2_REG_27__SCAN_IN), .ZN(
        n20785) );
  NAND4_X1 U23762 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A4(P3_D_C_N_REG_SCAN_IN), .ZN(
        n20784) );
  NAND4_X1 U23763 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_EAX_REG_12__SCAN_IN), .A3(P1_EBX_REG_18__SCAN_IN), .A4(
        P1_REIP_REG_30__SCAN_IN), .ZN(n20783) );
  NAND4_X1 U23764 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_15__3__SCAN_IN), .A3(P1_INSTQUEUE_REG_9__6__SCAN_IN), 
        .A4(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n20782) );
  NOR4_X1 U23765 ( .A1(n20785), .A2(n20784), .A3(n20783), .A4(n20782), .ZN(
        n20813) );
  NAND4_X1 U23766 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .A3(P3_INSTQUEUE_REG_14__2__SCAN_IN), 
        .A4(P3_UWORD_REG_2__SCAN_IN), .ZN(n20789) );
  NAND4_X1 U23767 ( .A1(READY22_REG_SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_LWORD_REG_14__SCAN_IN), .A4(P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(
        n20788) );
  NAND4_X1 U23768 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .A4(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n20787) );
  NAND4_X1 U23769 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_1__2__SCAN_IN), .A3(P3_INSTQUEUE_REG_0__6__SCAN_IN), 
        .A4(P3_REIP_REG_20__SCAN_IN), .ZN(n20786) );
  NOR4_X1 U23770 ( .A1(n20789), .A2(n20788), .A3(n20787), .A4(n20786), .ZN(
        n20812) );
  NOR4_X1 U23771 ( .A1(P1_BYTEENABLE_REG_1__SCAN_IN), .A2(
        P3_ADDRESS_REG_14__SCAN_IN), .A3(P3_ADDRESS_REG_8__SCAN_IN), .A4(
        P3_LWORD_REG_10__SCAN_IN), .ZN(n20793) );
  NOR4_X1 U23772 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(P3_DATAO_REG_17__SCAN_IN), .A3(P3_UWORD_REG_1__SCAN_IN), .A4(P1_LWORD_REG_14__SCAN_IN), .ZN(n20792) );
  NOR4_X1 U23773 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P1_EAX_REG_2__SCAN_IN), .A3(P1_EAX_REG_7__SCAN_IN), .A4(
        P2_READREQUEST_REG_SCAN_IN), .ZN(n20791) );
  NOR4_X1 U23774 ( .A1(DATAI_0_), .A2(P3_LWORD_REG_9__SCAN_IN), .A3(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A4(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(
        n20790) );
  NAND4_X1 U23775 ( .A1(n20793), .A2(n20792), .A3(n20791), .A4(n20790), .ZN(
        n20810) );
  INV_X1 U23776 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n21045) );
  NOR4_X1 U23777 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_10__3__SCAN_IN), .A3(P2_INSTQUEUE_REG_8__3__SCAN_IN), 
        .A4(n21045), .ZN(n20798) );
  NOR4_X1 U23778 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_7__5__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), 
        .A4(P1_DATAO_REG_7__SCAN_IN), .ZN(n20797) );
  NOR4_X1 U23779 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_10__4__SCAN_IN), .A3(P2_INSTQUEUE_REG_13__4__SCAN_IN), 
        .A4(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20794) );
  NAND3_X1 U23780 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20794), .A3(
        P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n20795) );
  NOR3_X1 U23781 ( .A1(n20795), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A3(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20796) );
  NAND3_X1 U23782 ( .A1(n20798), .A2(n20797), .A3(n20796), .ZN(n20809) );
  NOR4_X1 U23783 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A3(P3_EBX_REG_16__SCAN_IN), .A4(
        P3_EBX_REG_9__SCAN_IN), .ZN(n20802) );
  NOR4_X1 U23784 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(
        P3_EBX_REG_19__SCAN_IN), .A3(P3_EBX_REG_13__SCAN_IN), .A4(
        P3_EBX_REG_0__SCAN_IN), .ZN(n20801) );
  NOR4_X1 U23785 ( .A1(P2_EAX_REG_28__SCAN_IN), .A2(BUF2_REG_30__SCAN_IN), 
        .A3(P1_STATE2_REG_1__SCAN_IN), .A4(BUF1_REG_19__SCAN_IN), .ZN(n20800)
         );
  NOR4_X1 U23786 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(P2_REIP_REG_8__SCAN_IN), .A4(
        P3_EBX_REG_25__SCAN_IN), .ZN(n20799) );
  NAND4_X1 U23787 ( .A1(n20802), .A2(n20801), .A3(n20800), .A4(n20799), .ZN(
        n20808) );
  NOR4_X1 U23788 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A3(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A4(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20806) );
  NOR4_X1 U23789 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(BUF1_REG_14__SCAN_IN), 
        .A3(P2_LWORD_REG_5__SCAN_IN), .A4(P2_UWORD_REG_4__SCAN_IN), .ZN(n20805) );
  NOR4_X1 U23790 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .A3(P3_INSTQUEUE_REG_0__1__SCAN_IN), 
        .A4(P3_EAX_REG_22__SCAN_IN), .ZN(n20804) );
  NOR4_X1 U23791 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A4(P3_EAX_REG_5__SCAN_IN), .ZN(
        n20803) );
  NAND4_X1 U23792 ( .A1(n20806), .A2(n20805), .A3(n20804), .A4(n20803), .ZN(
        n20807) );
  NOR4_X1 U23793 ( .A1(n20810), .A2(n20809), .A3(n20808), .A4(n20807), .ZN(
        n20811) );
  NAND4_X1 U23794 ( .A1(n20814), .A2(n20813), .A3(n20812), .A4(n20811), .ZN(
        n21091) );
  AOI22_X1 U23795 ( .A1(n20817), .A2(keyinput17), .B1(keyinput125), .B2(n20816), .ZN(n20815) );
  OAI221_X1 U23796 ( .B1(n20817), .B2(keyinput17), .C1(n20816), .C2(
        keyinput125), .A(n20815), .ZN(n20828) );
  AOI22_X1 U23797 ( .A1(n20819), .A2(keyinput4), .B1(n12045), .B2(keyinput116), 
        .ZN(n20818) );
  OAI221_X1 U23798 ( .B1(n20819), .B2(keyinput4), .C1(n12045), .C2(keyinput116), .A(n20818), .ZN(n20827) );
  AOI22_X1 U23799 ( .A1(n20822), .A2(keyinput88), .B1(n20821), .B2(keyinput74), 
        .ZN(n20820) );
  OAI221_X1 U23800 ( .B1(n20822), .B2(keyinput88), .C1(n20821), .C2(keyinput74), .A(n20820), .ZN(n20826) );
  AOI22_X1 U23801 ( .A1(n14685), .A2(keyinput108), .B1(keyinput72), .B2(n20824), .ZN(n20823) );
  OAI221_X1 U23802 ( .B1(n14685), .B2(keyinput108), .C1(n20824), .C2(
        keyinput72), .A(n20823), .ZN(n20825) );
  NOR4_X1 U23803 ( .A1(n20828), .A2(n20827), .A3(n20826), .A4(n20825), .ZN(
        n20881) );
  AOI22_X1 U23804 ( .A1(n13344), .A2(keyinput25), .B1(keyinput113), .B2(n20830), .ZN(n20829) );
  OAI221_X1 U23805 ( .B1(n13344), .B2(keyinput25), .C1(n20830), .C2(
        keyinput113), .A(n20829), .ZN(n20833) );
  INV_X1 U23806 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n20831) );
  XNOR2_X1 U23807 ( .A(n20831), .B(keyinput43), .ZN(n20832) );
  NOR2_X1 U23808 ( .A1(n20833), .A2(n20832), .ZN(n20845) );
  AOI22_X1 U23809 ( .A1(n20836), .A2(keyinput61), .B1(n20835), .B2(keyinput10), 
        .ZN(n20834) );
  OAI221_X1 U23810 ( .B1(n20836), .B2(keyinput61), .C1(n20835), .C2(keyinput10), .A(n20834), .ZN(n20837) );
  INV_X1 U23811 ( .A(n20837), .ZN(n20844) );
  AOI22_X1 U23812 ( .A1(n20840), .A2(keyinput86), .B1(keyinput127), .B2(n20839), .ZN(n20838) );
  OAI221_X1 U23813 ( .B1(n20840), .B2(keyinput86), .C1(n20839), .C2(
        keyinput127), .A(n20838), .ZN(n20841) );
  INV_X1 U23814 ( .A(n20841), .ZN(n20843) );
  XNOR2_X1 U23815 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B(keyinput90), .ZN(
        n20842) );
  AND4_X1 U23816 ( .A1(n20845), .A2(n20844), .A3(n20843), .A4(n20842), .ZN(
        n20880) );
  AOI22_X1 U23817 ( .A1(n20848), .A2(keyinput98), .B1(n20847), .B2(keyinput111), .ZN(n20846) );
  OAI221_X1 U23818 ( .B1(n20848), .B2(keyinput98), .C1(n20847), .C2(
        keyinput111), .A(n20846), .ZN(n20861) );
  AOI22_X1 U23819 ( .A1(n20851), .A2(keyinput68), .B1(keyinput6), .B2(n20850), 
        .ZN(n20849) );
  OAI221_X1 U23820 ( .B1(n20851), .B2(keyinput68), .C1(n20850), .C2(keyinput6), 
        .A(n20849), .ZN(n20860) );
  AOI22_X1 U23821 ( .A1(n20854), .A2(keyinput38), .B1(n20853), .B2(keyinput14), 
        .ZN(n20852) );
  OAI221_X1 U23822 ( .B1(n20854), .B2(keyinput38), .C1(n20853), .C2(keyinput14), .A(n20852), .ZN(n20859) );
  AOI22_X1 U23823 ( .A1(n20857), .A2(keyinput55), .B1(keyinput71), .B2(n20856), 
        .ZN(n20855) );
  OAI221_X1 U23824 ( .B1(n20857), .B2(keyinput55), .C1(n20856), .C2(keyinput71), .A(n20855), .ZN(n20858) );
  NOR4_X1 U23825 ( .A1(n20861), .A2(n20860), .A3(n20859), .A4(n20858), .ZN(
        n20879) );
  INV_X1 U23826 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n20863) );
  AOI22_X1 U23827 ( .A1(n20864), .A2(keyinput59), .B1(keyinput21), .B2(n20863), 
        .ZN(n20862) );
  OAI221_X1 U23828 ( .B1(n20864), .B2(keyinput59), .C1(n20863), .C2(keyinput21), .A(n20862), .ZN(n20877) );
  AOI22_X1 U23829 ( .A1(n20867), .A2(keyinput94), .B1(keyinput79), .B2(n20866), 
        .ZN(n20865) );
  OAI221_X1 U23830 ( .B1(n20867), .B2(keyinput94), .C1(n20866), .C2(keyinput79), .A(n20865), .ZN(n20876) );
  AOI22_X1 U23831 ( .A1(n20870), .A2(keyinput28), .B1(n20869), .B2(keyinput84), 
        .ZN(n20868) );
  OAI221_X1 U23832 ( .B1(n20870), .B2(keyinput28), .C1(n20869), .C2(keyinput84), .A(n20868), .ZN(n20875) );
  AOI22_X1 U23833 ( .A1(n20873), .A2(keyinput12), .B1(n20872), .B2(keyinput92), 
        .ZN(n20871) );
  OAI221_X1 U23834 ( .B1(n20873), .B2(keyinput12), .C1(n20872), .C2(keyinput92), .A(n20871), .ZN(n20874) );
  NOR4_X1 U23835 ( .A1(n20877), .A2(n20876), .A3(n20875), .A4(n20874), .ZN(
        n20878) );
  NAND4_X1 U23836 ( .A1(n20881), .A2(n20880), .A3(n20879), .A4(n20878), .ZN(
        n21076) );
  INV_X1 U23837 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n20884) );
  AOI22_X1 U23838 ( .A1(n20884), .A2(keyinput67), .B1(keyinput1), .B2(n20883), 
        .ZN(n20882) );
  OAI221_X1 U23839 ( .B1(n20884), .B2(keyinput67), .C1(n20883), .C2(keyinput1), 
        .A(n20882), .ZN(n20897) );
  AOI22_X1 U23840 ( .A1(n20887), .A2(keyinput54), .B1(n20886), .B2(keyinput101), .ZN(n20885) );
  OAI221_X1 U23841 ( .B1(n20887), .B2(keyinput54), .C1(n20886), .C2(
        keyinput101), .A(n20885), .ZN(n20896) );
  AOI22_X1 U23842 ( .A1(n20890), .A2(keyinput0), .B1(n20889), .B2(keyinput83), 
        .ZN(n20888) );
  OAI221_X1 U23843 ( .B1(n20890), .B2(keyinput0), .C1(n20889), .C2(keyinput83), 
        .A(n20888), .ZN(n20895) );
  INV_X1 U23844 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n20893) );
  AOI22_X1 U23845 ( .A1(n20893), .A2(keyinput118), .B1(keyinput35), .B2(n20892), .ZN(n20891) );
  OAI221_X1 U23846 ( .B1(n20893), .B2(keyinput118), .C1(n20892), .C2(
        keyinput35), .A(n20891), .ZN(n20894) );
  NOR4_X1 U23847 ( .A1(n20897), .A2(n20896), .A3(n20895), .A4(n20894), .ZN(
        n20948) );
  INV_X1 U23848 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n20899) );
  AOI22_X1 U23849 ( .A1(n20900), .A2(keyinput62), .B1(n20899), .B2(keyinput97), 
        .ZN(n20898) );
  OAI221_X1 U23850 ( .B1(n20900), .B2(keyinput62), .C1(n20899), .C2(keyinput97), .A(n20898), .ZN(n20913) );
  AOI22_X1 U23851 ( .A1(n20903), .A2(keyinput119), .B1(keyinput66), .B2(n20902), .ZN(n20901) );
  OAI221_X1 U23852 ( .B1(n20903), .B2(keyinput119), .C1(n20902), .C2(
        keyinput66), .A(n20901), .ZN(n20912) );
  INV_X1 U23853 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n20906) );
  AOI22_X1 U23854 ( .A1(n20906), .A2(keyinput96), .B1(keyinput9), .B2(n20905), 
        .ZN(n20904) );
  OAI221_X1 U23855 ( .B1(n20906), .B2(keyinput96), .C1(n20905), .C2(keyinput9), 
        .A(n20904), .ZN(n20911) );
  AOI22_X1 U23856 ( .A1(n20909), .A2(keyinput33), .B1(n20908), .B2(keyinput75), 
        .ZN(n20907) );
  OAI221_X1 U23857 ( .B1(n20909), .B2(keyinput33), .C1(n20908), .C2(keyinput75), .A(n20907), .ZN(n20910) );
  NOR4_X1 U23858 ( .A1(n20913), .A2(n20912), .A3(n20911), .A4(n20910), .ZN(
        n20947) );
  INV_X1 U23859 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n20916) );
  AOI22_X1 U23860 ( .A1(n20916), .A2(keyinput120), .B1(keyinput122), .B2(
        n20915), .ZN(n20914) );
  OAI221_X1 U23861 ( .B1(n20916), .B2(keyinput120), .C1(n20915), .C2(
        keyinput122), .A(n20914), .ZN(n20928) );
  AOI22_X1 U23862 ( .A1(n20918), .A2(keyinput80), .B1(n10824), .B2(keyinput112), .ZN(n20917) );
  OAI221_X1 U23863 ( .B1(n20918), .B2(keyinput80), .C1(n10824), .C2(
        keyinput112), .A(n20917), .ZN(n20927) );
  AOI22_X1 U23864 ( .A1(n20921), .A2(keyinput22), .B1(keyinput110), .B2(n20920), .ZN(n20919) );
  OAI221_X1 U23865 ( .B1(n20921), .B2(keyinput22), .C1(n20920), .C2(
        keyinput110), .A(n20919), .ZN(n20926) );
  AOI22_X1 U23866 ( .A1(n20924), .A2(keyinput44), .B1(n20923), .B2(keyinput13), 
        .ZN(n20922) );
  OAI221_X1 U23867 ( .B1(n20924), .B2(keyinput44), .C1(n20923), .C2(keyinput13), .A(n20922), .ZN(n20925) );
  NOR4_X1 U23868 ( .A1(n20928), .A2(n20927), .A3(n20926), .A4(n20925), .ZN(
        n20946) );
  AOI22_X1 U23869 ( .A1(n20931), .A2(keyinput106), .B1(keyinput117), .B2(
        n20930), .ZN(n20929) );
  OAI221_X1 U23870 ( .B1(n20931), .B2(keyinput106), .C1(n20930), .C2(
        keyinput117), .A(n20929), .ZN(n20944) );
  AOI22_X1 U23871 ( .A1(n20934), .A2(keyinput63), .B1(n20933), .B2(keyinput42), 
        .ZN(n20932) );
  OAI221_X1 U23872 ( .B1(n20934), .B2(keyinput63), .C1(n20933), .C2(keyinput42), .A(n20932), .ZN(n20938) );
  XNOR2_X1 U23873 ( .A(n20935), .B(keyinput65), .ZN(n20937) );
  XOR2_X1 U23874 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B(keyinput26), .Z(
        n20936) );
  OR3_X1 U23875 ( .A1(n20938), .A2(n20937), .A3(n20936), .ZN(n20943) );
  INV_X1 U23876 ( .A(DATAI_0_), .ZN(n20941) );
  AOI22_X1 U23877 ( .A1(n20941), .A2(keyinput76), .B1(keyinput20), .B2(n20940), 
        .ZN(n20939) );
  OAI221_X1 U23878 ( .B1(n20941), .B2(keyinput76), .C1(n20940), .C2(keyinput20), .A(n20939), .ZN(n20942) );
  NOR3_X1 U23879 ( .A1(n20944), .A2(n20943), .A3(n20942), .ZN(n20945) );
  NAND4_X1 U23880 ( .A1(n20948), .A2(n20947), .A3(n20946), .A4(n20945), .ZN(
        n21075) );
  INV_X1 U23881 ( .A(P3_D_C_N_REG_SCAN_IN), .ZN(n20950) );
  AOI22_X1 U23882 ( .A1(n20951), .A2(keyinput39), .B1(keyinput60), .B2(n20950), 
        .ZN(n20949) );
  OAI221_X1 U23883 ( .B1(n20951), .B2(keyinput39), .C1(n20950), .C2(keyinput60), .A(n20949), .ZN(n20963) );
  AOI22_X1 U23884 ( .A1(n20954), .A2(keyinput124), .B1(n20953), .B2(keyinput3), 
        .ZN(n20952) );
  OAI221_X1 U23885 ( .B1(n20954), .B2(keyinput124), .C1(n20953), .C2(keyinput3), .A(n20952), .ZN(n20962) );
  AOI22_X1 U23886 ( .A1(n20957), .A2(keyinput100), .B1(keyinput109), .B2(
        n20956), .ZN(n20955) );
  OAI221_X1 U23887 ( .B1(n20957), .B2(keyinput100), .C1(n20956), .C2(
        keyinput109), .A(n20955), .ZN(n20961) );
  AOI22_X1 U23888 ( .A1(n10731), .A2(keyinput89), .B1(keyinput52), .B2(n20959), 
        .ZN(n20958) );
  OAI221_X1 U23889 ( .B1(n10731), .B2(keyinput89), .C1(n20959), .C2(keyinput52), .A(n20958), .ZN(n20960) );
  NOR4_X1 U23890 ( .A1(n20963), .A2(n20962), .A3(n20961), .A4(n20960), .ZN(
        n21010) );
  AOI22_X1 U23891 ( .A1(n10814), .A2(keyinput49), .B1(keyinput18), .B2(n11556), 
        .ZN(n20964) );
  OAI221_X1 U23892 ( .B1(n10814), .B2(keyinput49), .C1(n11556), .C2(keyinput18), .A(n20964), .ZN(n20977) );
  AOI22_X1 U23893 ( .A1(n20967), .A2(keyinput115), .B1(n20966), .B2(keyinput53), .ZN(n20965) );
  OAI221_X1 U23894 ( .B1(n20967), .B2(keyinput115), .C1(n20966), .C2(
        keyinput53), .A(n20965), .ZN(n20976) );
  INV_X1 U23895 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n20969) );
  AOI22_X1 U23896 ( .A1(n20970), .A2(keyinput36), .B1(n20969), .B2(keyinput16), 
        .ZN(n20968) );
  OAI221_X1 U23897 ( .B1(n20970), .B2(keyinput36), .C1(n20969), .C2(keyinput16), .A(n20968), .ZN(n20975) );
  AOI22_X1 U23898 ( .A1(n20973), .A2(keyinput32), .B1(keyinput70), .B2(n20972), 
        .ZN(n20971) );
  OAI221_X1 U23899 ( .B1(n20973), .B2(keyinput32), .C1(n20972), .C2(keyinput70), .A(n20971), .ZN(n20974) );
  NOR4_X1 U23900 ( .A1(n20977), .A2(n20976), .A3(n20975), .A4(n20974), .ZN(
        n21009) );
  INV_X1 U23901 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n20980) );
  AOI22_X1 U23902 ( .A1(n20980), .A2(keyinput77), .B1(keyinput40), .B2(n20979), 
        .ZN(n20978) );
  OAI221_X1 U23903 ( .B1(n20980), .B2(keyinput77), .C1(n20979), .C2(keyinput40), .A(n20978), .ZN(n20984) );
  XOR2_X1 U23904 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B(keyinput47), .Z(
        n20983) );
  XNOR2_X1 U23905 ( .A(n20981), .B(keyinput104), .ZN(n20982) );
  OR3_X1 U23906 ( .A1(n20984), .A2(n20983), .A3(n20982), .ZN(n20993) );
  AOI22_X1 U23907 ( .A1(n20987), .A2(keyinput103), .B1(n20986), .B2(keyinput93), .ZN(n20985) );
  OAI221_X1 U23908 ( .B1(n20987), .B2(keyinput103), .C1(n20986), .C2(
        keyinput93), .A(n20985), .ZN(n20992) );
  INV_X1 U23909 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n20990) );
  AOI22_X1 U23910 ( .A1(n20990), .A2(keyinput11), .B1(n20989), .B2(keyinput27), 
        .ZN(n20988) );
  OAI221_X1 U23911 ( .B1(n20990), .B2(keyinput11), .C1(n20989), .C2(keyinput27), .A(n20988), .ZN(n20991) );
  NOR3_X1 U23912 ( .A1(n20993), .A2(n20992), .A3(n20991), .ZN(n21008) );
  INV_X1 U23913 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20995) );
  AOI22_X1 U23914 ( .A1(n9862), .A2(keyinput37), .B1(keyinput29), .B2(n20995), 
        .ZN(n20994) );
  OAI221_X1 U23915 ( .B1(n9862), .B2(keyinput37), .C1(n20995), .C2(keyinput29), 
        .A(n20994), .ZN(n21006) );
  AOI22_X1 U23916 ( .A1(n20998), .A2(keyinput69), .B1(keyinput64), .B2(n20997), 
        .ZN(n20996) );
  OAI221_X1 U23917 ( .B1(n20998), .B2(keyinput69), .C1(n20997), .C2(keyinput64), .A(n20996), .ZN(n21005) );
  INV_X1 U23918 ( .A(DATAI_4_), .ZN(n21000) );
  AOI22_X1 U23919 ( .A1(n12062), .A2(keyinput31), .B1(keyinput57), .B2(n21000), 
        .ZN(n20999) );
  OAI221_X1 U23920 ( .B1(n12062), .B2(keyinput31), .C1(n21000), .C2(keyinput57), .A(n20999), .ZN(n21004) );
  INV_X1 U23921 ( .A(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n21002) );
  AOI22_X1 U23922 ( .A1(n10799), .A2(keyinput19), .B1(keyinput46), .B2(n21002), 
        .ZN(n21001) );
  OAI221_X1 U23923 ( .B1(n10799), .B2(keyinput19), .C1(n21002), .C2(keyinput46), .A(n21001), .ZN(n21003) );
  NOR4_X1 U23924 ( .A1(n21006), .A2(n21005), .A3(n21004), .A4(n21003), .ZN(
        n21007) );
  NAND4_X1 U23925 ( .A1(n21010), .A2(n21009), .A3(n21008), .A4(n21007), .ZN(
        n21074) );
  AOI22_X1 U23926 ( .A1(n21013), .A2(keyinput81), .B1(keyinput102), .B2(n21012), .ZN(n21011) );
  OAI221_X1 U23927 ( .B1(n21013), .B2(keyinput81), .C1(n21012), .C2(
        keyinput102), .A(n21011), .ZN(n21023) );
  AOI22_X1 U23928 ( .A1(n21015), .A2(keyinput2), .B1(n13709), .B2(keyinput24), 
        .ZN(n21014) );
  OAI221_X1 U23929 ( .B1(n21015), .B2(keyinput2), .C1(n13709), .C2(keyinput24), 
        .A(n21014), .ZN(n21022) );
  AOI22_X1 U23930 ( .A1(n11020), .A2(keyinput73), .B1(keyinput99), .B2(n11917), 
        .ZN(n21016) );
  OAI221_X1 U23931 ( .B1(n11020), .B2(keyinput73), .C1(n11917), .C2(keyinput99), .A(n21016), .ZN(n21021) );
  INV_X1 U23932 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n21019) );
  AOI22_X1 U23933 ( .A1(n21019), .A2(keyinput56), .B1(keyinput45), .B2(n21018), 
        .ZN(n21017) );
  OAI221_X1 U23934 ( .B1(n21019), .B2(keyinput56), .C1(n21018), .C2(keyinput45), .A(n21017), .ZN(n21020) );
  NOR4_X1 U23935 ( .A1(n21023), .A2(n21022), .A3(n21021), .A4(n21020), .ZN(
        n21072) );
  AOI22_X1 U23936 ( .A1(n21026), .A2(keyinput107), .B1(keyinput78), .B2(n21025), .ZN(n21024) );
  OAI221_X1 U23937 ( .B1(n21026), .B2(keyinput107), .C1(n21025), .C2(
        keyinput78), .A(n21024), .ZN(n21039) );
  AOI22_X1 U23938 ( .A1(n21029), .A2(keyinput23), .B1(keyinput41), .B2(n21028), 
        .ZN(n21027) );
  OAI221_X1 U23939 ( .B1(n21029), .B2(keyinput23), .C1(n21028), .C2(keyinput41), .A(n21027), .ZN(n21038) );
  INV_X1 U23940 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n21032) );
  INV_X1 U23941 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n21031) );
  AOI22_X1 U23942 ( .A1(n21032), .A2(keyinput82), .B1(keyinput5), .B2(n21031), 
        .ZN(n21030) );
  OAI221_X1 U23943 ( .B1(n21032), .B2(keyinput82), .C1(n21031), .C2(keyinput5), 
        .A(n21030), .ZN(n21037) );
  AOI22_X1 U23944 ( .A1(n21035), .A2(keyinput121), .B1(keyinput123), .B2(
        n21034), .ZN(n21033) );
  OAI221_X1 U23945 ( .B1(n21035), .B2(keyinput121), .C1(n21034), .C2(
        keyinput123), .A(n21033), .ZN(n21036) );
  NOR4_X1 U23946 ( .A1(n21039), .A2(n21038), .A3(n21037), .A4(n21036), .ZN(
        n21071) );
  AOI22_X1 U23947 ( .A1(n15122), .A2(keyinput91), .B1(n10939), .B2(keyinput105), .ZN(n21040) );
  OAI221_X1 U23948 ( .B1(n15122), .B2(keyinput91), .C1(n10939), .C2(
        keyinput105), .A(n21040), .ZN(n21053) );
  INV_X1 U23949 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n21042) );
  AOI22_X1 U23950 ( .A1(n21043), .A2(keyinput7), .B1(n21042), .B2(keyinput48), 
        .ZN(n21041) );
  OAI221_X1 U23951 ( .B1(n21043), .B2(keyinput7), .C1(n21042), .C2(keyinput48), 
        .A(n21041), .ZN(n21052) );
  AOI22_X1 U23952 ( .A1(n21046), .A2(keyinput30), .B1(n21045), .B2(keyinput95), 
        .ZN(n21044) );
  OAI221_X1 U23953 ( .B1(n21046), .B2(keyinput30), .C1(n21045), .C2(keyinput95), .A(n21044), .ZN(n21051) );
  AOI22_X1 U23954 ( .A1(n21049), .A2(keyinput87), .B1(n21048), .B2(keyinput51), 
        .ZN(n21047) );
  OAI221_X1 U23955 ( .B1(n21049), .B2(keyinput87), .C1(n21048), .C2(keyinput51), .A(n21047), .ZN(n21050) );
  NOR4_X1 U23956 ( .A1(n21053), .A2(n21052), .A3(n21051), .A4(n21050), .ZN(
        n21070) );
  AOI22_X1 U23957 ( .A1(n21056), .A2(keyinput126), .B1(n21055), .B2(keyinput50), .ZN(n21054) );
  OAI221_X1 U23958 ( .B1(n21056), .B2(keyinput126), .C1(n21055), .C2(
        keyinput50), .A(n21054), .ZN(n21068) );
  INV_X1 U23959 ( .A(READY22_REG_SCAN_IN), .ZN(n21058) );
  AOI22_X1 U23960 ( .A1(n21059), .A2(keyinput8), .B1(keyinput15), .B2(n21058), 
        .ZN(n21057) );
  OAI221_X1 U23961 ( .B1(n21059), .B2(keyinput8), .C1(n21058), .C2(keyinput15), 
        .A(n21057), .ZN(n21067) );
  INV_X1 U23962 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n21061) );
  AOI22_X1 U23963 ( .A1(n21061), .A2(keyinput85), .B1(keyinput114), .B2(n14507), .ZN(n21060) );
  OAI221_X1 U23964 ( .B1(n21061), .B2(keyinput85), .C1(n14507), .C2(
        keyinput114), .A(n21060), .ZN(n21066) );
  AOI22_X1 U23965 ( .A1(n21064), .A2(keyinput58), .B1(n21063), .B2(keyinput34), 
        .ZN(n21062) );
  OAI221_X1 U23966 ( .B1(n21064), .B2(keyinput58), .C1(n21063), .C2(keyinput34), .A(n21062), .ZN(n21065) );
  NOR4_X1 U23967 ( .A1(n21068), .A2(n21067), .A3(n21066), .A4(n21065), .ZN(
        n21069) );
  NAND4_X1 U23968 ( .A1(n21072), .A2(n21071), .A3(n21070), .A4(n21069), .ZN(
        n21073) );
  NOR4_X1 U23969 ( .A1(n21076), .A2(n21075), .A3(n21074), .A4(n21073), .ZN(
        n21089) );
  AOI22_X1 U23970 ( .A1(n21080), .A2(n21079), .B1(n21078), .B2(n21077), .ZN(
        n21085) );
  AOI22_X1 U23971 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n21083), .B1(
        n21082), .B2(n21081), .ZN(n21084) );
  OAI211_X1 U23972 ( .C1(n21087), .C2(n21086), .A(n21085), .B(n21084), .ZN(
        n21088) );
  XOR2_X1 U23973 ( .A(n21089), .B(n21088), .Z(n21090) );
  XNOR2_X1 U23974 ( .A(n21091), .B(n21090), .ZN(P2_U3093) );
  INV_X1 U11279 ( .A(n10204), .ZN(n10596) );
  NAND2_X2 U11286 ( .A1(n10161), .A2(n10162), .ZN(n10558) );
  BUF_X1 U11239 ( .A(n14301), .Z(n9707) );
  NAND2_X1 U11248 ( .A1(n10241), .A2(n10240), .ZN(n10247) );
  BUF_X2 U11158 ( .A(n11654), .Z(n13069) );
  BUF_X2 U11160 ( .A(n12403), .Z(n17048) );
  BUF_X2 U11164 ( .A(n12543), .Z(n16740) );
  NAND2_X1 U11175 ( .A1(n11393), .A2(n11392), .ZN(n11402) );
  CLKBUF_X1 U11198 ( .A(n9721), .Z(n13073) );
  CLKBUF_X1 U11206 ( .A(n10353), .Z(n14300) );
  CLKBUF_X1 U11210 ( .A(n10382), .Z(n14293) );
  CLKBUF_X1 U11250 ( .A(n12224), .Z(n13633) );
  CLKBUF_X1 U11267 ( .A(n10684), .Z(n10701) );
  CLKBUF_X1 U11269 ( .A(n15408), .Z(n16031) );
  CLKBUF_X1 U11283 ( .A(n15438), .Z(n9727) );
  AND3_X1 U11461 ( .A1(n10195), .A2(n10212), .A3(n10208), .ZN(n10176) );
  CLKBUF_X2 U11526 ( .A(n14495), .Z(n11771) );
  NAND4_X1 U11607 ( .A1(n11261), .A2(n11260), .A3(n11259), .A4(n11258), .ZN(
        n11271) );
  CLKBUF_X1 U11608 ( .A(n12213), .Z(n13548) );
  CLKBUF_X1 U11636 ( .A(n14970), .Z(n9766) );
  BUF_X2 U12388 ( .A(n10204), .Z(n9763) );
  CLKBUF_X1 U12439 ( .A(n10212), .Z(n13724) );
  CLKBUF_X1 U12796 ( .A(n11929), .Z(n20089) );
  CLKBUF_X1 U12890 ( .A(n16336), .Z(n16345) );
endmodule

