

module b21_C_SARLock_k_128_7 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4409, n4410, n4411, n4413, n4414, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10230;

  AOI21_X1 U4915 ( .B1(n9310), .B2(n9471), .A(n4725), .ZN(n4724) );
  INV_X1 U4916 ( .A(n7705), .ZN(n8538) );
  NAND2_X1 U4917 ( .A1(n6781), .A2(n6780), .ZN(n7002) );
  INV_X1 U4918 ( .A(n7674), .ZN(n7665) );
  NAND4_X1 U4919 ( .A1(n5784), .A2(n5783), .A3(n5782), .A4(n5781), .ZN(n6057)
         );
  CLKBUF_X1 U4920 ( .A(n7370), .Z(n4416) );
  AND4_X1 U4921 ( .A1(n5199), .A2(n5198), .A3(n5197), .A4(n5196), .ZN(n6424)
         );
  CLKBUF_X2 U4922 ( .A(n5223), .Z(n7674) );
  INV_X2 U4923 ( .A(n7314), .ZN(n7324) );
  NAND2_X1 U4926 ( .A1(n5130), .A2(n5129), .ZN(n7214) );
  INV_X4 U4927 ( .A(n9281), .ZN(n4419) );
  OAI211_X1 U4931 ( .C1(n6513), .C2(n8099), .A(n5316), .B(n5315), .ZN(n7062)
         );
  OR2_X1 U4932 ( .A1(n9322), .A2(n9097), .ZN(n7467) );
  CLKBUF_X2 U4933 ( .A(n6348), .Z(n7450) );
  OAI21_X1 U4934 ( .B1(n7448), .B2(n7223), .A(n7222), .ZN(n7226) );
  NAND2_X1 U4936 ( .A1(n8528), .A2(n7835), .ZN(n7705) );
  CLKBUF_X2 U4937 ( .A(n6394), .Z(n8004) );
  INV_X1 U4938 ( .A(n7998), .ZN(n8005) );
  INV_X1 U4939 ( .A(n7370), .ZN(n7456) );
  NAND2_X1 U4940 ( .A1(n7498), .A2(n7408), .ZN(n6231) );
  AND2_X1 U4941 ( .A1(n7612), .A2(n8214), .ZN(n9115) );
  OAI21_X1 U4942 ( .B1(n5502), .B2(n4878), .A(n4875), .ZN(n5534) );
  NAND2_X1 U4943 ( .A1(n5417), .A2(n5416), .ZN(n8848) );
  AND4_X1 U4944 ( .A1(n5216), .A2(n5215), .A3(n5214), .A4(n5213), .ZN(n6487)
         );
  INV_X1 U4945 ( .A(n8546), .ZN(n7711) );
  NAND2_X1 U4946 ( .A1(n5151), .A2(n5150), .ZN(n8883) );
  NAND2_X1 U4947 ( .A1(n7012), .A2(n7011), .ZN(n8914) );
  XNOR2_X1 U4948 ( .A(n5653), .B(n5652), .ZN(n7242) );
  NOR2_X1 U4949 ( .A1(n5794), .A2(n5793), .ZN(n9529) );
  AOI211_X1 U4950 ( .C1(n9727), .C2(n8782), .A(n8518), .B(n8517), .ZN(n8519)
         );
  INV_X1 U4951 ( .A(n5140), .ZN(n5702) );
  AOI211_X1 U4952 ( .C1(n9650), .C2(n9318), .A(n8223), .B(n8222), .ZN(n8224)
         );
  NAND2_X1 U4953 ( .A1(n5771), .A2(n4961), .ZN(n9419) );
  NOR2_X2 U4954 ( .A1(n6586), .A2(n8892), .ZN(n4730) );
  NOR2_X2 U4955 ( .A1(n6057), .A2(n6194), .ZN(n6187) );
  NAND2_X4 U4956 ( .A1(n5146), .A2(n6834), .ZN(n5200) );
  NAND3_X2 U4957 ( .A1(n5190), .A2(n5189), .A3(n5188), .ZN(n6275) );
  OAI211_X4 U4958 ( .C1(n7674), .C2(n5845), .A(n4672), .B(n4671), .ZN(n6270)
         );
  AND2_X4 U4959 ( .A1(n4654), .A2(n4653), .ZN(n7229) );
  INV_X4 U4960 ( .A(n7229), .ZN(n5844) );
  INV_X4 U4961 ( .A(n7229), .ZN(n7220) );
  AND2_X1 U4962 ( .A1(n5168), .A2(n8232), .ZN(n4409) );
  CLKBUF_X1 U4963 ( .A(n5212), .Z(n4410) );
  OAI222_X1 U4964 ( .A1(P2_U3152), .A2(n8232), .B1(n8236), .B2(n8234), .C1(
        n8233), .C2(n8881), .ZN(P2_U3328) );
  BUF_X2 U4965 ( .A(n6319), .Z(n4411) );
  NOR4_X2 U4966 ( .A1(n7493), .A2(n9095), .A3(n9129), .A4(n7492), .ZN(n7495)
         );
  INV_X1 U4967 ( .A(n10230), .ZN(n4413) );
  AND2_X1 U4970 ( .A1(n9419), .A2(n5772), .ZN(n7370) );
  AND4_X1 U4971 ( .A1(n4436), .A2(n7853), .A3(n7852), .A4(n7851), .ZN(n7858)
         );
  AND2_X1 U4972 ( .A1(n8853), .A2(n7191), .ZN(n8712) );
  AOI21_X1 U4973 ( .B1(n4752), .B2(n7697), .A(n4750), .ZN(n4749) );
  NAND2_X2 U4974 ( .A1(n7796), .A2(n7797), .ZN(n8711) );
  OAI21_X1 U4975 ( .B1(n6634), .B2(n6633), .A(n5301), .ZN(n6773) );
  INV_X1 U4976 ( .A(n6886), .ZN(n9783) );
  NAND2_X2 U4977 ( .A1(n7746), .A2(n6977), .ZN(n7685) );
  INV_X1 U4978 ( .A(n6501), .ZN(n4677) );
  NAND2_X1 U4979 ( .A1(n6226), .A2(n8930), .ZN(n7498) );
  NAND2_X1 U4980 ( .A1(n6487), .A2(n4421), .ZN(n7745) );
  BUF_X1 U4981 ( .A(n6924), .Z(n4421) );
  INV_X1 U4982 ( .A(n4411), .ZN(n7885) );
  INV_X1 U4983 ( .A(n9053), .ZN(n6226) );
  AND4_X2 U4984 ( .A1(n5180), .A2(n5179), .A3(n5178), .A4(n5177), .ZN(n6271)
         );
  INV_X2 U4985 ( .A(n5195), .ZN(n5393) );
  INV_X1 U4986 ( .A(n5195), .ZN(n4418) );
  INV_X1 U4987 ( .A(n7728), .ZN(n6680) );
  INV_X1 U4988 ( .A(n9419), .ZN(n5773) );
  AND2_X1 U4989 ( .A1(n8232), .A2(n8227), .ZN(n5212) );
  NAND2_X1 U4990 ( .A1(n5152), .A2(n8883), .ZN(n8227) );
  MUX2_X1 U4991 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5149), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5152) );
  MUX2_X1 U4992 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5128), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5130) );
  OR2_X1 U4993 ( .A1(n4674), .A2(n5355), .ZN(n4439) );
  INV_X1 U4994 ( .A(n4932), .ZN(n4728) );
  AND2_X1 U4995 ( .A1(n5793), .A2(n5748), .ZN(n4727) );
  NOR2_X1 U4996 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5740) );
  AOI21_X1 U4997 ( .B1(n8220), .B2(n9296), .A(n4511), .ZN(n9320) );
  AND2_X1 U4998 ( .A1(n8246), .A2(n8247), .ZN(n8301) );
  NAND2_X1 U4999 ( .A1(n4776), .A2(n8538), .ZN(n8541) );
  INV_X1 U5000 ( .A(n7521), .ZN(n9311) );
  NAND2_X1 U5001 ( .A1(n7676), .A2(n7675), .ZN(n8761) );
  NAND2_X1 U5002 ( .A1(n7234), .A2(n7233), .ZN(n7521) );
  AOI21_X1 U5003 ( .B1(n4777), .B2(n7705), .A(n4775), .ZN(n4774) );
  OAI21_X1 U5004 ( .B1(n9106), .B2(n8187), .A(n4942), .ZN(n9092) );
  NAND2_X1 U5005 ( .A1(n8603), .A2(n8602), .ZN(n8601) );
  OR2_X1 U5006 ( .A1(n8787), .A2(n8275), .ZN(n7839) );
  NAND2_X1 U5007 ( .A1(n5641), .A2(n5640), .ZN(n8781) );
  XNOR2_X1 U5008 ( .A(n7217), .B(n7216), .ZN(n8235) );
  NAND2_X1 U5009 ( .A1(n7258), .A2(n7257), .ZN(n9332) );
  OAI21_X1 U5010 ( .B1(n8380), .B2(n8813), .A(n7196), .ZN(n8581) );
  NAND2_X1 U5011 ( .A1(n4845), .A2(n5654), .ZN(n7217) );
  OR2_X1 U5012 ( .A1(n8792), .A2(n8561), .ZN(n8528) );
  OR2_X1 U5013 ( .A1(n8796), .A2(n8570), .ZN(n7198) );
  NAND2_X1 U5014 ( .A1(n5614), .A2(n5613), .ZN(n5634) );
  NAND2_X1 U5015 ( .A1(n5565), .A2(n5114), .ZN(n5591) );
  NAND2_X1 U5016 ( .A1(n5113), .A2(n5112), .ZN(n5565) );
  OR2_X1 U5017 ( .A1(n9218), .A2(n9368), .ZN(n9184) );
  OAI22_X1 U5018 ( .A1(n8712), .A2(n4822), .B1(n4823), .B2(n7193), .ZN(n8683)
         );
  NAND2_X1 U5019 ( .A1(n7037), .A2(n7486), .ZN(n7036) );
  AND2_X1 U5020 ( .A1(n7015), .A2(n7387), .ZN(n7037) );
  NAND2_X1 U5021 ( .A1(n4611), .A2(n4612), .ZN(n9452) );
  OAI21_X1 U5022 ( .B1(n7114), .B2(n7698), .A(n7115), .ZN(n7116) );
  NAND2_X1 U5023 ( .A1(n7320), .A2(n7319), .ZN(n9377) );
  AND2_X1 U5024 ( .A1(n7694), .A2(n7056), .ZN(n7094) );
  NAND2_X1 U5025 ( .A1(n5088), .A2(n5087), .ZN(n5502) );
  NAND2_X1 U5026 ( .A1(n9731), .A2(n9730), .ZN(n9729) );
  NAND2_X1 U5027 ( .A1(n5484), .A2(n5085), .ZN(n5088) );
  OR2_X1 U5028 ( .A1(n8914), .A2(n9033), .ZN(n8195) );
  NAND2_X1 U5029 ( .A1(n7384), .A2(n7383), .ZN(n9391) );
  AND2_X1 U5030 ( .A1(n7695), .A2(n7123), .ZN(n7124) );
  AND2_X1 U5031 ( .A1(n7768), .A2(n7771), .ZN(n7692) );
  NAND2_X1 U5032 ( .A1(n5079), .A2(n5078), .ZN(n5463) );
  OR2_X1 U5033 ( .A1(n6376), .A2(n7479), .ZN(n6562) );
  NAND2_X1 U5034 ( .A1(n5369), .A2(n5368), .ZN(n8855) );
  NAND2_X1 U5035 ( .A1(n6932), .A2(n6931), .ZN(n7386) );
  NAND2_X1 U5036 ( .A1(n6693), .A2(n6692), .ZN(n6859) );
  NAND2_X1 U5037 ( .A1(n5365), .A2(n4992), .ZN(n5063) );
  NAND2_X1 U5038 ( .A1(n6647), .A2(n6646), .ZN(n9649) );
  AND2_X1 U5039 ( .A1(n7759), .A2(n7753), .ZN(n8735) );
  NAND2_X1 U5040 ( .A1(n5335), .A2(n4438), .ZN(n5047) );
  OAI21_X2 U5041 ( .B1(n5313), .B2(n4871), .A(n4868), .ZN(n5335) );
  OR2_X1 U5042 ( .A1(n5314), .A2(n6354), .ZN(n5296) );
  NAND2_X1 U5043 ( .A1(n6186), .A2(n5787), .ZN(n7407) );
  NAND2_X1 U5044 ( .A1(n7723), .A2(n7745), .ZN(n7734) );
  NAND2_X1 U5045 ( .A1(n5026), .A2(n5025), .ZN(n5294) );
  INV_X1 U5046 ( .A(n6185), .ZN(n7473) );
  AND2_X1 U5047 ( .A1(n4605), .A2(n4604), .ZN(n6225) );
  INV_X2 U5048 ( .A(n7683), .ZN(n6450) );
  AND4_X1 U5049 ( .A1(n5255), .A2(n5254), .A3(n5253), .A4(n5252), .ZN(n6875)
         );
  AND4_X1 U5050 ( .A1(n5235), .A2(n5234), .A3(n5233), .A4(n5232), .ZN(n6872)
         );
  AND2_X2 U5051 ( .A1(n5878), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NAND4_X1 U5052 ( .A1(n5814), .A2(n5813), .A3(n5812), .A4(n5811), .ZN(n9053)
         );
  AND3_X1 U5053 ( .A1(n4953), .A2(n4954), .A3(n4949), .ZN(n4952) );
  NAND4_X1 U5054 ( .A1(n5791), .A2(n5790), .A3(n5789), .A4(n5788), .ZN(n9054)
         );
  OAI211_X1 U5055 ( .C1(n6513), .C2(n9444), .A(n5207), .B(n5206), .ZN(n6319)
         );
  NAND2_X2 U5056 ( .A1(n5702), .A2(n6680), .ZN(n9763) );
  AOI21_X1 U5057 ( .B1(n4856), .B2(n4437), .A(n4855), .ZN(n4854) );
  NAND2_X1 U5058 ( .A1(n6513), .A2(n5844), .ZN(n5223) );
  CLKBUF_X3 U5059 ( .A(n5211), .Z(n5644) );
  AND2_X2 U5060 ( .A1(n5772), .A2(n5773), .ZN(n7459) );
  NAND2_X2 U5061 ( .A1(n4780), .A2(n8227), .ZN(n5195) );
  NAND2_X1 U5062 ( .A1(n5010), .A2(n5009), .ZN(n5221) );
  NAND2_X4 U5063 ( .A1(n5721), .A2(n7214), .ZN(n6513) );
  NAND2_X1 U5064 ( .A1(n4997), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5675) );
  XNOR2_X1 U5065 ( .A(n5142), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7728) );
  INV_X2 U5066 ( .A(n6105), .ZN(n7382) );
  NAND2_X1 U5067 ( .A1(n6105), .A2(n5844), .ZN(n6644) );
  INV_X1 U5068 ( .A(n5772), .ZN(n8229) );
  OR2_X1 U5069 ( .A1(n5141), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n4997) );
  XNOR2_X1 U5070 ( .A(n5769), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U5071 ( .A1(n8883), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5153) );
  CLKBUF_X1 U5072 ( .A(n5809), .Z(n9536) );
  OR2_X1 U5073 ( .A1(n5151), .A2(n5126), .ZN(n5149) );
  NAND2_X1 U5074 ( .A1(n4961), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5769) );
  NOR2_X1 U5075 ( .A1(n5485), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5134) );
  XNOR2_X1 U5076 ( .A(n5764), .B(n5768), .ZN(n5809) );
  NAND2_X1 U5077 ( .A1(n5767), .A2(n5766), .ZN(n9532) );
  NAND2_X2 U5078 ( .A1(n5844), .A2(P1_U3084), .ZN(n9424) );
  NAND2_X2 U5079 ( .A1(n7229), .A2(P2_U3152), .ZN(n8236) );
  AND2_X1 U5080 ( .A1(n4818), .A2(n5125), .ZN(n4673) );
  AND2_X1 U5081 ( .A1(n4981), .A2(n4837), .ZN(n4836) );
  NAND4_X1 U5082 ( .A1(n4443), .A2(n4931), .A3(n5741), .A4(n5740), .ZN(n4932)
         );
  AND3_X1 U5083 ( .A1(n4427), .A2(n4424), .A3(n4486), .ZN(n4726) );
  AND4_X1 U5084 ( .A1(n4927), .A2(n10122), .A3(n5895), .A4(n5729), .ZN(n4424)
         );
  AND2_X1 U5085 ( .A1(n5739), .A2(n5734), .ZN(n4931) );
  AND4_X1 U5086 ( .A1(n5733), .A2(n5732), .A3(n5731), .A4(n5730), .ZN(n4427)
         );
  AND2_X1 U5087 ( .A1(n5119), .A2(n4838), .ZN(n4837) );
  AND2_X1 U5088 ( .A1(n5118), .A2(n4819), .ZN(n4818) );
  INV_X4 U5089 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U5090 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5895) );
  NOR2_X1 U5091 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5115) );
  INV_X1 U5092 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5734) );
  NOR2_X1 U5093 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5667) );
  NOR2_X1 U5094 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5731) );
  NOR2_X1 U5095 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5732) );
  INV_X1 U5096 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10122) );
  NOR2_X1 U5097 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4927) );
  NOR2_X1 U5098 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5133) );
  INV_X4 U5099 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U5100 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4657) );
  INV_X1 U5101 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6221) );
  NOR2_X1 U5102 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5741) );
  NOR2_X1 U5103 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4991) );
  NOR3_X1 U5104 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .A3(
        P2_IR_REG_10__SCAN_IN), .ZN(n5118) );
  INV_X1 U5105 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5729) );
  NOR2_X1 U5106 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5116) );
  OR2_X1 U5107 ( .A1(n5222), .A2(n5853), .ZN(n4672) );
  OAI211_X2 U5108 ( .C1(n7220), .C2(P1_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n5002), .ZN(n5003) );
  NAND2_X2 U5109 ( .A1(n7089), .A2(n7782), .ZN(n7110) );
  AND2_X1 U5110 ( .A1(n6105), .A2(n7229), .ZN(n6348) );
  OAI21_X2 U5111 ( .B1(n8555), .B2(n4831), .A(n4828), .ZN(n8521) );
  INV_X1 U5112 ( .A(n7229), .ZN(n4420) );
  AND2_X4 U5113 ( .A1(n5168), .A2(n8232), .ZN(n5248) );
  XNOR2_X2 U5114 ( .A(n5153), .B(n8880), .ZN(n8232) );
  NOR2_X1 U5115 ( .A1(n7581), .A2(n7580), .ZN(n7586) );
  NAND2_X1 U5116 ( .A1(n5069), .A2(n5068), .ZN(n5072) );
  OR2_X1 U5117 ( .A1(n7873), .A2(n7668), .ZN(n7849) );
  OR2_X1 U5118 ( .A1(n8776), .A2(n8494), .ZN(n7847) );
  NOR2_X1 U5119 ( .A1(n8590), .A2(n4765), .ZN(n4764) );
  INV_X1 U5120 ( .A(n7820), .ZN(n4765) );
  OR2_X1 U5121 ( .A1(n8818), .A2(n8257), .ZN(n7816) );
  AND2_X1 U5122 ( .A1(n4991), .A2(n4781), .ZN(n4981) );
  NOR2_X1 U5123 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n4781) );
  NAND2_X1 U5124 ( .A1(n8813), .A2(n8380), .ZN(n7195) );
  INV_X1 U5125 ( .A(n7792), .ZN(n4753) );
  NAND2_X1 U5126 ( .A1(n7534), .A2(n4706), .ZN(n4705) );
  AOI21_X1 U5127 ( .B1(n7533), .B2(n7627), .A(n7535), .ZN(n4707) );
  NAND2_X1 U5128 ( .A1(n4644), .A2(n4643), .ZN(n7819) );
  NOR2_X1 U5129 ( .A1(n7808), .A2(n8636), .ZN(n4643) );
  NAND2_X1 U5130 ( .A1(n4646), .A2(n4645), .ZN(n4644) );
  AND2_X1 U5131 ( .A1(n7552), .A2(n7554), .ZN(n4712) );
  NAND2_X1 U5132 ( .A1(n4710), .A2(n4709), .ZN(n4708) );
  INV_X1 U5133 ( .A(n9289), .ZN(n4709) );
  INV_X1 U5134 ( .A(n7568), .ZN(n4710) );
  NOR2_X1 U5135 ( .A1(n7585), .A2(n4706), .ZN(n4722) );
  NAND2_X1 U5136 ( .A1(n8192), .A2(n9089), .ZN(n4874) );
  INV_X1 U5137 ( .A(n5040), .ZN(n4869) );
  INV_X1 U5138 ( .A(n8255), .ZN(n5513) );
  AND2_X1 U5139 ( .A1(n7161), .A2(n7156), .ZN(n5406) );
  OAI21_X1 U5140 ( .B1(n7858), .B2(n7857), .A(n4449), .ZN(n4667) );
  OAI21_X1 U5141 ( .B1(n7858), .B2(n7855), .A(n4476), .ZN(n4666) );
  NOR2_X1 U5142 ( .A1(n8232), .A2(n8227), .ZN(n5211) );
  AOI21_X1 U5143 ( .B1(n4811), .B2(n4809), .A(n4432), .ZN(n4807) );
  NAND2_X1 U5144 ( .A1(n7052), .A2(n7051), .ZN(n9721) );
  NAND2_X1 U5145 ( .A1(n6271), .A2(n6270), .ZN(n7739) );
  AND2_X1 U5146 ( .A1(n6267), .A2(n6266), .ZN(n6832) );
  OR2_X1 U5147 ( .A1(n4883), .A2(n4542), .ZN(n4543) );
  NOR2_X1 U5148 ( .A1(n4542), .A2(n4885), .ZN(n4547) );
  NAND2_X1 U5149 ( .A1(n4928), .A2(n8005), .ZN(n6049) );
  INV_X1 U5150 ( .A(n6048), .ZN(n4928) );
  INV_X1 U5151 ( .A(n6003), .ZN(n4578) );
  AND2_X1 U5152 ( .A1(n9372), .A2(n9206), .ZN(n8203) );
  NOR2_X1 U5153 ( .A1(n9383), .A2(n9388), .ZN(n4741) );
  INV_X1 U5154 ( .A(n6668), .ZN(n4524) );
  XNOR2_X1 U5155 ( .A(n7226), .B(n7225), .ZN(n7235) );
  NAND2_X1 U5156 ( .A1(n4844), .A2(n4843), .ZN(n7448) );
  AOI21_X1 U5157 ( .B1(n4846), .B2(n4848), .A(n4506), .ZN(n4843) );
  NAND2_X1 U5158 ( .A1(n5545), .A2(n5104), .ZN(n5549) );
  AND2_X1 U5159 ( .A1(n5096), .A2(n5095), .ZN(n5517) );
  INV_X1 U5160 ( .A(n5066), .ZN(n4858) );
  INV_X1 U5161 ( .A(n4863), .ZN(n4862) );
  OAI21_X1 U5162 ( .B1(n4866), .B2(n4440), .A(n5057), .ZN(n4863) );
  NAND2_X1 U5163 ( .A1(n5246), .A2(n5245), .ZN(n6441) );
  OAI21_X1 U5164 ( .B1(n8490), .B2(n7669), .A(n7850), .ZN(n7672) );
  INV_X1 U5165 ( .A(n8232), .ZN(n4780) );
  NAND2_X1 U5166 ( .A1(n4771), .A2(n4769), .ZN(n7208) );
  AOI21_X1 U5167 ( .B1(n4772), .B2(n4778), .A(n4770), .ZN(n4769) );
  AND2_X1 U5168 ( .A1(n4774), .A2(n8512), .ZN(n4772) );
  NAND2_X1 U5169 ( .A1(n4766), .A2(n4763), .ZN(n8567) );
  NOR2_X1 U5170 ( .A1(n8577), .A2(n7205), .ZN(n4763) );
  AND2_X1 U5171 ( .A1(n8818), .A2(n8604), .ZN(n7194) );
  INV_X1 U5172 ( .A(n7796), .ZN(n4750) );
  INV_X1 U5173 ( .A(n5314), .ZN(n7673) );
  NAND2_X1 U5175 ( .A1(n6513), .A2(n7229), .ZN(n5222) );
  INV_X1 U5176 ( .A(n9753), .ZN(n7869) );
  NAND2_X1 U5177 ( .A1(n4442), .A2(n4836), .ZN(n4674) );
  NAND2_X1 U5178 ( .A1(n5135), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5138) );
  OR2_X1 U5179 ( .A1(n9006), .A2(n9005), .ZN(n4541) );
  OAI21_X1 U5180 ( .B1(n8010), .B2(n4894), .A(n4892), .ZN(n4891) );
  OAI21_X1 U5181 ( .B1(n8010), .B2(n8003), .A(n4894), .ZN(n4892) );
  INV_X1 U5182 ( .A(n7969), .ZN(n4914) );
  INV_X1 U5183 ( .A(n7459), .ZN(n7434) );
  NAND2_X1 U5184 ( .A1(n8229), .A2(n9419), .ZN(n7314) );
  OAI21_X1 U5185 ( .B1(n9529), .B2(n5912), .A(n4568), .ZN(n9528) );
  NAND2_X1 U5186 ( .A1(n9529), .A2(n5912), .ZN(n4568) );
  NAND2_X1 U5187 ( .A1(n9564), .A2(n9563), .ZN(n4566) );
  AOI21_X1 U5188 ( .B1(n4939), .B2(n8187), .A(n4479), .ZN(n4937) );
  NAND2_X1 U5189 ( .A1(n9106), .A2(n4939), .ZN(n4936) );
  NAND2_X1 U5190 ( .A1(n9117), .A2(n9291), .ZN(n4802) );
  AOI21_X1 U5191 ( .B1(n4623), .B2(n4625), .A(n4957), .ZN(n4622) );
  INV_X1 U5192 ( .A(n4625), .ZN(n4624) );
  AND2_X1 U5193 ( .A1(n9362), .A2(n9177), .ZN(n4957) );
  AOI21_X1 U5194 ( .B1(n4590), .B2(n7469), .A(n4589), .ZN(n4588) );
  OAI22_X1 U5195 ( .A1(n7035), .A2(n7009), .B1(n7386), .B2(n9043), .ZN(n8173)
         );
  INV_X1 U5196 ( .A(n6644), .ZN(n7449) );
  INV_X1 U5197 ( .A(n9296), .ZN(n9459) );
  NAND2_X1 U5198 ( .A1(n8238), .A2(n5651), .ZN(n4967) );
  XNOR2_X1 U5199 ( .A(n9313), .B(n9311), .ZN(n9310) );
  NAND2_X1 U5200 ( .A1(n4702), .A2(n4706), .ZN(n4701) );
  NAND2_X1 U5201 ( .A1(n4698), .A2(n7627), .ZN(n4697) );
  NAND2_X1 U5202 ( .A1(n4703), .A2(n7537), .ZN(n4702) );
  OAI21_X1 U5203 ( .B1(n7819), .B2(n7818), .A(n4642), .ZN(n4641) );
  AND2_X1 U5204 ( .A1(n7817), .A2(n7816), .ZN(n4642) );
  NOR3_X1 U5205 ( .A1(n7573), .A2(n7572), .A3(n9269), .ZN(n7577) );
  AOI21_X1 U5206 ( .B1(n4711), .B2(n7569), .A(n4708), .ZN(n7573) );
  OAI21_X1 U5207 ( .B1(n7841), .B2(n7840), .A(n4473), .ZN(n4651) );
  INV_X1 U5208 ( .A(n7590), .ZN(n7593) );
  NAND2_X1 U5209 ( .A1(n4648), .A2(n4647), .ZN(n7853) );
  INV_X1 U5210 ( .A(n7848), .ZN(n4647) );
  INV_X1 U5211 ( .A(n6873), .ZN(n4817) );
  OAI21_X1 U5212 ( .B1(n7685), .B2(n4817), .A(n7690), .ZN(n4816) );
  NAND2_X1 U5213 ( .A1(n5054), .A2(n5053), .ZN(n5057) );
  INV_X1 U5214 ( .A(SI_12_), .ZN(n5053) );
  INV_X1 U5215 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5041) );
  INV_X1 U5216 ( .A(n5430), .ZN(n4971) );
  INV_X1 U5217 ( .A(n7174), .ZN(n5425) );
  NAND2_X1 U5218 ( .A1(n7175), .A2(n5430), .ZN(n4970) );
  NAND2_X1 U5219 ( .A1(n8556), .A2(n7198), .ZN(n4832) );
  AND2_X1 U5220 ( .A1(n8824), .A2(n8624), .ZN(n7818) );
  NAND2_X1 U5221 ( .A1(n8649), .A2(n8669), .ZN(n4812) );
  OR2_X1 U5222 ( .A1(n8828), .A2(n8669), .ZN(n7807) );
  OAI21_X1 U5223 ( .B1(n8711), .B2(n4825), .A(n8702), .ZN(n4824) );
  NAND2_X1 U5224 ( .A1(n4481), .A2(n4749), .ZN(n4744) );
  NAND2_X1 U5225 ( .A1(n4749), .A2(n7801), .ZN(n4748) );
  NAND2_X1 U5226 ( .A1(n4690), .A2(n9811), .ZN(n4689) );
  INV_X1 U5227 ( .A(n4691), .ZN(n4690) );
  OAI21_X1 U5228 ( .B1(n6881), .B2(n4835), .A(n4833), .ZN(n9719) );
  AOI21_X1 U5229 ( .B1(n4834), .B2(n8735), .A(n4470), .ZN(n4833) );
  NAND2_X1 U5230 ( .A1(n6424), .A2(n4411), .ZN(n7742) );
  NAND2_X1 U5231 ( .A1(n8391), .A2(n7885), .ZN(n7731) );
  INV_X1 U5232 ( .A(n6270), .ZN(n6282) );
  AND2_X1 U5233 ( .A1(n5140), .A2(n7728), .ZN(n6512) );
  AND2_X1 U5234 ( .A1(n4429), .A2(n4695), .ZN(n4694) );
  NOR2_X1 U5235 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5123) );
  NAND2_X1 U5236 ( .A1(n5676), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5699) );
  INV_X1 U5237 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n4838) );
  INV_X1 U5238 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5117) );
  INV_X1 U5239 ( .A(n6398), .ZN(n4548) );
  NOR2_X1 U5240 ( .A1(n7945), .A2(n4538), .ZN(n4537) );
  INV_X1 U5241 ( .A(n4540), .ZN(n4538) );
  NOR2_X1 U5242 ( .A1(n4721), .A2(n7622), .ZN(n4720) );
  AND2_X1 U5243 ( .A1(n7625), .A2(n4850), .ZN(n4849) );
  NAND2_X1 U5244 ( .A1(n7622), .A2(n4706), .ZN(n4850) );
  NAND2_X1 U5245 ( .A1(n7629), .A2(n7628), .ZN(n4852) );
  NAND2_X1 U5246 ( .A1(n7524), .A2(n7627), .ZN(n4851) );
  NOR2_X1 U5247 ( .A1(n8192), .A2(n9089), .ZN(n7622) );
  INV_X1 U5248 ( .A(n4874), .ZN(n7623) );
  NOR2_X1 U5249 ( .A1(n4795), .A2(n8213), .ZN(n4794) );
  INV_X1 U5250 ( .A(n4796), .ZN(n4795) );
  OR2_X1 U5251 ( .A1(n9337), .A2(n9141), .ZN(n9113) );
  NOR2_X1 U5252 ( .A1(n9354), .A2(n9362), .ZN(n4735) );
  AND2_X1 U5253 ( .A1(n9354), .A2(n9191), .ZN(n8209) );
  NOR2_X1 U5254 ( .A1(n4629), .A2(n8184), .ZN(n4628) );
  INV_X1 U5255 ( .A(n8182), .ZN(n4629) );
  INV_X1 U5256 ( .A(n9377), .ZN(n4740) );
  OR2_X1 U5257 ( .A1(n7002), .A2(n6816), .ZN(n7557) );
  NAND2_X1 U5258 ( .A1(n4610), .A2(n4609), .ZN(n9457) );
  OR2_X1 U5259 ( .A1(n9649), .A2(n9047), .ZN(n6683) );
  INV_X1 U5260 ( .A(n6665), .ZN(n4616) );
  INV_X1 U5261 ( .A(n7481), .ZN(n4617) );
  NAND2_X1 U5262 ( .A1(n9053), .A2(n6225), .ZN(n7408) );
  AND2_X1 U5263 ( .A1(n6846), .A2(n7661), .ZN(n7627) );
  AND2_X1 U5264 ( .A1(n5654), .A2(n5639), .ZN(n5652) );
  AND2_X1 U5265 ( .A1(n4929), .A2(n4490), .ZN(n4561) );
  NAND2_X1 U5266 ( .A1(n5549), .A2(n5105), .ZN(n5113) );
  NAND2_X1 U5267 ( .A1(n5753), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5757) );
  AOI21_X1 U5268 ( .B1(n4879), .B2(n4877), .A(n4876), .ZN(n4875) );
  INV_X1 U5269 ( .A(n4879), .ZN(n4878) );
  INV_X1 U5270 ( .A(n5096), .ZN(n4876) );
  INV_X1 U5271 ( .A(n5462), .ZN(n5084) );
  INV_X1 U5272 ( .A(n6200), .ZN(n4930) );
  AND2_X1 U5273 ( .A1(n5078), .A2(n5077), .ZN(n5431) );
  INV_X1 U5274 ( .A(n4857), .ZN(n4856) );
  OAI21_X1 U5275 ( .B1(n4860), .B2(n4437), .A(n5072), .ZN(n4857) );
  NAND2_X1 U5276 ( .A1(n5065), .A2(SI_14_), .ZN(n5066) );
  NOR2_X1 U5277 ( .A1(n5067), .A2(n4861), .ZN(n4860) );
  INV_X1 U5278 ( .A(n5062), .ZN(n4861) );
  INV_X1 U5279 ( .A(n5412), .ZN(n5067) );
  NAND2_X1 U5280 ( .A1(n5072), .A2(n5071), .ZN(n5447) );
  NOR2_X1 U5281 ( .A1(n5051), .A2(n4867), .ZN(n4866) );
  INV_X1 U5282 ( .A(n5046), .ZN(n4867) );
  INV_X1 U5283 ( .A(n5382), .ZN(n5051) );
  XNOR2_X1 U5284 ( .A(n5048), .B(SI_11_), .ZN(n5382) );
  INV_X1 U5285 ( .A(n4872), .ZN(n4871) );
  AOI21_X1 U5286 ( .B1(n4872), .B2(n4870), .A(n4869), .ZN(n4868) );
  AND2_X1 U5287 ( .A1(n4873), .A2(n4993), .ZN(n4872) );
  NAND2_X1 U5288 ( .A1(n5205), .A2(n5204), .ZN(n5010) );
  NAND2_X1 U5289 ( .A1(n6970), .A2(n6969), .ZN(n6968) );
  AND2_X1 U5290 ( .A1(n8313), .A2(n5516), .ZN(n4985) );
  NAND2_X1 U5291 ( .A1(n5513), .A2(n5512), .ZN(n8253) );
  NAND2_X1 U5292 ( .A1(n5406), .A2(n4461), .ZN(n5403) );
  INV_X1 U5293 ( .A(n6991), .ZN(n4979) );
  OR2_X1 U5294 ( .A1(n5392), .A2(n5359), .ZN(n5371) );
  NAND2_X1 U5295 ( .A1(n6441), .A2(n4460), .ZN(n4988) );
  OR2_X1 U5296 ( .A1(n5629), .A2(n8349), .ZN(n8351) );
  INV_X1 U5297 ( .A(n7861), .ZN(n7864) );
  OR2_X1 U5298 ( .A1(n5195), .A2(n6507), .ZN(n5177) );
  AOI21_X1 U5299 ( .B1(n8039), .B2(P2_REG1_REG_7__SCAN_IN), .A(n9870), .ZN(
        n8091) );
  NOR3_X1 U5300 ( .A1(n8522), .A2(n4678), .A3(n8481), .ZN(n8480) );
  NAND2_X1 U5301 ( .A1(n4680), .A2(n4679), .ZN(n4678) );
  INV_X1 U5302 ( .A(n4681), .ZN(n4680) );
  AND2_X1 U5303 ( .A1(n5665), .A2(n5664), .ZN(n8494) );
  OR2_X1 U5304 ( .A1(n7199), .A2(n5722), .ZN(n5665) );
  AND3_X1 U5305 ( .A1(n5647), .A2(n5646), .A3(n5645), .ZN(n8357) );
  NAND2_X1 U5306 ( .A1(n7847), .A2(n7846), .ZN(n8486) );
  INV_X1 U5307 ( .A(n7837), .ZN(n4775) );
  OR2_X1 U5308 ( .A1(n8555), .A2(n8556), .ZN(n8553) );
  NOR2_X1 U5309 ( .A1(n8622), .A2(n7204), .ZN(n8603) );
  AOI21_X1 U5310 ( .B1(n4807), .B2(n4808), .A(n4474), .ZN(n4805) );
  NAND2_X1 U5311 ( .A1(n4468), .A2(n4812), .ZN(n4809) );
  NAND2_X1 U5312 ( .A1(n8664), .A2(n7715), .ZN(n8651) );
  NOR2_X1 U5313 ( .A1(n8670), .A2(n8828), .ZN(n8646) );
  NAND2_X1 U5314 ( .A1(n4814), .A2(n8680), .ZN(n4813) );
  AOI21_X1 U5315 ( .B1(n8683), .B2(n8682), .A(n4826), .ZN(n8662) );
  AND2_X1 U5316 ( .A1(n8838), .A2(n8705), .ZN(n4826) );
  NAND2_X1 U5317 ( .A1(n8662), .A2(n8661), .ZN(n8660) );
  INV_X1 U5318 ( .A(n7202), .ZN(n4755) );
  NAND2_X1 U5319 ( .A1(n8712), .A2(n8711), .ZN(n8710) );
  NOR2_X1 U5320 ( .A1(n7118), .A2(n8855), .ZN(n8714) );
  AND2_X1 U5321 ( .A1(n4452), .A2(n7053), .ZN(n4841) );
  AND4_X1 U5322 ( .A1(n5376), .A2(n5375), .A3(n5374), .A4(n5373), .ZN(n7176)
         );
  AND2_X1 U5323 ( .A1(n7046), .A2(n7768), .ZN(n4767) );
  OR2_X1 U5324 ( .A1(n6274), .A2(n5721), .ZN(n9734) );
  NAND2_X1 U5325 ( .A1(n6489), .A2(n6488), .ZN(n6490) );
  AND2_X1 U5326 ( .A1(n7731), .A2(n7742), .ZN(n7687) );
  NAND2_X1 U5327 ( .A1(n6322), .A2(n7739), .ZN(n7733) );
  NAND2_X1 U5328 ( .A1(n6449), .A2(n6282), .ZN(n7730) );
  NAND4_X1 U5329 ( .A1(n7733), .A2(n7742), .A3(n7731), .A4(n7730), .ZN(n6428)
         );
  OR2_X1 U5330 ( .A1(n9787), .A2(n7728), .ZN(n6268) );
  NAND2_X1 U5331 ( .A1(n6881), .A2(n6880), .ZN(n9777) );
  NAND2_X1 U5332 ( .A1(n6509), .A2(n9760), .ZN(n9753) );
  AND2_X1 U5333 ( .A1(n5682), .A2(n4439), .ZN(n5696) );
  NAND2_X1 U5334 ( .A1(n5138), .A2(n5137), .ZN(n5143) );
  INV_X1 U5335 ( .A(n5236), .ZN(n4974) );
  AND2_X1 U5336 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n6357) );
  INV_X1 U5337 ( .A(n4884), .ZN(n4883) );
  OAI21_X1 U5338 ( .B1(n6397), .B2(n4885), .A(n6606), .ZN(n4884) );
  NAND2_X1 U5339 ( .A1(n4548), .A2(n6400), .ZN(n4549) );
  NAND2_X1 U5340 ( .A1(n4919), .A2(n4918), .ZN(n4917) );
  NAND2_X1 U5341 ( .A1(n4898), .A2(n4896), .ZN(n6936) );
  NOR2_X1 U5342 ( .A1(n6787), .A2(n4897), .ZN(n4896) );
  INV_X1 U5343 ( .A(n4900), .ZN(n4897) );
  AND2_X1 U5344 ( .A1(n4906), .A2(n7981), .ZN(n4903) );
  NAND2_X1 U5345 ( .A1(n4916), .A2(n4907), .ZN(n4906) );
  OAI21_X1 U5346 ( .B1(n6293), .B2(n6294), .A(n6295), .ZN(n6395) );
  OR2_X1 U5347 ( .A1(n9008), .A2(n4536), .ZN(n4533) );
  INV_X1 U5348 ( .A(n4537), .ZN(n4536) );
  NAND2_X1 U5349 ( .A1(n6942), .A2(n4920), .ZN(n7904) );
  NOR2_X1 U5350 ( .A1(n6953), .A2(n4921), .ZN(n4920) );
  INV_X1 U5351 ( .A(n6941), .ZN(n4921) );
  NAND2_X1 U5352 ( .A1(n4882), .A2(n6051), .ZN(n6075) );
  NAND2_X1 U5353 ( .A1(n9025), .A2(n9028), .ZN(n4550) );
  AND2_X1 U5354 ( .A1(n8971), .A2(n4925), .ZN(n4924) );
  OR2_X1 U5355 ( .A1(n8963), .A2(n4926), .ZN(n4925) );
  INV_X1 U5356 ( .A(n7929), .ZN(n4926) );
  AND2_X1 U5357 ( .A1(n4903), .A2(n4445), .ZN(n4560) );
  NAND2_X1 U5358 ( .A1(n4559), .A2(n4445), .ZN(n4558) );
  INV_X1 U5359 ( .A(n8954), .ZN(n4559) );
  AND2_X1 U5360 ( .A1(n4556), .A2(n9017), .ZN(n4555) );
  OR2_X1 U5361 ( .A1(n4560), .A2(n4557), .ZN(n4556) );
  INV_X1 U5362 ( .A(n4558), .ZN(n4557) );
  NOR2_X1 U5363 ( .A1(n8977), .A2(n4909), .ZN(n4908) );
  INV_X1 U5364 ( .A(n4911), .ZN(n4909) );
  NAND2_X1 U5365 ( .A1(n4551), .A2(n7921), .ZN(n9026) );
  NAND2_X1 U5366 ( .A1(n5935), .A2(n5934), .ZN(n4569) );
  AND2_X1 U5367 ( .A1(n9568), .A2(n9567), .ZN(n9570) );
  AND2_X1 U5368 ( .A1(n4566), .A2(n4492), .ZN(n9577) );
  NOR2_X1 U5369 ( .A1(n4577), .A2(n4494), .ZN(n4576) );
  NOR2_X1 U5370 ( .A1(n6001), .A2(n4578), .ZN(n4577) );
  OR2_X1 U5371 ( .A1(n6000), .A2(n4578), .ZN(n4575) );
  OR2_X1 U5372 ( .A1(n6023), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6137) );
  NOR2_X1 U5373 ( .A1(n6719), .A2(n4580), .ZN(n6720) );
  AND2_X1 U5374 ( .A1(n6930), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4580) );
  NAND2_X1 U5375 ( .A1(n6725), .A2(n4516), .ZN(n9620) );
  OR2_X1 U5376 ( .A1(n6930), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4516) );
  OR2_X1 U5377 ( .A1(n6908), .A2(n6907), .ZN(n4565) );
  AND2_X1 U5378 ( .A1(n9322), .A2(n9041), .ZN(n4941) );
  NOR2_X1 U5379 ( .A1(n7622), .A2(n7623), .ZN(n8218) );
  NAND2_X1 U5380 ( .A1(n9121), .A2(n8186), .ZN(n9106) );
  NAND2_X1 U5381 ( .A1(n4797), .A2(n4799), .ZN(n4796) );
  NAND2_X1 U5382 ( .A1(n8211), .A2(n4798), .ZN(n4797) );
  NAND2_X1 U5383 ( .A1(n9155), .A2(n8209), .ZN(n4798) );
  NAND2_X1 U5384 ( .A1(n9160), .A2(n4448), .ZN(n4789) );
  NAND2_X1 U5385 ( .A1(n9122), .A2(n9129), .ZN(n9121) );
  AOI21_X1 U5386 ( .B1(n4956), .B2(n4955), .A(n4466), .ZN(n9150) );
  NAND2_X1 U5387 ( .A1(n9173), .A2(n9191), .ZN(n4955) );
  OR2_X1 U5388 ( .A1(n9368), .A2(n9228), .ZN(n4630) );
  AND2_X1 U5389 ( .A1(n4482), .A2(n8178), .ZN(n4944) );
  AOI21_X1 U5390 ( .B1(n4588), .B2(n4591), .A(n4587), .ZN(n4586) );
  INV_X1 U5391 ( .A(n9226), .ZN(n4587) );
  NAND2_X1 U5392 ( .A1(n9250), .A2(n8201), .ZN(n4593) );
  AND2_X1 U5393 ( .A1(n7582), .A2(n8202), .ZN(n9238) );
  OR2_X1 U5394 ( .A1(n7469), .A2(n8200), .ZN(n9251) );
  NAND2_X1 U5395 ( .A1(n9265), .A2(n9269), .ZN(n4621) );
  NAND2_X1 U5396 ( .A1(n7036), .A2(n7392), .ZN(n7016) );
  AOI21_X1 U5397 ( .B1(n9452), .B2(n7004), .A(n4469), .ZN(n7035) );
  NOR2_X1 U5398 ( .A1(n4451), .A2(n4608), .ZN(n4607) );
  INV_X1 U5399 ( .A(n4609), .ZN(n4608) );
  AOI21_X1 U5400 ( .B1(n4787), .B2(n4786), .A(n4785), .ZN(n4784) );
  INV_X1 U5401 ( .A(n7389), .ZN(n4785) );
  INV_X1 U5402 ( .A(n7013), .ZN(n4787) );
  NOR2_X1 U5403 ( .A1(n7547), .A2(n4788), .ZN(n4786) );
  OR2_X1 U5404 ( .A1(n6695), .A2(n6694), .ZN(n6704) );
  OR2_X1 U5405 ( .A1(n6564), .A2(n6563), .ZN(n6654) );
  NAND2_X1 U5406 ( .A1(n9457), .A2(n7547), .ZN(n9453) );
  NAND2_X1 U5407 ( .A1(n4618), .A2(n4617), .ZN(n6666) );
  INV_X1 U5408 ( .A(n6560), .ZN(n4618) );
  NAND2_X1 U5409 ( .A1(n6406), .A2(n4946), .ZN(n6584) );
  AND2_X1 U5410 ( .A1(n7535), .A2(n6346), .ZN(n4946) );
  NAND2_X1 U5411 ( .A1(n6225), .A2(n4508), .ZN(n6238) );
  NAND2_X1 U5412 ( .A1(n4948), .A2(n4636), .ZN(n4635) );
  NAND2_X1 U5413 ( .A1(n4952), .A2(n4951), .ZN(n4948) );
  OR2_X1 U5414 ( .A1(n7631), .A2(n7643), .ZN(n9462) );
  NAND2_X1 U5415 ( .A1(n5802), .A2(n5801), .ZN(n9296) );
  INV_X1 U5416 ( .A(n9462), .ZN(n9293) );
  INV_X1 U5417 ( .A(n8192), .ZN(n9317) );
  OR3_X1 U5418 ( .A1(n7187), .A2(n7071), .A3(n7169), .ZN(n6123) );
  XNOR2_X1 U5419 ( .A(n7448), .B(n7447), .ZN(n8225) );
  XNOR2_X1 U5420 ( .A(n5608), .B(n5607), .ZN(n7266) );
  OAI21_X1 U5421 ( .B1(n5502), .B2(n5501), .A(n5092), .ZN(n5518) );
  INV_X1 U5422 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5728) );
  NOR2_X2 U5423 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5775) );
  XNOR2_X1 U5424 ( .A(n5003), .B(SI_1_), .ZN(n5176) );
  NAND3_X1 U5425 ( .A1(n4842), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4653) );
  INV_X1 U5426 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4842) );
  NAND2_X1 U5427 ( .A1(n4967), .A2(n5712), .ZN(n4966) );
  INV_X1 U5428 ( .A(n8600), .ZN(n8813) );
  AND4_X1 U5429 ( .A1(n5423), .A2(n5422), .A3(n5421), .A4(n5420), .ZN(n8371)
         );
  NAND2_X1 U5430 ( .A1(n5551), .A2(n5550), .ZN(n8808) );
  INV_X1 U5431 ( .A(n8374), .ZN(n8348) );
  NAND2_X1 U5432 ( .A1(n6448), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8368) );
  INV_X1 U5433 ( .A(n4998), .ZN(n4761) );
  AND3_X1 U5434 ( .A1(n5725), .A2(n5724), .A3(n5723), .ZN(n7668) );
  AND4_X1 U5435 ( .A1(n5578), .A2(n5577), .A3(n5576), .A4(n5575), .ZN(n8591)
         );
  NAND2_X1 U5436 ( .A1(n4522), .A2(n8478), .ZN(n4521) );
  OR2_X1 U5437 ( .A1(n8479), .A2(n4656), .ZN(n4522) );
  INV_X1 U5438 ( .A(n6838), .ZN(n6833) );
  NAND2_X1 U5439 ( .A1(n9008), .A2(n4541), .ZN(n4539) );
  NOR2_X1 U5440 ( .A1(n4431), .A2(n9038), .ZN(n4887) );
  INV_X1 U5441 ( .A(n8010), .ZN(n4890) );
  NAND2_X1 U5442 ( .A1(n4891), .A2(n4893), .ZN(n4889) );
  NAND2_X1 U5443 ( .A1(n8010), .A2(n8003), .ZN(n4893) );
  NAND2_X1 U5444 ( .A1(n7312), .A2(n7311), .ZN(n9383) );
  INV_X1 U5445 ( .A(n9332), .ZN(n9112) );
  INV_X1 U5446 ( .A(n6846), .ZN(n7646) );
  NAND2_X1 U5447 ( .A1(n7255), .A2(n7254), .ZN(n9117) );
  NAND2_X1 U5448 ( .A1(n7265), .A2(n7264), .ZN(n9130) );
  OR2_X1 U5449 ( .A1(n9019), .A2(n7434), .ZN(n7265) );
  NAND2_X1 U5450 ( .A1(n9526), .A2(n5919), .ZN(n5917) );
  NOR2_X1 U5451 ( .A1(n6727), .A2(n6726), .ZN(n6910) );
  OAI21_X1 U5452 ( .B1(n9311), .B2(n9691), .A(n9314), .ZN(n4725) );
  NAND2_X1 U5453 ( .A1(n4704), .A2(n4450), .ZN(n4703) );
  NAND2_X1 U5454 ( .A1(n4699), .A2(n7538), .ZN(n4698) );
  NAND2_X1 U5455 ( .A1(n4704), .A2(n4700), .ZN(n4699) );
  INV_X1 U5456 ( .A(n7539), .ZN(n4700) );
  NAND2_X1 U5457 ( .A1(n7806), .A2(n7805), .ZN(n4646) );
  NOR2_X1 U5458 ( .A1(n4661), .A2(n8577), .ZN(n4660) );
  NAND2_X1 U5459 ( .A1(n4641), .A2(n4453), .ZN(n7823) );
  INV_X1 U5460 ( .A(n8528), .ZN(n4665) );
  NAND2_X1 U5461 ( .A1(n4770), .A2(n7859), .ZN(n4652) );
  NAND2_X1 U5462 ( .A1(n4650), .A2(n4649), .ZN(n4648) );
  INV_X1 U5463 ( .A(n7845), .ZN(n4649) );
  NAND2_X1 U5464 ( .A1(n4651), .A2(n7846), .ZN(n4650) );
  NAND2_X1 U5465 ( .A1(n8728), .A2(n8735), .ZN(n6893) );
  NOR2_X1 U5466 ( .A1(n8217), .A2(n4706), .ZN(n4721) );
  OR2_X1 U5467 ( .A1(n9328), .A2(n7427), .ZN(n7615) );
  INV_X1 U5468 ( .A(n5654), .ZN(n4848) );
  INV_X1 U5469 ( .A(n4847), .ZN(n4846) );
  OAI21_X1 U5470 ( .B1(n5652), .B2(n4848), .A(n7216), .ZN(n4847) );
  AND2_X1 U5471 ( .A1(n4880), .A2(n5517), .ZN(n4879) );
  NAND2_X1 U5472 ( .A1(n5501), .A2(n5092), .ZN(n4880) );
  INV_X1 U5473 ( .A(n5092), .ZN(n4877) );
  INV_X1 U5474 ( .A(n5431), .ZN(n4855) );
  INV_X1 U5475 ( .A(n5050), .ZN(n4864) );
  NAND2_X1 U5476 ( .A1(n5311), .A2(n5035), .ZN(n4873) );
  INV_X1 U5477 ( .A(n5035), .ZN(n4870) );
  NAND2_X1 U5478 ( .A1(n5037), .A2(n5036), .ZN(n5040) );
  NAND2_X1 U5479 ( .A1(n8485), .A2(n8770), .ZN(n4681) );
  INV_X1 U5480 ( .A(n4809), .ZN(n4808) );
  OR2_X1 U5481 ( .A1(n8835), .A2(n8680), .ZN(n7715) );
  NOR2_X1 U5482 ( .A1(n8843), .A2(n8848), .ZN(n4685) );
  NAND2_X1 U5483 ( .A1(n9802), .A2(n9795), .ZN(n4691) );
  NAND2_X1 U5484 ( .A1(n7074), .A2(n7692), .ZN(n4768) );
  INV_X1 U5485 ( .A(n7685), .ZN(n6495) );
  OAI21_X1 U5486 ( .B1(n6490), .B2(n4817), .A(n4815), .ZN(n6877) );
  INV_X1 U5487 ( .A(n4816), .ZN(n4815) );
  INV_X1 U5488 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4980) );
  INV_X1 U5489 ( .A(n5355), .ZN(n5120) );
  AND2_X1 U5490 ( .A1(n4820), .A2(n4821), .ZN(n5325) );
  NOR2_X1 U5491 ( .A1(n5236), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5256) );
  INV_X1 U5492 ( .A(n4912), .ZN(n4907) );
  NAND2_X1 U5493 ( .A1(n8944), .A2(n7964), .ZN(n7970) );
  NAND2_X1 U5494 ( .A1(n4874), .A2(n7467), .ZN(n7619) );
  NOR2_X1 U5495 ( .A1(n5932), .A2(n4572), .ZN(n4571) );
  INV_X1 U5496 ( .A(n5929), .ZN(n4572) );
  AND2_X1 U5497 ( .A1(n7615), .A2(n7616), .ZN(n8188) );
  AND2_X1 U5498 ( .A1(n7423), .A2(n9138), .ZN(n8211) );
  OR2_X1 U5499 ( .A1(n7360), .A2(n8955), .ZN(n7270) );
  AND2_X1 U5500 ( .A1(n9345), .A2(n8956), .ZN(n7605) );
  AND2_X1 U5501 ( .A1(n4735), .A2(n4734), .ZN(n4733) );
  INV_X1 U5502 ( .A(n4628), .ZN(n4623) );
  OR2_X1 U5503 ( .A1(n9362), .A2(n9207), .ZN(n7596) );
  NOR2_X1 U5504 ( .A1(n4472), .A2(n4620), .ZN(n4619) );
  INV_X1 U5505 ( .A(n8177), .ZN(n4620) );
  OR2_X1 U5506 ( .A1(n6957), .A2(n8910), .ZN(n7020) );
  OR2_X1 U5507 ( .A1(n6800), .A2(n6799), .ZN(n6957) );
  NAND2_X1 U5508 ( .A1(n6702), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6800) );
  INV_X1 U5509 ( .A(n6704), .ZN(n6702) );
  AND2_X1 U5510 ( .A1(n6711), .A2(n7388), .ZN(n4609) );
  AND2_X1 U5511 ( .A1(n9473), .A2(n9479), .ZN(n6714) );
  NAND2_X1 U5512 ( .A1(n7411), .A2(n4583), .ZN(n4582) );
  NOR2_X1 U5513 ( .A1(n9194), .A2(n4626), .ZN(n4625) );
  INV_X1 U5514 ( .A(n4630), .ZN(n4626) );
  INV_X1 U5515 ( .A(n9184), .ZN(n9208) );
  NAND2_X1 U5516 ( .A1(n4730), .A2(n4729), .ZN(n6670) );
  NAND2_X1 U5517 ( .A1(n5766), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U5518 ( .A1(n9415), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4595) );
  NAND2_X1 U5519 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5763), .ZN(n4596) );
  AND2_X1 U5520 ( .A1(n5633), .A2(n5612), .ZN(n5613) );
  INV_X1 U5521 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5739) );
  AND2_X1 U5522 ( .A1(n5736), .A2(n5734), .ZN(n4929) );
  INV_X1 U5523 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U5524 ( .A1(n5032), .A2(n9949), .ZN(n5035) );
  INV_X1 U5525 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U5526 ( .A1(n4420), .A2(n5001), .ZN(n5002) );
  NAND2_X1 U5527 ( .A1(n5425), .A2(n5424), .ZN(n7172) );
  OR2_X1 U5528 ( .A1(n5553), .A2(n5163), .ZN(n5572) );
  AOI21_X1 U5529 ( .B1(n4985), .B2(n8256), .A(n4983), .ZN(n4982) );
  INV_X1 U5530 ( .A(n4985), .ZN(n4984) );
  INV_X1 U5531 ( .A(n5532), .ZN(n4983) );
  INV_X1 U5532 ( .A(n5580), .ZN(n5570) );
  OR2_X1 U5533 ( .A1(n5582), .A2(n8570), .ZN(n5579) );
  NAND2_X1 U5534 ( .A1(n4969), .A2(n4458), .ZN(n8294) );
  NAND2_X1 U5535 ( .A1(n4447), .A2(n4971), .ZN(n4968) );
  OR2_X1 U5536 ( .A1(n5441), .A2(n8366), .ZN(n5469) );
  NOR2_X1 U5537 ( .A1(n4464), .A2(n4425), .ZN(n4975) );
  INV_X1 U5538 ( .A(n6969), .ZN(n4976) );
  NAND2_X1 U5539 ( .A1(n6968), .A2(n4977), .ZN(n7147) );
  OR2_X1 U5540 ( .A1(n5489), .A2(n8343), .ZN(n5506) );
  NAND2_X1 U5541 ( .A1(n7172), .A2(n5430), .ZN(n8282) );
  NOR2_X1 U5542 ( .A1(n5713), .A2(n9753), .ZN(n5720) );
  OR2_X2 U5543 ( .A1(n9763), .A2(n5714), .ZN(n7683) );
  AND3_X1 U5544 ( .A1(n5624), .A2(n5623), .A3(n5622), .ZN(n8275) );
  INV_X1 U5545 ( .A(n5644), .ZN(n5722) );
  AND4_X1 U5546 ( .A1(n5526), .A2(n5525), .A3(n5524), .A4(n5523), .ZN(n8257)
         );
  AND4_X1 U5547 ( .A1(n5269), .A2(n5268), .A3(n5267), .A4(n5266), .ZN(n6878)
         );
  OR2_X1 U5548 ( .A1(n5195), .A2(n5194), .ZN(n5197) );
  INV_X1 U5549 ( .A(n8227), .ZN(n5168) );
  AND2_X1 U5550 ( .A1(n6543), .A2(n6544), .ZN(n8017) );
  AOI21_X1 U5551 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n8044), .A(n8017), .ZN(
        n8103) );
  AOI21_X1 U5552 ( .B1(n8036), .B2(P2_REG1_REG_9__SCAN_IN), .A(n8077), .ZN(
        n8067) );
  AOI21_X1 U5553 ( .B1(n8167), .B2(P2_REG1_REG_11__SCAN_IN), .A(n8163), .ZN(
        n8027) );
  NOR2_X1 U5554 ( .A1(n8415), .A2(n8414), .ZN(n8417) );
  AOI21_X1 U5555 ( .B1(n8455), .B2(P2_REG1_REG_17__SCAN_IN), .A(n8454), .ZN(
        n8456) );
  NAND2_X1 U5556 ( .A1(n7671), .A2(n7670), .ZN(n8481) );
  NAND2_X1 U5557 ( .A1(n7667), .A2(n7666), .ZN(n7873) );
  NOR2_X1 U5558 ( .A1(n4682), .A2(n8776), .ZN(n8498) );
  INV_X1 U5559 ( .A(n8486), .ZN(n7207) );
  NAND2_X1 U5560 ( .A1(n8538), .A2(n8537), .ZN(n4779) );
  NOR2_X1 U5561 ( .A1(n8792), .A2(n4693), .ZN(n4692) );
  INV_X1 U5562 ( .A(n4694), .ZN(n4693) );
  OR2_X1 U5563 ( .A1(n8543), .A2(n8787), .ZN(n8522) );
  INV_X1 U5564 ( .A(n8529), .ZN(n8520) );
  AOI21_X1 U5565 ( .B1(n4830), .B2(n4829), .A(n4475), .ZN(n4828) );
  INV_X1 U5566 ( .A(n7198), .ZN(n4829) );
  OR2_X1 U5567 ( .A1(n8559), .A2(n8537), .ZN(n4776) );
  NAND2_X1 U5568 ( .A1(n8612), .A2(n4429), .ZN(n8572) );
  NAND2_X1 U5569 ( .A1(n8612), .A2(n4426), .ZN(n8582) );
  INV_X1 U5570 ( .A(n7818), .ZN(n8619) );
  AND2_X1 U5571 ( .A1(n8631), .A2(n8616), .ZN(n8612) );
  AND2_X1 U5572 ( .A1(n8646), .A2(n8635), .ZN(n8631) );
  NAND2_X1 U5573 ( .A1(n8651), .A2(n4468), .ZN(n8650) );
  NAND2_X1 U5574 ( .A1(n8714), .A2(n4683), .ZN(n8670) );
  AND2_X1 U5575 ( .A1(n4428), .A2(n4814), .ZN(n4683) );
  NAND2_X1 U5576 ( .A1(n4756), .A2(n7804), .ZN(n8665) );
  NOR2_X1 U5577 ( .A1(n4747), .A2(n7203), .ZN(n4743) );
  NAND2_X1 U5578 ( .A1(n7192), .A2(n4827), .ZN(n4822) );
  INV_X1 U5579 ( .A(n4824), .ZN(n4823) );
  NAND2_X1 U5580 ( .A1(n8714), .A2(n4428), .ZN(n8687) );
  NAND2_X1 U5581 ( .A1(n4745), .A2(n4434), .ZN(n8679) );
  AND4_X1 U5582 ( .A1(n5446), .A2(n5445), .A3(n5444), .A4(n5443), .ZN(n8681)
         );
  NAND2_X1 U5583 ( .A1(n8714), .A2(n4685), .ZN(n8696) );
  AND2_X1 U5584 ( .A1(n8714), .A2(n8719), .ZN(n8715) );
  NOR2_X1 U5585 ( .A1(n4689), .A2(n9816), .ZN(n4687) );
  NAND2_X1 U5586 ( .A1(n7129), .A2(n7774), .ZN(n7089) );
  NOR2_X1 U5587 ( .A1(n9724), .A2(n4691), .ZN(n7134) );
  AND4_X1 U5588 ( .A1(n5397), .A2(n5396), .A3(n5395), .A4(n5394), .ZN(n7130)
         );
  NAND2_X1 U5589 ( .A1(n9721), .A2(n7053), .ZN(n7113) );
  NOR2_X1 U5590 ( .A1(n9724), .A2(n7080), .ZN(n7136) );
  NAND2_X1 U5591 ( .A1(n9729), .A2(n7765), .ZN(n7074) );
  NAND2_X1 U5592 ( .A1(n8737), .A2(n9783), .ZN(n9723) );
  AND4_X1 U5593 ( .A1(n5290), .A2(n5289), .A3(n5288), .A4(n5287), .ZN(n9735)
         );
  AND4_X1 U5594 ( .A1(n5324), .A2(n5323), .A3(n5322), .A4(n5321), .ZN(n9733)
         );
  NAND2_X1 U5595 ( .A1(n4676), .A2(n9770), .ZN(n8738) );
  NOR2_X1 U5596 ( .A1(n8738), .A2(n9773), .ZN(n8737) );
  NAND2_X1 U5597 ( .A1(n8389), .A2(n4677), .ZN(n6977) );
  NAND2_X1 U5598 ( .A1(n6318), .A2(n6317), .ZN(n6321) );
  AND3_X1 U5599 ( .A1(n6832), .A2(n6831), .A3(n6830), .ZN(n6838) );
  NOR2_X1 U5600 ( .A1(n6325), .A2(n4411), .ZN(n6431) );
  NAND2_X1 U5601 ( .A1(n7688), .A2(n6272), .ZN(n6318) );
  NAND2_X1 U5602 ( .A1(n7730), .A2(n7739), .ZN(n7688) );
  NAND2_X1 U5603 ( .A1(n5488), .A2(n5487), .ZN(n8828) );
  INV_X1 U5604 ( .A(n9820), .ZN(n9774) );
  AND3_X1 U5605 ( .A1(n6269), .A2(n6832), .A3(n6268), .ZN(n6290) );
  OR2_X1 U5606 ( .A1(n7144), .A2(n5679), .ZN(n5683) );
  INV_X1 U5607 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5147) );
  INV_X1 U5608 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5125) );
  OR2_X1 U5609 ( .A1(n5699), .A2(n5698), .ZN(n5700) );
  AND2_X1 U5610 ( .A1(n5116), .A2(n5237), .ZN(n4973) );
  NAND2_X1 U5611 ( .A1(n6115), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6361) );
  NAND2_X1 U5612 ( .A1(n9006), .A2(n9005), .ZN(n4540) );
  AND2_X1 U5613 ( .A1(n4487), .A2(n4895), .ZN(n4894) );
  NAND2_X1 U5614 ( .A1(n8003), .A2(n4493), .ZN(n4895) );
  NAND2_X1 U5615 ( .A1(n4491), .A2(n8963), .ZN(n8962) );
  INV_X1 U5616 ( .A(n7343), .ZN(n7249) );
  OR2_X1 U5617 ( .A1(n7358), .A2(n7357), .ZN(n7360) );
  OR2_X1 U5618 ( .A1(n7974), .A2(n4913), .ZN(n4912) );
  NAND2_X1 U5619 ( .A1(n7974), .A2(n4913), .ZN(n4911) );
  NAND2_X1 U5620 ( .A1(n6641), .A2(n4902), .ZN(n4900) );
  NOR2_X1 U5621 ( .A1(n4901), .A2(n4545), .ZN(n4544) );
  INV_X1 U5622 ( .A(n6615), .ZN(n4545) );
  NOR2_X1 U5623 ( .A1(n6641), .A2(n4902), .ZN(n4901) );
  NAND2_X1 U5624 ( .A1(n5964), .A2(n6048), .ZN(n6050) );
  INV_X1 U5625 ( .A(n7333), .ZN(n7247) );
  AOI21_X1 U5626 ( .B1(n4537), .B2(n4535), .A(n4480), .ZN(n4534) );
  INV_X1 U5627 ( .A(n4541), .ZN(n4535) );
  NAND2_X1 U5628 ( .A1(n4533), .A2(n4532), .ZN(n8984) );
  AND2_X1 U5629 ( .A1(n4534), .A2(n4496), .ZN(n4532) );
  OR2_X1 U5630 ( .A1(n7292), .A2(n7280), .ZN(n7301) );
  NAND2_X1 U5631 ( .A1(n7248), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n7343) );
  INV_X1 U5632 ( .A(n7301), .ZN(n7248) );
  OR2_X1 U5633 ( .A1(n6395), .A2(n4531), .ZN(n6397) );
  INV_X1 U5634 ( .A(n6396), .ZN(n4531) );
  NAND2_X1 U5635 ( .A1(n4851), .A2(n4852), .ZN(n4717) );
  NAND2_X1 U5636 ( .A1(n4719), .A2(n4849), .ZN(n4718) );
  NAND2_X1 U5637 ( .A1(n4417), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4954) );
  NAND2_X1 U5638 ( .A1(n7459), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4953) );
  NAND2_X1 U5639 ( .A1(n4413), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4949) );
  NAND2_X1 U5640 ( .A1(n9527), .A2(n9528), .ZN(n9526) );
  AOI21_X1 U5641 ( .B1(n9540), .B2(n5908), .A(n5907), .ZN(n5924) );
  NAND2_X1 U5642 ( .A1(n5930), .A2(n4571), .ZN(n9546) );
  NOR2_X1 U5643 ( .A1(n5926), .A2(n5925), .ZN(n5988) );
  NOR2_X1 U5644 ( .A1(n6015), .A2(n4567), .ZN(n9564) );
  AND2_X1 U5645 ( .A1(n6349), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4567) );
  NOR2_X1 U5646 ( .A1(n5989), .A2(n9570), .ZN(n9584) );
  NAND2_X1 U5647 ( .A1(n9604), .A2(n4512), .ZN(n6164) );
  OR2_X1 U5648 ( .A1(n9603), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4512) );
  NAND2_X1 U5649 ( .A1(n6164), .A2(n6165), .ZN(n6258) );
  NOR2_X1 U5650 ( .A1(n4574), .A2(n4579), .ZN(n4573) );
  INV_X1 U5651 ( .A(n9608), .ZN(n4579) );
  INV_X1 U5652 ( .A(n4576), .ZN(n4574) );
  NAND2_X1 U5653 ( .A1(n6259), .A2(n6260), .ZN(n6725) );
  NOR2_X1 U5654 ( .A1(n6252), .A2(n4581), .ZN(n6255) );
  AND2_X1 U5655 ( .A1(n6779), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4581) );
  NOR2_X1 U5656 ( .A1(n6255), .A2(n6254), .ZN(n6719) );
  XNOR2_X1 U5657 ( .A(n4514), .B(n4513), .ZN(n7657) );
  INV_X1 U5658 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n4513) );
  NAND2_X1 U5659 ( .A1(n9637), .A2(n4515), .ZN(n4514) );
  OR2_X1 U5660 ( .A1(n9636), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n4515) );
  NAND2_X1 U5661 ( .A1(n7237), .A2(n7236), .ZN(n9075) );
  NOR2_X1 U5662 ( .A1(n9080), .A2(n9317), .ZN(n9073) );
  NOR2_X1 U5663 ( .A1(n9107), .A2(n9328), .ZN(n9100) );
  OAI21_X1 U5664 ( .B1(n4789), .B2(n8215), .A(n4790), .ZN(n9094) );
  AOI21_X1 U5665 ( .B1(n4792), .B2(n4793), .A(n4791), .ZN(n4790) );
  INV_X1 U5666 ( .A(n4794), .ZN(n4792) );
  INV_X1 U5667 ( .A(n8188), .ZN(n9095) );
  NOR2_X1 U5668 ( .A1(n9348), .A2(n4634), .ZN(n9122) );
  AND2_X1 U5669 ( .A1(n9345), .A2(n9161), .ZN(n4634) );
  NAND2_X1 U5670 ( .A1(n9208), .A2(n4731), .ZN(n9135) );
  NOR2_X1 U5671 ( .A1(n9345), .A2(n4732), .ZN(n4731) );
  INV_X1 U5672 ( .A(n4733), .ZN(n4732) );
  NOR2_X1 U5673 ( .A1(n8210), .A2(n7605), .ZN(n9144) );
  OAI21_X1 U5674 ( .B1(n9160), .B2(n8209), .A(n9155), .ZN(n9158) );
  NAND2_X1 U5675 ( .A1(n9208), .A2(n4735), .ZN(n9168) );
  NAND2_X1 U5676 ( .A1(n9208), .A2(n8949), .ZN(n9182) );
  AND2_X1 U5677 ( .A1(n7596), .A2(n8206), .ZN(n9194) );
  NAND2_X1 U5678 ( .A1(n8183), .A2(n4628), .ZN(n4627) );
  NOR2_X1 U5679 ( .A1(n9372), .A2(n4739), .ZN(n4737) );
  NAND2_X1 U5680 ( .A1(n4945), .A2(n8178), .ZN(n9233) );
  OR2_X1 U5681 ( .A1(n9233), .A2(n9238), .ZN(n9234) );
  OR2_X1 U5682 ( .A1(n7374), .A2(n8972), .ZN(n7322) );
  NAND2_X1 U5683 ( .A1(n9284), .A2(n9279), .ZN(n9273) );
  NAND2_X1 U5684 ( .A1(n9284), .A2(n4741), .ZN(n9255) );
  NAND2_X1 U5685 ( .A1(n7018), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7372) );
  INV_X1 U5686 ( .A(n7020), .ZN(n7018) );
  NAND2_X1 U5687 ( .A1(n7245), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7374) );
  INV_X1 U5688 ( .A(n7372), .ZN(n7245) );
  AND2_X1 U5689 ( .A1(n7896), .A2(n9288), .ZN(n9284) );
  NAND2_X1 U5690 ( .A1(n4526), .A2(n4525), .ZN(n8196) );
  AND2_X1 U5691 ( .A1(n6714), .A2(n6761), .ZN(n6822) );
  INV_X1 U5692 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6694) );
  INV_X1 U5693 ( .A(n6654), .ZN(n6652) );
  NOR2_X1 U5694 ( .A1(n6670), .A2(n9649), .ZN(n9473) );
  INV_X1 U5695 ( .A(n4613), .ZN(n4612) );
  NAND2_X1 U5696 ( .A1(n6560), .A2(n4615), .ZN(n4611) );
  OAI21_X1 U5697 ( .B1(n4617), .B2(n4614), .A(n6683), .ZN(n4613) );
  NAND2_X1 U5698 ( .A1(n6562), .A2(n7538), .ZN(n6668) );
  NAND2_X1 U5699 ( .A1(n7646), .A2(n9243), .ZN(n4563) );
  NOR2_X1 U5700 ( .A1(n6238), .A2(n6239), .ZN(n6410) );
  NAND2_X1 U5701 ( .A1(n6209), .A2(n6208), .ZN(n6210) );
  NOR2_X1 U5702 ( .A1(n7400), .A2(n6179), .ZN(n6192) );
  AND2_X1 U5703 ( .A1(n4627), .A2(n4625), .ZN(n9365) );
  INV_X1 U5704 ( .A(n9692), .ZN(n9471) );
  NAND2_X1 U5705 ( .A1(n4610), .A2(n7388), .ZN(n6710) );
  NAND2_X1 U5706 ( .A1(n6666), .A2(n6665), .ZN(n6685) );
  INV_X1 U5707 ( .A(n9691), .ZN(n9392) );
  NAND2_X1 U5708 ( .A1(n7450), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4604) );
  INV_X1 U5709 ( .A(n4606), .ZN(n4605) );
  OAI21_X1 U5710 ( .B1(n6644), .B2(n6089), .A(n6088), .ZN(n4606) );
  NAND2_X1 U5711 ( .A1(n6183), .A2(n5803), .ZN(n5805) );
  AND2_X1 U5712 ( .A1(n7627), .A2(n6678), .ZN(n9697) );
  XNOR2_X1 U5713 ( .A(n7235), .B(SI_30_), .ZN(n8228) );
  NOR2_X1 U5714 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n4716) );
  NAND2_X1 U5715 ( .A1(n5653), .A2(n5652), .ZN(n4845) );
  INV_X1 U5716 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5748) );
  INV_X1 U5717 ( .A(n5113), .ZN(n5564) );
  NAND2_X1 U5718 ( .A1(n4930), .A2(n5734), .ZN(n6205) );
  OAI21_X1 U5719 ( .B1(n5063), .B2(n4437), .A(n4856), .ZN(n5432) );
  NAND2_X1 U5720 ( .A1(n4859), .A2(n5066), .ZN(n5448) );
  NAND2_X1 U5721 ( .A1(n5063), .A2(n4860), .ZN(n4859) );
  NAND2_X1 U5722 ( .A1(n4865), .A2(n5050), .ZN(n5354) );
  NAND2_X1 U5723 ( .A1(n5047), .A2(n4866), .ZN(n4865) );
  NAND2_X1 U5724 ( .A1(n5047), .A2(n5046), .ZN(n5383) );
  OR2_X1 U5725 ( .A1(n5872), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5873) );
  XNOR2_X1 U5726 ( .A(n5028), .B(SI_7_), .ZN(n5293) );
  NAND2_X1 U5727 ( .A1(n5022), .A2(n5021), .ZN(n5275) );
  XNOR2_X1 U5728 ( .A(n5023), .B(SI_6_), .ZN(n5274) );
  AND2_X1 U5729 ( .A1(n5793), .A2(n5729), .ZN(n5849) );
  INV_X1 U5730 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5850) );
  OR2_X1 U5731 ( .A1(n5697), .A2(n7069), .ZN(n6509) );
  AND2_X1 U5732 ( .A1(n8351), .A2(n5631), .ZN(n5632) );
  NAND2_X1 U5733 ( .A1(n6968), .A2(n5334), .ZN(n6992) );
  NAND2_X1 U5734 ( .A1(n5504), .A2(n5503), .ZN(n8824) );
  NAND2_X1 U5735 ( .A1(n4963), .A2(n5193), .ZN(n7888) );
  INV_X1 U5736 ( .A(n4964), .ZN(n4963) );
  AND2_X1 U5737 ( .A1(n5193), .A2(n5185), .ZN(n7890) );
  NAND2_X1 U5738 ( .A1(n6441), .A2(n5247), .ZN(n6467) );
  AND4_X1 U5739 ( .A1(n5348), .A2(n5347), .A3(n5346), .A4(n5345), .ZN(n7075)
         );
  NAND2_X1 U5740 ( .A1(n5520), .A2(n5519), .ZN(n8818) );
  NAND2_X1 U5741 ( .A1(n8253), .A2(n4985), .ZN(n8312) );
  AND2_X1 U5742 ( .A1(n8253), .A2(n5516), .ZN(n8314) );
  AND4_X1 U5743 ( .A1(n5364), .A2(n5363), .A3(n5362), .A4(n5361), .ZN(n7163)
         );
  AND2_X1 U5744 ( .A1(n5411), .A2(n5381), .ZN(n7161) );
  XNOR2_X1 U5745 ( .A(n5561), .B(n5559), .ZN(n8321) );
  INV_X1 U5746 ( .A(n8278), .ZN(n8358) );
  NOR2_X1 U5747 ( .A1(n4989), .A2(n4987), .ZN(n4986) );
  INV_X1 U5748 ( .A(n6627), .ZN(n4987) );
  OR2_X1 U5749 ( .A1(n8278), .A2(n9734), .ZN(n8370) );
  INV_X1 U5750 ( .A(n8376), .ZN(n8353) );
  AND3_X1 U5751 ( .A1(n6068), .A2(n6067), .A3(n6066), .ZN(n7876) );
  AND4_X1 U5752 ( .A1(n5494), .A2(n5493), .A3(n5492), .A4(n5491), .ZN(n8669)
         );
  INV_X1 U5753 ( .A(n9735), .ZN(n8732) );
  INV_X1 U5754 ( .A(n6424), .ZN(n8391) );
  INV_X1 U5755 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5001) );
  NAND2_X1 U5756 ( .A1(n4418), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5189) );
  INV_X1 U5757 ( .A(n9869), .ZN(n9714) );
  INV_X1 U5758 ( .A(n8479), .ZN(n9875) );
  OR2_X1 U5759 ( .A1(n7063), .A2(n9820), .ZN(n8499) );
  INV_X1 U5760 ( .A(n7873), .ZN(n8770) );
  NAND2_X1 U5761 ( .A1(n8485), .A2(n8494), .ZN(n4529) );
  NAND2_X1 U5762 ( .A1(n8553), .A2(n7198), .ZN(n8536) );
  NAND2_X1 U5763 ( .A1(n8578), .A2(n8577), .ZN(n8801) );
  AND2_X1 U5764 ( .A1(n4762), .A2(n7824), .ZN(n8568) );
  NAND2_X1 U5765 ( .A1(n8601), .A2(n7820), .ZN(n8589) );
  AND2_X1 U5766 ( .A1(n5536), .A2(n5535), .ZN(n8600) );
  NAND2_X1 U5767 ( .A1(n4806), .A2(n4809), .ZN(n8630) );
  NAND2_X1 U5768 ( .A1(n8660), .A2(n4810), .ZN(n4806) );
  NAND2_X1 U5769 ( .A1(n8660), .A2(n4813), .ZN(n8645) );
  NAND2_X1 U5770 ( .A1(n4746), .A2(n4749), .ZN(n8703) );
  NAND2_X1 U5771 ( .A1(n7202), .A2(n4752), .ZN(n4746) );
  NAND2_X1 U5772 ( .A1(n8710), .A2(n7192), .ZN(n8695) );
  NAND2_X1 U5773 ( .A1(n4754), .A2(n7792), .ZN(n8721) );
  NAND2_X1 U5774 ( .A1(n4755), .A2(n7789), .ZN(n4754) );
  NAND2_X1 U5775 ( .A1(n9749), .A2(n6841), .ZN(n9747) );
  NAND3_X1 U5776 ( .A1(n4839), .A2(n7697), .A3(n4840), .ZN(n8853) );
  AND2_X1 U5777 ( .A1(n4840), .A2(n4839), .ZN(n7117) );
  NAND2_X1 U5778 ( .A1(n9777), .A2(n4834), .ZN(n7050) );
  AND2_X1 U5779 ( .A1(n9777), .A2(n6882), .ZN(n5000) );
  OR2_X1 U5780 ( .A1(n6296), .A2(n5314), .ZN(n4668) );
  NOR2_X1 U5781 ( .A1(n4456), .A2(n4670), .ZN(n4669) );
  NOR2_X1 U5782 ( .A1(n6513), .A2(n6548), .ZN(n4670) );
  NAND2_X1 U5783 ( .A1(n6874), .A2(n6873), .ZN(n6988) );
  AND2_X1 U5784 ( .A1(n7733), .A2(n7730), .ZN(n6323) );
  OR2_X1 U5785 ( .A1(n6513), .A2(n9427), .ZN(n4671) );
  INV_X1 U5786 ( .A(n8727), .ZN(n8751) );
  NAND2_X1 U5787 ( .A1(n7869), .A2(n5704), .ZN(n9743) );
  INV_X1 U5788 ( .A(n9747), .ZN(n8749) );
  INV_X1 U5789 ( .A(n8499), .ZN(n9727) );
  AND2_X2 U5790 ( .A1(n6290), .A2(n6289), .ZN(n9839) );
  AND2_X2 U5791 ( .A1(n6290), .A2(n6831), .ZN(n9826) );
  NOR2_X1 U5792 ( .A1(n9753), .A2(n9752), .ZN(n9754) );
  AND2_X1 U5793 ( .A1(n7185), .A2(n7069), .ZN(n9756) );
  AND2_X1 U5794 ( .A1(n6142), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9760) );
  INV_X1 U5795 ( .A(n9754), .ZN(n9757) );
  XNOR2_X1 U5796 ( .A(n5678), .B(n5677), .ZN(n7069) );
  NAND2_X1 U5797 ( .A1(n5701), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5678) );
  XNOR2_X1 U5798 ( .A(n5145), .B(n5144), .ZN(n7860) );
  INV_X1 U5799 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10084) );
  INV_X1 U5800 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6204) );
  INV_X1 U5801 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10140) );
  INV_X1 U5802 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10001) );
  INV_X1 U5803 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9996) );
  INV_X1 U5804 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10174) );
  INV_X1 U5805 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5888) );
  INV_X1 U5806 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5877) );
  INV_X1 U5807 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n5869) );
  INV_X1 U5808 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5862) );
  INV_X1 U5809 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10109) );
  INV_X1 U5810 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U5811 ( .A1(n8888), .A2(n8889), .ZN(n8887) );
  NAND2_X1 U5812 ( .A1(n4549), .A2(n4883), .ZN(n8888) );
  AOI21_X1 U5813 ( .B1(n4555), .B2(n4557), .A(n4493), .ZN(n4553) );
  NAND2_X1 U5814 ( .A1(n4917), .A2(n7974), .ZN(n8918) );
  INV_X1 U5815 ( .A(n7974), .ZN(n4910) );
  NAND2_X1 U5816 ( .A1(n6618), .A2(n6617), .ZN(n6642) );
  NAND2_X1 U5817 ( .A1(n4899), .A2(n4902), .ZN(n6643) );
  INV_X1 U5818 ( .A(n6618), .ZN(n4899) );
  NAND2_X1 U5819 ( .A1(n8984), .A2(n8987), .ZN(n8945) );
  INV_X1 U5820 ( .A(n9130), .ZN(n9096) );
  NAND2_X1 U5821 ( .A1(n7268), .A2(n7267), .ZN(n9337) );
  NAND2_X1 U5822 ( .A1(n8962), .A2(n7929), .ZN(n8970) );
  NAND2_X1 U5823 ( .A1(n8926), .A2(n6096), .ZN(n6293) );
  NAND2_X1 U5824 ( .A1(n4898), .A2(n4900), .ZN(n6788) );
  NAND2_X1 U5825 ( .A1(n4533), .A2(n4534), .ZN(n8986) );
  NAND2_X1 U5826 ( .A1(n7290), .A2(n7289), .ZN(n9368) );
  NAND2_X1 U5827 ( .A1(n6942), .A2(n6941), .ZN(n6952) );
  INV_X1 U5828 ( .A(n9177), .ZN(n9207) );
  INV_X1 U5829 ( .A(n4918), .ZN(n8998) );
  NAND2_X1 U5830 ( .A1(n7300), .A2(n7299), .ZN(n9354) );
  NAND2_X1 U5831 ( .A1(n4881), .A2(n6076), .ZN(n6148) );
  NAND2_X1 U5832 ( .A1(n4923), .A2(n4922), .ZN(n9008) );
  AOI21_X1 U5833 ( .B1(n4924), .B2(n4926), .A(n4467), .ZN(n4922) );
  NAND2_X1 U5834 ( .A1(n6399), .A2(n6400), .ZN(n6607) );
  NAND2_X1 U5835 ( .A1(n6398), .A2(n6397), .ZN(n6399) );
  NAND2_X1 U5836 ( .A1(n4554), .A2(n4558), .ZN(n9018) );
  INV_X1 U5837 ( .A(n8978), .ZN(n9034) );
  NAND2_X1 U5838 ( .A1(n4570), .A2(n4569), .ZN(n5997) );
  NAND2_X1 U5839 ( .A1(n4570), .A2(n4462), .ZN(n6017) );
  INV_X1 U5840 ( .A(n4566), .ZN(n9566) );
  AOI21_X1 U5841 ( .B1(n9577), .B2(n9575), .A(n4497), .ZN(n9597) );
  NAND2_X1 U5842 ( .A1(n6000), .A2(n6001), .ZN(n6002) );
  XNOR2_X1 U5843 ( .A(n6720), .B(n9615), .ZN(n9618) );
  NOR2_X1 U5844 ( .A1(n6910), .A2(n6911), .ZN(n6913) );
  NOR2_X1 U5845 ( .A1(n6904), .A2(n6905), .ZN(n6908) );
  INV_X1 U5846 ( .A(n4565), .ZN(n7650) );
  NOR2_X1 U5847 ( .A1(n9058), .A2(n9057), .ZN(n9056) );
  AND2_X1 U5848 ( .A1(n4565), .A2(n4564), .ZN(n9058) );
  NAND2_X1 U5849 ( .A1(n7655), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4564) );
  INV_X1 U5850 ( .A(n9075), .ZN(n9316) );
  INV_X1 U5851 ( .A(n8221), .ZN(n4511) );
  AND2_X1 U5852 ( .A1(n7452), .A2(n7451), .ZN(n8192) );
  INV_X1 U5853 ( .A(n4940), .ZN(n8189) );
  AOI21_X1 U5854 ( .B1(n4934), .B2(n4938), .A(n4941), .ZN(n4933) );
  NAND2_X1 U5855 ( .A1(n4633), .A2(n4465), .ZN(n9326) );
  NAND2_X1 U5856 ( .A1(n9079), .A2(n9088), .ZN(n4633) );
  NAND2_X1 U5857 ( .A1(n4936), .A2(n4937), .ZN(n9079) );
  AOI21_X1 U5858 ( .B1(n9090), .B2(n9296), .A(n4801), .ZN(n9325) );
  NAND2_X1 U5859 ( .A1(n4803), .A2(n4802), .ZN(n4801) );
  NAND2_X1 U5860 ( .A1(n9089), .A2(n9293), .ZN(n4803) );
  AOI21_X1 U5861 ( .B1(n9333), .B2(n9650), .A(n9120), .ZN(n4599) );
  AND2_X1 U5862 ( .A1(n4603), .A2(n4601), .ZN(n9335) );
  AOI21_X1 U5863 ( .B1(n9117), .B2(n9293), .A(n4602), .ZN(n4601) );
  NAND2_X1 U5864 ( .A1(n9119), .A2(n9296), .ZN(n4603) );
  NOR2_X1 U5865 ( .A1(n9141), .A2(n9464), .ZN(n4602) );
  NAND2_X1 U5866 ( .A1(n4789), .A2(n4796), .ZN(n9128) );
  INV_X1 U5867 ( .A(n4956), .ZN(n9167) );
  OAI21_X1 U5868 ( .B1(n9250), .B2(n4591), .A(n4588), .ZN(n9225) );
  NAND2_X1 U5869 ( .A1(n4593), .A2(n4590), .ZN(n9237) );
  NAND2_X1 U5870 ( .A1(n4621), .A2(n8177), .ZN(n9249) );
  NAND2_X1 U5871 ( .A1(n4783), .A2(n4784), .ZN(n6819) );
  NAND2_X1 U5872 ( .A1(n9453), .A2(n9460), .ZN(n6818) );
  OR2_X1 U5873 ( .A1(n4419), .A2(n5966), .ZN(n9656) );
  AND2_X1 U5874 ( .A1(n6406), .A2(n6346), .ZN(n6585) );
  NAND2_X1 U5875 ( .A1(n5839), .A2(n9258), .ZN(n9281) );
  INV_X1 U5876 ( .A(n9258), .ZN(n9652) );
  INV_X1 U5877 ( .A(n9656), .ZN(n9469) );
  AND2_X1 U5878 ( .A1(n6998), .A2(n5833), .ZN(n7641) );
  AND2_X1 U5879 ( .A1(n4959), .A2(n5763), .ZN(n4958) );
  AND2_X1 U5880 ( .A1(n5768), .A2(n4960), .ZN(n4959) );
  INV_X1 U5881 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4960) );
  XNOR2_X1 U5882 ( .A(n5756), .B(n5755), .ZN(n6846) );
  INV_X1 U5883 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10056) );
  INV_X1 U5884 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6202) );
  INV_X1 U5885 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6141) );
  INV_X1 U5886 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6061) );
  INV_X1 U5887 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10204) );
  INV_X1 U5888 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5876) );
  INV_X1 U5889 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5858) );
  INV_X1 U5890 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10108) );
  NAND2_X1 U5891 ( .A1(n4640), .A2(n5014), .ZN(n5240) );
  NAND2_X1 U5892 ( .A1(n5221), .A2(n5220), .ZN(n4640) );
  NOR2_X1 U5893 ( .A1(n5775), .A2(n9415), .ZN(n5792) );
  INV_X1 U5894 ( .A(n5775), .ZN(n5776) );
  NOR2_X1 U5895 ( .A1(n9510), .A2(n10209), .ZN(n9868) );
  AOI21_X1 U5896 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9866), .ZN(n9865) );
  NOR2_X1 U5897 ( .A1(n9865), .A2(n9864), .ZN(n9863) );
  OAI211_X1 U5898 ( .C1(n4967), .C2(n5711), .A(n4966), .B(n5710), .ZN(n4965)
         );
  AOI21_X1 U5899 ( .B1(n4760), .B2(n4761), .A(n4759), .ZN(n4758) );
  INV_X1 U5900 ( .A(n7872), .ZN(n4759) );
  NAND2_X1 U5901 ( .A1(n4523), .A2(n4520), .ZN(P2_U3264) );
  NAND2_X1 U5902 ( .A1(n8477), .A2(n7711), .ZN(n4523) );
  AOI21_X1 U5903 ( .B1(n8476), .B2(n8546), .A(n4521), .ZN(n4520) );
  NAND2_X1 U5904 ( .A1(n4889), .A2(n9015), .ZN(n4888) );
  NAND2_X1 U5905 ( .A1(n4519), .A2(n4517), .ZN(P1_U3260) );
  AOI21_X1 U5906 ( .B1(n7663), .B2(n9243), .A(n4518), .ZN(n4517) );
  NAND2_X1 U5907 ( .A1(n7662), .A2(n7661), .ZN(n4519) );
  OAI21_X1 U5908 ( .B1(n9627), .B2(n4657), .A(n8939), .ZN(n4518) );
  OAI21_X1 U5909 ( .B1(n9325), .B2(n4419), .A(n4800), .ZN(P1_U3263) );
  INV_X1 U5910 ( .A(n4631), .ZN(n4800) );
  OAI21_X1 U5911 ( .B1(n9326), .B2(n9308), .A(n4632), .ZN(n4631) );
  AOI21_X1 U5912 ( .B1(n9323), .B2(n9650), .A(n9091), .ZN(n4632) );
  NAND2_X1 U5913 ( .A1(n4600), .A2(n4597), .ZN(P1_U3265) );
  OR2_X1 U5914 ( .A1(n9335), .A2(n4419), .ZN(n4600) );
  INV_X1 U5915 ( .A(n4598), .ZN(n4597) );
  OAI21_X1 U5916 ( .B1(n9336), .B2(n9308), .A(n4599), .ZN(n4598) );
  INV_X1 U5917 ( .A(n4724), .ZN(n9398) );
  INV_X1 U5918 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n4723) );
  INV_X2 U5920 ( .A(n5200), .ZN(n5208) );
  INV_X1 U5921 ( .A(n4414), .ZN(n6097) );
  INV_X1 U5922 ( .A(n8889), .ZN(n4542) );
  INV_X1 U5923 ( .A(n4972), .ZN(n4821) );
  NOR2_X1 U5924 ( .A1(n8188), .A2(n4943), .ZN(n4939) );
  NAND2_X1 U5925 ( .A1(n5656), .A2(n5655), .ZN(n8776) );
  INV_X1 U5926 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U5927 ( .A1(n7146), .A2(n5403), .ZN(n4425) );
  AND2_X1 U5928 ( .A1(n8587), .A2(n8600), .ZN(n4426) );
  AND2_X1 U5929 ( .A1(n4563), .A2(n5954), .ZN(n7998) );
  AND2_X1 U5930 ( .A1(n4685), .A2(n4684), .ZN(n4428) );
  AND2_X1 U5931 ( .A1(n4426), .A2(n4696), .ZN(n4429) );
  INV_X1 U5932 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9415) );
  AND2_X1 U5933 ( .A1(n7626), .A2(n7529), .ZN(n4430) );
  NAND2_X1 U5934 ( .A1(n7329), .A2(n7328), .ZN(n9372) );
  AND2_X1 U5935 ( .A1(n4891), .A2(n4471), .ZN(n4431) );
  INV_X1 U5936 ( .A(n8735), .ZN(n6880) );
  NAND2_X1 U5937 ( .A1(n5454), .A2(n5453), .ZN(n8843) );
  NOR2_X1 U5938 ( .A1(n8824), .A2(n8652), .ZN(n4432) );
  INV_X1 U5939 ( .A(n6225), .ZN(n8930) );
  AND2_X1 U5940 ( .A1(n5804), .A2(n5803), .ZN(n4433) );
  INV_X1 U5941 ( .A(n9118), .ZN(n9141) );
  OR2_X1 U5942 ( .A1(n8808), .A2(n8248), .ZN(n7824) );
  NAND2_X1 U5943 ( .A1(n4669), .A2(n4668), .ZN(n6987) );
  INV_X1 U5944 ( .A(n6987), .ZN(n9770) );
  AND2_X1 U5945 ( .A1(n4744), .A2(n7800), .ZN(n4434) );
  AND2_X1 U5946 ( .A1(n5414), .A2(n4503), .ZN(n4435) );
  NOR2_X1 U5947 ( .A1(n6142), .A2(P2_U3152), .ZN(n7867) );
  NAND2_X1 U5948 ( .A1(n4915), .A2(n4914), .ZN(n4918) );
  OR2_X1 U5949 ( .A1(n8481), .A2(n8492), .ZN(n4436) );
  OR2_X1 U5950 ( .A1(n5447), .A2(n4858), .ZN(n4437) );
  AND2_X1 U5951 ( .A1(n5046), .A2(n5045), .ZN(n4438) );
  NAND2_X1 U5952 ( .A1(n8650), .A2(n4999), .ZN(n8617) );
  INV_X1 U5953 ( .A(n9460), .ZN(n4788) );
  INV_X1 U5954 ( .A(n4591), .ZN(n4590) );
  NAND2_X1 U5955 ( .A1(n9238), .A2(n4592), .ZN(n4591) );
  OR2_X1 U5956 ( .A1(n5353), .A2(n4864), .ZN(n4440) );
  INV_X1 U5957 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4562) );
  NOR2_X1 U5958 ( .A1(n6200), .A2(n4932), .ZN(n5743) );
  INV_X1 U5959 ( .A(n8200), .ZN(n4592) );
  AND2_X1 U5960 ( .A1(n8520), .A2(n8528), .ZN(n4441) );
  AND4_X1 U5961 ( .A1(n5124), .A2(n5123), .A3(n5667), .A4(n5122), .ZN(n4442)
         );
  AND3_X1 U5962 ( .A1(n6221), .A2(n5799), .A3(n4562), .ZN(n4443) );
  OR2_X1 U5963 ( .A1(n6297), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4444) );
  NAND2_X1 U5964 ( .A1(n7987), .A2(n7986), .ZN(n4445) );
  AND2_X1 U5965 ( .A1(n4905), .A2(n4912), .ZN(n4446) );
  AND2_X1 U5966 ( .A1(n5455), .A2(n4970), .ZN(n4447) );
  INV_X1 U5967 ( .A(n8661), .ZN(n4645) );
  NOR2_X1 U5968 ( .A1(n9345), .A2(n8956), .ZN(n8210) );
  INV_X1 U5969 ( .A(n8210), .ZN(n4799) );
  AND2_X1 U5970 ( .A1(n4799), .A2(n9155), .ZN(n4448) );
  INV_X1 U5971 ( .A(n4778), .ZN(n4777) );
  NAND2_X1 U5972 ( .A1(n4441), .A2(n4779), .ZN(n4778) );
  NAND2_X1 U5973 ( .A1(n7198), .A2(n7197), .ZN(n8556) );
  INV_X1 U5974 ( .A(n8556), .ZN(n4661) );
  INV_X1 U5975 ( .A(n8202), .ZN(n4589) );
  INV_X1 U5976 ( .A(n8214), .ZN(n4791) );
  AND2_X1 U5977 ( .A1(n7856), .A2(n7859), .ZN(n4449) );
  AND2_X1 U5978 ( .A1(n7538), .A2(n7536), .ZN(n4450) );
  OR2_X1 U5979 ( .A1(n7013), .A2(n4788), .ZN(n4451) );
  NOR2_X1 U5980 ( .A1(n8522), .A2(n8781), .ZN(n8509) );
  INV_X1 U5981 ( .A(n8509), .ZN(n4682) );
  XNOR2_X1 U5982 ( .A(n8387), .B(n7062), .ZN(n9730) );
  AND2_X1 U5983 ( .A1(n7760), .A2(n7761), .ZN(n7757) );
  INV_X1 U5984 ( .A(n8977), .ZN(n4916) );
  NOR2_X1 U5985 ( .A1(n7112), .A2(n7698), .ZN(n4452) );
  AND2_X1 U5986 ( .A1(n7820), .A2(n7821), .ZN(n4453) );
  AND2_X1 U5987 ( .A1(n4784), .A2(n4782), .ZN(n4454) );
  NAND2_X1 U5988 ( .A1(n8994), .A2(n8997), .ZN(n4919) );
  OR2_X1 U5989 ( .A1(n4682), .A2(n4681), .ZN(n4455) );
  NAND2_X1 U5990 ( .A1(n5568), .A2(n5567), .ZN(n8803) );
  INV_X1 U5991 ( .A(n8803), .ZN(n4696) );
  NAND2_X1 U5992 ( .A1(n4974), .A2(n4973), .ZN(n5291) );
  NOR2_X1 U5993 ( .A1(n7674), .A2(n10109), .ZN(n4456) );
  NAND2_X1 U5994 ( .A1(n7353), .A2(n7352), .ZN(n9349) );
  INV_X1 U5995 ( .A(n9349), .ZN(n4734) );
  AND3_X1 U5996 ( .A1(n8283), .A2(n5458), .A3(n8284), .ZN(n4457) );
  NAND2_X1 U5997 ( .A1(n7279), .A2(n7278), .ZN(n9362) );
  NAND2_X1 U5998 ( .A1(n7369), .A2(n7368), .ZN(n9388) );
  NAND2_X1 U5999 ( .A1(n7356), .A2(n7355), .ZN(n9345) );
  AND2_X1 U6000 ( .A1(n7467), .A2(n8217), .ZN(n9088) );
  NAND2_X1 U6001 ( .A1(n5598), .A2(n5597), .ZN(n8792) );
  AND2_X1 U6002 ( .A1(n4968), .A2(n5461), .ZN(n4458) );
  OR2_X1 U6003 ( .A1(n7583), .A2(n7584), .ZN(n4459) );
  AND2_X1 U6004 ( .A1(n4990), .A2(n5247), .ZN(n4460) );
  NAND2_X1 U6005 ( .A1(n7148), .A2(n7158), .ZN(n4461) );
  AND2_X1 U6006 ( .A1(n4569), .A2(n4444), .ZN(n4462) );
  INV_X1 U6007 ( .A(n4615), .ZN(n4614) );
  NOR2_X1 U6008 ( .A1(n6684), .A2(n4616), .ZN(n4615) );
  AND2_X1 U6009 ( .A1(n4596), .A2(n4595), .ZN(n4463) );
  AND2_X1 U6010 ( .A1(n4977), .A2(n4976), .ZN(n4464) );
  INV_X1 U6011 ( .A(n4939), .ZN(n4938) );
  INV_X1 U6012 ( .A(n7193), .ZN(n4827) );
  NAND2_X1 U6013 ( .A1(n4936), .A2(n4934), .ZN(n4465) );
  AND2_X1 U6014 ( .A1(n9354), .A2(n9162), .ZN(n4466) );
  AND2_X1 U6015 ( .A1(n7936), .A2(n7935), .ZN(n4467) );
  AND2_X1 U6016 ( .A1(n7807), .A2(n7809), .ZN(n4468) );
  NOR2_X1 U6017 ( .A1(n7008), .A2(n7007), .ZN(n4469) );
  INV_X1 U6018 ( .A(n7471), .ZN(n4525) );
  INV_X1 U6019 ( .A(n4943), .ZN(n4942) );
  NOR2_X1 U6020 ( .A1(n9096), .A2(n9112), .ZN(n4943) );
  AND2_X1 U6021 ( .A1(n9735), .A2(n9783), .ZN(n4470) );
  NAND2_X1 U6022 ( .A1(n4890), .A2(n4894), .ZN(n4471) );
  OR2_X1 U6023 ( .A1(n8781), .A2(n8357), .ZN(n7843) );
  INV_X1 U6024 ( .A(n7843), .ZN(n4770) );
  AND2_X1 U6025 ( .A1(n9383), .A2(n9239), .ZN(n4472) );
  AND2_X1 U6026 ( .A1(n7847), .A2(n4652), .ZN(n4473) );
  NOR2_X1 U6027 ( .A1(n8635), .A2(n8624), .ZN(n4474) );
  NOR2_X1 U6028 ( .A1(n8792), .A2(n8379), .ZN(n4475) );
  INV_X1 U6029 ( .A(n6400), .ZN(n4885) );
  AND2_X1 U6030 ( .A1(n7854), .A2(n7842), .ZN(n4476) );
  NAND3_X1 U6031 ( .A1(n4919), .A2(n4918), .A3(n4910), .ZN(n4477) );
  OR2_X1 U6032 ( .A1(n5797), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n4478) );
  INV_X1 U6033 ( .A(n4739), .ZN(n4738) );
  NAND2_X1 U6034 ( .A1(n4741), .A2(n4740), .ZN(n4739) );
  INV_X1 U6035 ( .A(n8215), .ZN(n4793) );
  NOR2_X1 U6036 ( .A1(n9328), .A2(n9117), .ZN(n4479) );
  INV_X1 U6037 ( .A(n4835), .ZN(n4834) );
  NAND2_X1 U6038 ( .A1(n6891), .A2(n6882), .ZN(n4835) );
  AND2_X1 U6039 ( .A1(n7947), .A2(n7946), .ZN(n4480) );
  INV_X1 U6040 ( .A(n4831), .ZN(n4830) );
  NAND2_X1 U6041 ( .A1(n7705), .A2(n4832), .ZN(n4831) );
  INV_X1 U6042 ( .A(n8776), .ZN(n8485) );
  INV_X1 U6043 ( .A(n4811), .ZN(n4810) );
  NAND2_X1 U6044 ( .A1(n4812), .A2(n4813), .ZN(n4811) );
  INV_X1 U6045 ( .A(n7192), .ZN(n4825) );
  AND2_X1 U6046 ( .A1(n4751), .A2(n7801), .ZN(n4481) );
  INV_X1 U6047 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5799) );
  AND2_X1 U6048 ( .A1(n7849), .A2(n7850), .ZN(n8488) );
  NOR2_X1 U6049 ( .A1(n9238), .A2(n8181), .ZN(n4482) );
  AND2_X1 U6050 ( .A1(n4789), .A2(n4794), .ZN(n4483) );
  INV_X1 U6051 ( .A(n8512), .ZN(n8507) );
  AND2_X1 U6052 ( .A1(n8618), .A2(n8619), .ZN(n4484) );
  AND2_X1 U6053 ( .A1(n5935), .A2(n4571), .ZN(n4485) );
  AND2_X1 U6054 ( .A1(n5750), .A2(n5745), .ZN(n4486) );
  NAND2_X1 U6055 ( .A1(n8002), .A2(n8897), .ZN(n4487) );
  AND2_X1 U6056 ( .A1(n5014), .A2(n5009), .ZN(n4488) );
  AND2_X1 U6057 ( .A1(n4744), .A2(n4743), .ZN(n4489) );
  AND2_X1 U6058 ( .A1(n5799), .A2(n4562), .ZN(n4490) );
  INV_X1 U6059 ( .A(n4978), .ZN(n4977) );
  NAND2_X1 U6060 ( .A1(n4979), .A2(n5334), .ZN(n4978) );
  INV_X1 U6061 ( .A(n4935), .ZN(n4934) );
  NAND2_X1 U6062 ( .A1(n4937), .A2(n7493), .ZN(n4935) );
  NAND2_X1 U6063 ( .A1(n6276), .A2(n6869), .ZN(n6322) );
  NAND2_X1 U6064 ( .A1(n4524), .A2(n7540), .ZN(n4610) );
  NAND2_X1 U6065 ( .A1(n5132), .A2(n5131), .ZN(n8796) );
  INV_X1 U6066 ( .A(n8796), .ZN(n4695) );
  INV_X1 U6067 ( .A(n7627), .ZN(n4706) );
  INV_X1 U6068 ( .A(n8919), .ZN(n4913) );
  INV_X1 U6069 ( .A(n8781), .ZN(n4679) );
  AND4_X1 U6070 ( .A1(n5540), .A2(n5539), .A3(n5538), .A4(n5537), .ZN(n8623)
         );
  INV_X1 U6071 ( .A(n8623), .ZN(n8380) );
  AND4_X1 U6072 ( .A1(n5474), .A2(n5473), .A3(n5472), .A4(n5471), .ZN(n8680)
         );
  NAND2_X1 U6073 ( .A1(n8183), .A2(n8182), .ZN(n9201) );
  NAND2_X1 U6074 ( .A1(n4539), .A2(n4540), .ZN(n8935) );
  INV_X1 U6075 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4819) );
  AND2_X1 U6076 ( .A1(n4550), .A2(n9026), .ZN(n4491) );
  OR2_X1 U6077 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n9562), .ZN(n4492) );
  AND2_X1 U6078 ( .A1(n7992), .A2(n7994), .ZN(n4493) );
  AND2_X1 U6079 ( .A1(n6687), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4494) );
  NAND2_X1 U6080 ( .A1(n5120), .A2(n4836), .ZN(n5485) );
  NAND2_X1 U6081 ( .A1(n4768), .A2(n7768), .ZN(n7128) );
  NAND2_X1 U6082 ( .A1(n4821), .A2(n4974), .ZN(n5309) );
  NAND2_X1 U6083 ( .A1(n5120), .A2(n5119), .ZN(n5366) );
  NAND2_X1 U6084 ( .A1(n5414), .A2(n4991), .ZN(n5433) );
  INV_X1 U6085 ( .A(n4752), .ZN(n4751) );
  NOR2_X1 U6086 ( .A1(n8711), .A2(n4753), .ZN(n4752) );
  NAND2_X1 U6087 ( .A1(n9208), .A2(n4733), .ZN(n4736) );
  NAND2_X1 U6088 ( .A1(n9284), .A2(n4738), .ZN(n4742) );
  NAND2_X1 U6089 ( .A1(n8612), .A2(n4694), .ZN(n4495) );
  NAND2_X1 U6090 ( .A1(n7953), .A2(n7954), .ZN(n4496) );
  AND2_X1 U6091 ( .A1(n5120), .A2(n4837), .ZN(n5414) );
  AND2_X1 U6092 ( .A1(n9580), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4497) );
  OR2_X1 U6093 ( .A1(n8302), .A2(n8306), .ZN(n4498) );
  NOR2_X1 U6094 ( .A1(n5726), .A2(n5727), .ZN(n4499) );
  AND2_X1 U6095 ( .A1(n4593), .A2(n4592), .ZN(n4500) );
  AND2_X1 U6096 ( .A1(n5760), .A2(n5759), .ZN(n5807) );
  NAND2_X1 U6097 ( .A1(n5466), .A2(n5465), .ZN(n8835) );
  INV_X1 U6098 ( .A(n8835), .ZN(n4814) );
  AND2_X1 U6099 ( .A1(n7531), .A2(n7536), .ZN(n7411) );
  INV_X1 U6100 ( .A(n7411), .ZN(n4584) );
  INV_X1 U6101 ( .A(n7499), .ZN(n4583) );
  NAND2_X1 U6102 ( .A1(n5436), .A2(n5435), .ZN(n8838) );
  INV_X1 U6103 ( .A(n8838), .ZN(n4684) );
  OR2_X1 U6104 ( .A1(n9671), .A2(n4723), .ZN(n4501) );
  OR2_X1 U6105 ( .A1(n9724), .A2(n4689), .ZN(n4502) );
  AND2_X1 U6106 ( .A1(n4991), .A2(n4980), .ZN(n4503) );
  INV_X1 U6107 ( .A(n4730), .ZN(n6577) );
  AND2_X1 U6108 ( .A1(n4575), .A2(n4576), .ZN(n4504) );
  INV_X1 U6109 ( .A(n7800), .ZN(n4747) );
  NAND2_X1 U6110 ( .A1(n6002), .A2(n6003), .ZN(n4505) );
  INV_X1 U6111 ( .A(n5263), .ZN(n4989) );
  NAND2_X1 U6112 ( .A1(n4947), .A2(n6345), .ZN(n6406) );
  AND2_X1 U6113 ( .A1(n7219), .A2(n9998), .ZN(n4506) );
  AND2_X1 U6114 ( .A1(n4988), .A2(n5263), .ZN(n4507) );
  XNOR2_X1 U6115 ( .A(n5127), .B(n5147), .ZN(n5721) );
  INV_X1 U6116 ( .A(n7400), .ZN(n4636) );
  AND2_X1 U6117 ( .A1(n9674), .A2(n6192), .ZN(n4508) );
  INV_X1 U6118 ( .A(n9464), .ZN(n9291) );
  INV_X1 U6119 ( .A(n6271), .ZN(n6449) );
  NAND2_X1 U6120 ( .A1(n6559), .A2(n6558), .ZN(n9690) );
  INV_X1 U6121 ( .A(n9690), .ZN(n4729) );
  NAND2_X1 U6122 ( .A1(n5358), .A2(n5357), .ZN(n9816) );
  INV_X1 U6123 ( .A(n9816), .ZN(n4688) );
  NAND2_X1 U6124 ( .A1(n5965), .A2(n5953), .ZN(n9038) );
  AND2_X1 U6125 ( .A1(n7683), .A2(n7682), .ZN(n4509) );
  NAND2_X1 U6126 ( .A1(n6432), .A2(n4677), .ZN(n6983) );
  INV_X1 U6127 ( .A(n6983), .ZN(n4676) );
  INV_X1 U6128 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5449) );
  INV_X1 U6129 ( .A(n9243), .ZN(n7661) );
  NAND2_X1 U6130 ( .A1(n5139), .A2(n5143), .ZN(n8546) );
  AND2_X1 U6131 ( .A1(n5930), .A2(n5929), .ZN(n4510) );
  INV_X1 U6132 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4656) );
  NAND2_X1 U6133 ( .A1(n5010), .A2(n4488), .ZN(n4639) );
  OAI22_X2 U6134 ( .A1(n8508), .A2(n8512), .B1(n8781), .B2(n8378), .ZN(n8487)
         );
  NAND2_X1 U6135 ( .A1(n4745), .A2(n4489), .ZN(n4756) );
  NAND2_X1 U6136 ( .A1(n4773), .A2(n4774), .ZN(n8513) );
  NAND3_X1 U6137 ( .A1(n4639), .A2(n4638), .A3(n5239), .ZN(n4527) );
  INV_X1 U6138 ( .A(n7016), .ZN(n4526) );
  NOR2_X2 U6139 ( .A1(n9175), .A2(n8208), .ZN(n9160) );
  INV_X1 U6140 ( .A(n7485), .ZN(n4782) );
  NOR2_X1 U6141 ( .A1(n9094), .A2(n9095), .ZN(n9093) );
  NAND2_X1 U6142 ( .A1(n8265), .A2(n5544), .ZN(n5561) );
  NAND2_X1 U6143 ( .A1(n8240), .A2(n8239), .ZN(n8238) );
  NAND2_X1 U6144 ( .A1(n4527), .A2(n5017), .ZN(n5258) );
  NAND2_X1 U6145 ( .A1(n4962), .A2(n5627), .ZN(n8352) );
  NAND2_X1 U6146 ( .A1(n4965), .A2(n4499), .ZN(P2_U3222) );
  AND3_X2 U6147 ( .A1(n4726), .A2(n4727), .A3(n4728), .ZN(n5765) );
  NAND2_X1 U6148 ( .A1(n4783), .A2(n4454), .ZN(n7015) );
  NOR2_X1 U6149 ( .A1(n9320), .A2(n4419), .ZN(n8222) );
  OAI211_X1 U6150 ( .C1(n6373), .C2(n4584), .A(n4582), .B(n6375), .ZN(n6376)
         );
  XNOR2_X1 U6151 ( .A(n4528), .B(n8489), .ZN(n8769) );
  NAND2_X1 U6152 ( .A1(n4530), .A2(n4529), .ZN(n4528) );
  NAND2_X1 U6153 ( .A1(n8487), .A2(n8486), .ZN(n4530) );
  XNOR2_X2 U6154 ( .A(n5335), .B(n4438), .ZN(n6686) );
  INV_X1 U6155 ( .A(n7116), .ZN(n4840) );
  NAND2_X1 U6156 ( .A1(n4548), .A2(n4547), .ZN(n4546) );
  NAND3_X1 U6157 ( .A1(n4546), .A2(n6615), .A3(n4543), .ZN(n6618) );
  NAND3_X1 U6158 ( .A1(n4546), .A2(n4544), .A3(n4543), .ZN(n4898) );
  NAND3_X1 U6159 ( .A1(n4550), .A2(n9026), .A3(n4924), .ZN(n4923) );
  NAND2_X1 U6160 ( .A1(n7919), .A2(n8907), .ZN(n4551) );
  NAND3_X1 U6161 ( .A1(n7919), .A2(n8907), .A3(n7920), .ZN(n9025) );
  NAND2_X1 U6162 ( .A1(n4904), .A2(n4555), .ZN(n4552) );
  OAI21_X1 U6163 ( .B1(n4904), .B2(n4557), .A(n4555), .ZN(n9016) );
  NAND2_X1 U6164 ( .A1(n4904), .A2(n4560), .ZN(n4554) );
  NAND2_X1 U6165 ( .A1(n4552), .A2(n4553), .ZN(n8900) );
  NAND2_X1 U6166 ( .A1(n4904), .A2(n4903), .ZN(n8953) );
  NAND2_X1 U6167 ( .A1(n4930), .A2(n4561), .ZN(n5753) );
  NAND2_X1 U6168 ( .A1(n4930), .A2(n4929), .ZN(n5797) );
  XNOR2_X1 U6169 ( .A(n6047), .B(n7998), .ZN(n6052) );
  NAND2_X1 U6170 ( .A1(n5930), .A2(n4485), .ZN(n4570) );
  NAND2_X1 U6171 ( .A1(n4575), .A2(n4573), .ZN(n9607) );
  NAND2_X1 U6172 ( .A1(n6373), .A2(n7499), .ZN(n7532) );
  NAND2_X1 U6173 ( .A1(n9250), .A2(n4588), .ZN(n4585) );
  NAND2_X1 U6174 ( .A1(n4585), .A2(n4586), .ZN(n9224) );
  NAND2_X1 U6175 ( .A1(n4594), .A2(n4463), .ZN(n5767) );
  NAND4_X1 U6176 ( .A1(n4726), .A2(n4728), .A3(n4727), .A4(
        P1_IR_REG_27__SCAN_IN), .ZN(n4594) );
  NAND2_X1 U6177 ( .A1(n4610), .A2(n4607), .ZN(n4783) );
  NAND2_X1 U6178 ( .A1(n4433), .A2(n6183), .ZN(n6209) );
  NAND2_X1 U6179 ( .A1(n4621), .A2(n4619), .ZN(n4945) );
  NAND4_X1 U6180 ( .A1(n4726), .A2(n4728), .A3(n5763), .A4(n4727), .ZN(n5766)
         );
  OAI21_X1 U6181 ( .B1(n8183), .B2(n4624), .A(n4622), .ZN(n4956) );
  NAND2_X1 U6182 ( .A1(n4627), .A2(n4630), .ZN(n9195) );
  NAND2_X1 U6183 ( .A1(n4950), .A2(n4635), .ZN(n6185) );
  NAND2_X1 U6184 ( .A1(n5014), .A2(n4637), .ZN(n4638) );
  INV_X1 U6185 ( .A(n5220), .ZN(n4637) );
  NAND3_X1 U6186 ( .A1(n4657), .A2(n4656), .A3(n4655), .ZN(n4654) );
  INV_X2 U6187 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4655) );
  NAND4_X1 U6188 ( .A1(n4663), .A2(n7839), .A3(n4662), .A4(n4658), .ZN(n7838)
         );
  NAND3_X1 U6189 ( .A1(n4659), .A2(n7842), .A3(n4664), .ZN(n4658) );
  INV_X1 U6190 ( .A(n7828), .ZN(n4659) );
  NAND3_X1 U6191 ( .A1(n7835), .A2(n7833), .A3(n7859), .ZN(n4662) );
  NAND4_X1 U6192 ( .A1(n4664), .A2(n7826), .A3(n7827), .A4(n4660), .ZN(n4663)
         );
  NOR2_X1 U6193 ( .A1(n7834), .A2(n4665), .ZN(n4664) );
  NAND3_X1 U6194 ( .A1(n7860), .A2(n4667), .A3(n4666), .ZN(n7861) );
  XNOR2_X1 U6195 ( .A(n5258), .B(n5257), .ZN(n6296) );
  NAND2_X1 U6196 ( .A1(n4818), .A2(n4675), .ZN(n5355) );
  NOR2_X2 U6197 ( .A1(n4972), .A2(n5236), .ZN(n4675) );
  AND4_X2 U6198 ( .A1(n4442), .A2(n4675), .A3(n4836), .A4(n4673), .ZN(n5148)
         );
  INV_X1 U6199 ( .A(n9724), .ZN(n4686) );
  NAND2_X1 U6200 ( .A1(n4686), .A2(n4687), .ZN(n7118) );
  NAND2_X1 U6201 ( .A1(n8612), .A2(n4692), .ZN(n8543) );
  NAND2_X1 U6202 ( .A1(n4701), .A2(n4697), .ZN(n7546) );
  NAND2_X1 U6203 ( .A1(n4707), .A2(n4705), .ZN(n4704) );
  NAND4_X1 U6204 ( .A1(n4714), .A2(n7553), .A3(n4713), .A4(n4712), .ZN(n4711)
         );
  NAND3_X1 U6205 ( .A1(n7548), .A2(n7627), .A3(n7547), .ZN(n4713) );
  NAND4_X1 U6206 ( .A1(n7543), .A2(n6711), .A3(n9460), .A4(n4706), .ZN(n4714)
         );
  NAND2_X1 U6207 ( .A1(n4715), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U6208 ( .A1(n5765), .A2(n4716), .ZN(n4715) );
  AOI21_X2 U6209 ( .B1(n4718), .B2(n4430), .A(n4717), .ZN(n7635) );
  NAND3_X1 U6210 ( .A1(n7621), .A2(n7620), .A3(n4720), .ZN(n4719) );
  OAI21_X1 U6211 ( .B1(n7586), .B2(n4459), .A(n4722), .ZN(n7590) );
  OAI21_X1 U6212 ( .B1(n4724), .B2(n9698), .A(n4501), .ZN(P1_U3522) );
  NAND4_X1 U6213 ( .A1(n4728), .A2(n4727), .A3(n4427), .A4(n4424), .ZN(n5762)
         );
  INV_X1 U6214 ( .A(n4736), .ZN(n9151) );
  NAND2_X1 U6215 ( .A1(n9284), .A2(n4737), .ZN(n9218) );
  INV_X1 U6216 ( .A(n4742), .ZN(n9242) );
  OR2_X2 U6217 ( .A1(n7202), .A2(n4748), .ZN(n4745) );
  NAND2_X1 U6218 ( .A1(n4757), .A2(n4758), .ZN(P2_U3244) );
  NAND2_X1 U6219 ( .A1(n7684), .A2(n4760), .ZN(n4757) );
  AOI21_X2 U6220 ( .B1(n4998), .B2(n4509), .A(n7871), .ZN(n4760) );
  NAND2_X1 U6221 ( .A1(n8601), .A2(n4764), .ZN(n4766) );
  CLKBUF_X1 U6222 ( .A(n4766), .Z(n4762) );
  INV_X1 U6223 ( .A(n4762), .ZN(n8588) );
  NAND2_X1 U6224 ( .A1(n4768), .A2(n4767), .ZN(n7129) );
  OR2_X1 U6225 ( .A1(n8559), .A2(n4778), .ZN(n4773) );
  NAND2_X1 U6226 ( .A1(n8559), .A2(n4772), .ZN(n4771) );
  AND2_X2 U6227 ( .A1(n8617), .A2(n4484), .ZN(n8622) );
  AND2_X2 U6228 ( .A1(n5148), .A2(n5147), .ZN(n5151) );
  AOI21_X2 U6229 ( .B1(n7532), .B2(n7531), .A(n7530), .ZN(n7533) );
  NAND2_X1 U6230 ( .A1(n6211), .A2(n7402), .ZN(n6232) );
  NAND2_X1 U6231 ( .A1(n7473), .A2(n6187), .ZN(n6186) );
  NAND2_X1 U6232 ( .A1(n7208), .A2(n7207), .ZN(n7664) );
  AOI21_X2 U6233 ( .B1(n7110), .B2(n7783), .A(n7109), .ZN(n7202) );
  NOR2_X2 U6234 ( .A1(n8560), .A2(n4661), .ZN(n8559) );
  NAND2_X1 U6235 ( .A1(n6496), .A2(n6495), .ZN(n6887) );
  OAI211_X2 U6236 ( .C1(n6513), .C2(n9882), .A(n5296), .B(n5295), .ZN(n6886)
         );
  INV_X1 U6237 ( .A(n7757), .ZN(n6891) );
  NAND2_X1 U6238 ( .A1(n8660), .A2(n4807), .ZN(n4804) );
  NAND2_X1 U6239 ( .A1(n4804), .A2(n4805), .ZN(n8611) );
  NAND2_X1 U6240 ( .A1(n6490), .A2(n7685), .ZN(n6874) );
  NOR2_X1 U6241 ( .A1(n5236), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n4820) );
  NAND2_X1 U6242 ( .A1(n9721), .A2(n4841), .ZN(n4839) );
  AOI21_X2 U6243 ( .B1(n5099), .B2(n5533), .A(n4995), .ZN(n5545) );
  NAND2_X1 U6244 ( .A1(n5653), .A2(n4846), .ZN(n4844) );
  NAND2_X1 U6245 ( .A1(n5063), .A2(n4856), .ZN(n4853) );
  NAND2_X1 U6246 ( .A1(n4853), .A2(n4854), .ZN(n5079) );
  NAND2_X1 U6247 ( .A1(n5063), .A2(n5062), .ZN(n5413) );
  OAI21_X2 U6248 ( .B1(n5047), .B2(n4440), .A(n4862), .ZN(n5365) );
  OAI21_X1 U6249 ( .B1(n5313), .B2(n5311), .A(n5035), .ZN(n5326) );
  NAND2_X1 U6250 ( .A1(n6075), .A2(n6074), .ZN(n4881) );
  INV_X1 U6251 ( .A(n6053), .ZN(n4882) );
  NAND2_X1 U6252 ( .A1(n9016), .A2(n4887), .ZN(n4886) );
  OAI211_X1 U6253 ( .C1(n9016), .C2(n4888), .A(n4886), .B(n8016), .ZN(P1_U3218) );
  INV_X1 U6254 ( .A(n6617), .ZN(n4902) );
  INV_X1 U6255 ( .A(n7970), .ZN(n4915) );
  NAND3_X1 U6256 ( .A1(n4919), .A2(n4908), .A3(n4918), .ZN(n4904) );
  NAND3_X1 U6257 ( .A1(n4919), .A2(n4918), .A3(n4911), .ZN(n4905) );
  NAND2_X1 U6258 ( .A1(n7904), .A2(n7903), .ZN(n7913) );
  INV_X1 U6259 ( .A(n7913), .ZN(n7916) );
  NAND3_X1 U6260 ( .A1(n4424), .A2(n4427), .A3(n5793), .ZN(n6200) );
  OAI21_X1 U6261 ( .B1(n9106), .B2(n4935), .A(n4933), .ZN(n4940) );
  NAND2_X1 U6262 ( .A1(n4945), .A2(n4944), .ZN(n8183) );
  INV_X1 U6263 ( .A(n6408), .ZN(n4947) );
  NAND2_X1 U6264 ( .A1(n4952), .A2(n4951), .ZN(n9055) );
  NAND3_X1 U6265 ( .A1(n7400), .A2(n4952), .A3(n4951), .ZN(n4950) );
  NAND2_X1 U6266 ( .A1(n7324), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4951) );
  NAND2_X1 U6267 ( .A1(n5765), .A2(n4958), .ZN(n4961) );
  NAND3_X1 U6268 ( .A1(n5585), .A2(n4498), .A3(n5584), .ZN(n4962) );
  OAI211_X1 U6269 ( .C1(n4962), .C2(n8272), .A(n8350), .B(n8353), .ZN(n8281)
         );
  NAND2_X1 U6270 ( .A1(n4962), .A2(n8272), .ZN(n8350) );
  NAND2_X1 U6271 ( .A1(n4964), .A2(n5193), .ZN(n7880) );
  NAND2_X1 U6272 ( .A1(n7889), .A2(n5185), .ZN(n4964) );
  OAI22_X1 U6273 ( .A1(n7880), .A2(n7881), .B1(n5210), .B2(n5209), .ZN(n6335)
         );
  NAND2_X1 U6274 ( .A1(n5425), .A2(n4447), .ZN(n4969) );
  NAND3_X1 U6275 ( .A1(n5116), .A2(n5117), .A3(n5237), .ZN(n4972) );
  OAI21_X1 U6276 ( .B1(n6970), .B2(n4978), .A(n4975), .ZN(n5410) );
  OAI21_X2 U6277 ( .B1(n5513), .B2(n4984), .A(n4982), .ZN(n8267) );
  NAND2_X1 U6278 ( .A1(n4988), .A2(n4986), .ZN(n6626) );
  INV_X1 U6279 ( .A(n6466), .ZN(n4990) );
  INV_X1 U6280 ( .A(n5534), .ZN(n5099) );
  MUX2_X2 U6281 ( .A(n7640), .B(n7639), .S(n7638), .Z(n7649) );
  INV_X1 U6282 ( .A(n4423), .ZN(n5662) );
  NOR2_X1 U6283 ( .A1(n4997), .A2(n5668), .ZN(n5672) );
  OR2_X1 U6284 ( .A1(n9763), .A2(n7709), .ZN(n9820) );
  NAND2_X1 U6285 ( .A1(n4436), .A2(n7672), .ZN(n7678) );
  INV_X1 U6286 ( .A(n9730), .ZN(n7051) );
  AND2_X1 U6287 ( .A1(n5062), .A2(n5061), .ZN(n4992) );
  NAND2_X1 U6288 ( .A1(n6040), .A2(n6031), .ZN(n9698) );
  AND2_X1 U6289 ( .A1(n5040), .A2(n5039), .ZN(n4993) );
  OR2_X1 U6290 ( .A1(n6859), .A2(n9045), .ZN(n4994) );
  INV_X1 U6291 ( .A(n9745), .ZN(n9749) );
  AND2_X1 U6292 ( .A1(n7500), .A2(n6374), .ZN(n7476) );
  AND2_X1 U6293 ( .A1(n5098), .A2(SI_21_), .ZN(n4995) );
  AND2_X1 U6294 ( .A1(n5579), .A2(n8247), .ZN(n4996) );
  AND2_X1 U6295 ( .A1(n7863), .A2(n7682), .ZN(n8620) );
  INV_X1 U6296 ( .A(n7542), .ZN(n6711) );
  AND2_X1 U6297 ( .A1(n7866), .A2(n7865), .ZN(n4998) );
  AND2_X1 U6298 ( .A1(n8638), .A2(n7807), .ZN(n4999) );
  INV_X1 U6299 ( .A(n7857), .ZN(n7677) );
  INV_X1 U6300 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5119) );
  NOR2_X1 U6301 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n5122) );
  INV_X1 U6302 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10027) );
  OR2_X1 U6303 ( .A1(n5418), .A2(n7179), .ZN(n5441) );
  NAND2_X1 U6304 ( .A1(n5675), .A2(n5674), .ZN(n5676) );
  INV_X1 U6305 ( .A(n7270), .ZN(n7250) );
  INV_X1 U6306 ( .A(n7322), .ZN(n7246) );
  INV_X1 U6307 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6563) );
  INV_X1 U6308 ( .A(n7476), .ZN(n6345) );
  INV_X1 U6309 ( .A(n5483), .ZN(n5085) );
  INV_X1 U6310 ( .A(SI_13_), .ZN(n10011) );
  INV_X1 U6311 ( .A(SI_8_), .ZN(n9949) );
  INV_X1 U6312 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5284) );
  OR2_X1 U6313 ( .A1(n5302), .A2(n10027), .ZN(n5343) );
  INV_X1 U6314 ( .A(n6443), .ZN(n5245) );
  OR2_X1 U6315 ( .A1(n5599), .A2(n8276), .ZN(n5620) );
  AND2_X1 U6316 ( .A1(n7786), .A2(n7787), .ZN(n7698) );
  OR2_X1 U6317 ( .A1(n9723), .A2(n7062), .ZN(n9724) );
  AOI21_X1 U6318 ( .B1(n9752), .B2(n9758), .A(n9759), .ZN(n6830) );
  INV_X1 U6319 ( .A(n5414), .ZN(n5415) );
  INV_X1 U6320 ( .A(n7993), .ZN(n7994) );
  OR3_X1 U6321 ( .A1(n7432), .A2(n7431), .A3(n7430), .ZN(n7453) );
  NAND2_X1 U6322 ( .A1(n7250), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7432) );
  NAND2_X1 U6323 ( .A1(n7249), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7358) );
  NAND2_X1 U6324 ( .A1(n7247), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n7292) );
  NAND2_X1 U6325 ( .A1(n6379), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6564) );
  INV_X1 U6326 ( .A(n9194), .ZN(n9189) );
  NAND2_X1 U6327 ( .A1(n7246), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7331) );
  OR2_X1 U6328 ( .A1(n7040), .A2(n7386), .ZN(n7028) );
  AND2_X1 U6329 ( .A1(n5821), .A2(n5864), .ZN(n5949) );
  OAI21_X2 U6330 ( .B1(n5608), .B2(n5607), .A(n5606), .ZN(n5614) );
  INV_X1 U6331 ( .A(n5546), .ZN(n5104) );
  OR2_X1 U6332 ( .A1(n5285), .A2(n5284), .ZN(n5302) );
  OR2_X1 U6333 ( .A1(n5642), .A2(n10144), .ZN(n5658) );
  NAND2_X1 U6334 ( .A1(n8246), .A2(n4996), .ZN(n5585) );
  INV_X1 U6335 ( .A(n8293), .ZN(n5480) );
  INV_X1 U6336 ( .A(n8379), .ZN(n8561) );
  OR2_X1 U6337 ( .A1(n5521), .A2(n10059), .ZN(n5553) );
  INV_X1 U6338 ( .A(n8652), .ZN(n8624) );
  INV_X1 U6339 ( .A(n6513), .ZN(n6143) );
  NAND2_X1 U6340 ( .A1(n7839), .A2(n7837), .ZN(n8529) );
  INV_X1 U6341 ( .A(n8808), .ZN(n8587) );
  OR2_X1 U6342 ( .A1(n7113), .A2(n7692), .ZN(n7125) );
  INV_X1 U6343 ( .A(n8731), .ZN(n9732) );
  INV_X1 U6344 ( .A(n7687), .ZN(n6320) );
  INV_X1 U6345 ( .A(n7054), .ZN(n9802) );
  INV_X1 U6346 ( .A(n9810), .ZN(n9815) );
  NAND2_X1 U6347 ( .A1(n5699), .A2(n5698), .ZN(n5701) );
  INV_X1 U6348 ( .A(n9041), .ZN(n9097) );
  OR2_X1 U6349 ( .A1(n7980), .A2(n7979), .ZN(n7981) );
  INV_X1 U6350 ( .A(n9029), .ZN(n9010) );
  AND2_X1 U6351 ( .A1(n7270), .A2(n7269), .ZN(n9125) );
  OR2_X1 U6352 ( .A1(n7331), .A2(n7330), .ZN(n7333) );
  AND2_X1 U6353 ( .A1(n6032), .A2(n7638), .ZN(n6127) );
  OR2_X1 U6354 ( .A1(n9337), .A2(n9118), .ZN(n8186) );
  INV_X1 U6355 ( .A(n9162), .ZN(n9191) );
  INV_X1 U6356 ( .A(n9239), .ZN(n9271) );
  NAND2_X1 U6357 ( .A1(n6652), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6695) );
  AND2_X1 U6358 ( .A1(n7388), .A2(n7540), .ZN(n7481) );
  OR2_X1 U6359 ( .A1(n6034), .A2(n7638), .ZN(n9692) );
  AND2_X1 U6360 ( .A1(n5658), .A2(n5643), .ZN(n8510) );
  OR2_X1 U6361 ( .A1(n8278), .A2(n9732), .ZN(n8369) );
  INV_X1 U6362 ( .A(n8368), .ZN(n8345) );
  NAND2_X1 U6363 ( .A1(n5705), .A2(n9743), .ZN(n8374) );
  AND4_X1 U6364 ( .A1(n5558), .A2(n5557), .A3(n5556), .A4(n5555), .ZN(n8248)
         );
  AND4_X1 U6365 ( .A1(n5440), .A2(n5439), .A3(n5438), .A4(n5437), .ZN(n8666)
         );
  INV_X1 U6366 ( .A(n9883), .ZN(n9433) );
  INV_X1 U6367 ( .A(n8474), .ZN(n9877) );
  INV_X1 U6368 ( .A(n9734), .ZN(n8729) );
  INV_X1 U6369 ( .A(n8620), .ZN(n9737) );
  INV_X1 U6370 ( .A(n9743), .ZN(n8752) );
  AND2_X1 U6371 ( .A1(n5685), .A2(n5684), .ZN(n6289) );
  OR2_X1 U6372 ( .A1(n9763), .A2(n7868), .ZN(n9810) );
  AND2_X1 U6373 ( .A1(n8655), .A2(n8654), .ZN(n8831) );
  INV_X1 U6374 ( .A(n9822), .ZN(n9764) );
  INV_X1 U6375 ( .A(n6289), .ZN(n6831) );
  AND2_X1 U6376 ( .A1(n5683), .A2(n5696), .ZN(n9752) );
  AND2_X1 U6377 ( .A1(n5673), .A2(n5680), .ZN(n7144) );
  INV_X1 U6378 ( .A(n9038), .ZN(n9015) );
  OR2_X1 U6379 ( .A1(n8011), .A2(n7434), .ZN(n7440) );
  OR2_X1 U6380 ( .A1(n9137), .A2(n7434), .ZN(n7365) );
  INV_X1 U6381 ( .A(n9629), .ZN(n9623) );
  INV_X1 U6382 ( .A(n9060), .ZN(n9641) );
  INV_X1 U6383 ( .A(n6127), .ZN(n5966) );
  OR2_X1 U6384 ( .A1(n8208), .A2(n8209), .ZN(n9174) );
  NOR2_X1 U6385 ( .A1(n7583), .A2(n8203), .ZN(n9226) );
  NAND2_X1 U6386 ( .A1(n9697), .A2(n5836), .ZN(n9258) );
  OR2_X1 U6387 ( .A1(n6034), .A2(n5955), .ZN(n9691) );
  AND2_X1 U6388 ( .A1(n6574), .A2(n6409), .ZN(n9396) );
  AND3_X1 U6389 ( .A1(n6028), .A2(n6027), .A3(n6026), .ZN(n6040) );
  INV_X1 U6390 ( .A(n7641), .ZN(n6029) );
  INV_X1 U6391 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5750) );
  AND2_X1 U6392 ( .A1(n5902), .A2(n6023), .ZN(n6687) );
  INV_X1 U6393 ( .A(n9760), .ZN(n5752) );
  NAND2_X1 U6394 ( .A1(n5720), .A2(n5709), .ZN(n8376) );
  OR2_X1 U6395 ( .A1(n5603), .A2(n5602), .ZN(n8379) );
  INV_X2 U6396 ( .A(P2_U3966), .ZN(n8392) );
  NAND2_X1 U6397 ( .A1(n6526), .A2(n5721), .ZN(n9883) );
  OR2_X1 U6398 ( .A1(n9710), .A2(n5721), .ZN(n8474) );
  AND2_X1 U6399 ( .A1(n6146), .A2(n6145), .ZN(n8479) );
  INV_X1 U6400 ( .A(n9749), .ZN(n8656) );
  INV_X1 U6401 ( .A(n9749), .ZN(n8754) );
  AND2_X1 U6402 ( .A1(n6833), .A2(n9743), .ZN(n9745) );
  NAND2_X1 U6403 ( .A1(n9749), .A2(n6835), .ZN(n8727) );
  INV_X1 U6404 ( .A(n9839), .ZN(n9837) );
  INV_X1 U6405 ( .A(n9826), .ZN(n9824) );
  INV_X1 U6406 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10081) );
  OR2_X1 U6407 ( .A1(n6056), .A2(n7643), .ZN(n9009) );
  INV_X1 U6408 ( .A(n9036), .ZN(n9024) );
  NAND2_X1 U6409 ( .A1(n7440), .A2(n7439), .ZN(n9041) );
  NAND2_X1 U6410 ( .A1(n7276), .A2(n7275), .ZN(n9118) );
  OR2_X1 U6411 ( .A1(n7317), .A2(n7316), .ZN(n9239) );
  OR2_X1 U6412 ( .A1(P1_U3083), .A2(n5878), .ZN(n9627) );
  OR2_X1 U6413 ( .A1(n4419), .A2(n6369), .ZN(n9308) );
  NAND2_X1 U6414 ( .A1(n6040), .A2(n6039), .ZN(n9707) );
  INV_X1 U6415 ( .A(n9664), .ZN(n9663) );
  INV_X1 U6416 ( .A(n5807), .ZN(n7630) );
  INV_X1 U6417 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10026) );
  INV_X1 U6418 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5972) );
  NOR2_X1 U6419 ( .A1(n10211), .A2(n10210), .ZN(n10209) );
  NOR2_X1 U6420 ( .A1(n9868), .A2(n9867), .ZN(n9866) );
  NOR2_X2 U6421 ( .A1(n6509), .A2(n5752), .ZN(P2_U3966) );
  MUX2_X1 U6422 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n7220), .Z(n5175) );
  NAND2_X1 U6423 ( .A1(n5176), .A2(n5175), .ZN(n5006) );
  INV_X1 U6424 ( .A(n5003), .ZN(n5004) );
  NAND2_X1 U6425 ( .A1(n5004), .A2(SI_1_), .ZN(n5005) );
  NAND2_X1 U6426 ( .A1(n5006), .A2(n5005), .ZN(n5205) );
  MUX2_X1 U6427 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n7220), .Z(n5008) );
  INV_X1 U6428 ( .A(SI_2_), .ZN(n5007) );
  XNOR2_X1 U6429 ( .A(n5008), .B(n5007), .ZN(n5204) );
  NAND2_X1 U6430 ( .A1(n5008), .A2(SI_2_), .ZN(n5009) );
  INV_X1 U6431 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5861) );
  INV_X1 U6432 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5011) );
  MUX2_X1 U6433 ( .A(n5861), .B(n5011), .S(n5844), .Z(n5012) );
  XNOR2_X1 U6434 ( .A(n5012), .B(SI_3_), .ZN(n5220) );
  INV_X1 U6435 ( .A(n5012), .ZN(n5013) );
  NAND2_X1 U6436 ( .A1(n5013), .A2(SI_3_), .ZN(n5014) );
  MUX2_X1 U6437 ( .A(n5860), .B(n10108), .S(n7220), .Z(n5015) );
  XNOR2_X1 U6438 ( .A(n5015), .B(SI_4_), .ZN(n5239) );
  INV_X1 U6439 ( .A(n5015), .ZN(n5016) );
  NAND2_X1 U6440 ( .A1(n5016), .A2(SI_4_), .ZN(n5017) );
  INV_X1 U6441 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5018) );
  MUX2_X1 U6442 ( .A(n10109), .B(n5018), .S(n5844), .Z(n5019) );
  XNOR2_X1 U6443 ( .A(n5019), .B(SI_5_), .ZN(n5257) );
  NAND2_X1 U6444 ( .A1(n5258), .A2(n5257), .ZN(n5022) );
  INV_X1 U6445 ( .A(n5019), .ZN(n5020) );
  NAND2_X1 U6446 ( .A1(n5020), .A2(SI_5_), .ZN(n5021) );
  MUX2_X1 U6447 ( .A(n5862), .B(n5858), .S(n5844), .Z(n5023) );
  NAND2_X1 U6448 ( .A1(n5275), .A2(n5274), .ZN(n5026) );
  INV_X1 U6449 ( .A(n5023), .ZN(n5024) );
  NAND2_X1 U6450 ( .A1(n5024), .A2(SI_6_), .ZN(n5025) );
  MUX2_X1 U6451 ( .A(n5869), .B(n5027), .S(n7220), .Z(n5028) );
  NAND2_X1 U6452 ( .A1(n5294), .A2(n5293), .ZN(n5031) );
  INV_X1 U6453 ( .A(n5028), .ZN(n5029) );
  NAND2_X1 U6454 ( .A1(n5029), .A2(SI_7_), .ZN(n5030) );
  NAND2_X2 U6455 ( .A1(n5031), .A2(n5030), .ZN(n5313) );
  MUX2_X1 U6456 ( .A(n5877), .B(n5876), .S(n7220), .Z(n5032) );
  INV_X1 U6457 ( .A(n5032), .ZN(n5033) );
  NAND2_X1 U6458 ( .A1(n5033), .A2(SI_8_), .ZN(n5034) );
  NAND2_X1 U6459 ( .A1(n5035), .A2(n5034), .ZN(n5311) );
  MUX2_X1 U6460 ( .A(n5888), .B(n10204), .S(n7220), .Z(n5037) );
  INV_X1 U6461 ( .A(SI_9_), .ZN(n5036) );
  INV_X1 U6462 ( .A(n5037), .ZN(n5038) );
  NAND2_X1 U6463 ( .A1(n5038), .A2(SI_9_), .ZN(n5039) );
  MUX2_X1 U6464 ( .A(n10174), .B(n5041), .S(n7220), .Z(n5043) );
  INV_X1 U6465 ( .A(SI_10_), .ZN(n5042) );
  NAND2_X1 U6466 ( .A1(n5043), .A2(n5042), .ZN(n5046) );
  INV_X1 U6467 ( .A(n5043), .ZN(n5044) );
  NAND2_X1 U6468 ( .A1(n5044), .A2(SI_10_), .ZN(n5045) );
  MUX2_X1 U6469 ( .A(n9996), .B(n5972), .S(n7220), .Z(n5048) );
  INV_X1 U6470 ( .A(n5048), .ZN(n5049) );
  NAND2_X1 U6471 ( .A1(n5049), .A2(SI_11_), .ZN(n5050) );
  INV_X1 U6472 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5052) );
  MUX2_X1 U6473 ( .A(n10001), .B(n5052), .S(n5844), .Z(n5054) );
  INV_X1 U6474 ( .A(n5054), .ZN(n5055) );
  NAND2_X1 U6475 ( .A1(n5055), .A2(SI_12_), .ZN(n5056) );
  NAND2_X1 U6476 ( .A1(n5057), .A2(n5056), .ZN(n5353) );
  INV_X1 U6477 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5058) );
  MUX2_X1 U6478 ( .A(n10081), .B(n5058), .S(n5844), .Z(n5059) );
  NAND2_X1 U6479 ( .A1(n5059), .A2(n10011), .ZN(n5062) );
  INV_X1 U6480 ( .A(n5059), .ZN(n5060) );
  NAND2_X1 U6481 ( .A1(n5060), .A2(SI_13_), .ZN(n5061) );
  MUX2_X1 U6482 ( .A(n10140), .B(n6141), .S(n5844), .Z(n5064) );
  XNOR2_X1 U6483 ( .A(n5064), .B(SI_14_), .ZN(n5412) );
  INV_X1 U6484 ( .A(n5064), .ZN(n5065) );
  MUX2_X1 U6485 ( .A(n6204), .B(n6202), .S(n7220), .Z(n5069) );
  INV_X1 U6486 ( .A(SI_15_), .ZN(n5068) );
  INV_X1 U6487 ( .A(n5069), .ZN(n5070) );
  NAND2_X1 U6488 ( .A1(n5070), .A2(SI_15_), .ZN(n5071) );
  INV_X1 U6489 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5073) );
  MUX2_X1 U6490 ( .A(n5073), .B(n10026), .S(n7220), .Z(n5075) );
  INV_X1 U6491 ( .A(SI_16_), .ZN(n5074) );
  NAND2_X1 U6492 ( .A1(n5075), .A2(n5074), .ZN(n5078) );
  INV_X1 U6493 ( .A(n5075), .ZN(n5076) );
  NAND2_X1 U6494 ( .A1(n5076), .A2(SI_16_), .ZN(n5077) );
  INV_X1 U6495 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5080) );
  MUX2_X1 U6496 ( .A(n10084), .B(n5080), .S(n5844), .Z(n5081) );
  XNOR2_X1 U6497 ( .A(n5081), .B(SI_17_), .ZN(n5462) );
  INV_X1 U6498 ( .A(n5081), .ZN(n5082) );
  NAND2_X1 U6499 ( .A1(n5082), .A2(SI_17_), .ZN(n5083) );
  OAI21_X2 U6500 ( .B1(n5463), .B2(n5084), .A(n5083), .ZN(n5484) );
  MUX2_X1 U6501 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5844), .Z(n5086) );
  XNOR2_X1 U6502 ( .A(n5086), .B(SI_18_), .ZN(n5483) );
  NAND2_X1 U6503 ( .A1(n5086), .A2(SI_18_), .ZN(n5087) );
  INV_X1 U6504 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6554) );
  INV_X1 U6505 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6552) );
  MUX2_X1 U6506 ( .A(n6554), .B(n6552), .S(n7220), .Z(n5089) );
  INV_X1 U6507 ( .A(SI_19_), .ZN(n10168) );
  NAND2_X1 U6508 ( .A1(n5089), .A2(n10168), .ZN(n5092) );
  INV_X1 U6509 ( .A(n5089), .ZN(n5090) );
  NAND2_X1 U6510 ( .A1(n5090), .A2(SI_19_), .ZN(n5091) );
  NAND2_X1 U6511 ( .A1(n5092), .A2(n5091), .ZN(n5501) );
  INV_X1 U6512 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6640) );
  INV_X1 U6513 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6679) );
  MUX2_X1 U6514 ( .A(n6640), .B(n6679), .S(n7220), .Z(n5093) );
  INV_X1 U6515 ( .A(SI_20_), .ZN(n9971) );
  NAND2_X1 U6516 ( .A1(n5093), .A2(n9971), .ZN(n5096) );
  INV_X1 U6517 ( .A(n5093), .ZN(n5094) );
  NAND2_X1 U6518 ( .A1(n5094), .A2(SI_20_), .ZN(n5095) );
  INV_X1 U6519 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6681) );
  MUX2_X1 U6520 ( .A(n6681), .B(n10056), .S(n7220), .Z(n5097) );
  XNOR2_X1 U6521 ( .A(n5097), .B(SI_21_), .ZN(n5533) );
  INV_X1 U6522 ( .A(n5097), .ZN(n5098) );
  INV_X1 U6523 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7887) );
  INV_X1 U6524 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n6847) );
  MUX2_X1 U6525 ( .A(n7887), .B(n6847), .S(n5844), .Z(n5101) );
  INV_X1 U6526 ( .A(SI_22_), .ZN(n5100) );
  NAND2_X1 U6527 ( .A1(n5101), .A2(n5100), .ZN(n5105) );
  INV_X1 U6528 ( .A(n5101), .ZN(n5102) );
  NAND2_X1 U6529 ( .A1(n5102), .A2(SI_22_), .ZN(n5103) );
  NAND2_X1 U6530 ( .A1(n5105), .A2(n5103), .ZN(n5546) );
  INV_X1 U6531 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5107) );
  INV_X1 U6532 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5106) );
  MUX2_X1 U6533 ( .A(n5107), .B(n5106), .S(n5844), .Z(n5109) );
  INV_X1 U6534 ( .A(SI_23_), .ZN(n5108) );
  NAND2_X1 U6535 ( .A1(n5109), .A2(n5108), .ZN(n5114) );
  INV_X1 U6536 ( .A(n5109), .ZN(n5110) );
  NAND2_X1 U6537 ( .A1(n5110), .A2(SI_23_), .ZN(n5111) );
  NAND2_X1 U6538 ( .A1(n5114), .A2(n5111), .ZN(n5563) );
  INV_X1 U6539 ( .A(n5563), .ZN(n5112) );
  INV_X1 U6540 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7068) );
  INV_X1 U6541 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10167) );
  MUX2_X1 U6542 ( .A(n7068), .B(n10167), .S(n4420), .Z(n5587) );
  XNOR2_X1 U6543 ( .A(n5587), .B(SI_24_), .ZN(n5586) );
  XNOR2_X1 U6544 ( .A(n5591), .B(n5586), .ZN(n7354) );
  NOR2_X2 U6545 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5201) );
  NAND2_X1 U6546 ( .A1(n5201), .A2(n5115), .ZN(n5236) );
  INV_X1 U6547 ( .A(n5133), .ZN(n5121) );
  NOR2_X1 U6548 ( .A1(n5121), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n5124) );
  INV_X1 U6549 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5126) );
  OR2_X1 U6550 ( .A1(n5148), .A2(n5126), .ZN(n5127) );
  NAND2_X1 U6551 ( .A1(n4439), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5128) );
  INV_X1 U6552 ( .A(n5148), .ZN(n5129) );
  NAND2_X1 U6553 ( .A1(n7354), .A2(n7673), .ZN(n5132) );
  NAND2_X1 U6554 ( .A1(n7665), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5131) );
  NAND2_X1 U6555 ( .A1(n5134), .A2(n5133), .ZN(n5141) );
  XNOR2_X2 U6556 ( .A(n5675), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5140) );
  INV_X1 U6557 ( .A(n5134), .ZN(n5135) );
  INV_X1 U6558 ( .A(n5138), .ZN(n5136) );
  NAND2_X1 U6559 ( .A1(n5136), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n5139) );
  INV_X1 U6560 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U6561 ( .A1(n5140), .A2(n7711), .ZN(n7863) );
  NAND2_X1 U6562 ( .A1(n5141), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5142) );
  NAND3_X1 U6563 ( .A1(n7863), .A2(n9763), .A3(n6680), .ZN(n5146) );
  NAND2_X1 U6564 ( .A1(n5143), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5145) );
  INV_X1 U6565 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U6566 ( .A1(n7860), .A2(n7728), .ZN(n6834) );
  XNOR2_X1 U6567 ( .A(n8796), .B(n5200), .ZN(n5582) );
  INV_X1 U6568 ( .A(n5582), .ZN(n8302) );
  INV_X1 U6569 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5150) );
  INV_X1 U6570 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8880) );
  INV_X1 U6571 ( .A(n5248), .ZN(n5467) );
  NAND2_X1 U6572 ( .A1(n4409), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U6573 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5250) );
  INV_X1 U6574 ( .A(n5250), .ZN(n5154) );
  NAND2_X1 U6575 ( .A1(n5154), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5264) );
  INV_X1 U6576 ( .A(n5264), .ZN(n5155) );
  NAND2_X1 U6577 ( .A1(n5155), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5285) );
  INV_X1 U6578 ( .A(n5343), .ZN(n5157) );
  AND2_X1 U6579 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n5156) );
  NAND2_X1 U6580 ( .A1(n5157), .A2(n5156), .ZN(n5390) );
  INV_X1 U6581 ( .A(n5390), .ZN(n5158) );
  NAND2_X1 U6582 ( .A1(n5158), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5392) );
  INV_X1 U6583 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5359) );
  INV_X1 U6584 ( .A(n5371), .ZN(n5159) );
  NAND2_X1 U6585 ( .A1(n5159), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5418) );
  INV_X1 U6586 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7179) );
  INV_X1 U6587 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8366) );
  INV_X1 U6588 ( .A(n5469), .ZN(n5161) );
  AND2_X1 U6589 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n5160) );
  NAND2_X1 U6590 ( .A1(n5161), .A2(n5160), .ZN(n5489) );
  INV_X1 U6591 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8343) );
  INV_X1 U6592 ( .A(n5506), .ZN(n5162) );
  NAND2_X1 U6593 ( .A1(n5162), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5521) );
  INV_X1 U6594 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10059) );
  NAND2_X1 U6595 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n5163) );
  INV_X1 U6596 ( .A(n5572), .ZN(n5164) );
  NAND2_X1 U6597 ( .A1(n5164), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5574) );
  INV_X1 U6598 ( .A(n5574), .ZN(n5165) );
  NAND2_X1 U6599 ( .A1(n5165), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5599) );
  INV_X1 U6600 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6601 ( .A1(n5574), .A2(n5166), .ZN(n5167) );
  AND2_X1 U6602 ( .A1(n5599), .A2(n5167), .ZN(n8557) );
  NAND2_X1 U6603 ( .A1(n5644), .A2(n8557), .ZN(n5171) );
  NAND2_X1 U6604 ( .A1(n4423), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6605 ( .A1(n5393), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5169) );
  NAND4_X1 U6606 ( .A1(n5172), .A2(n5171), .A3(n5170), .A4(n5169), .ZN(n8570)
         );
  INV_X1 U6607 ( .A(n8570), .ZN(n8274) );
  NAND2_X1 U6608 ( .A1(n7860), .A2(n8546), .ZN(n5714) );
  NOR2_X1 U6609 ( .A1(n8274), .A2(n6450), .ZN(n5583) );
  INV_X1 U6610 ( .A(n5583), .ZN(n8306) );
  INV_X1 U6611 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U6612 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5173) );
  XNOR2_X1 U6613 ( .A(n5174), .B(n5173), .ZN(n9427) );
  XNOR2_X1 U6614 ( .A(n5176), .B(n5175), .ZN(n5853) );
  INV_X1 U6615 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5845) );
  XNOR2_X1 U6616 ( .A(n6270), .B(n5200), .ZN(n5182) );
  NAND2_X1 U6617 ( .A1(n5248), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5180) );
  NAND2_X1 U6618 ( .A1(n5211), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5179) );
  NAND2_X1 U6619 ( .A1(n4410), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5178) );
  INV_X1 U6620 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6507) );
  NOR2_X1 U6621 ( .A1(n6271), .A2(n6450), .ZN(n5181) );
  NAND2_X1 U6622 ( .A1(n5182), .A2(n5181), .ZN(n5185) );
  INV_X1 U6623 ( .A(n5181), .ZN(n5184) );
  INV_X1 U6624 ( .A(n5182), .ZN(n5183) );
  NAND2_X1 U6625 ( .A1(n5184), .A2(n5183), .ZN(n5193) );
  NAND2_X1 U6626 ( .A1(n5212), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6627 ( .A1(n5211), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5186) );
  AND2_X1 U6628 ( .A1(n5187), .A2(n5186), .ZN(n5190) );
  NAND2_X1 U6629 ( .A1(n4409), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5188) );
  NAND2_X1 U6630 ( .A1(n6275), .A2(n7683), .ZN(n5192) );
  NAND2_X1 U6631 ( .A1(n7229), .A2(SI_0_), .ZN(n5191) );
  XNOR2_X1 U6632 ( .A(n5191), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8886) );
  MUX2_X1 U6633 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8886), .S(n6513), .Z(n6869) );
  MUX2_X1 U6634 ( .A(n5569), .B(n5192), .S(n6869), .Z(n7889) );
  NAND2_X1 U6635 ( .A1(n5248), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U6636 ( .A1(n5211), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5198) );
  INV_X1 U6637 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6638 ( .A1(n4410), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5196) );
  OR2_X1 U6639 ( .A1(n6424), .A2(n6450), .ZN(n5209) );
  OR2_X1 U6640 ( .A1(n5201), .A2(n5126), .ZN(n5203) );
  INV_X1 U6641 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5202) );
  NAND2_X1 U6642 ( .A1(n5203), .A2(n5202), .ZN(n5217) );
  OAI21_X1 U6643 ( .B1(n5203), .B2(n5202), .A(n5217), .ZN(n9444) );
  XNOR2_X1 U6644 ( .A(n5205), .B(n5204), .ZN(n5859) );
  OR2_X1 U6645 ( .A1(n5222), .A2(n5859), .ZN(n5207) );
  INV_X1 U6646 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10154) );
  OR2_X1 U6647 ( .A1(n5223), .A2(n10154), .ZN(n5206) );
  XNOR2_X1 U6648 ( .A(n5208), .B(n4411), .ZN(n5210) );
  XNOR2_X1 U6649 ( .A(n5209), .B(n5210), .ZN(n7881) );
  NAND2_X1 U6650 ( .A1(n5248), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5216) );
  INV_X1 U6651 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10012) );
  NAND2_X1 U6652 ( .A1(n5211), .A2(n10012), .ZN(n5215) );
  NAND2_X1 U6653 ( .A1(n4422), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6654 ( .A1(n4418), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5213) );
  OR2_X1 U6655 ( .A1(n6487), .A2(n6450), .ZN(n5226) );
  NAND2_X1 U6656 ( .A1(n5217), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5219) );
  INV_X1 U6657 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5218) );
  XNOR2_X1 U6658 ( .A(n5219), .B(n5218), .ZN(n6533) );
  XNOR2_X1 U6659 ( .A(n5221), .B(n5220), .ZN(n6089) );
  OR2_X1 U6660 ( .A1(n5222), .A2(n6089), .ZN(n5225) );
  OR2_X1 U6661 ( .A1(n5223), .A2(n5861), .ZN(n5224) );
  OAI211_X1 U6662 ( .C1(n6513), .C2(n6533), .A(n5225), .B(n5224), .ZN(n6924)
         );
  XNOR2_X1 U6663 ( .A(n4421), .B(n5569), .ZN(n5227) );
  XNOR2_X1 U6664 ( .A(n5226), .B(n5227), .ZN(n6334) );
  NAND2_X1 U6665 ( .A1(n6335), .A2(n6334), .ZN(n5230) );
  INV_X1 U6666 ( .A(n5226), .ZN(n5228) );
  NAND2_X1 U6667 ( .A1(n5228), .A2(n5227), .ZN(n5229) );
  NAND2_X1 U6668 ( .A1(n5230), .A2(n5229), .ZN(n6444) );
  INV_X1 U6669 ( .A(n6444), .ZN(n5246) );
  NAND2_X1 U6670 ( .A1(n5248), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5235) );
  INV_X1 U6671 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8400) );
  NAND2_X1 U6672 ( .A1(n10012), .A2(n8400), .ZN(n5231) );
  AND2_X1 U6673 ( .A1(n5231), .A2(n5250), .ZN(n6839) );
  NAND2_X1 U6674 ( .A1(n5644), .A2(n6839), .ZN(n5234) );
  NAND2_X1 U6675 ( .A1(n4422), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U6676 ( .A1(n5393), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5232) );
  OR2_X1 U6677 ( .A1(n6872), .A2(n6450), .ZN(n5244) );
  NAND2_X1 U6678 ( .A1(n5236), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5238) );
  INV_X1 U6679 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5237) );
  XNOR2_X1 U6680 ( .A(n5238), .B(n5237), .ZN(n8402) );
  XNOR2_X1 U6681 ( .A(n5240), .B(n5239), .ZN(n6102) );
  OR2_X1 U6682 ( .A1(n5314), .A2(n6102), .ZN(n5242) );
  OR2_X1 U6683 ( .A1(n5223), .A2(n5860), .ZN(n5241) );
  OAI211_X1 U6684 ( .C1(n6513), .C2(n8402), .A(n5242), .B(n5241), .ZN(n6501)
         );
  XNOR2_X1 U6685 ( .A(n5208), .B(n6501), .ZN(n5243) );
  NAND2_X1 U6686 ( .A1(n5244), .A2(n5243), .ZN(n5247) );
  OAI21_X1 U6687 ( .B1(n5244), .B2(n5243), .A(n5247), .ZN(n6443) );
  NAND2_X1 U6688 ( .A1(n5248), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5255) );
  INV_X1 U6689 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6690 ( .A1(n5250), .A2(n5249), .ZN(n5251) );
  AND2_X1 U6691 ( .A1(n5264), .A2(n5251), .ZN(n6981) );
  NAND2_X1 U6692 ( .A1(n5644), .A2(n6981), .ZN(n5254) );
  NAND2_X1 U6693 ( .A1(n5393), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U6694 ( .A1(n4422), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5252) );
  OR2_X1 U6695 ( .A1(n6875), .A2(n6450), .ZN(n5259) );
  OR2_X1 U6696 ( .A1(n5256), .A2(n5126), .ZN(n5271) );
  XNOR2_X1 U6697 ( .A(n5271), .B(P2_IR_REG_5__SCAN_IN), .ZN(n8044) );
  INV_X1 U6698 ( .A(n8044), .ZN(n6548) );
  XNOR2_X1 U6699 ( .A(n5208), .B(n6987), .ZN(n5260) );
  XNOR2_X1 U6700 ( .A(n5259), .B(n5260), .ZN(n6466) );
  INV_X1 U6701 ( .A(n5259), .ZN(n5262) );
  INV_X1 U6702 ( .A(n5260), .ZN(n5261) );
  NAND2_X1 U6703 ( .A1(n5262), .A2(n5261), .ZN(n5263) );
  NAND2_X1 U6704 ( .A1(n5248), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5269) );
  INV_X1 U6705 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10063) );
  NAND2_X1 U6706 ( .A1(n5264), .A2(n10063), .ZN(n5265) );
  AND2_X1 U6707 ( .A1(n5285), .A2(n5265), .ZN(n8734) );
  NAND2_X1 U6708 ( .A1(n5644), .A2(n8734), .ZN(n5268) );
  NAND2_X1 U6709 ( .A1(n4422), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U6710 ( .A1(n5393), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5266) );
  NOR2_X1 U6711 ( .A1(n6878), .A2(n6450), .ZN(n5278) );
  INV_X1 U6712 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6713 ( .A1(n5271), .A2(n5270), .ZN(n5272) );
  NAND2_X1 U6714 ( .A1(n5272), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5273) );
  XNOR2_X1 U6715 ( .A(n5273), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8041) );
  INV_X1 U6716 ( .A(n8041), .ZN(n8111) );
  XNOR2_X1 U6717 ( .A(n5275), .B(n5274), .ZN(n6347) );
  OR2_X1 U6718 ( .A1(n5314), .A2(n6347), .ZN(n5277) );
  OR2_X1 U6719 ( .A1(n7674), .A2(n5862), .ZN(n5276) );
  OAI211_X1 U6720 ( .C1(n6513), .C2(n8111), .A(n5277), .B(n5276), .ZN(n9773)
         );
  XNOR2_X1 U6721 ( .A(n9773), .B(n5569), .ZN(n5279) );
  NAND2_X1 U6722 ( .A1(n5278), .A2(n5279), .ZN(n5282) );
  INV_X1 U6723 ( .A(n5278), .ZN(n5281) );
  INV_X1 U6724 ( .A(n5279), .ZN(n5280) );
  NAND2_X1 U6725 ( .A1(n5281), .A2(n5280), .ZN(n5283) );
  AND2_X1 U6726 ( .A1(n5282), .A2(n5283), .ZN(n6627) );
  NAND2_X1 U6727 ( .A1(n6626), .A2(n5283), .ZN(n6634) );
  NAND2_X1 U6728 ( .A1(n5248), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6729 ( .A1(n5285), .A2(n5284), .ZN(n5286) );
  AND2_X1 U6730 ( .A1(n5302), .A2(n5286), .ZN(n6883) );
  NAND2_X1 U6731 ( .A1(n5644), .A2(n6883), .ZN(n5289) );
  NAND2_X1 U6732 ( .A1(n5393), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5288) );
  NAND2_X1 U6733 ( .A1(n4422), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5287) );
  OR2_X1 U6734 ( .A1(n9735), .A2(n6450), .ZN(n5297) );
  NAND2_X1 U6735 ( .A1(n5291), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5292) );
  XNOR2_X1 U6736 ( .A(n5292), .B(P2_IR_REG_7__SCAN_IN), .ZN(n8039) );
  INV_X1 U6737 ( .A(n8039), .ZN(n9882) );
  XNOR2_X1 U6738 ( .A(n5294), .B(n5293), .ZN(n6354) );
  OR2_X1 U6739 ( .A1(n7674), .A2(n5869), .ZN(n5295) );
  XNOR2_X1 U6740 ( .A(n5208), .B(n6886), .ZN(n5298) );
  XNOR2_X1 U6741 ( .A(n5297), .B(n5298), .ZN(n6633) );
  INV_X1 U6742 ( .A(n5297), .ZN(n5300) );
  INV_X1 U6743 ( .A(n5298), .ZN(n5299) );
  NAND2_X1 U6744 ( .A1(n5300), .A2(n5299), .ZN(n5301) );
  NAND2_X1 U6745 ( .A1(n5302), .A2(n10027), .ZN(n5303) );
  NAND2_X1 U6746 ( .A1(n5343), .A2(n5303), .ZN(n9742) );
  INV_X1 U6747 ( .A(n9742), .ZN(n5304) );
  NAND2_X1 U6748 ( .A1(n5644), .A2(n5304), .ZN(n5308) );
  NAND2_X1 U6749 ( .A1(n5248), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U6750 ( .A1(n5393), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6751 ( .A1(n4423), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5305) );
  NAND4_X1 U6752 ( .A1(n5308), .A2(n5307), .A3(n5306), .A4(n5305), .ZN(n8387)
         );
  NAND2_X1 U6753 ( .A1(n8387), .A2(n7683), .ZN(n5319) );
  NAND2_X1 U6754 ( .A1(n5309), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5310) );
  XNOR2_X1 U6755 ( .A(n5310), .B(n4819), .ZN(n8099) );
  INV_X1 U6756 ( .A(n5311), .ZN(n5312) );
  XNOR2_X1 U6757 ( .A(n5313), .B(n5312), .ZN(n6557) );
  OR2_X1 U6758 ( .A1(n5314), .A2(n6557), .ZN(n5316) );
  OR2_X1 U6759 ( .A1(n7674), .A2(n5877), .ZN(n5315) );
  XNOR2_X1 U6760 ( .A(n7062), .B(n5200), .ZN(n5317) );
  XNOR2_X1 U6761 ( .A(n5319), .B(n5317), .ZN(n6772) );
  INV_X1 U6762 ( .A(n5317), .ZN(n5318) );
  NOR2_X1 U6763 ( .A1(n5319), .A2(n5318), .ZN(n5320) );
  AOI21_X1 U6764 ( .B1(n6773), .B2(n6772), .A(n5320), .ZN(n6970) );
  NAND2_X1 U6765 ( .A1(n5248), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5324) );
  XNOR2_X1 U6766 ( .A(n5343), .B(P2_REG3_REG_9__SCAN_IN), .ZN(n7083) );
  NAND2_X1 U6767 ( .A1(n5644), .A2(n7083), .ZN(n5323) );
  NAND2_X1 U6768 ( .A1(n5393), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6769 ( .A1(n4410), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5321) );
  NOR2_X1 U6770 ( .A1(n9733), .A2(n6450), .ZN(n5329) );
  OR2_X1 U6771 ( .A1(n5325), .A2(n5126), .ZN(n5337) );
  XNOR2_X1 U6772 ( .A(n5337), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8036) );
  AOI22_X1 U6773 ( .A1(n7665), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6143), .B2(
        n8036), .ZN(n5328) );
  XNOR2_X1 U6774 ( .A(n5326), .B(n4993), .ZN(n6645) );
  NAND2_X1 U6775 ( .A1(n6645), .A2(n7673), .ZN(n5327) );
  NAND2_X1 U6776 ( .A1(n5328), .A2(n5327), .ZN(n7080) );
  XNOR2_X1 U6777 ( .A(n7080), .B(n5569), .ZN(n5330) );
  NAND2_X1 U6778 ( .A1(n5329), .A2(n5330), .ZN(n5333) );
  INV_X1 U6779 ( .A(n5329), .ZN(n5332) );
  INV_X1 U6780 ( .A(n5330), .ZN(n5331) );
  NAND2_X1 U6781 ( .A1(n5332), .A2(n5331), .ZN(n5334) );
  AND2_X1 U6782 ( .A1(n5333), .A2(n5334), .ZN(n6969) );
  NAND2_X1 U6783 ( .A1(n6686), .A2(n7673), .ZN(n5340) );
  INV_X1 U6784 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6785 ( .A1(n5337), .A2(n5336), .ZN(n5338) );
  NAND2_X1 U6786 ( .A1(n5338), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5385) );
  XNOR2_X1 U6787 ( .A(n5385), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8033) );
  AOI22_X1 U6788 ( .A1(n7665), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6143), .B2(
        n8033), .ZN(n5339) );
  NAND2_X1 U6789 ( .A1(n5340), .A2(n5339), .ZN(n7054) );
  XNOR2_X1 U6790 ( .A(n7054), .B(n5208), .ZN(n5350) );
  NAND2_X1 U6791 ( .A1(n5248), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5348) );
  INV_X1 U6792 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5342) );
  INV_X1 U6793 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5341) );
  OAI21_X1 U6794 ( .B1(n5343), .B2(n5342), .A(n5341), .ZN(n5344) );
  AND2_X1 U6795 ( .A1(n5390), .A2(n5344), .ZN(n7137) );
  NAND2_X1 U6796 ( .A1(n5644), .A2(n7137), .ZN(n5347) );
  NAND2_X1 U6797 ( .A1(n5393), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6798 ( .A1(n4422), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5345) );
  OR2_X1 U6799 ( .A1(n7075), .A2(n6450), .ZN(n5349) );
  XNOR2_X1 U6800 ( .A(n5350), .B(n5349), .ZN(n6991) );
  INV_X1 U6801 ( .A(n5349), .ZN(n5352) );
  INV_X1 U6802 ( .A(n5350), .ZN(n5351) );
  NAND2_X1 U6803 ( .A1(n5352), .A2(n5351), .ZN(n7146) );
  XNOR2_X1 U6804 ( .A(n5354), .B(n5353), .ZN(n6778) );
  NAND2_X1 U6805 ( .A1(n6778), .A2(n7673), .ZN(n5358) );
  NAND2_X1 U6806 ( .A1(n5355), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5356) );
  XNOR2_X1 U6807 ( .A(n5356), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8122) );
  AOI22_X1 U6808 ( .A1(n7665), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6143), .B2(
        n8122), .ZN(n5357) );
  XNOR2_X1 U6809 ( .A(n9816), .B(n5208), .ZN(n5399) );
  NAND2_X1 U6810 ( .A1(n5248), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U6811 ( .A1(n5392), .A2(n5359), .ZN(n5360) );
  AND2_X1 U6812 ( .A1(n5371), .A2(n5360), .ZN(n7102) );
  NAND2_X1 U6813 ( .A1(n5644), .A2(n7102), .ZN(n5363) );
  NAND2_X1 U6814 ( .A1(n4423), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6815 ( .A1(n5393), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5361) );
  OR2_X1 U6816 ( .A1(n7163), .A2(n6450), .ZN(n5400) );
  NAND2_X1 U6817 ( .A1(n5399), .A2(n5400), .ZN(n7156) );
  XNOR2_X1 U6818 ( .A(n5365), .B(n4992), .ZN(n6929) );
  NAND2_X1 U6819 ( .A1(n6929), .A2(n7673), .ZN(n5369) );
  NAND2_X1 U6820 ( .A1(n5366), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5367) );
  XNOR2_X1 U6821 ( .A(n5367), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8123) );
  AOI22_X1 U6822 ( .A1(n7665), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6143), .B2(
        n8123), .ZN(n5368) );
  XNOR2_X1 U6823 ( .A(n8855), .B(n5569), .ZN(n5377) );
  NAND2_X1 U6824 ( .A1(n5248), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5376) );
  INV_X1 U6825 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6826 ( .A1(n5371), .A2(n5370), .ZN(n5372) );
  AND2_X1 U6827 ( .A1(n5418), .A2(n5372), .ZN(n7165) );
  NAND2_X1 U6828 ( .A1(n5644), .A2(n7165), .ZN(n5375) );
  NAND2_X1 U6829 ( .A1(n4423), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6830 ( .A1(n5393), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5373) );
  NOR2_X1 U6831 ( .A1(n7176), .A2(n6450), .ZN(n5378) );
  NAND2_X1 U6832 ( .A1(n5377), .A2(n5378), .ZN(n5411) );
  INV_X1 U6833 ( .A(n5377), .ZN(n5380) );
  INV_X1 U6834 ( .A(n5378), .ZN(n5379) );
  NAND2_X1 U6835 ( .A1(n5380), .A2(n5379), .ZN(n5381) );
  XNOR2_X1 U6836 ( .A(n5383), .B(n5382), .ZN(n6691) );
  NAND2_X1 U6837 ( .A1(n6691), .A2(n7673), .ZN(n5389) );
  INV_X1 U6838 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6839 ( .A1(n5385), .A2(n5384), .ZN(n5386) );
  NAND2_X1 U6840 ( .A1(n5386), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5387) );
  XNOR2_X1 U6841 ( .A(n5387), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8167) );
  AOI22_X1 U6842 ( .A1(n7665), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6143), .B2(
        n8167), .ZN(n5388) );
  NAND2_X1 U6843 ( .A1(n5389), .A2(n5388), .ZN(n8334) );
  XNOR2_X1 U6844 ( .A(n8334), .B(n5208), .ZN(n5405) );
  INV_X1 U6845 ( .A(n5405), .ZN(n5398) );
  NAND2_X1 U6846 ( .A1(n5248), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5397) );
  INV_X1 U6847 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9953) );
  NAND2_X1 U6848 ( .A1(n5390), .A2(n9953), .ZN(n5391) );
  AND2_X1 U6849 ( .A1(n5392), .A2(n5391), .ZN(n7061) );
  NAND2_X1 U6850 ( .A1(n5644), .A2(n7061), .ZN(n5396) );
  NAND2_X1 U6851 ( .A1(n5393), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U6852 ( .A1(n4423), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5394) );
  NOR2_X1 U6853 ( .A1(n7130), .A2(n6450), .ZN(n5404) );
  NAND2_X1 U6854 ( .A1(n5398), .A2(n5404), .ZN(n7148) );
  INV_X1 U6855 ( .A(n5399), .ZN(n5402) );
  INV_X1 U6856 ( .A(n5400), .ZN(n5401) );
  NAND2_X1 U6857 ( .A1(n5402), .A2(n5401), .ZN(n7158) );
  INV_X1 U6858 ( .A(n5403), .ZN(n5408) );
  XNOR2_X1 U6859 ( .A(n5405), .B(n5404), .ZN(n8330) );
  AND2_X1 U6860 ( .A1(n8330), .A2(n5406), .ZN(n5407) );
  OR2_X1 U6861 ( .A1(n5408), .A2(n5407), .ZN(n5409) );
  NAND2_X1 U6862 ( .A1(n5410), .A2(n5409), .ZN(n7160) );
  NAND2_X1 U6863 ( .A1(n7160), .A2(n5411), .ZN(n7174) );
  XNOR2_X1 U6864 ( .A(n5413), .B(n5412), .ZN(n7010) );
  NAND2_X1 U6865 ( .A1(n7010), .A2(n7673), .ZN(n5417) );
  NAND2_X1 U6866 ( .A1(n5415), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5450) );
  XNOR2_X1 U6867 ( .A(n5450), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8124) );
  AOI22_X1 U6868 ( .A1(n7665), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6143), .B2(
        n8124), .ZN(n5416) );
  XNOR2_X1 U6869 ( .A(n8848), .B(n5200), .ZN(n5426) );
  NAND2_X1 U6870 ( .A1(n5248), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U6871 ( .A1(n5418), .A2(n7179), .ZN(n5419) );
  AND2_X1 U6872 ( .A1(n5441), .A2(n5419), .ZN(n8717) );
  NAND2_X1 U6873 ( .A1(n5644), .A2(n8717), .ZN(n5422) );
  NAND2_X1 U6874 ( .A1(n4423), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U6875 ( .A1(n5393), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5420) );
  NOR2_X1 U6876 ( .A1(n8371), .A2(n6450), .ZN(n5427) );
  XNOR2_X1 U6877 ( .A(n5426), .B(n5427), .ZN(n7175) );
  INV_X1 U6878 ( .A(n7175), .ZN(n5424) );
  INV_X1 U6879 ( .A(n5426), .ZN(n5429) );
  INV_X1 U6880 ( .A(n5427), .ZN(n5428) );
  NAND2_X1 U6881 ( .A1(n5429), .A2(n5428), .ZN(n5430) );
  XNOR2_X1 U6882 ( .A(n5432), .B(n5431), .ZN(n7367) );
  NAND2_X1 U6883 ( .A1(n7367), .A2(n7673), .ZN(n5436) );
  NAND2_X1 U6884 ( .A1(n5433), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5434) );
  XNOR2_X1 U6885 ( .A(n5434), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8439) );
  AOI22_X1 U6886 ( .A1(n7665), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6143), .B2(
        n8439), .ZN(n5435) );
  XNOR2_X1 U6887 ( .A(n8838), .B(n5200), .ZN(n8285) );
  NAND2_X1 U6888 ( .A1(n5248), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5440) );
  XNOR2_X1 U6889 ( .A(n5469), .B(P2_REG3_REG_16__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U6890 ( .A1(n5644), .A2(n8689), .ZN(n5439) );
  NAND2_X1 U6891 ( .A1(n4423), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5438) );
  NAND2_X1 U6892 ( .A1(n5393), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5437) );
  NOR2_X1 U6893 ( .A1(n8666), .A2(n6450), .ZN(n5457) );
  NAND2_X1 U6894 ( .A1(n5248), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U6895 ( .A1(n5441), .A2(n8366), .ZN(n5442) );
  AND2_X1 U6896 ( .A1(n5469), .A2(n5442), .ZN(n8699) );
  NAND2_X1 U6897 ( .A1(n5644), .A2(n8699), .ZN(n5445) );
  NAND2_X1 U6898 ( .A1(n4423), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U6899 ( .A1(n5393), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5443) );
  NOR2_X1 U6900 ( .A1(n8681), .A2(n6450), .ZN(n8364) );
  XNOR2_X1 U6901 ( .A(n5448), .B(n5447), .ZN(n7379) );
  NAND2_X1 U6902 ( .A1(n7379), .A2(n7673), .ZN(n5454) );
  NAND2_X1 U6903 ( .A1(n5450), .A2(n5449), .ZN(n5451) );
  NAND2_X1 U6904 ( .A1(n5451), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5452) );
  XNOR2_X1 U6905 ( .A(n5452), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8422) );
  AOI22_X1 U6906 ( .A1(n7665), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6143), .B2(
        n8422), .ZN(n5453) );
  XNOR2_X1 U6907 ( .A(n8843), .B(n5200), .ZN(n5456) );
  AOI22_X1 U6908 ( .A1(n8285), .A2(n5457), .B1(n8364), .B2(n5456), .ZN(n5455)
         );
  INV_X1 U6909 ( .A(n8285), .ZN(n5460) );
  OAI21_X1 U6910 ( .B1(n5456), .B2(n8364), .A(n5457), .ZN(n5459) );
  INV_X1 U6911 ( .A(n5456), .ZN(n8283) );
  INV_X1 U6912 ( .A(n8364), .ZN(n5458) );
  INV_X1 U6913 ( .A(n5457), .ZN(n8284) );
  AOI21_X1 U6914 ( .B1(n5460), .B2(n5459), .A(n4457), .ZN(n5461) );
  INV_X1 U6915 ( .A(n8294), .ZN(n5481) );
  XNOR2_X1 U6916 ( .A(n5463), .B(n5462), .ZN(n7310) );
  NAND2_X1 U6917 ( .A1(n7310), .A2(n7673), .ZN(n5466) );
  OR2_X1 U6918 ( .A1(n4435), .A2(n5126), .ZN(n5464) );
  XNOR2_X1 U6919 ( .A(n5464), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8455) );
  AOI22_X1 U6920 ( .A1(n7665), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6143), .B2(
        n8455), .ZN(n5465) );
  XNOR2_X1 U6921 ( .A(n8835), .B(n5200), .ZN(n5475) );
  NAND2_X1 U6922 ( .A1(n4409), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5474) );
  INV_X1 U6923 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5468) );
  INV_X1 U6924 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9951) );
  OAI21_X1 U6925 ( .B1(n5469), .B2(n5468), .A(n9951), .ZN(n5470) );
  AND2_X1 U6926 ( .A1(n5489), .A2(n5470), .ZN(n8673) );
  NAND2_X1 U6927 ( .A1(n5644), .A2(n8673), .ZN(n5473) );
  NAND2_X1 U6928 ( .A1(n4423), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6929 ( .A1(n5393), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5471) );
  NOR2_X1 U6930 ( .A1(n8680), .A2(n6450), .ZN(n5476) );
  NAND2_X1 U6931 ( .A1(n5475), .A2(n5476), .ZN(n5482) );
  INV_X1 U6932 ( .A(n5475), .ZN(n5478) );
  INV_X1 U6933 ( .A(n5476), .ZN(n5477) );
  NAND2_X1 U6934 ( .A1(n5478), .A2(n5477), .ZN(n5479) );
  NAND2_X1 U6935 ( .A1(n5482), .A2(n5479), .ZN(n8293) );
  NAND2_X1 U6936 ( .A1(n5481), .A2(n5480), .ZN(n8295) );
  NAND2_X1 U6937 ( .A1(n8295), .A2(n5482), .ZN(n8342) );
  XNOR2_X1 U6938 ( .A(n5484), .B(n5483), .ZN(n7318) );
  NAND2_X1 U6939 ( .A1(n7318), .A2(n7673), .ZN(n5488) );
  NAND2_X1 U6940 ( .A1(n5485), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5486) );
  XNOR2_X1 U6941 ( .A(n5486), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8468) );
  AOI22_X1 U6942 ( .A1(n7665), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6143), .B2(
        n8468), .ZN(n5487) );
  XNOR2_X1 U6943 ( .A(n8828), .B(n5200), .ZN(n5495) );
  NAND2_X1 U6944 ( .A1(n4409), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U6945 ( .A1(n5489), .A2(n8343), .ZN(n5490) );
  AND2_X1 U6946 ( .A1(n5506), .A2(n5490), .ZN(n8647) );
  NAND2_X1 U6947 ( .A1(n5644), .A2(n8647), .ZN(n5493) );
  NAND2_X1 U6948 ( .A1(n4423), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U6949 ( .A1(n5393), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5491) );
  NOR2_X1 U6950 ( .A1(n8669), .A2(n6450), .ZN(n5496) );
  NAND2_X1 U6951 ( .A1(n5495), .A2(n5496), .ZN(n5500) );
  INV_X1 U6952 ( .A(n5495), .ZN(n5498) );
  INV_X1 U6953 ( .A(n5496), .ZN(n5497) );
  NAND2_X1 U6954 ( .A1(n5498), .A2(n5497), .ZN(n5499) );
  AND2_X1 U6955 ( .A1(n5500), .A2(n5499), .ZN(n8341) );
  NAND2_X1 U6956 ( .A1(n8342), .A2(n8341), .ZN(n8340) );
  NAND2_X1 U6957 ( .A1(n8340), .A2(n5500), .ZN(n8255) );
  XNOR2_X1 U6958 ( .A(n5502), .B(n5501), .ZN(n7327) );
  NAND2_X1 U6959 ( .A1(n7327), .A2(n7673), .ZN(n5504) );
  AOI22_X1 U6960 ( .A1(n7665), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7711), .B2(
        n6143), .ZN(n5503) );
  XNOR2_X1 U6961 ( .A(n8824), .B(n5208), .ZN(n5515) );
  NAND2_X1 U6962 ( .A1(n5248), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5511) );
  INV_X1 U6963 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U6964 ( .A1(n5506), .A2(n5505), .ZN(n5507) );
  AND2_X1 U6965 ( .A1(n5521), .A2(n5507), .ZN(n8633) );
  NAND2_X1 U6966 ( .A1(n5644), .A2(n8633), .ZN(n5510) );
  NAND2_X1 U6967 ( .A1(n4423), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U6968 ( .A1(n5393), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5508) );
  NAND4_X1 U6969 ( .A1(n5511), .A2(n5510), .A3(n5509), .A4(n5508), .ZN(n8652)
         );
  NAND2_X1 U6970 ( .A1(n8652), .A2(n7683), .ZN(n5514) );
  XNOR2_X1 U6971 ( .A(n5515), .B(n5514), .ZN(n8256) );
  INV_X1 U6972 ( .A(n8256), .ZN(n5512) );
  NAND2_X1 U6973 ( .A1(n5515), .A2(n5514), .ZN(n5516) );
  XNOR2_X1 U6974 ( .A(n5518), .B(n5517), .ZN(n7288) );
  NAND2_X1 U6975 ( .A1(n7288), .A2(n7673), .ZN(n5520) );
  NAND2_X1 U6976 ( .A1(n7665), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5519) );
  XNOR2_X1 U6977 ( .A(n8818), .B(n5200), .ZN(n5527) );
  NAND2_X1 U6978 ( .A1(n5248), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U6979 ( .A1(n5521), .A2(n10059), .ZN(n5522) );
  AND2_X1 U6980 ( .A1(n5553), .A2(n5522), .ZN(n8614) );
  NAND2_X1 U6981 ( .A1(n5644), .A2(n8614), .ZN(n5525) );
  NAND2_X1 U6982 ( .A1(n4423), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U6983 ( .A1(n5393), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5523) );
  NOR2_X1 U6984 ( .A1(n8257), .A2(n6450), .ZN(n5528) );
  NAND2_X1 U6985 ( .A1(n5527), .A2(n5528), .ZN(n5532) );
  INV_X1 U6986 ( .A(n5527), .ZN(n5530) );
  INV_X1 U6987 ( .A(n5528), .ZN(n5529) );
  NAND2_X1 U6988 ( .A1(n5530), .A2(n5529), .ZN(n5531) );
  AND2_X1 U6989 ( .A1(n5532), .A2(n5531), .ZN(n8313) );
  XNOR2_X1 U6990 ( .A(n5534), .B(n5533), .ZN(n7277) );
  NAND2_X1 U6991 ( .A1(n7277), .A2(n7673), .ZN(n5536) );
  NAND2_X1 U6992 ( .A1(n7665), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5535) );
  XNOR2_X1 U6993 ( .A(n8600), .B(n5200), .ZN(n5541) );
  NAND2_X1 U6994 ( .A1(n5248), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5540) );
  XNOR2_X1 U6995 ( .A(n5553), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U6996 ( .A1(n5644), .A2(n8598), .ZN(n5539) );
  NAND2_X1 U6997 ( .A1(n4423), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U6998 ( .A1(n5393), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5537) );
  NOR2_X1 U6999 ( .A1(n8623), .A2(n6450), .ZN(n5542) );
  XNOR2_X1 U7000 ( .A(n5541), .B(n5542), .ZN(n8266) );
  NAND2_X1 U7001 ( .A1(n8267), .A2(n8266), .ZN(n8265) );
  INV_X1 U7002 ( .A(n5541), .ZN(n5543) );
  NAND2_X1 U7003 ( .A1(n5543), .A2(n5542), .ZN(n5544) );
  INV_X1 U7004 ( .A(n5545), .ZN(n5547) );
  NAND2_X1 U7005 ( .A1(n5547), .A2(n5546), .ZN(n5548) );
  NAND2_X1 U7006 ( .A1(n5549), .A2(n5548), .ZN(n7298) );
  NAND2_X1 U7007 ( .A1(n7298), .A2(n7673), .ZN(n5551) );
  NAND2_X1 U7008 ( .A1(n7665), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5550) );
  XNOR2_X1 U7009 ( .A(n8808), .B(n5208), .ZN(n5559) );
  NAND2_X1 U7010 ( .A1(n4409), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5558) );
  INV_X1 U7011 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5552) );
  INV_X1 U7012 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8323) );
  OAI21_X1 U7013 ( .B1(n5553), .B2(n5552), .A(n8323), .ZN(n5554) );
  AND2_X1 U7014 ( .A1(n5572), .A2(n5554), .ZN(n8585) );
  NAND2_X1 U7015 ( .A1(n5644), .A2(n8585), .ZN(n5557) );
  NAND2_X1 U7016 ( .A1(n4423), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7017 ( .A1(n5393), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5555) );
  OR2_X1 U7018 ( .A1(n8248), .A2(n6450), .ZN(n8322) );
  INV_X1 U7019 ( .A(n5559), .ZN(n5560) );
  NOR2_X1 U7020 ( .A1(n5561), .A2(n5560), .ZN(n5562) );
  AOI21_X2 U7021 ( .B1(n8321), .B2(n8322), .A(n5562), .ZN(n5581) );
  NAND2_X1 U7022 ( .A1(n5564), .A2(n5563), .ZN(n5566) );
  NAND2_X1 U7023 ( .A1(n5566), .A2(n5565), .ZN(n7351) );
  NAND2_X1 U7024 ( .A1(n7351), .A2(n7673), .ZN(n5568) );
  NAND2_X1 U7025 ( .A1(n7665), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5567) );
  XNOR2_X1 U7026 ( .A(n8803), .B(n5200), .ZN(n5580) );
  XNOR2_X2 U7027 ( .A(n5581), .B(n5570), .ZN(n8246) );
  NAND2_X1 U7028 ( .A1(n5248), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5578) );
  INV_X1 U7029 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U7030 ( .A1(n5572), .A2(n5571), .ZN(n5573) );
  AND2_X1 U7031 ( .A1(n5574), .A2(n5573), .ZN(n8574) );
  NAND2_X1 U7032 ( .A1(n5644), .A2(n8574), .ZN(n5577) );
  NAND2_X1 U7033 ( .A1(n4423), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7034 ( .A1(n5393), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5575) );
  NOR2_X1 U7035 ( .A1(n8591), .A2(n6450), .ZN(n8247) );
  AND2_X1 U7036 ( .A1(n5581), .A2(n5580), .ZN(n8300) );
  OAI21_X1 U7037 ( .B1(n5583), .B2(n5582), .A(n8300), .ZN(n5584) );
  INV_X1 U7038 ( .A(n5586), .ZN(n5590) );
  INV_X1 U7039 ( .A(n5587), .ZN(n5588) );
  NAND2_X1 U7040 ( .A1(n5588), .A2(SI_24_), .ZN(n5589) );
  OAI21_X2 U7041 ( .B1(n5591), .B2(n5590), .A(n5589), .ZN(n5608) );
  INV_X1 U7042 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n5592) );
  INV_X1 U7043 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7171) );
  MUX2_X1 U7044 ( .A(n5592), .B(n7171), .S(n5844), .Z(n5594) );
  INV_X1 U7045 ( .A(SI_25_), .ZN(n5593) );
  NAND2_X1 U7046 ( .A1(n5594), .A2(n5593), .ZN(n5606) );
  INV_X1 U7047 ( .A(n5594), .ZN(n5595) );
  NAND2_X1 U7048 ( .A1(n5595), .A2(SI_25_), .ZN(n5596) );
  NAND2_X1 U7049 ( .A1(n5606), .A2(n5596), .ZN(n5607) );
  NAND2_X1 U7050 ( .A1(n7266), .A2(n7673), .ZN(n5598) );
  NAND2_X1 U7051 ( .A1(n7665), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5597) );
  XNOR2_X1 U7052 ( .A(n8792), .B(n5208), .ZN(n5605) );
  INV_X1 U7053 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8276) );
  NAND2_X1 U7054 ( .A1(n5599), .A2(n8276), .ZN(n5600) );
  NAND2_X1 U7055 ( .A1(n5620), .A2(n5600), .ZN(n8273) );
  INV_X1 U7056 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8548) );
  OAI22_X1 U7057 ( .A1(n8273), .A2(n5722), .B1(n5195), .B2(n8548), .ZN(n5603)
         );
  INV_X1 U7058 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n10033) );
  INV_X1 U7059 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n5601) );
  OAI22_X1 U7060 ( .A1(n5662), .A2(n10033), .B1(n5467), .B2(n5601), .ZN(n5602)
         );
  NAND2_X1 U7061 ( .A1(n8379), .A2(n7683), .ZN(n5604) );
  NOR2_X1 U7062 ( .A1(n5605), .A2(n5604), .ZN(n5628) );
  AOI21_X1 U7063 ( .B1(n5605), .B2(n5604), .A(n5628), .ZN(n8272) );
  INV_X1 U7064 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7186) );
  INV_X1 U7065 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9983) );
  MUX2_X1 U7066 ( .A(n7186), .B(n9983), .S(n4420), .Z(n5610) );
  INV_X1 U7067 ( .A(SI_26_), .ZN(n5609) );
  NAND2_X1 U7068 ( .A1(n5610), .A2(n5609), .ZN(n5633) );
  INV_X1 U7069 ( .A(n5610), .ZN(n5611) );
  NAND2_X1 U7070 ( .A1(n5611), .A2(SI_26_), .ZN(n5612) );
  OR2_X1 U7071 ( .A1(n5614), .A2(n5613), .ZN(n5615) );
  NAND2_X1 U7072 ( .A1(n5634), .A2(n5615), .ZN(n7256) );
  NAND2_X1 U7073 ( .A1(n7256), .A2(n7673), .ZN(n5617) );
  NAND2_X1 U7074 ( .A1(n7665), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5616) );
  NAND2_X2 U7075 ( .A1(n5617), .A2(n5616), .ZN(n8787) );
  XNOR2_X1 U7076 ( .A(n8787), .B(n5208), .ZN(n5626) );
  INV_X1 U7077 ( .A(n5620), .ZN(n5618) );
  NAND2_X1 U7078 ( .A1(n5618), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5642) );
  INV_X1 U7079 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U7080 ( .A1(n5620), .A2(n5619), .ZN(n5621) );
  NAND2_X1 U7081 ( .A1(n5642), .A2(n5621), .ZN(n8524) );
  OR2_X1 U7082 ( .A1(n8524), .A2(n5722), .ZN(n5624) );
  AOI22_X1 U7083 ( .A1(n4409), .A2(P2_REG1_REG_26__SCAN_IN), .B1(n4423), .B2(
        P2_REG0_REG_26__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U7084 ( .A1(n5393), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5622) );
  INV_X1 U7085 ( .A(n8275), .ZN(n8514) );
  NAND2_X1 U7086 ( .A1(n8514), .A2(n7683), .ZN(n5625) );
  NOR2_X1 U7087 ( .A1(n5626), .A2(n5625), .ZN(n5630) );
  AOI21_X1 U7088 ( .B1(n5626), .B2(n5625), .A(n5630), .ZN(n8355) );
  AND2_X1 U7089 ( .A1(n8272), .A2(n8355), .ZN(n5627) );
  INV_X1 U7090 ( .A(n8355), .ZN(n5629) );
  INV_X1 U7091 ( .A(n5628), .ZN(n8349) );
  INV_X1 U7092 ( .A(n5630), .ZN(n5631) );
  NAND2_X1 U7093 ( .A1(n8352), .A2(n5632), .ZN(n8240) );
  NAND2_X2 U7094 ( .A1(n5634), .A2(n5633), .ZN(n5653) );
  INV_X1 U7095 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n10091) );
  INV_X1 U7096 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5635) );
  MUX2_X1 U7097 ( .A(n10091), .B(n5635), .S(n7220), .Z(n5637) );
  INV_X1 U7098 ( .A(SI_27_), .ZN(n5636) );
  NAND2_X1 U7099 ( .A1(n5637), .A2(n5636), .ZN(n5654) );
  INV_X1 U7100 ( .A(n5637), .ZN(n5638) );
  NAND2_X1 U7101 ( .A1(n5638), .A2(SI_27_), .ZN(n5639) );
  NAND2_X1 U7102 ( .A1(n7242), .A2(n7673), .ZN(n5641) );
  OR2_X1 U7103 ( .A1(n7674), .A2(n10091), .ZN(n5640) );
  XNOR2_X1 U7104 ( .A(n8781), .B(n5208), .ZN(n5649) );
  INV_X1 U7105 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U7106 ( .A1(n5642), .A2(n10144), .ZN(n5643) );
  NAND2_X1 U7107 ( .A1(n8510), .A2(n5644), .ZN(n5647) );
  AOI22_X1 U7108 ( .A1(n5248), .A2(P2_REG1_REG_27__SCAN_IN), .B1(n4423), .B2(
        P2_REG0_REG_27__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U7109 ( .A1(n5393), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5645) );
  INV_X1 U7110 ( .A(n8357), .ZN(n8378) );
  NAND2_X1 U7111 ( .A1(n8378), .A2(n7683), .ZN(n5648) );
  NOR2_X1 U7112 ( .A1(n5649), .A2(n5648), .ZN(n5650) );
  AOI21_X1 U7113 ( .B1(n5649), .B2(n5648), .A(n5650), .ZN(n8239) );
  INV_X1 U7114 ( .A(n5650), .ZN(n5651) );
  MUX2_X1 U7115 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n4420), .Z(n7218) );
  INV_X1 U7116 ( .A(SI_28_), .ZN(n9998) );
  XNOR2_X1 U7117 ( .A(n7218), .B(n9998), .ZN(n7216) );
  NAND2_X1 U7118 ( .A1(n8235), .A2(n7673), .ZN(n5656) );
  INV_X1 U7119 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10185) );
  OR2_X1 U7120 ( .A1(n7674), .A2(n10185), .ZN(n5655) );
  INV_X1 U7121 ( .A(n5658), .ZN(n5657) );
  NAND2_X1 U7122 ( .A1(n5657), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8500) );
  INV_X1 U7123 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U7124 ( .A1(n5658), .A2(n5719), .ZN(n5659) );
  NAND2_X1 U7125 ( .A1(n8500), .A2(n5659), .ZN(n7199) );
  INV_X1 U7126 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10112) );
  NAND2_X1 U7127 ( .A1(n4409), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7128 ( .A1(n5393), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5660) );
  OAI211_X1 U7129 ( .C1(n5662), .C2(n10112), .A(n5661), .B(n5660), .ZN(n5663)
         );
  INV_X1 U7130 ( .A(n5663), .ZN(n5664) );
  NOR2_X1 U7131 ( .A1(n8494), .A2(n6450), .ZN(n5666) );
  XNOR2_X1 U7132 ( .A(n5666), .B(n5208), .ZN(n5708) );
  INV_X1 U7133 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7134 ( .A1(n5667), .A2(n5677), .ZN(n5668) );
  NOR2_X1 U7135 ( .A1(n5672), .A2(n5126), .ZN(n5669) );
  MUX2_X1 U7136 ( .A(n5126), .B(n5669), .S(P2_IR_REG_25__SCAN_IN), .Z(n5670)
         );
  INV_X1 U7137 ( .A(n5670), .ZN(n5673) );
  INV_X1 U7138 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U7139 ( .A1(n5672), .A2(n5671), .ZN(n5680) );
  INV_X1 U7140 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5674) );
  INV_X1 U7141 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5698) );
  XOR2_X1 U7142 ( .A(n7069), .B(P2_B_REG_SCAN_IN), .Z(n5679) );
  NAND2_X1 U7143 ( .A1(n5680), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5681) );
  MUX2_X1 U7144 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5681), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5682) );
  INV_X1 U7145 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9758) );
  NOR2_X1 U7146 ( .A1(n7144), .A2(n5696), .ZN(n9759) );
  INV_X1 U7147 ( .A(n5696), .ZN(n7185) );
  INV_X1 U7148 ( .A(n9756), .ZN(n5685) );
  INV_X1 U7149 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9755) );
  NAND2_X1 U7150 ( .A1(n9752), .A2(n9755), .ZN(n5684) );
  NOR4_X1 U7151 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n5689) );
  NOR4_X1 U7152 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n5688) );
  NOR4_X1 U7153 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5687) );
  NOR4_X1 U7154 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5686) );
  NAND4_X1 U7155 ( .A1(n5689), .A2(n5688), .A3(n5687), .A4(n5686), .ZN(n5695)
         );
  NOR2_X1 U7156 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n5693) );
  NOR4_X1 U7157 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n5692) );
  NOR4_X1 U7158 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n5691) );
  NOR4_X1 U7159 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5690) );
  NAND4_X1 U7160 ( .A1(n5693), .A2(n5692), .A3(n5691), .A4(n5690), .ZN(n5694)
         );
  OAI21_X1 U7161 ( .B1(n5695), .B2(n5694), .A(n9752), .ZN(n6266) );
  NAND3_X1 U7162 ( .A1(n6830), .A2(n6289), .A3(n6266), .ZN(n5713) );
  NAND2_X1 U7163 ( .A1(n7144), .A2(n5696), .ZN(n5697) );
  NAND2_X1 U7164 ( .A1(n5701), .A2(n5700), .ZN(n6142) );
  NOR2_X1 U7165 ( .A1(n9763), .A2(n7860), .ZN(n6841) );
  NAND2_X1 U7166 ( .A1(n5720), .A2(n6841), .ZN(n5705) );
  AND2_X1 U7167 ( .A1(n7860), .A2(n7711), .ZN(n5703) );
  NAND2_X1 U7168 ( .A1(n5702), .A2(n5703), .ZN(n9787) );
  INV_X1 U7169 ( .A(n6268), .ZN(n5704) );
  NAND3_X1 U7170 ( .A1(n8776), .A2(n8348), .A3(n5708), .ZN(n5706) );
  OAI21_X1 U7171 ( .B1(n8776), .B2(n5708), .A(n5706), .ZN(n5712) );
  NOR3_X1 U7172 ( .A1(n8485), .A2(n8374), .A3(n5708), .ZN(n5707) );
  AOI21_X1 U7173 ( .B1(n8485), .B2(n5708), .A(n5707), .ZN(n5711) );
  INV_X1 U7174 ( .A(n6512), .ZN(n6274) );
  INV_X1 U7175 ( .A(n5714), .ZN(n7868) );
  AND2_X1 U7176 ( .A1(n6274), .A2(n9810), .ZN(n5709) );
  OAI21_X1 U7177 ( .B1(n8485), .B2(n8348), .A(n8376), .ZN(n5710) );
  NAND2_X1 U7178 ( .A1(n5713), .A2(n6268), .ZN(n5718) );
  AND2_X1 U7179 ( .A1(n6512), .A2(n5714), .ZN(n6265) );
  INV_X1 U7180 ( .A(n6142), .ZN(n5715) );
  NOR2_X1 U7181 ( .A1(n6265), .A2(n5715), .ZN(n5716) );
  AND2_X1 U7182 ( .A1(n6509), .A2(n5716), .ZN(n5717) );
  NAND2_X1 U7183 ( .A1(n5718), .A2(n5717), .ZN(n6448) );
  OAI22_X1 U7184 ( .A1(n8368), .A2(n7199), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5719), .ZN(n5727) );
  NAND2_X1 U7185 ( .A1(n5720), .A2(n7868), .ZN(n8278) );
  AND2_X1 U7186 ( .A1(n6512), .A2(n5721), .ZN(n8731) );
  OR2_X1 U7187 ( .A1(n8500), .A2(n5722), .ZN(n5725) );
  AOI22_X1 U7188 ( .A1(P2_REG1_REG_29__SCAN_IN), .A2(n4409), .B1(n4423), .B2(
        P2_REG0_REG_29__SCAN_IN), .ZN(n5724) );
  NAND2_X1 U7189 ( .A1(n5393), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5723) );
  OAI22_X1 U7190 ( .A1(n8357), .A2(n8370), .B1(n8369), .B2(n7668), .ZN(n5726)
         );
  AND2_X2 U7191 ( .A1(n5775), .A2(n5728), .ZN(n5793) );
  NOR2_X1 U7192 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5733) );
  INV_X1 U7193 ( .A(n5741), .ZN(n5735) );
  NOR2_X1 U7194 ( .A1(n5735), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5736) );
  INV_X1 U7195 ( .A(n5753), .ZN(n5737) );
  AOI21_X1 U7196 ( .B1(n5737), .B2(n5740), .A(n9415), .ZN(n5738) );
  MUX2_X1 U7197 ( .A(n9415), .B(n5738), .S(P1_IR_REG_23__SCAN_IN), .Z(n5742)
         );
  OR2_X1 U7198 ( .A1(n5742), .A2(n5743), .ZN(n6998) );
  NAND2_X1 U7199 ( .A1(n5762), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U7200 ( .A1(n5751), .A2(n5750), .ZN(n5744) );
  NAND2_X1 U7201 ( .A1(n5744), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5746) );
  INV_X1 U7202 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5745) );
  XNOR2_X1 U7203 ( .A(n5746), .B(n5745), .ZN(n7187) );
  INV_X1 U7204 ( .A(n5743), .ZN(n5747) );
  NAND2_X1 U7205 ( .A1(n5747), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5749) );
  XNOR2_X1 U7206 ( .A(n5749), .B(n5748), .ZN(n7071) );
  XNOR2_X1 U7207 ( .A(n5751), .B(n5750), .ZN(n7169) );
  INV_X1 U7208 ( .A(n6123), .ZN(n5961) );
  AND2_X1 U7209 ( .A1(n6998), .A2(n5961), .ZN(n5878) );
  INV_X1 U7210 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U7211 ( .A1(n5757), .A2(n5754), .ZN(n5759) );
  NAND2_X1 U7212 ( .A1(n5759), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5756) );
  INV_X1 U7213 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5755) );
  INV_X1 U7214 ( .A(n5757), .ZN(n5758) );
  NAND2_X1 U7215 ( .A1(n5758), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n5760) );
  NAND2_X1 U7216 ( .A1(n7646), .A2(n5807), .ZN(n7631) );
  NAND2_X1 U7217 ( .A1(n7631), .A2(n6123), .ZN(n5761) );
  NAND2_X1 U7218 ( .A1(n5761), .A2(n6998), .ZN(n5904) );
  INV_X1 U7219 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5763) );
  NAND2_X2 U7220 ( .A1(n5809), .A2(n9532), .ZN(n6105) );
  NAND2_X1 U7221 ( .A1(n5904), .A2(n6105), .ZN(n5883) );
  NAND2_X1 U7222 ( .A1(n5883), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  MUX2_X1 U7223 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5770), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5771) );
  NAND2_X1 U7224 ( .A1(n6348), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U7225 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5774) );
  MUX2_X1 U7226 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5774), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5777) );
  NAND2_X1 U7227 ( .A1(n5777), .A2(n5776), .ZN(n5980) );
  INV_X1 U7228 ( .A(n5980), .ZN(n5778) );
  NAND2_X1 U7229 ( .A1(n7382), .A2(n5778), .ZN(n5779) );
  OAI211_X2 U7230 ( .C1(n6644), .C2(n5853), .A(n5780), .B(n5779), .ZN(n7400)
         );
  NAND2_X1 U7231 ( .A1(n7459), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U7232 ( .A1(n7324), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U7233 ( .A1(n4416), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U7234 ( .A1(n4414), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5781) );
  INV_X1 U7235 ( .A(SI_0_), .ZN(n5785) );
  NOR2_X1 U7236 ( .A1(n7229), .A2(n5785), .ZN(n5786) );
  XNOR2_X1 U7237 ( .A(n5786), .B(n5001), .ZN(n9426) );
  MUX2_X1 U7238 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9426), .S(n6105), .Z(n6179) );
  INV_X1 U7239 ( .A(n6179), .ZN(n6194) );
  INV_X1 U7240 ( .A(n9055), .ZN(n7401) );
  NAND2_X1 U7241 ( .A1(n7401), .A2(n7400), .ZN(n5787) );
  NAND2_X1 U7242 ( .A1(n7459), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U7243 ( .A1(n7324), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U7244 ( .A1(n4417), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U7245 ( .A1(n4414), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U7246 ( .A1(n6348), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5796) );
  MUX2_X1 U7247 ( .A(n9415), .B(n5792), .S(P1_IR_REG_2__SCAN_IN), .Z(n5794) );
  NAND2_X1 U7248 ( .A1(n7382), .A2(n9529), .ZN(n5795) );
  OAI211_X1 U7249 ( .C1(n6644), .C2(n5859), .A(n5796), .B(n5795), .ZN(n7404)
         );
  XNOR2_X1 U7250 ( .A(n9054), .B(n7404), .ZN(n7472) );
  XNOR2_X1 U7251 ( .A(n7407), .B(n5804), .ZN(n5817) );
  NAND2_X1 U7252 ( .A1(n5797), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5798) );
  XNOR2_X2 U7253 ( .A(n5798), .B(n4562), .ZN(n9243) );
  OR2_X1 U7254 ( .A1(n6846), .A2(n9243), .ZN(n5802) );
  NAND2_X1 U7255 ( .A1(n4478), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5800) );
  XNOR2_X1 U7256 ( .A(n5800), .B(n5799), .ZN(n6678) );
  INV_X1 U7257 ( .A(n6678), .ZN(n7638) );
  NAND2_X1 U7258 ( .A1(n5807), .A2(n7638), .ZN(n5801) );
  AND2_X1 U7259 ( .A1(n6057), .A2(n6179), .ZN(n6184) );
  NAND2_X1 U7260 ( .A1(n6185), .A2(n6184), .ZN(n6183) );
  NAND2_X1 U7261 ( .A1(n9055), .A2(n7400), .ZN(n5803) );
  INV_X1 U7262 ( .A(n7472), .ZN(n5804) );
  NAND2_X1 U7263 ( .A1(n5805), .A2(n7472), .ZN(n5806) );
  NAND2_X1 U7264 ( .A1(n6209), .A2(n5806), .ZN(n9677) );
  NAND2_X1 U7265 ( .A1(n5807), .A2(n6678), .ZN(n5954) );
  INV_X1 U7266 ( .A(n5954), .ZN(n5957) );
  AND3_X1 U7267 ( .A1(n5957), .A2(n7646), .A3(n9243), .ZN(n7644) );
  NOR2_X1 U7268 ( .A1(n7644), .A2(n7661), .ZN(n5808) );
  NAND2_X1 U7269 ( .A1(n5808), .A2(n8005), .ZN(n6574) );
  INV_X1 U7270 ( .A(n6574), .ZN(n9648) );
  NAND2_X1 U7271 ( .A1(n9677), .A2(n9648), .ZN(n5816) );
  INV_X1 U7272 ( .A(n9536), .ZN(n7643) );
  NAND2_X1 U7273 ( .A1(n7324), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7274 ( .A1(n4416), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7275 ( .A1(n4414), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5812) );
  INV_X1 U7276 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U7277 ( .A1(n7459), .A2(n5810), .ZN(n5811) );
  OR2_X1 U7278 ( .A1(n7631), .A2(n9536), .ZN(n9464) );
  AOI22_X1 U7279 ( .A1(n9293), .A2(n9053), .B1(n9055), .B2(n9291), .ZN(n5815)
         );
  OAI211_X1 U7280 ( .C1(n5817), .C2(n9459), .A(n5816), .B(n5815), .ZN(n9675)
         );
  NAND2_X1 U7281 ( .A1(n7169), .A2(P1_B_REG_SCAN_IN), .ZN(n5818) );
  MUX2_X1 U7282 ( .A(P1_B_REG_SCAN_IN), .B(n5818), .S(n7071), .Z(n5820) );
  INV_X1 U7283 ( .A(n7187), .ZN(n5819) );
  NAND2_X1 U7284 ( .A1(n5820), .A2(n5819), .ZN(n5863) );
  OR2_X1 U7285 ( .A1(n5863), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U7286 ( .A1(n7187), .A2(n7071), .ZN(n5864) );
  INV_X1 U7287 ( .A(n5949), .ZN(n6037) );
  AND2_X1 U7288 ( .A1(n6678), .A2(n9243), .ZN(n5955) );
  OR2_X1 U7289 ( .A1(n7631), .A2(n5955), .ZN(n6124) );
  NAND2_X1 U7290 ( .A1(n6037), .A2(n6124), .ZN(n6030) );
  INV_X1 U7291 ( .A(n6030), .ZN(n5835) );
  OR2_X1 U7292 ( .A1(n5863), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U7293 ( .A1(n7187), .A2(n7169), .ZN(n5870) );
  AND2_X1 U7294 ( .A1(n5822), .A2(n5870), .ZN(n6025) );
  NOR4_X1 U7295 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5831) );
  NOR4_X1 U7296 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5830) );
  INV_X1 U7297 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10137) );
  INV_X1 U7298 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10181) );
  INV_X1 U7299 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10094) );
  INV_X1 U7300 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10123) );
  NAND4_X1 U7301 ( .A1(n10137), .A2(n10181), .A3(n10094), .A4(n10123), .ZN(
        n5828) );
  NOR4_X1 U7302 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5826) );
  NOR4_X1 U7303 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5825) );
  NOR4_X1 U7304 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5824) );
  NOR4_X1 U7305 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5823) );
  NAND4_X1 U7306 ( .A1(n5826), .A2(n5825), .A3(n5824), .A4(n5823), .ZN(n5827)
         );
  NOR4_X1 U7307 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5828), .A4(n5827), .ZN(n5829) );
  AND3_X1 U7308 ( .A1(n5831), .A2(n5830), .A3(n5829), .ZN(n5832) );
  OR2_X1 U7309 ( .A1(n5863), .A2(n5832), .ZN(n6027) );
  AND2_X1 U7310 ( .A1(n6025), .A2(n6027), .ZN(n5950) );
  AND2_X1 U7311 ( .A1(n6123), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5833) );
  AND2_X1 U7312 ( .A1(n5950), .A2(n7641), .ZN(n5834) );
  NAND2_X1 U7313 ( .A1(n5835), .A2(n5834), .ZN(n5839) );
  NOR2_X1 U7314 ( .A1(n6029), .A2(n5807), .ZN(n5836) );
  MUX2_X1 U7315 ( .A(n9675), .B(P1_REG2_REG_2__SCAN_IN), .S(n4419), .Z(n5843)
         );
  INV_X1 U7316 ( .A(n9677), .ZN(n5838) );
  OR2_X1 U7317 ( .A1(n5954), .A2(n9243), .ZN(n5837) );
  OR2_X1 U7318 ( .A1(n4419), .A2(n5837), .ZN(n6583) );
  NOR2_X1 U7319 ( .A1(n5838), .A2(n6583), .ZN(n5842) );
  NOR2_X1 U7320 ( .A1(n5839), .A2(n7661), .ZN(n9475) );
  INV_X1 U7321 ( .A(n9475), .ZN(n7031) );
  NAND2_X1 U7322 ( .A1(n6846), .A2(n7630), .ZN(n6034) );
  NOR2_X2 U7323 ( .A1(n7031), .A2(n9692), .ZN(n9650) );
  INV_X1 U7324 ( .A(n9650), .ZN(n6591) );
  INV_X1 U7325 ( .A(n7404), .ZN(n9674) );
  NOR2_X1 U7326 ( .A1(n6192), .A2(n9674), .ZN(n9672) );
  NOR3_X1 U7327 ( .A1(n6591), .A2(n4508), .A3(n9672), .ZN(n5841) );
  INV_X1 U7328 ( .A(n6034), .ZN(n6032) );
  INV_X1 U7329 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6150) );
  OAI22_X1 U7330 ( .A1(n9656), .A2(n9674), .B1(n9258), .B2(n6150), .ZN(n5840)
         );
  OR4_X1 U7331 ( .A1(n5843), .A2(n5842), .A3(n5841), .A4(n5840), .ZN(P1_U3289)
         );
  NAND2_X1 U7332 ( .A1(n7220), .A2(P2_U3152), .ZN(n8237) );
  INV_X1 U7333 ( .A(n8237), .ZN(n7143) );
  INV_X1 U7334 ( .A(n7143), .ZN(n8881) );
  OAI222_X1 U7335 ( .A1(n8881), .A2(n5845), .B1(n8236), .B2(n5853), .C1(n9427), 
        .C2(P2_U3152), .ZN(P2_U3357) );
  NAND2_X1 U7336 ( .A1(n5849), .A2(n5850), .ZN(n5898) );
  NAND2_X1 U7337 ( .A1(n5898), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5867) );
  XNOR2_X1 U7338 ( .A(n5867), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U7339 ( .A1(n7229), .A2(P1_U3084), .ZN(n8231) );
  INV_X1 U7340 ( .A(n8231), .ZN(n9421) );
  AOI22_X1 U7341 ( .A1(n6297), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9421), .ZN(n5846) );
  OAI21_X1 U7342 ( .B1(n6296), .B2(n9424), .A(n5846), .ZN(P1_U3348) );
  OR2_X1 U7343 ( .A1(n5793), .A2(n9415), .ZN(n5847) );
  XNOR2_X1 U7344 ( .A(n5847), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6087) );
  AOI22_X1 U7345 ( .A1(n6087), .A2(P1_STATE_REG_SCAN_IN), .B1(n9421), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n5848) );
  OAI21_X1 U7346 ( .B1(n6089), .B2(n9424), .A(n5848), .ZN(P1_U3350) );
  OR2_X1 U7347 ( .A1(n5849), .A2(n9415), .ZN(n5851) );
  XNOR2_X1 U7348 ( .A(n5851), .B(n5850), .ZN(n9545) );
  OAI222_X1 U7349 ( .A1(n8231), .A2(n10108), .B1(n9424), .B2(n6102), .C1(
        P1_U3084), .C2(n9545), .ZN(P1_U3349) );
  INV_X1 U7350 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5852) );
  OAI222_X1 U7351 ( .A1(P1_U3084), .A2(n5980), .B1(n9424), .B2(n5853), .C1(
        n5852), .C2(n8231), .ZN(P1_U3352) );
  INV_X1 U7352 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9981) );
  INV_X1 U7353 ( .A(n9529), .ZN(n5854) );
  OAI222_X1 U7354 ( .A1(n8231), .A2(n9981), .B1(n9424), .B2(n5859), .C1(
        P1_U3084), .C2(n5854), .ZN(P1_U3351) );
  INV_X1 U7355 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U7356 ( .A1(n5867), .A2(n5855), .ZN(n5856) );
  NAND2_X1 U7357 ( .A1(n5856), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5857) );
  XNOR2_X1 U7358 ( .A(n5857), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6349) );
  INV_X1 U7359 ( .A(n6349), .ZN(n6014) );
  OAI222_X1 U7360 ( .A1(n8231), .A2(n5858), .B1(n9424), .B2(n6347), .C1(
        P1_U3084), .C2(n6014), .ZN(P1_U3347) );
  OAI222_X1 U7361 ( .A1(n8881), .A2(n10154), .B1(n8236), .B2(n5859), .C1(
        P2_U3152), .C2(n9444), .ZN(P2_U3356) );
  OAI222_X1 U7362 ( .A1(n8881), .A2(n5860), .B1(n8236), .B2(n6102), .C1(
        P2_U3152), .C2(n8402), .ZN(P2_U3354) );
  OAI222_X1 U7363 ( .A1(n8881), .A2(n10109), .B1(n8236), .B2(n6296), .C1(
        P2_U3152), .C2(n6548), .ZN(P2_U3353) );
  OAI222_X1 U7364 ( .A1(n8881), .A2(n5861), .B1(n8236), .B2(n6089), .C1(
        P2_U3152), .C2(n6533), .ZN(P2_U3355) );
  OAI222_X1 U7365 ( .A1(n8881), .A2(n5862), .B1(n8236), .B2(n6347), .C1(
        P2_U3152), .C2(n8111), .ZN(P2_U3352) );
  NAND2_X1 U7366 ( .A1(n7641), .A2(n5863), .ZN(n9664) );
  INV_X1 U7367 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10111) );
  INV_X1 U7368 ( .A(n5864), .ZN(n5865) );
  AOI22_X1 U7369 ( .A1(n9664), .A2(n10111), .B1(n5865), .B2(n7641), .ZN(
        P1_U3440) );
  NOR2_X1 U7370 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5896) );
  OR2_X1 U7371 ( .A1(n5896), .A2(n9415), .ZN(n5866) );
  NAND2_X1 U7372 ( .A1(n5867), .A2(n5866), .ZN(n5872) );
  INV_X1 U7373 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5893) );
  XNOR2_X1 U7374 ( .A(n5872), .B(n5893), .ZN(n9562) );
  AOI22_X1 U7375 ( .A1(n9562), .A2(P1_STATE_REG_SCAN_IN), .B1(n9421), .B2(
        P2_DATAO_REG_7__SCAN_IN), .ZN(n5868) );
  OAI21_X1 U7376 ( .B1(n6354), .B2(n9424), .A(n5868), .ZN(P1_U3346) );
  OAI222_X1 U7377 ( .A1(n8881), .A2(n5869), .B1(n8236), .B2(n6354), .C1(
        P2_U3152), .C2(n9882), .ZN(P2_U3351) );
  OAI22_X1 U7378 ( .A1(n9663), .A2(P1_D_REG_1__SCAN_IN), .B1(n6029), .B2(n5870), .ZN(n5871) );
  INV_X1 U7379 ( .A(n5871), .ZN(P1_U3441) );
  NAND2_X1 U7380 ( .A1(n5873), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7381 ( .A1(n5874), .A2(n5895), .ZN(n5889) );
  OR2_X1 U7382 ( .A1(n5874), .A2(n5895), .ZN(n5875) );
  NAND2_X1 U7383 ( .A1(n5889), .A2(n5875), .ZN(n9582) );
  OAI222_X1 U7384 ( .A1(n8231), .A2(n5876), .B1(n9424), .B2(n6557), .C1(
        P1_U3084), .C2(n9582), .ZN(P1_U3345) );
  OAI222_X1 U7385 ( .A1(n8881), .A2(n5877), .B1(n8236), .B2(n6557), .C1(
        P2_U3152), .C2(n8099), .ZN(P2_U3350) );
  NOR2_X1 U7386 ( .A1(n9532), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5879) );
  INV_X1 U7387 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5974) );
  OAI21_X1 U7388 ( .B1(n9536), .B2(n5879), .A(n5974), .ZN(n9535) );
  INV_X1 U7389 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6043) );
  INV_X1 U7390 ( .A(n9532), .ZN(n7642) );
  NAND2_X1 U7391 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9534) );
  NAND2_X1 U7392 ( .A1(n7642), .A2(n9534), .ZN(n5880) );
  OAI211_X1 U7393 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n6043), .A(n7643), .B(n5880), .ZN(n5881) );
  NAND3_X1 U7394 ( .A1(n9535), .A2(P1_STATE_REG_SCAN_IN), .A3(n5881), .ZN(
        n5882) );
  NOR2_X1 U7395 ( .A1(n5883), .A2(n5882), .ZN(n5886) );
  OR2_X1 U7396 ( .A1(n9536), .A2(P1_U3084), .ZN(n9422) );
  NOR2_X1 U7397 ( .A1(n9422), .A2(n7642), .ZN(n5884) );
  NAND2_X1 U7398 ( .A1(n5904), .A2(n5884), .ZN(n9060) );
  AND3_X1 U7399 ( .A1(n9641), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6043), .ZN(n5885) );
  AOI211_X1 U7400 ( .C1(P1_REG3_REG_0__SCAN_IN), .C2(P1_U3084), .A(n5886), .B(
        n5885), .ZN(n5887) );
  OAI21_X1 U7401 ( .B1(n9627), .B2(n9844), .A(n5887), .ZN(P1_U3241) );
  INV_X1 U7402 ( .A(n6645), .ZN(n5892) );
  INV_X1 U7403 ( .A(n8036), .ZN(n8087) );
  OAI222_X1 U7404 ( .A1(n8881), .A2(n5888), .B1(n8236), .B2(n5892), .C1(n8087), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  NAND2_X1 U7405 ( .A1(n5889), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5890) );
  XNOR2_X1 U7406 ( .A(n5890), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9599) );
  INV_X1 U7407 ( .A(n9599), .ZN(n5891) );
  OAI222_X1 U7408 ( .A1(n8231), .A2(n10204), .B1(n9424), .B2(n5892), .C1(n5891), .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U7409 ( .A(n6686), .ZN(n5970) );
  INV_X1 U7410 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5894) );
  NAND4_X1 U7411 ( .A1(n5896), .A2(n5895), .A3(n5894), .A4(n5893), .ZN(n5897)
         );
  NOR2_X1 U7412 ( .A1(n5898), .A2(n5897), .ZN(n5901) );
  OR2_X1 U7413 ( .A1(n5901), .A2(n9415), .ZN(n5899) );
  MUX2_X1 U7414 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5899), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5902) );
  INV_X1 U7415 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7416 ( .A1(n5901), .A2(n5900), .ZN(n6023) );
  AOI22_X1 U7417 ( .A1(n6687), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9421), .ZN(n5903) );
  OAI21_X1 U7418 ( .B1(n5970), .B2(n9424), .A(n5903), .ZN(P1_U3343) );
  INV_X1 U7419 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n5923) );
  NOR2_X1 U7420 ( .A1(n9532), .A2(P1_U3084), .ZN(n7189) );
  NAND2_X1 U7421 ( .A1(n5904), .A2(n7189), .ZN(n7659) );
  INV_X1 U7422 ( .A(n7659), .ZN(n5905) );
  AND2_X1 U7423 ( .A1(n5905), .A2(n9536), .ZN(n9635) );
  AND2_X1 U7424 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3084), .ZN(n5911) );
  INV_X1 U7425 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5906) );
  MUX2_X1 U7426 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n5906), .S(n9529), .Z(n9541)
         );
  INV_X1 U7427 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9700) );
  MUX2_X1 U7428 ( .A(n9700), .B(P1_REG1_REG_1__SCAN_IN), .S(n5980), .Z(n5976)
         );
  NAND3_X1 U7429 ( .A1(n5976), .A2(P1_REG1_REG_0__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n5975) );
  OAI21_X1 U7430 ( .B1(n9700), .B2(n5980), .A(n5975), .ZN(n9542) );
  NAND2_X1 U7431 ( .A1(n9541), .A2(n9542), .ZN(n9540) );
  NAND2_X1 U7432 ( .A1(n9529), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5908) );
  INV_X1 U7433 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6217) );
  MUX2_X1 U7434 ( .A(n6217), .B(P1_REG1_REG_3__SCAN_IN), .S(n6087), .Z(n5907)
         );
  AND3_X1 U7435 ( .A1(n9540), .A2(n5908), .A3(n5907), .ZN(n5909) );
  NOR3_X1 U7436 ( .A1(n9060), .A2(n5924), .A3(n5909), .ZN(n5910) );
  AOI211_X1 U7437 ( .C1(n9635), .C2(n6087), .A(n5911), .B(n5910), .ZN(n5922)
         );
  OR2_X1 U7438 ( .A1(n7659), .A2(n9536), .ZN(n9629) );
  INV_X1 U7439 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5912) );
  INV_X1 U7440 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5914) );
  MUX2_X1 U7441 ( .A(n5914), .B(P1_REG2_REG_1__SCAN_IN), .S(n5980), .Z(n5983)
         );
  AND2_X1 U7442 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n5913) );
  NAND2_X1 U7443 ( .A1(n5983), .A2(n5913), .ZN(n5982) );
  OAI21_X1 U7444 ( .B1(n5914), .B2(n5980), .A(n5982), .ZN(n9527) );
  NAND2_X1 U7445 ( .A1(n9529), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5919) );
  INV_X1 U7446 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5915) );
  MUX2_X1 U7447 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n5915), .S(n6087), .Z(n5916)
         );
  NAND2_X1 U7448 ( .A1(n5917), .A2(n5916), .ZN(n5930) );
  MUX2_X1 U7449 ( .A(n5915), .B(P1_REG2_REG_3__SCAN_IN), .S(n6087), .Z(n5918)
         );
  NAND3_X1 U7450 ( .A1(n9526), .A2(n5919), .A3(n5918), .ZN(n5920) );
  NAND3_X1 U7451 ( .A1(n9623), .A2(n5930), .A3(n5920), .ZN(n5921) );
  OAI211_X1 U7452 ( .C1(n5923), .C2(n9627), .A(n5922), .B(n5921), .ZN(P1_U3244) );
  INV_X1 U7453 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n5940) );
  AND2_X1 U7454 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3084), .ZN(n5928) );
  INV_X1 U7455 ( .A(n9545), .ZN(n9549) );
  AOI21_X1 U7456 ( .B1(n6087), .B2(P1_REG1_REG_3__SCAN_IN), .A(n5924), .ZN(
        n9555) );
  INV_X1 U7457 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10032) );
  MUX2_X1 U7458 ( .A(n10032), .B(P1_REG1_REG_4__SCAN_IN), .S(n9545), .Z(n9556)
         );
  NAND2_X1 U7459 ( .A1(n9555), .A2(n9556), .ZN(n9554) );
  OAI21_X1 U7460 ( .B1(n9549), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9554), .ZN(
        n5926) );
  INV_X1 U7461 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6423) );
  MUX2_X1 U7462 ( .A(n6423), .B(P1_REG1_REG_5__SCAN_IN), .S(n6297), .Z(n5925)
         );
  AOI211_X1 U7463 ( .C1(n5926), .C2(n5925), .A(n9060), .B(n5988), .ZN(n5927)
         );
  AOI211_X1 U7464 ( .C1(n9635), .C2(n6297), .A(n5928), .B(n5927), .ZN(n5939)
         );
  NAND2_X1 U7465 ( .A1(n6087), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5929) );
  INV_X1 U7466 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5931) );
  MUX2_X1 U7467 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n5931), .S(n9545), .Z(n5932)
         );
  AND2_X1 U7468 ( .A1(n9545), .A2(n5931), .ZN(n5934) );
  INV_X1 U7469 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5933) );
  MUX2_X1 U7470 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n5933), .S(n6297), .Z(n5935)
         );
  INV_X1 U7471 ( .A(n9546), .ZN(n5936) );
  NOR3_X1 U7472 ( .A1(n5936), .A2(n5935), .A3(n5934), .ZN(n5937) );
  OAI21_X1 U7473 ( .B1(n5997), .B2(n5937), .A(n9623), .ZN(n5938) );
  OAI211_X1 U7474 ( .C1(n5940), .C2(n9627), .A(n5939), .B(n5938), .ZN(P1_U3246) );
  INV_X1 U7475 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5942) );
  NAND2_X1 U7476 ( .A1(n6057), .A2(P1_U4006), .ZN(n5941) );
  OAI21_X1 U7477 ( .B1(P1_U4006), .B2(n5942), .A(n5941), .ZN(P1_U3555) );
  INV_X1 U7478 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7479 ( .A1(n4414), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7480 ( .A1(n4416), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7481 ( .A1(n7324), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5944) );
  NAND3_X1 U7482 ( .A1(n5946), .A2(n5945), .A3(n5944), .ZN(n7899) );
  NAND2_X1 U7483 ( .A1(n7899), .A2(P1_U4006), .ZN(n5947) );
  OAI21_X1 U7484 ( .B1(P1_U4006), .B2(n5948), .A(n5947), .ZN(P1_U3586) );
  NAND2_X1 U7485 ( .A1(n5950), .A2(n5949), .ZN(n6128) );
  INV_X1 U7486 ( .A(n6128), .ZN(n5951) );
  AND2_X1 U7487 ( .A1(n5951), .A2(n7641), .ZN(n5965) );
  NAND2_X1 U7488 ( .A1(n5965), .A2(n7644), .ZN(n6056) );
  AOI21_X1 U7489 ( .B1(n9392), .B2(n5966), .A(n5951), .ZN(n5952) );
  NAND2_X1 U7490 ( .A1(n6124), .A2(n7641), .ZN(n6038) );
  NOR2_X1 U7491 ( .A1(n5952), .A2(n6038), .ZN(n6151) );
  INV_X1 U7492 ( .A(n6151), .ZN(n6055) );
  AND2_X1 U7493 ( .A1(n9691), .A2(n7631), .ZN(n5953) );
  AND2_X1 U7494 ( .A1(n5954), .A2(n6123), .ZN(n6077) );
  NAND2_X1 U7495 ( .A1(n6846), .A2(n5955), .ZN(n5956) );
  AND2_X2 U7496 ( .A1(n6077), .A2(n5956), .ZN(n8007) );
  NAND2_X1 U7497 ( .A1(n6057), .A2(n8007), .ZN(n5960) );
  AND2_X2 U7498 ( .A1(n5957), .A2(n6123), .ZN(n6394) );
  NOR2_X1 U7499 ( .A1(n6123), .A2(n5974), .ZN(n5958) );
  AOI21_X1 U7500 ( .B1(n6179), .B2(n6394), .A(n5958), .ZN(n5959) );
  AND2_X1 U7501 ( .A1(n5960), .A2(n5959), .ZN(n5964) );
  NAND2_X1 U7502 ( .A1(n6057), .A2(n6394), .ZN(n5963) );
  AOI22_X1 U7503 ( .A1(n6179), .A2(n6077), .B1(n5961), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7504 ( .A1(n5963), .A2(n5962), .ZN(n6048) );
  OAI21_X1 U7505 ( .B1(n5964), .B2(n6048), .A(n6050), .ZN(n9533) );
  AOI22_X1 U7506 ( .A1(n6055), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9015), .B2(
        n9533), .ZN(n5969) );
  INV_X1 U7507 ( .A(n5965), .ZN(n5967) );
  OAI21_X2 U7508 ( .B1(n5967), .B2(n5966), .A(n9258), .ZN(n9036) );
  NAND2_X1 U7509 ( .A1(n9036), .A2(n6179), .ZN(n5968) );
  OAI211_X1 U7510 ( .C1(n7401), .C2(n9009), .A(n5969), .B(n5968), .ZN(P1_U3230) );
  INV_X1 U7511 ( .A(n8033), .ZN(n8075) );
  OAI222_X1 U7512 ( .A1(n8237), .A2(n10174), .B1(n8236), .B2(n5970), .C1(n8075), .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7513 ( .A(n6691), .ZN(n5973) );
  NAND2_X1 U7514 ( .A1(n6023), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5971) );
  XNOR2_X1 U7515 ( .A(n5971), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9603) );
  INV_X1 U7516 ( .A(n9603), .ZN(n6171) );
  OAI222_X1 U7517 ( .A1(n8231), .A2(n5972), .B1(n9424), .B2(n5973), .C1(n6171), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U7518 ( .A(n8167), .ZN(n8056) );
  OAI222_X1 U7519 ( .A1(n8237), .A2(n9996), .B1(n8236), .B2(n5973), .C1(n8056), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U7520 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n5986) );
  INV_X1 U7521 ( .A(n9635), .ZN(n9069) );
  NAND2_X1 U7522 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P1_U3084), .ZN(n5979) );
  NOR2_X1 U7523 ( .A1(n5974), .A2(n6043), .ZN(n5977) );
  OAI211_X1 U7524 ( .C1(n5977), .C2(n5976), .A(n9641), .B(n5975), .ZN(n5978)
         );
  OAI211_X1 U7525 ( .C1(n9069), .C2(n5980), .A(n5979), .B(n5978), .ZN(n5981)
         );
  INV_X1 U7526 ( .A(n5981), .ZN(n5985) );
  OAI211_X1 U7527 ( .C1(n5913), .C2(n5983), .A(n9623), .B(n5982), .ZN(n5984)
         );
  OAI211_X1 U7528 ( .C1(n5986), .C2(n9627), .A(n5985), .B(n5984), .ZN(P1_U3242) );
  NOR2_X1 U7529 ( .A1(n9599), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5987) );
  AOI21_X1 U7530 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9599), .A(n5987), .ZN(
        n9591) );
  NOR2_X1 U7531 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n9562), .ZN(n5989) );
  AOI21_X1 U7532 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n6297), .A(n5988), .ZN(
        n6012) );
  INV_X1 U7533 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9705) );
  MUX2_X1 U7534 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n9705), .S(n6349), .Z(n6011)
         );
  NAND2_X1 U7535 ( .A1(n6012), .A2(n6011), .ZN(n6010) );
  OAI21_X1 U7536 ( .B1(n6349), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6010), .ZN(
        n9568) );
  INV_X1 U7537 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6478) );
  MUX2_X1 U7538 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6478), .S(n9562), .Z(n9567)
         );
  INV_X1 U7539 ( .A(n9584), .ZN(n5990) );
  INV_X1 U7540 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9708) );
  OAI21_X1 U7541 ( .B1(n5990), .B2(n9708), .A(n9582), .ZN(n5991) );
  OAI21_X1 U7542 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9584), .A(n5991), .ZN(
        n9590) );
  NAND2_X1 U7543 ( .A1(n9591), .A2(n9590), .ZN(n9589) );
  OAI21_X1 U7544 ( .B1(n9599), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9589), .ZN(
        n5994) );
  INV_X1 U7545 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5992) );
  MUX2_X1 U7546 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n5992), .S(n6687), .Z(n5993)
         );
  NAND2_X1 U7547 ( .A1(n5994), .A2(n5993), .ZN(n6163) );
  OAI21_X1 U7548 ( .B1(n5994), .B2(n5993), .A(n6163), .ZN(n6008) );
  INV_X1 U7549 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U7550 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6767) );
  INV_X1 U7551 ( .A(n6767), .ZN(n5995) );
  AOI21_X1 U7552 ( .B1(n9635), .B2(n6687), .A(n5995), .ZN(n6005) );
  INV_X1 U7553 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5996) );
  XNOR2_X1 U7554 ( .A(n6687), .B(n5996), .ZN(n6003) );
  NAND2_X1 U7555 ( .A1(n9599), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6001) );
  INV_X1 U7556 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5998) );
  MUX2_X1 U7557 ( .A(n5998), .B(P1_REG2_REG_6__SCAN_IN), .S(n6349), .Z(n6016)
         );
  NOR2_X1 U7558 ( .A1(n6017), .A2(n6016), .ZN(n6015) );
  INV_X1 U7559 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5999) );
  MUX2_X1 U7560 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n5999), .S(n9562), .Z(n9563)
         );
  NAND2_X1 U7561 ( .A1(n9582), .A2(n6576), .ZN(n9575) );
  INV_X1 U7562 ( .A(n9582), .ZN(n9580) );
  OAI21_X1 U7563 ( .B1(n9599), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6001), .ZN(
        n9596) );
  NOR2_X1 U7564 ( .A1(n9597), .A2(n9596), .ZN(n9595) );
  INV_X1 U7565 ( .A(n9595), .ZN(n6000) );
  OAI211_X1 U7566 ( .C1(n6003), .C2(n6002), .A(n9623), .B(n4505), .ZN(n6004)
         );
  OAI211_X1 U7567 ( .C1(n6006), .C2(n9627), .A(n6005), .B(n6004), .ZN(n6007)
         );
  AOI21_X1 U7568 ( .B1(n6008), .B2(n9641), .A(n6007), .ZN(n6009) );
  INV_X1 U7569 ( .A(n6009), .ZN(P1_U3251) );
  INV_X1 U7570 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6022) );
  OAI21_X1 U7571 ( .B1(n6012), .B2(n6011), .A(n6010), .ZN(n6020) );
  NAND2_X1 U7572 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3084), .ZN(n6013) );
  OAI21_X1 U7573 ( .B1(n9069), .B2(n6014), .A(n6013), .ZN(n6019) );
  AOI211_X1 U7574 ( .C1(n6017), .C2(n6016), .A(n6015), .B(n9629), .ZN(n6018)
         );
  AOI211_X1 U7575 ( .C1(n9641), .C2(n6020), .A(n6019), .B(n6018), .ZN(n6021)
         );
  OAI21_X1 U7576 ( .B1(n9627), .B2(n6022), .A(n6021), .ZN(P1_U3247) );
  INV_X1 U7577 ( .A(n6778), .ZN(n6044) );
  NAND2_X1 U7578 ( .A1(n6137), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6062) );
  XNOR2_X1 U7579 ( .A(n6062), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6779) );
  AOI22_X1 U7580 ( .A1(n6779), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9421), .ZN(n6024) );
  OAI21_X1 U7581 ( .B1(n6044), .B2(n9424), .A(n6024), .ZN(P1_U3341) );
  NAND2_X1 U7582 ( .A1(n9697), .A2(n7630), .ZN(n6028) );
  INV_X1 U7583 ( .A(n6025), .ZN(n6026) );
  NOR2_X1 U7584 ( .A1(n6030), .A2(n6029), .ZN(n6031) );
  INV_X2 U7585 ( .A(n9698), .ZN(n9671) );
  INV_X1 U7586 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6036) );
  INV_X1 U7587 ( .A(n6057), .ZN(n6188) );
  NOR2_X1 U7588 ( .A1(n6188), .A2(n6179), .ZN(n7398) );
  NOR2_X1 U7589 ( .A1(n7398), .A2(n6187), .ZN(n7475) );
  NOR3_X1 U7590 ( .A1(n7475), .A2(n6032), .A3(n7644), .ZN(n6033) );
  AOI21_X1 U7591 ( .B1(n9293), .B2(n9055), .A(n6033), .ZN(n6182) );
  OAI21_X1 U7592 ( .B1(n6194), .B2(n6034), .A(n6182), .ZN(n6041) );
  NAND2_X1 U7593 ( .A1(n6041), .A2(n9671), .ZN(n6035) );
  OAI21_X1 U7594 ( .B1(n9671), .B2(n6036), .A(n6035), .ZN(P1_U3454) );
  NOR2_X1 U7595 ( .A1(n6038), .A2(n6037), .ZN(n6039) );
  INV_X2 U7596 ( .A(n9707), .ZN(n9702) );
  NAND2_X1 U7597 ( .A1(n6041), .A2(n9702), .ZN(n6042) );
  OAI21_X1 U7598 ( .B1(n9702), .B2(n6043), .A(n6042), .ZN(P1_U3523) );
  INV_X1 U7599 ( .A(n8122), .ZN(n8063) );
  OAI222_X1 U7600 ( .A1(n8237), .A2(n10001), .B1(n8236), .B2(n6044), .C1(
        P2_U3152), .C2(n8063), .ZN(P2_U3346) );
  NAND2_X1 U7601 ( .A1(n9055), .A2(n6394), .ZN(n6046) );
  NAND2_X1 U7602 ( .A1(n7400), .A2(n6077), .ZN(n6045) );
  NAND2_X1 U7603 ( .A1(n6046), .A2(n6045), .ZN(n6047) );
  INV_X1 U7604 ( .A(n6052), .ZN(n6051) );
  NAND2_X1 U7605 ( .A1(n6050), .A2(n6049), .ZN(n6053) );
  NAND2_X1 U7606 ( .A1(n6053), .A2(n6052), .ZN(n6076) );
  NAND2_X1 U7607 ( .A1(n6075), .A2(n6076), .ZN(n6054) );
  AOI22_X1 U7608 ( .A1(n9055), .A2(n8007), .B1(n8004), .B2(n7400), .ZN(n6074)
         );
  XNOR2_X1 U7609 ( .A(n6054), .B(n6074), .ZN(n6060) );
  AOI22_X1 U7610 ( .A1(n6055), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n7400), .B2(
        n9036), .ZN(n6059) );
  NOR2_X2 U7611 ( .A1(n6056), .A2(n9536), .ZN(n8978) );
  INV_X1 U7612 ( .A(n9009), .ZN(n9030) );
  AOI22_X1 U7613 ( .A1(n8978), .A2(n6057), .B1(n9030), .B2(n9054), .ZN(n6058)
         );
  OAI211_X1 U7614 ( .C1(n6060), .C2(n9038), .A(n6059), .B(n6058), .ZN(P1_U3220) );
  INV_X1 U7615 ( .A(n6929), .ZN(n6073) );
  NAND2_X1 U7616 ( .A1(n6062), .A2(n6061), .ZN(n6063) );
  NAND2_X1 U7617 ( .A1(n6063), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6064) );
  XNOR2_X1 U7618 ( .A(n6064), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6930) );
  AOI22_X1 U7619 ( .A1(n6930), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9421), .ZN(n6065) );
  OAI21_X1 U7620 ( .B1(n6073), .B2(n9424), .A(n6065), .ZN(P1_U3340) );
  INV_X1 U7621 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7622 ( .A1(n4409), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7623 ( .A1(n5393), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7624 ( .A1(n4423), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6066) );
  INV_X1 U7625 ( .A(n7876), .ZN(n6069) );
  NAND2_X1 U7626 ( .A1(n6069), .A2(P2_U3966), .ZN(n6070) );
  OAI21_X1 U7627 ( .B1(P2_U3966), .B2(n6071), .A(n6070), .ZN(P2_U3583) );
  NAND2_X1 U7628 ( .A1(n6275), .A2(P2_U3966), .ZN(n6072) );
  OAI21_X1 U7629 ( .B1(P2_U3966), .B2(n5001), .A(n6072), .ZN(P2_U3552) );
  INV_X1 U7630 ( .A(n8123), .ZN(n8150) );
  OAI222_X1 U7631 ( .A1(n8237), .A2(n10081), .B1(n8236), .B2(n6073), .C1(n8150), .C2(P2_U3152), .ZN(P2_U3345) );
  NAND2_X1 U7632 ( .A1(n9054), .A2(n6394), .ZN(n6079) );
  NAND2_X1 U7633 ( .A1(n7404), .A2(n6077), .ZN(n6078) );
  NAND2_X1 U7634 ( .A1(n6079), .A2(n6078), .ZN(n6080) );
  XNOR2_X1 U7635 ( .A(n6080), .B(n7998), .ZN(n6081) );
  AOI22_X1 U7636 ( .A1(n9054), .A2(n8007), .B1(n8004), .B2(n7404), .ZN(n6082)
         );
  NAND2_X1 U7637 ( .A1(n6081), .A2(n6082), .ZN(n6086) );
  INV_X1 U7638 ( .A(n6081), .ZN(n6084) );
  INV_X1 U7639 ( .A(n6082), .ZN(n6083) );
  NAND2_X1 U7640 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  AND2_X1 U7641 ( .A1(n6086), .A2(n6085), .ZN(n6149) );
  NAND2_X1 U7642 ( .A1(n6148), .A2(n6149), .ZN(n6147) );
  NAND2_X1 U7643 ( .A1(n6147), .A2(n6086), .ZN(n8927) );
  NAND2_X1 U7644 ( .A1(n9053), .A2(n6394), .ZN(n6091) );
  NAND2_X1 U7645 ( .A1(n7382), .A2(n6087), .ZN(n6088) );
  NAND2_X1 U7646 ( .A1(n8930), .A2(n6077), .ZN(n6090) );
  NAND2_X1 U7647 ( .A1(n6091), .A2(n6090), .ZN(n6092) );
  XNOR2_X1 U7648 ( .A(n6092), .B(n8005), .ZN(n6093) );
  AOI22_X1 U7649 ( .A1(n9053), .A2(n8007), .B1(n8004), .B2(n8930), .ZN(n6094)
         );
  XNOR2_X1 U7650 ( .A(n6093), .B(n6094), .ZN(n8928) );
  NAND2_X1 U7651 ( .A1(n8927), .A2(n8928), .ZN(n8926) );
  INV_X1 U7652 ( .A(n6093), .ZN(n6095) );
  NAND2_X1 U7653 ( .A1(n6095), .A2(n6094), .ZN(n6096) );
  NAND2_X1 U7654 ( .A1(n4414), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7655 ( .A1(n7324), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7656 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6117) );
  OAI21_X1 U7657 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n6117), .ZN(n6240) );
  INV_X1 U7658 ( .A(n6240), .ZN(n6131) );
  NAND2_X1 U7659 ( .A1(n7459), .A2(n6131), .ZN(n6099) );
  NAND2_X1 U7660 ( .A1(n4417), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6098) );
  NAND4_X1 U7661 ( .A1(n6101), .A2(n6100), .A3(n6099), .A4(n6098), .ZN(n9052)
         );
  NAND2_X1 U7662 ( .A1(n9052), .A2(n6394), .ZN(n6107) );
  OR2_X1 U7663 ( .A1(n6644), .A2(n6102), .ZN(n6104) );
  NAND2_X1 U7664 ( .A1(n7450), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6103) );
  OAI211_X1 U7665 ( .C1(n6105), .C2(n9545), .A(n6104), .B(n6103), .ZN(n6239)
         );
  NAND2_X1 U7666 ( .A1(n6239), .A2(n7995), .ZN(n6106) );
  NAND2_X1 U7667 ( .A1(n6107), .A2(n6106), .ZN(n6108) );
  XNOR2_X1 U7668 ( .A(n6108), .B(n7998), .ZN(n6109) );
  AOI22_X1 U7669 ( .A1(n9052), .A2(n8007), .B1(n8004), .B2(n6239), .ZN(n6110)
         );
  AND2_X1 U7670 ( .A1(n6109), .A2(n6110), .ZN(n6294) );
  INV_X1 U7671 ( .A(n6294), .ZN(n6113) );
  INV_X1 U7672 ( .A(n6109), .ZN(n6112) );
  INV_X1 U7673 ( .A(n6110), .ZN(n6111) );
  NAND2_X1 U7674 ( .A1(n6112), .A2(n6111), .ZN(n6295) );
  NAND2_X1 U7675 ( .A1(n6113), .A2(n6295), .ZN(n6114) );
  XNOR2_X1 U7676 ( .A(n6293), .B(n6114), .ZN(n6136) );
  NAND2_X1 U7677 ( .A1(n4414), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6122) );
  OR2_X1 U7678 ( .A1(n7456), .A2(n5933), .ZN(n6121) );
  NAND2_X1 U7679 ( .A1(n7324), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6120) );
  INV_X1 U7680 ( .A(n6117), .ZN(n6115) );
  INV_X1 U7681 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U7682 ( .A1(n6117), .A2(n6116), .ZN(n6118) );
  AND2_X1 U7683 ( .A1(n6361), .A2(n6118), .ZN(n6457) );
  NAND2_X1 U7684 ( .A1(n7459), .A2(n6457), .ZN(n6119) );
  NAND4_X1 U7685 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .ZN(n9051)
         );
  NAND3_X1 U7686 ( .A1(n6124), .A2(n6123), .A3(n6998), .ZN(n6125) );
  AOI21_X1 U7687 ( .B1(n6128), .B2(n9691), .A(n6125), .ZN(n6126) );
  OR2_X1 U7688 ( .A1(n6126), .A2(P1_U3084), .ZN(n6130) );
  NAND3_X1 U7689 ( .A1(n6128), .A2(n7641), .A3(n6127), .ZN(n6129) );
  NAND2_X1 U7690 ( .A1(n6130), .A2(n6129), .ZN(n9029) );
  AOI22_X1 U7691 ( .A1(n9030), .A2(n9051), .B1(n6131), .B2(n9029), .ZN(n6135)
         );
  NAND2_X1 U7692 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9560) );
  INV_X1 U7693 ( .A(n9560), .ZN(n6133) );
  INV_X1 U7694 ( .A(n6239), .ZN(n9679) );
  NOR2_X1 U7695 ( .A1(n9024), .A2(n9679), .ZN(n6132) );
  AOI211_X1 U7696 ( .C1(n8978), .C2(n9053), .A(n6133), .B(n6132), .ZN(n6134)
         );
  OAI211_X1 U7697 ( .C1(n6136), .C2(n9038), .A(n6135), .B(n6134), .ZN(P1_U3228) );
  INV_X1 U7698 ( .A(n7010), .ZN(n6140) );
  INV_X1 U7699 ( .A(n8124), .ZN(n8141) );
  OAI222_X1 U7700 ( .A1(n8881), .A2(n10140), .B1(n8236), .B2(n6140), .C1(n8141), .C2(P2_U3152), .ZN(P2_U3344) );
  OR3_X1 U7701 ( .A1(n6137), .A2(P1_IR_REG_13__SCAN_IN), .A3(
        P1_IR_REG_12__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7702 ( .A1(n6138), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6139) );
  XNOR2_X1 U7703 ( .A(n6139), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9615) );
  INV_X1 U7704 ( .A(n9615), .ZN(n6724) );
  OAI222_X1 U7705 ( .A1(n8231), .A2(n6141), .B1(n9424), .B2(n6140), .C1(n6724), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  NAND2_X1 U7706 ( .A1(n7869), .A2(n6512), .ZN(n6146) );
  INV_X1 U7707 ( .A(n7867), .ZN(n7871) );
  NAND2_X1 U7708 ( .A1(n9753), .A2(n7871), .ZN(n6144) );
  NAND2_X1 U7709 ( .A1(n6144), .A2(n6143), .ZN(n6145) );
  NOR2_X1 U7710 ( .A1(n9875), .A2(P2_U3966), .ZN(P2_U3151) );
  OAI21_X1 U7711 ( .B1(n6149), .B2(n6148), .A(n6147), .ZN(n6154) );
  OAI22_X1 U7712 ( .A1(n6151), .A2(n6150), .B1(n9024), .B2(n9674), .ZN(n6153)
         );
  OAI22_X1 U7713 ( .A1(n9034), .A2(n7401), .B1(n6226), .B2(n9009), .ZN(n6152)
         );
  AOI211_X1 U7714 ( .C1(n6154), .C2(n9015), .A(n6153), .B(n6152), .ZN(n6155)
         );
  INV_X1 U7715 ( .A(n6155), .ZN(P1_U3235) );
  NAND2_X1 U7716 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n8392), .ZN(n6156) );
  OAI21_X1 U7717 ( .B1(n8669), .B2(n8392), .A(n6156), .ZN(P2_U3570) );
  NAND2_X1 U7718 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n8392), .ZN(n6157) );
  OAI21_X1 U7719 ( .B1(n8591), .B2(n8392), .A(n6157), .ZN(P2_U3575) );
  NAND2_X1 U7720 ( .A1(n5248), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7721 ( .A1(n4423), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6159) );
  NAND2_X1 U7722 ( .A1(n5393), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6158) );
  AND3_X1 U7723 ( .A1(n6160), .A2(n6159), .A3(n6158), .ZN(n8492) );
  NAND2_X1 U7724 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n8392), .ZN(n6161) );
  OAI21_X1 U7725 ( .B1(n8492), .B2(n8392), .A(n6161), .ZN(P2_U3582) );
  INV_X1 U7726 ( .A(n9627), .ZN(n9640) );
  INV_X1 U7727 ( .A(n6779), .ZN(n6169) );
  INV_X1 U7728 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6703) );
  NOR2_X1 U7729 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6703), .ZN(n6808) );
  INV_X1 U7730 ( .A(n6808), .ZN(n6168) );
  INV_X1 U7731 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6162) );
  MUX2_X1 U7732 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6162), .S(n6779), .Z(n6165)
         );
  INV_X1 U7733 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6866) );
  AOI22_X1 U7734 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n9603), .B1(n6171), .B2(
        n6866), .ZN(n9605) );
  OAI21_X1 U7735 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n6687), .A(n6163), .ZN(
        n9606) );
  NAND2_X1 U7736 ( .A1(n9605), .A2(n9606), .ZN(n9604) );
  OAI21_X1 U7737 ( .B1(n6165), .B2(n6164), .A(n6258), .ZN(n6166) );
  NAND2_X1 U7738 ( .A1(n9641), .A2(n6166), .ZN(n6167) );
  OAI211_X1 U7739 ( .C1(n9069), .C2(n6169), .A(n6168), .B(n6167), .ZN(n6176)
         );
  INV_X1 U7740 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6170) );
  AOI22_X1 U7741 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n9603), .B1(n6171), .B2(
        n6170), .ZN(n9608) );
  OAI21_X1 U7742 ( .B1(n9603), .B2(P1_REG2_REG_11__SCAN_IN), .A(n9607), .ZN(
        n6174) );
  NAND2_X1 U7743 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6779), .ZN(n6172) );
  OAI21_X1 U7744 ( .B1(n6779), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6172), .ZN(
        n6173) );
  NOR2_X1 U7745 ( .A1(n6173), .A2(n6174), .ZN(n6252) );
  AOI211_X1 U7746 ( .C1(n6174), .C2(n6173), .A(n6252), .B(n9629), .ZN(n6175)
         );
  AOI211_X1 U7747 ( .C1(P1_ADDR_REG_12__SCAN_IN), .C2(n9640), .A(n6176), .B(
        n6175), .ZN(n6177) );
  INV_X1 U7748 ( .A(n6177), .ZN(P1_U3253) );
  NAND2_X1 U7749 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8392), .ZN(n6178) );
  OAI21_X1 U7750 ( .B1(n7668), .B2(n8392), .A(n6178), .ZN(P2_U3581) );
  AOI22_X1 U7751 ( .A1(n4419), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9652), .ZN(n6181) );
  OAI21_X1 U7752 ( .B1(n9650), .B2(n9469), .A(n6179), .ZN(n6180) );
  OAI211_X1 U7753 ( .C1(n6182), .C2(n4419), .A(n6181), .B(n6180), .ZN(P1_U3291) );
  OAI21_X1 U7754 ( .B1(n6185), .B2(n6184), .A(n6183), .ZN(n9665) );
  OAI21_X1 U7755 ( .B1(n7473), .B2(n6187), .A(n6186), .ZN(n6190) );
  INV_X1 U7756 ( .A(n9054), .ZN(n7405) );
  OAI22_X1 U7757 ( .A1(n6188), .A2(n9464), .B1(n7405), .B2(n9462), .ZN(n6189)
         );
  AOI21_X1 U7758 ( .B1(n6190), .B2(n9296), .A(n6189), .ZN(n6191) );
  OAI21_X1 U7759 ( .B1(n6574), .B2(n9665), .A(n6191), .ZN(n9667) );
  INV_X1 U7760 ( .A(n6192), .ZN(n6193) );
  OAI211_X1 U7761 ( .C1(n4636), .C2(n6194), .A(n6193), .B(n9471), .ZN(n9666)
         );
  INV_X1 U7762 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6195) );
  OAI22_X1 U7763 ( .A1(n9666), .A2(n7661), .B1(n9258), .B2(n6195), .ZN(n6196)
         );
  OAI21_X1 U7764 ( .B1(n9667), .B2(n6196), .A(n9281), .ZN(n6198) );
  AOI22_X1 U7765 ( .A1(n9469), .A2(n7400), .B1(n4419), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6197) );
  OAI211_X1 U7766 ( .C1(n9665), .C2(n6583), .A(n6198), .B(n6197), .ZN(P1_U3290) );
  INV_X1 U7767 ( .A(n7367), .ZN(n6207) );
  AOI22_X1 U7768 ( .A1(n8439), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n7143), .ZN(n6199) );
  OAI21_X1 U7769 ( .B1(n6207), .B2(n8236), .A(n6199), .ZN(P2_U3342) );
  INV_X1 U7770 ( .A(n7379), .ZN(n6203) );
  NAND2_X1 U7771 ( .A1(n6200), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6201) );
  XNOR2_X1 U7772 ( .A(n6201), .B(n5734), .ZN(n7380) );
  OAI222_X1 U7773 ( .A1(n8231), .A2(n6202), .B1(n9424), .B2(n6203), .C1(
        P1_U3084), .C2(n7380), .ZN(P1_U3338) );
  INV_X1 U7774 ( .A(n8422), .ZN(n8413) );
  OAI222_X1 U7775 ( .A1(n8881), .A2(n6204), .B1(n8236), .B2(n6203), .C1(
        P2_U3152), .C2(n8413), .ZN(P2_U3343) );
  NAND2_X1 U7776 ( .A1(n6205), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6222) );
  XNOR2_X1 U7777 ( .A(n6222), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7655) );
  INV_X1 U7778 ( .A(n7655), .ZN(n6206) );
  OAI222_X1 U7779 ( .A1(n8231), .A2(n10026), .B1(n9424), .B2(n6207), .C1(n6206), .C2(P1_U3084), .ZN(P1_U3337) );
  NAND2_X1 U7780 ( .A1(n7405), .A2(n9674), .ZN(n6208) );
  NAND2_X1 U7781 ( .A1(n6210), .A2(n6231), .ZN(n6228) );
  OAI21_X1 U7782 ( .B1(n6210), .B2(n6231), .A(n6228), .ZN(n6250) );
  OAI21_X1 U7783 ( .B1(n4508), .B2(n6225), .A(n6238), .ZN(n6246) );
  OAI22_X1 U7784 ( .A1(n6246), .A2(n9692), .B1(n6225), .B2(n9691), .ZN(n6215)
         );
  NAND2_X1 U7785 ( .A1(n7407), .A2(n7472), .ZN(n6211) );
  NAND2_X1 U7786 ( .A1(n7405), .A2(n7404), .ZN(n7402) );
  XNOR2_X1 U7787 ( .A(n6232), .B(n6231), .ZN(n6214) );
  NAND2_X1 U7788 ( .A1(n6250), .A2(n9648), .ZN(n6213) );
  AOI22_X1 U7789 ( .A1(n9291), .A2(n9054), .B1(n9052), .B2(n9293), .ZN(n6212)
         );
  OAI211_X1 U7790 ( .C1(n9459), .C2(n6214), .A(n6213), .B(n6212), .ZN(n6247)
         );
  AOI211_X1 U7791 ( .C1(n9697), .C2(n6250), .A(n6215), .B(n6247), .ZN(n6218)
         );
  OR2_X1 U7792 ( .A1(n6218), .A2(n9707), .ZN(n6216) );
  OAI21_X1 U7793 ( .B1(n9702), .B2(n6217), .A(n6216), .ZN(P1_U3526) );
  INV_X1 U7794 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6220) );
  OR2_X1 U7795 ( .A1(n6218), .A2(n9698), .ZN(n6219) );
  OAI21_X1 U7796 ( .B1(n9671), .B2(n6220), .A(n6219), .ZN(P1_U3463) );
  INV_X1 U7797 ( .A(n7310), .ZN(n6316) );
  NAND2_X1 U7798 ( .A1(n6222), .A2(n6221), .ZN(n6223) );
  NAND2_X1 U7799 ( .A1(n6223), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6480) );
  XNOR2_X1 U7800 ( .A(n6480), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9059) );
  AOI22_X1 U7801 ( .A1(n9059), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9421), .ZN(n6224) );
  OAI21_X1 U7802 ( .B1(n6316), .B2(n9424), .A(n6224), .ZN(P1_U3336) );
  NAND2_X1 U7803 ( .A1(n6226), .A2(n6225), .ZN(n6227) );
  NAND2_X1 U7804 ( .A1(n6228), .A2(n6227), .ZN(n6229) );
  INV_X1 U7805 ( .A(n9052), .ZN(n6341) );
  NAND2_X1 U7806 ( .A1(n6341), .A2(n6239), .ZN(n6413) );
  NAND2_X1 U7807 ( .A1(n9052), .A2(n9679), .ZN(n7499) );
  NAND2_X1 U7808 ( .A1(n6413), .A2(n7499), .ZN(n7477) );
  NAND2_X1 U7809 ( .A1(n6229), .A2(n7477), .ZN(n6343) );
  OR2_X1 U7810 ( .A1(n6229), .A2(n7477), .ZN(n6230) );
  NAND2_X1 U7811 ( .A1(n6343), .A2(n6230), .ZN(n9683) );
  INV_X1 U7812 ( .A(n9683), .ZN(n6244) );
  INV_X1 U7813 ( .A(n6231), .ZN(n7474) );
  NAND2_X1 U7814 ( .A1(n6232), .A2(n7474), .ZN(n6233) );
  NAND2_X1 U7815 ( .A1(n6233), .A2(n7498), .ZN(n6373) );
  XNOR2_X1 U7816 ( .A(n6373), .B(n7477), .ZN(n6236) );
  NAND2_X1 U7817 ( .A1(n9683), .A2(n9648), .ZN(n6235) );
  AOI22_X1 U7818 ( .A1(n9291), .A2(n9053), .B1(n9051), .B2(n9293), .ZN(n6234)
         );
  OAI211_X1 U7819 ( .C1(n9459), .C2(n6236), .A(n6235), .B(n6234), .ZN(n9681)
         );
  MUX2_X1 U7820 ( .A(n9681), .B(P1_REG2_REG_4__SCAN_IN), .S(n4419), .Z(n6237)
         );
  INV_X1 U7821 ( .A(n6237), .ZN(n6243) );
  AOI21_X1 U7822 ( .B1(n6239), .B2(n6238), .A(n6410), .ZN(n9678) );
  OAI22_X1 U7823 ( .A1(n9656), .A2(n9679), .B1(n6240), .B2(n9258), .ZN(n6241)
         );
  AOI21_X1 U7824 ( .B1(n9678), .B2(n9650), .A(n6241), .ZN(n6242) );
  OAI211_X1 U7825 ( .C1(n6244), .C2(n6583), .A(n6243), .B(n6242), .ZN(P1_U3287) );
  INV_X1 U7826 ( .A(n6583), .ZN(n9659) );
  AOI22_X1 U7827 ( .A1(n9469), .A2(n8930), .B1(n5810), .B2(n9652), .ZN(n6245)
         );
  OAI21_X1 U7828 ( .B1(n6591), .B2(n6246), .A(n6245), .ZN(n6249) );
  MUX2_X1 U7829 ( .A(n6247), .B(P1_REG2_REG_3__SCAN_IN), .S(n4419), .Z(n6248)
         );
  AOI211_X1 U7830 ( .C1(n9659), .C2(n6250), .A(n6249), .B(n6248), .ZN(n6251)
         );
  INV_X1 U7831 ( .A(n6251), .ZN(P1_U3288) );
  INV_X1 U7832 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6264) );
  NAND2_X1 U7833 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n6930), .ZN(n6253) );
  OAI21_X1 U7834 ( .B1(n6930), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6253), .ZN(
        n6254) );
  AOI211_X1 U7835 ( .C1(n6255), .C2(n6254), .A(n6719), .B(n9629), .ZN(n6256)
         );
  AOI21_X1 U7836 ( .B1(n9635), .B2(n6930), .A(n6256), .ZN(n6263) );
  INV_X1 U7837 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6257) );
  MUX2_X1 U7838 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6257), .S(n6930), .Z(n6260)
         );
  OAI21_X1 U7839 ( .B1(n6779), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6258), .ZN(
        n6259) );
  OAI21_X1 U7840 ( .B1(n6260), .B2(n6259), .A(n6725), .ZN(n6261) );
  AND2_X1 U7841 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6965) );
  AOI21_X1 U7842 ( .B1(n9641), .B2(n6261), .A(n6965), .ZN(n6262) );
  OAI211_X1 U7843 ( .C1(n9627), .C2(n6264), .A(n6263), .B(n6262), .ZN(P1_U3254) );
  INV_X1 U7844 ( .A(n6830), .ZN(n6269) );
  NOR2_X1 U7845 ( .A1(n9753), .A2(n6265), .ZN(n6267) );
  INV_X1 U7846 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7847 ( .A1(n6275), .A2(n6869), .ZN(n6272) );
  OAI21_X1 U7848 ( .B1(n7688), .B2(n6272), .A(n6318), .ZN(n8750) );
  INV_X1 U7849 ( .A(n8750), .ZN(n6286) );
  NAND2_X1 U7850 ( .A1(n5702), .A2(n6834), .ZN(n6273) );
  NAND3_X1 U7851 ( .A1(n6274), .A2(n8546), .A3(n6273), .ZN(n9740) );
  NAND2_X1 U7852 ( .A1(n9740), .A2(n9787), .ZN(n9822) );
  INV_X1 U7853 ( .A(n6275), .ZN(n6276) );
  XNOR2_X1 U7854 ( .A(n6322), .B(n7688), .ZN(n6277) );
  INV_X1 U7855 ( .A(n7860), .ZN(n7709) );
  NAND2_X1 U7856 ( .A1(n7709), .A2(n7728), .ZN(n7682) );
  NAND2_X1 U7857 ( .A1(n6277), .A2(n9737), .ZN(n6281) );
  OR2_X1 U7858 ( .A1(n6424), .A2(n9732), .ZN(n6279) );
  NAND2_X1 U7859 ( .A1(n6275), .A2(n8729), .ZN(n6278) );
  NAND2_X1 U7860 ( .A1(n6279), .A2(n6278), .ZN(n7891) );
  INV_X1 U7861 ( .A(n7891), .ZN(n6280) );
  NAND2_X1 U7862 ( .A1(n6281), .A2(n6280), .ZN(n8753) );
  INV_X1 U7863 ( .A(n8753), .ZN(n6285) );
  AOI21_X1 U7864 ( .B1(n6270), .B2(n6869), .A(n9820), .ZN(n6283) );
  INV_X1 U7865 ( .A(n6869), .ZN(n9762) );
  NAND2_X1 U7866 ( .A1(n6282), .A2(n9762), .ZN(n6325) );
  AND2_X1 U7867 ( .A1(n6283), .A2(n6325), .ZN(n8755) );
  AOI21_X1 U7868 ( .B1(n9815), .B2(n6270), .A(n8755), .ZN(n6284) );
  OAI211_X1 U7869 ( .C1(n6286), .C2(n9764), .A(n6285), .B(n6284), .ZN(n6291)
         );
  NAND2_X1 U7870 ( .A1(n6291), .A2(n9826), .ZN(n6287) );
  OAI21_X1 U7871 ( .B1(n9826), .B2(n6288), .A(n6287), .ZN(P2_U3454) );
  NAND2_X1 U7872 ( .A1(n6291), .A2(n9839), .ZN(n6292) );
  OAI21_X1 U7873 ( .B1(n9839), .B2(n6521), .A(n6292), .ZN(P2_U3521) );
  NAND2_X1 U7874 ( .A1(n9051), .A2(n6394), .ZN(n6301) );
  OR2_X1 U7875 ( .A1(n6296), .A2(n6644), .ZN(n6299) );
  AOI22_X1 U7876 ( .A1(n7450), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7382), .B2(
        n6297), .ZN(n6298) );
  NAND2_X1 U7877 ( .A1(n6299), .A2(n6298), .ZN(n6458) );
  NAND2_X1 U7878 ( .A1(n6458), .A2(n7995), .ZN(n6300) );
  NAND2_X1 U7879 ( .A1(n6301), .A2(n6300), .ZN(n6302) );
  XNOR2_X1 U7880 ( .A(n6302), .B(n7998), .ZN(n6396) );
  XNOR2_X1 U7881 ( .A(n6395), .B(n6396), .ZN(n6306) );
  NAND2_X1 U7882 ( .A1(n9051), .A2(n8007), .ZN(n6304) );
  NAND2_X1 U7883 ( .A1(n6458), .A2(n6394), .ZN(n6303) );
  AND2_X1 U7884 ( .A1(n6304), .A2(n6303), .ZN(n6305) );
  NAND2_X1 U7885 ( .A1(n6306), .A2(n6305), .ZN(n6398) );
  OAI21_X1 U7886 ( .B1(n6306), .B2(n6305), .A(n6398), .ZN(n6314) );
  INV_X1 U7887 ( .A(n6458), .ZN(n6412) );
  AOI22_X1 U7888 ( .A1(n8978), .A2(n9052), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3084), .ZN(n6312) );
  NAND2_X1 U7889 ( .A1(n7324), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U7890 ( .A1(n4416), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6309) );
  XNOR2_X1 U7891 ( .A(n6361), .B(P1_REG3_REG_6__SCAN_IN), .ZN(n6588) );
  NAND2_X1 U7892 ( .A1(n7459), .A2(n6588), .ZN(n6308) );
  NAND2_X1 U7893 ( .A1(n4414), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6307) );
  NAND4_X1 U7894 ( .A1(n6310), .A2(n6309), .A3(n6308), .A4(n6307), .ZN(n9050)
         );
  AOI22_X1 U7895 ( .A1(n9030), .A2(n9050), .B1(n6457), .B2(n9029), .ZN(n6311)
         );
  OAI211_X1 U7896 ( .C1(n6412), .C2(n9024), .A(n6312), .B(n6311), .ZN(n6313)
         );
  AOI21_X1 U7897 ( .B1(n6314), .B2(n9015), .A(n6313), .ZN(n6315) );
  INV_X1 U7898 ( .A(n6315), .ZN(P1_U3225) );
  INV_X1 U7899 ( .A(n8455), .ZN(n8438) );
  OAI222_X1 U7900 ( .A1(n8881), .A2(n10084), .B1(n8236), .B2(n6316), .C1(n8438), .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U7901 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6519) );
  NAND2_X1 U7902 ( .A1(n6271), .A2(n6282), .ZN(n6317) );
  NAND2_X1 U7903 ( .A1(n6321), .A2(n6320), .ZN(n6426) );
  OAI21_X1 U7904 ( .B1(n6321), .B2(n6320), .A(n6426), .ZN(n8743) );
  INV_X1 U7905 ( .A(n8743), .ZN(n6329) );
  OAI21_X1 U7906 ( .B1(n6323), .B2(n7687), .A(n6428), .ZN(n6324) );
  OAI22_X1 U7907 ( .A1(n6271), .A2(n9734), .B1(n6487), .B2(n9732), .ZN(n7879)
         );
  AOI21_X1 U7908 ( .B1(n6324), .B2(n9737), .A(n7879), .ZN(n8745) );
  NAND2_X1 U7909 ( .A1(n6325), .A2(n4411), .ZN(n6326) );
  NAND2_X1 U7910 ( .A1(n6326), .A2(n9774), .ZN(n6327) );
  NOR2_X1 U7911 ( .A1(n6431), .A2(n6327), .ZN(n8744) );
  AOI21_X1 U7912 ( .B1(n9815), .B2(n4411), .A(n8744), .ZN(n6328) );
  OAI211_X1 U7913 ( .C1(n6329), .C2(n9764), .A(n8745), .B(n6328), .ZN(n6331)
         );
  NAND2_X1 U7914 ( .A1(n6331), .A2(n9839), .ZN(n6330) );
  OAI21_X1 U7915 ( .B1(n9839), .B2(n6519), .A(n6330), .ZN(P2_U3522) );
  INV_X1 U7916 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6333) );
  NAND2_X1 U7917 ( .A1(n6331), .A2(n9826), .ZN(n6332) );
  OAI21_X1 U7918 ( .B1(n9826), .B2(n6333), .A(n6332), .ZN(P2_U3457) );
  XNOR2_X1 U7919 ( .A(n6335), .B(n6334), .ZN(n6340) );
  OR2_X1 U7920 ( .A1(n6872), .A2(n9732), .ZN(n6337) );
  OR2_X1 U7921 ( .A1(n6424), .A2(n9734), .ZN(n6336) );
  NAND2_X1 U7922 ( .A1(n6337), .A2(n6336), .ZN(n6429) );
  AOI22_X1 U7923 ( .A1(n8358), .A2(n6429), .B1(n8374), .B2(n4421), .ZN(n6339)
         );
  MUX2_X1 U7924 ( .A(n8368), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n6338) );
  OAI211_X1 U7925 ( .C1(n6340), .C2(n8376), .A(n6339), .B(n6338), .ZN(P2_U3220) );
  NAND2_X1 U7926 ( .A1(n6341), .A2(n9679), .ZN(n6342) );
  NAND2_X1 U7927 ( .A1(n6343), .A2(n6342), .ZN(n6408) );
  INV_X1 U7928 ( .A(n9051), .ZN(n6344) );
  NAND2_X1 U7929 ( .A1(n6344), .A2(n6458), .ZN(n7500) );
  NAND2_X1 U7930 ( .A1(n6412), .A2(n9051), .ZN(n6374) );
  NAND2_X1 U7931 ( .A1(n9051), .A2(n6458), .ZN(n6346) );
  INV_X1 U7932 ( .A(n9050), .ZN(n6352) );
  OR2_X1 U7933 ( .A1(n6347), .A2(n6644), .ZN(n6351) );
  AOI22_X1 U7934 ( .A1(n7450), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7382), .B2(
        n6349), .ZN(n6350) );
  NAND2_X1 U7935 ( .A1(n6351), .A2(n6350), .ZN(n6589) );
  OR2_X1 U7936 ( .A1(n6352), .A2(n6589), .ZN(n7413) );
  NAND2_X1 U7937 ( .A1(n6589), .A2(n6352), .ZN(n7536) );
  NAND2_X1 U7938 ( .A1(n7413), .A2(n7536), .ZN(n7535) );
  OR2_X1 U7939 ( .A1(n6589), .A2(n9050), .ZN(n6353) );
  NAND2_X1 U7940 ( .A1(n6584), .A2(n6353), .ZN(n6367) );
  OR2_X1 U7941 ( .A1(n6354), .A2(n6644), .ZN(n6356) );
  AOI22_X1 U7942 ( .A1(n7450), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7382), .B2(
        n9562), .ZN(n6355) );
  NAND2_X1 U7943 ( .A1(n6356), .A2(n6355), .ZN(n8892) );
  NAND2_X1 U7944 ( .A1(n7324), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6366) );
  OR2_X1 U7945 ( .A1(n7456), .A2(n5999), .ZN(n6365) );
  INV_X1 U7946 ( .A(n6361), .ZN(n6358) );
  NAND2_X1 U7947 ( .A1(n6358), .A2(n6357), .ZN(n6380) );
  INV_X1 U7948 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6360) );
  INV_X1 U7949 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6359) );
  OAI21_X1 U7950 ( .B1(n6361), .B2(n6360), .A(n6359), .ZN(n6362) );
  AND2_X1 U7951 ( .A1(n6380), .A2(n6362), .ZN(n8891) );
  NAND2_X1 U7952 ( .A1(n7459), .A2(n8891), .ZN(n6364) );
  NAND2_X1 U7953 ( .A1(n4414), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6363) );
  NAND4_X1 U7954 ( .A1(n6366), .A2(n6365), .A3(n6364), .A4(n6363), .ZN(n9049)
         );
  INV_X1 U7955 ( .A(n9049), .ZN(n6570) );
  OR2_X1 U7956 ( .A1(n8892), .A2(n6570), .ZN(n7537) );
  NAND2_X1 U7957 ( .A1(n8892), .A2(n6570), .ZN(n7538) );
  NAND2_X1 U7958 ( .A1(n7537), .A2(n7538), .ZN(n7479) );
  NAND2_X1 U7959 ( .A1(n6367), .A2(n7479), .ZN(n6556) );
  OAI21_X1 U7960 ( .B1(n6367), .B2(n7479), .A(n6556), .ZN(n6368) );
  INV_X1 U7961 ( .A(n6368), .ZN(n6474) );
  OR2_X1 U7962 ( .A1(n7998), .A2(n7644), .ZN(n6369) );
  AND2_X1 U7963 ( .A1(n6410), .A2(n6412), .ZN(n6587) );
  INV_X1 U7964 ( .A(n6589), .ZN(n9684) );
  NAND2_X1 U7965 ( .A1(n6587), .A2(n9684), .ZN(n6586) );
  AOI211_X1 U7966 ( .C1(n8892), .C2(n6586), .A(n9692), .B(n4730), .ZN(n6471)
         );
  INV_X1 U7967 ( .A(n8892), .ZN(n6371) );
  INV_X1 U7968 ( .A(n8891), .ZN(n6370) );
  OAI22_X1 U7969 ( .A1(n6371), .A2(n9656), .B1(n6370), .B2(n9258), .ZN(n6372)
         );
  AOI21_X1 U7970 ( .B1(n6471), .B2(n9475), .A(n6372), .ZN(n6390) );
  AND2_X1 U7971 ( .A1(n7500), .A2(n6413), .ZN(n7531) );
  INV_X1 U7972 ( .A(n6374), .ZN(n7530) );
  NAND2_X1 U7973 ( .A1(n7536), .A2(n7530), .ZN(n7503) );
  AND2_X1 U7974 ( .A1(n7503), .A2(n7413), .ZN(n6375) );
  NAND2_X1 U7975 ( .A1(n6376), .A2(n7479), .ZN(n6377) );
  NAND2_X1 U7976 ( .A1(n6562), .A2(n6377), .ZN(n6378) );
  NAND2_X1 U7977 ( .A1(n6378), .A2(n9296), .ZN(n6387) );
  NAND2_X1 U7978 ( .A1(n4414), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6385) );
  NAND2_X1 U7979 ( .A1(n7324), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6384) );
  INV_X1 U7980 ( .A(n6380), .ZN(n6379) );
  INV_X1 U7981 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6620) );
  NAND2_X1 U7982 ( .A1(n6380), .A2(n6620), .ZN(n6381) );
  AND2_X1 U7983 ( .A1(n6564), .A2(n6381), .ZN(n6575) );
  NAND2_X1 U7984 ( .A1(n7459), .A2(n6575), .ZN(n6383) );
  NAND2_X1 U7985 ( .A1(n4417), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6382) );
  NAND4_X1 U7986 ( .A1(n6385), .A2(n6384), .A3(n6383), .A4(n6382), .ZN(n9048)
         );
  AOI22_X1 U7987 ( .A1(n9291), .A2(n9050), .B1(n9048), .B2(n9293), .ZN(n6386)
         );
  NAND2_X1 U7988 ( .A1(n6387), .A2(n6386), .ZN(n6472) );
  MUX2_X1 U7989 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6472), .S(n9281), .Z(n6388)
         );
  INV_X1 U7990 ( .A(n6388), .ZN(n6389) );
  OAI211_X1 U7991 ( .C1(n6474), .C2(n9308), .A(n6390), .B(n6389), .ZN(P1_U3284) );
  NAND2_X1 U7992 ( .A1(n6589), .A2(n7995), .ZN(n6392) );
  NAND2_X1 U7993 ( .A1(n9050), .A2(n8004), .ZN(n6391) );
  NAND2_X1 U7994 ( .A1(n6392), .A2(n6391), .ZN(n6393) );
  XNOR2_X1 U7995 ( .A(n6393), .B(n8005), .ZN(n6603) );
  AOI22_X1 U7996 ( .A1(n6589), .A2(n8004), .B1(n8007), .B2(n9050), .ZN(n6604)
         );
  XNOR2_X1 U7997 ( .A(n6603), .B(n6604), .ZN(n6400) );
  OAI21_X1 U7998 ( .B1(n6400), .B2(n6399), .A(n6607), .ZN(n6404) );
  AOI22_X1 U7999 ( .A1(n8978), .A2(n9051), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3084), .ZN(n6402) );
  AOI22_X1 U8000 ( .A1(n9030), .A2(n9049), .B1(n6588), .B2(n9029), .ZN(n6401)
         );
  OAI211_X1 U8001 ( .C1(n9684), .C2(n9024), .A(n6402), .B(n6401), .ZN(n6403)
         );
  AOI21_X1 U8002 ( .B1(n6404), .B2(n9015), .A(n6403), .ZN(n6405) );
  INV_X1 U8003 ( .A(n6405), .ZN(P1_U3237) );
  INV_X1 U8004 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6420) );
  INV_X1 U8005 ( .A(n6406), .ZN(n6407) );
  AOI21_X1 U8006 ( .B1(n7476), .B2(n6408), .A(n6407), .ZN(n6464) );
  INV_X1 U8007 ( .A(n9697), .ZN(n6409) );
  INV_X1 U8008 ( .A(n9396), .ZN(n9521) );
  NOR2_X1 U8009 ( .A1(n6410), .A2(n6412), .ZN(n6411) );
  OR2_X1 U8010 ( .A1(n6587), .A2(n6411), .ZN(n6460) );
  OAI22_X1 U8011 ( .A1(n6460), .A2(n9692), .B1(n6412), .B2(n9691), .ZN(n6418)
         );
  NAND2_X1 U8012 ( .A1(n7532), .A2(n6413), .ZN(n6414) );
  NAND2_X1 U8013 ( .A1(n6414), .A2(n7476), .ZN(n6592) );
  OAI21_X1 U8014 ( .B1(n7476), .B2(n6414), .A(n6592), .ZN(n6415) );
  NAND2_X1 U8015 ( .A1(n6415), .A2(n9296), .ZN(n6417) );
  AOI22_X1 U8016 ( .A1(n9291), .A2(n9052), .B1(n9050), .B2(n9293), .ZN(n6416)
         );
  NAND2_X1 U8017 ( .A1(n6417), .A2(n6416), .ZN(n6461) );
  AOI211_X1 U8018 ( .C1(n6464), .C2(n9521), .A(n6418), .B(n6461), .ZN(n6421)
         );
  OR2_X1 U8019 ( .A1(n6421), .A2(n9698), .ZN(n6419) );
  OAI21_X1 U8020 ( .B1(n9671), .B2(n6420), .A(n6419), .ZN(P1_U3469) );
  OR2_X1 U8021 ( .A1(n6421), .A2(n9707), .ZN(n6422) );
  OAI21_X1 U8022 ( .B1(n9702), .B2(n6423), .A(n6422), .ZN(P1_U3528) );
  INV_X1 U8023 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U8024 ( .A1(n6424), .A2(n7885), .ZN(n6425) );
  NAND2_X1 U8025 ( .A1(n6426), .A2(n6425), .ZN(n6427) );
  INV_X1 U8026 ( .A(n6924), .ZN(n6486) );
  INV_X1 U8027 ( .A(n6487), .ZN(n8390) );
  NAND2_X1 U8028 ( .A1(n6486), .A2(n8390), .ZN(n7723) );
  NAND2_X1 U8029 ( .A1(n6427), .A2(n7734), .ZN(n6489) );
  OAI21_X1 U8030 ( .B1(n6427), .B2(n7734), .A(n6489), .ZN(n6925) );
  INV_X1 U8031 ( .A(n6925), .ZN(n6435) );
  NAND2_X1 U8032 ( .A1(n6428), .A2(n7742), .ZN(n6492) );
  INV_X1 U8033 ( .A(n7734), .ZN(n7686) );
  XNOR2_X1 U8034 ( .A(n6492), .B(n7686), .ZN(n6430) );
  AOI21_X1 U8035 ( .B1(n6430), .B2(n9737), .A(n6429), .ZN(n6928) );
  INV_X1 U8036 ( .A(n6431), .ZN(n6433) );
  NAND2_X1 U8037 ( .A1(n6431), .A2(n6486), .ZN(n6499) );
  INV_X1 U8038 ( .A(n6499), .ZN(n6432) );
  AOI211_X1 U8039 ( .C1(n4421), .C2(n6433), .A(n9820), .B(n6432), .ZN(n6920)
         );
  AOI21_X1 U8040 ( .B1(n9815), .B2(n4421), .A(n6920), .ZN(n6434) );
  OAI211_X1 U8041 ( .C1(n6435), .C2(n9764), .A(n6928), .B(n6434), .ZN(n6438)
         );
  NAND2_X1 U8042 ( .A1(n6438), .A2(n9839), .ZN(n6436) );
  OAI21_X1 U8043 ( .B1(n9839), .B2(n6437), .A(n6436), .ZN(P2_U3523) );
  INV_X1 U8044 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U8045 ( .A1(n6438), .A2(n9826), .ZN(n6439) );
  OAI21_X1 U8046 ( .B1(n9826), .B2(n6440), .A(n6439), .ZN(P2_U3460) );
  INV_X1 U8047 ( .A(n6441), .ZN(n6442) );
  AOI21_X1 U8048 ( .B1(n6444), .B2(n6443), .A(n6442), .ZN(n6447) );
  OAI22_X1 U8049 ( .A1(n6875), .A2(n9732), .B1(n6487), .B2(n9734), .ZN(n6497)
         );
  AOI22_X1 U8050 ( .A1(n8358), .A2(n6497), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n6446) );
  AOI22_X1 U8051 ( .A1(n6501), .A2(n8374), .B1(n8345), .B2(n6839), .ZN(n6445)
         );
  OAI211_X1 U8052 ( .C1(n6447), .C2(n8376), .A(n6446), .B(n6445), .ZN(P2_U3232) );
  OR2_X1 U8053 ( .A1(n6448), .A2(P2_U3152), .ZN(n7893) );
  INV_X1 U8054 ( .A(n7893), .ZN(n6456) );
  INV_X1 U8055 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6455) );
  INV_X1 U8056 ( .A(n8369), .ZN(n8315) );
  AOI22_X1 U8057 ( .A1(n8315), .A2(n6449), .B1(n6869), .B2(n8374), .ZN(n6454)
         );
  INV_X1 U8058 ( .A(n6322), .ZN(n6452) );
  NAND2_X1 U8059 ( .A1(n6275), .A2(n9762), .ZN(n7729) );
  INV_X1 U8060 ( .A(n7729), .ZN(n7738) );
  MUX2_X1 U8061 ( .A(n7738), .B(n6869), .S(n6450), .Z(n6451) );
  OAI21_X1 U8062 ( .B1(n6452), .B2(n6451), .A(n8353), .ZN(n6453) );
  OAI211_X1 U8063 ( .C1(n6456), .C2(n6455), .A(n6454), .B(n6453), .ZN(P2_U3234) );
  INV_X1 U8064 ( .A(n9308), .ZN(n9196) );
  AOI22_X1 U8065 ( .A1(n9469), .A2(n6458), .B1(n9652), .B2(n6457), .ZN(n6459)
         );
  OAI21_X1 U8066 ( .B1(n6460), .B2(n6591), .A(n6459), .ZN(n6463) );
  MUX2_X1 U8067 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6461), .S(n9281), .Z(n6462)
         );
  AOI211_X1 U8068 ( .C1(n9196), .C2(n6464), .A(n6463), .B(n6462), .ZN(n6465)
         );
  INV_X1 U8069 ( .A(n6465), .ZN(P1_U3286) );
  XNOR2_X1 U8070 ( .A(n6467), .B(n6466), .ZN(n6470) );
  OAI22_X1 U8071 ( .A1(n6872), .A2(n9734), .B1(n6878), .B2(n9732), .ZN(n6979)
         );
  AOI22_X1 U8072 ( .A1(n8358), .A2(n6979), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n6469) );
  AOI22_X1 U8073 ( .A1(n6987), .A2(n8374), .B1(n8345), .B2(n6981), .ZN(n6468)
         );
  OAI211_X1 U8074 ( .C1(n6470), .C2(n8376), .A(n6469), .B(n6468), .ZN(P2_U3229) );
  INV_X1 U8075 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10075) );
  AOI211_X1 U8076 ( .C1(n9392), .C2(n8892), .A(n6472), .B(n6471), .ZN(n6473)
         );
  OAI21_X1 U8077 ( .B1(n6474), .B2(n9396), .A(n6473), .ZN(n6476) );
  NAND2_X1 U8078 ( .A1(n6476), .A2(n9671), .ZN(n6475) );
  OAI21_X1 U8079 ( .B1(n9671), .B2(n10075), .A(n6475), .ZN(P1_U3475) );
  NAND2_X1 U8080 ( .A1(n6476), .A2(n9702), .ZN(n6477) );
  OAI21_X1 U8081 ( .B1(n9702), .B2(n6478), .A(n6477), .ZN(P1_U3530) );
  INV_X1 U8082 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6483) );
  INV_X1 U8083 ( .A(n7318), .ZN(n6484) );
  INV_X1 U8084 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U8085 ( .A1(n6480), .A2(n6479), .ZN(n6481) );
  NAND2_X1 U8086 ( .A1(n6481), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6482) );
  XNOR2_X1 U8087 ( .A(n6482), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9636) );
  INV_X1 U8088 ( .A(n9636), .ZN(n7653) );
  OAI222_X1 U8089 ( .A1(n8231), .A2(n6483), .B1(n9424), .B2(n6484), .C1(
        P1_U3084), .C2(n7653), .ZN(P1_U3335) );
  INV_X1 U8090 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6485) );
  INV_X1 U8091 ( .A(n8468), .ZN(n8453) );
  OAI222_X1 U8092 ( .A1(n8881), .A2(n6485), .B1(n8236), .B2(n6484), .C1(
        P2_U3152), .C2(n8453), .ZN(P2_U3340) );
  INV_X1 U8093 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6540) );
  NAND2_X1 U8094 ( .A1(n6487), .A2(n6486), .ZN(n6488) );
  NAND2_X1 U8095 ( .A1(n6872), .A2(n6501), .ZN(n7746) );
  INV_X1 U8096 ( .A(n6872), .ZN(n8389) );
  OAI21_X1 U8097 ( .B1(n6490), .B2(n7685), .A(n6874), .ZN(n6491) );
  INV_X1 U8098 ( .A(n6491), .ZN(n6837) );
  NAND2_X1 U8099 ( .A1(n6492), .A2(n7686), .ZN(n6493) );
  NAND2_X1 U8100 ( .A1(n6493), .A2(n7745), .ZN(n6494) );
  AOI21_X1 U8101 ( .B1(n6494), .B2(n7685), .A(n8620), .ZN(n6498) );
  INV_X1 U8102 ( .A(n6494), .ZN(n6496) );
  AOI21_X1 U8103 ( .B1(n6498), .B2(n6887), .A(n6497), .ZN(n6836) );
  AOI21_X1 U8104 ( .B1(n6499), .B2(n6501), .A(n9820), .ZN(n6500) );
  AND2_X1 U8105 ( .A1(n6500), .A2(n6983), .ZN(n6840) );
  AOI21_X1 U8106 ( .B1(n9815), .B2(n6501), .A(n6840), .ZN(n6502) );
  OAI211_X1 U8107 ( .C1(n6837), .C2(n9764), .A(n6836), .B(n6502), .ZN(n6504)
         );
  NAND2_X1 U8108 ( .A1(n6504), .A2(n9839), .ZN(n6503) );
  OAI21_X1 U8109 ( .B1(n9839), .B2(n6540), .A(n6503), .ZN(P2_U3524) );
  INV_X1 U8110 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U8111 ( .A1(n6504), .A2(n9826), .ZN(n6505) );
  OAI21_X1 U8112 ( .B1(n9826), .B2(n6506), .A(n6505), .ZN(P2_U3463) );
  INV_X1 U8113 ( .A(n9444), .ZN(n6522) );
  MUX2_X1 U8114 ( .A(n5194), .B(P2_REG2_REG_2__SCAN_IN), .S(n9444), .Z(n9447)
         );
  XNOR2_X1 U8115 ( .A(n9427), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n9435) );
  NAND3_X1 U8116 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9435), .ZN(n9434) );
  OAI21_X1 U8117 ( .B1(n9427), .B2(n6507), .A(n9434), .ZN(n9448) );
  NAND2_X1 U8118 ( .A1(n9447), .A2(n9448), .ZN(n9446) );
  INV_X1 U8119 ( .A(n9446), .ZN(n6508) );
  AOI21_X1 U8120 ( .B1(n6522), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6508), .ZN(
        n6516) );
  INV_X1 U8121 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6922) );
  MUX2_X1 U8122 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6922), .S(n6533), .Z(n6515)
         );
  NOR2_X1 U8123 ( .A1(n6516), .A2(n6515), .ZN(n8399) );
  INV_X1 U8124 ( .A(n6509), .ZN(n6510) );
  NAND2_X1 U8125 ( .A1(n6510), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6511) );
  OAI211_X1 U8126 ( .C1(n9753), .C2(n6512), .A(n6511), .B(n7871), .ZN(n6514)
         );
  NAND2_X1 U8127 ( .A1(n6514), .A2(n6513), .ZN(n6517) );
  NAND2_X1 U8128 ( .A1(n6517), .A2(n8392), .ZN(n6526) );
  INV_X1 U8129 ( .A(n7214), .ZN(n7874) );
  NAND2_X1 U8130 ( .A1(n6526), .A2(n7874), .ZN(n9710) );
  AOI211_X1 U8131 ( .C1(n6516), .C2(n6515), .A(n8399), .B(n8474), .ZN(n6532)
         );
  INV_X1 U8132 ( .A(n6517), .ZN(n6518) );
  NAND2_X1 U8133 ( .A1(n6518), .A2(n7214), .ZN(n9869) );
  XNOR2_X1 U8134 ( .A(n6533), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n6525) );
  MUX2_X1 U8135 ( .A(n6519), .B(P2_REG1_REG_2__SCAN_IN), .S(n9444), .Z(n9442)
         );
  INV_X1 U8136 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U8137 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9430) );
  MUX2_X1 U8138 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6521), .S(n9427), .Z(n9429)
         );
  NOR2_X1 U8139 ( .A1(n9430), .A2(n9429), .ZN(n9428) );
  INV_X1 U8140 ( .A(n9428), .ZN(n6520) );
  OAI21_X1 U8141 ( .B1(n9427), .B2(n6521), .A(n6520), .ZN(n9441) );
  NAND2_X1 U8142 ( .A1(n9442), .A2(n9441), .ZN(n9440) );
  NAND2_X1 U8143 ( .A1(n6522), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U8144 ( .A1(n9440), .A2(n6523), .ZN(n6524) );
  NAND2_X1 U8145 ( .A1(n6524), .A2(n6525), .ZN(n6539) );
  OAI21_X1 U8146 ( .B1(n6525), .B2(n6524), .A(n6539), .ZN(n6530) );
  INV_X1 U8147 ( .A(n6533), .ZN(n6537) );
  NAND2_X1 U8148 ( .A1(n9433), .A2(n6537), .ZN(n6529) );
  NOR2_X1 U8149 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10012), .ZN(n6527) );
  AOI21_X1 U8150 ( .B1(n9875), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6527), .ZN(
        n6528) );
  OAI211_X1 U8151 ( .C1(n9869), .C2(n6530), .A(n6529), .B(n6528), .ZN(n6531)
         );
  OR2_X1 U8152 ( .A1(n6532), .A2(n6531), .ZN(P2_U3248) );
  INV_X1 U8153 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n8394) );
  NOR2_X1 U8154 ( .A1(n6533), .A2(n6922), .ZN(n8393) );
  MUX2_X1 U8155 ( .A(n8394), .B(P2_REG2_REG_4__SCAN_IN), .S(n8402), .Z(n6534)
         );
  OAI21_X1 U8156 ( .B1(n8399), .B2(n8393), .A(n6534), .ZN(n8397) );
  OAI21_X1 U8157 ( .B1(n8394), .B2(n8402), .A(n8397), .ZN(n8047) );
  INV_X1 U8158 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9985) );
  MUX2_X1 U8159 ( .A(n9985), .B(P2_REG2_REG_5__SCAN_IN), .S(n8044), .Z(n8045)
         );
  XNOR2_X1 U8160 ( .A(n8047), .B(n8045), .ZN(n6550) );
  OR2_X1 U8161 ( .A1(n8044), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U8162 ( .A1(n8044), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6535) );
  AND2_X1 U8163 ( .A1(n6536), .A2(n6535), .ZN(n6544) );
  NAND2_X1 U8164 ( .A1(n6537), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U8165 ( .A1(n6539), .A2(n6538), .ZN(n8405) );
  MUX2_X1 U8166 ( .A(n6540), .B(P2_REG1_REG_4__SCAN_IN), .S(n8402), .Z(n8406)
         );
  NAND2_X1 U8167 ( .A1(n8405), .A2(n8406), .ZN(n8404) );
  OR2_X1 U8168 ( .A1(n8402), .A2(n6540), .ZN(n6541) );
  NAND2_X1 U8169 ( .A1(n8404), .A2(n6541), .ZN(n6543) );
  INV_X1 U8170 ( .A(n8017), .ZN(n6542) );
  OAI211_X1 U8171 ( .C1(n6544), .C2(n6543), .A(n9714), .B(n6542), .ZN(n6547)
         );
  AND2_X1 U8172 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6545) );
  AOI21_X1 U8173 ( .B1(n9875), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6545), .ZN(
        n6546) );
  OAI211_X1 U8174 ( .C1(n9883), .C2(n6548), .A(n6547), .B(n6546), .ZN(n6549)
         );
  AOI21_X1 U8175 ( .B1(n9877), .B2(n6550), .A(n6549), .ZN(n6551) );
  INV_X1 U8176 ( .A(n6551), .ZN(P2_U3250) );
  INV_X1 U8177 ( .A(n7327), .ZN(n6553) );
  OAI222_X1 U8178 ( .A1(n8231), .A2(n6552), .B1(n9424), .B2(n6553), .C1(n9243), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OAI222_X1 U8179 ( .A1(n8237), .A2(n6554), .B1(n8236), .B2(n6553), .C1(
        P2_U3152), .C2(n8546), .ZN(P2_U3339) );
  OR2_X1 U8180 ( .A1(n8892), .A2(n9049), .ZN(n6555) );
  NAND2_X1 U8181 ( .A1(n6556), .A2(n6555), .ZN(n6560) );
  OR2_X1 U8182 ( .A1(n6557), .A2(n6644), .ZN(n6559) );
  AOI22_X1 U8183 ( .A1(n7450), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7382), .B2(
        n9580), .ZN(n6558) );
  INV_X1 U8184 ( .A(n9048), .ZN(n6661) );
  OR2_X1 U8185 ( .A1(n9690), .A2(n6661), .ZN(n7388) );
  NAND2_X1 U8186 ( .A1(n9690), .A2(n6661), .ZN(n7540) );
  NAND2_X1 U8187 ( .A1(n6560), .A2(n7481), .ZN(n6561) );
  NAND2_X1 U8188 ( .A1(n6666), .A2(n6561), .ZN(n9689) );
  XNOR2_X1 U8189 ( .A(n6668), .B(n7481), .ZN(n6572) );
  NAND2_X1 U8190 ( .A1(n6564), .A2(n6563), .ZN(n6565) );
  AND2_X1 U8191 ( .A1(n6654), .A2(n6565), .ZN(n9653) );
  NAND2_X1 U8192 ( .A1(n7459), .A2(n9653), .ZN(n6569) );
  NAND2_X1 U8193 ( .A1(n7324), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6568) );
  NAND2_X1 U8194 ( .A1(n4416), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U8195 ( .A1(n4414), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6566) );
  NAND4_X1 U8196 ( .A1(n6569), .A2(n6568), .A3(n6567), .A4(n6566), .ZN(n9047)
         );
  INV_X1 U8197 ( .A(n9047), .ZN(n9465) );
  OAI22_X1 U8198 ( .A1(n6570), .A2(n9464), .B1(n9465), .B2(n9462), .ZN(n6571)
         );
  AOI21_X1 U8199 ( .B1(n6572), .B2(n9296), .A(n6571), .ZN(n6573) );
  OAI21_X1 U8200 ( .B1(n9689), .B2(n6574), .A(n6573), .ZN(n9694) );
  NAND2_X1 U8201 ( .A1(n9694), .A2(n9281), .ZN(n6582) );
  INV_X1 U8202 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6576) );
  INV_X1 U8203 ( .A(n6575), .ZN(n6621) );
  OAI22_X1 U8204 ( .A1(n9281), .A2(n6576), .B1(n6621), .B2(n9258), .ZN(n6580)
         );
  NAND2_X1 U8205 ( .A1(n6577), .A2(n9690), .ZN(n6578) );
  NAND2_X1 U8206 ( .A1(n6670), .A2(n6578), .ZN(n9693) );
  NOR2_X1 U8207 ( .A1(n9693), .A2(n6591), .ZN(n6579) );
  AOI211_X1 U8208 ( .C1(n9469), .C2(n9690), .A(n6580), .B(n6579), .ZN(n6581)
         );
  OAI211_X1 U8209 ( .C1(n9689), .C2(n6583), .A(n6582), .B(n6581), .ZN(P1_U3283) );
  OAI21_X1 U8210 ( .B1(n6585), .B2(n7535), .A(n6584), .ZN(n9688) );
  OAI21_X1 U8211 ( .B1(n6587), .B2(n9684), .A(n6586), .ZN(n9685) );
  AOI22_X1 U8212 ( .A1(n9469), .A2(n6589), .B1(n9652), .B2(n6588), .ZN(n6590)
         );
  OAI21_X1 U8213 ( .B1(n9685), .B2(n6591), .A(n6590), .ZN(n6598) );
  NAND2_X1 U8214 ( .A1(n6592), .A2(n7500), .ZN(n6593) );
  XNOR2_X1 U8215 ( .A(n6593), .B(n7535), .ZN(n6596) );
  NAND2_X1 U8216 ( .A1(n9688), .A2(n9648), .ZN(n6595) );
  AOI22_X1 U8217 ( .A1(n9293), .A2(n9049), .B1(n9051), .B2(n9291), .ZN(n6594)
         );
  OAI211_X1 U8218 ( .C1(n9459), .C2(n6596), .A(n6595), .B(n6594), .ZN(n9686)
         );
  MUX2_X1 U8219 ( .A(n9686), .B(P1_REG2_REG_6__SCAN_IN), .S(n4419), .Z(n6597)
         );
  AOI211_X1 U8220 ( .C1(n9659), .C2(n9688), .A(n6598), .B(n6597), .ZN(n6599)
         );
  INV_X1 U8221 ( .A(n6599), .ZN(P1_U3285) );
  NAND2_X1 U8222 ( .A1(n9690), .A2(n7995), .ZN(n6601) );
  NAND2_X1 U8223 ( .A1(n9048), .A2(n8004), .ZN(n6600) );
  NAND2_X1 U8224 ( .A1(n6601), .A2(n6600), .ZN(n6602) );
  XNOR2_X1 U8225 ( .A(n6602), .B(n8005), .ZN(n6641) );
  INV_X1 U8226 ( .A(n6603), .ZN(n6605) );
  NAND2_X1 U8227 ( .A1(n6605), .A2(n6604), .ZN(n6606) );
  NAND2_X1 U8228 ( .A1(n8892), .A2(n6077), .ZN(n6609) );
  NAND2_X1 U8229 ( .A1(n9049), .A2(n6394), .ZN(n6608) );
  NAND2_X1 U8230 ( .A1(n6609), .A2(n6608), .ZN(n6610) );
  XNOR2_X1 U8231 ( .A(n6610), .B(n8005), .ZN(n6612) );
  AND2_X1 U8232 ( .A1(n9049), .A2(n8007), .ZN(n6611) );
  AOI21_X1 U8233 ( .B1(n8892), .B2(n8004), .A(n6611), .ZN(n6613) );
  XNOR2_X1 U8234 ( .A(n6612), .B(n6613), .ZN(n8889) );
  INV_X1 U8235 ( .A(n6612), .ZN(n6614) );
  NAND2_X1 U8236 ( .A1(n6614), .A2(n6613), .ZN(n6615) );
  AND2_X1 U8237 ( .A1(n9048), .A2(n8007), .ZN(n6616) );
  AOI21_X1 U8238 ( .B1(n9690), .B2(n8004), .A(n6616), .ZN(n6617) );
  NAND2_X1 U8239 ( .A1(n6643), .A2(n6642), .ZN(n6619) );
  XOR2_X1 U8240 ( .A(n6641), .B(n6619), .Z(n6625) );
  NOR2_X1 U8241 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6620), .ZN(n9579) );
  OAI22_X1 U8242 ( .A1(n9010), .A2(n6621), .B1(n9009), .B2(n9465), .ZN(n6622)
         );
  AOI211_X1 U8243 ( .C1(n8978), .C2(n9049), .A(n9579), .B(n6622), .ZN(n6624)
         );
  NAND2_X1 U8244 ( .A1(n9690), .A2(n9036), .ZN(n6623) );
  OAI211_X1 U8245 ( .C1(n6625), .C2(n9038), .A(n6624), .B(n6623), .ZN(P1_U3219) );
  OAI21_X1 U8246 ( .B1(n6627), .B2(n4507), .A(n6626), .ZN(n6631) );
  INV_X1 U8247 ( .A(n9773), .ZN(n6879) );
  OAI22_X1 U8248 ( .A1(n8348), .A2(n6879), .B1(n8369), .B2(n9735), .ZN(n6630)
         );
  NAND2_X1 U8249 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8100) );
  NAND2_X1 U8250 ( .A1(n8345), .A2(n8734), .ZN(n6628) );
  OAI211_X1 U8251 ( .C1(n8370), .C2(n6875), .A(n8100), .B(n6628), .ZN(n6629)
         );
  AOI211_X1 U8252 ( .C1(n6631), .C2(n8353), .A(n6630), .B(n6629), .ZN(n6632)
         );
  INV_X1 U8253 ( .A(n6632), .ZN(P2_U3241) );
  XNOR2_X1 U8254 ( .A(n6634), .B(n6633), .ZN(n6639) );
  OR2_X1 U8255 ( .A1(n6878), .A2(n9734), .ZN(n6636) );
  NAND2_X1 U8256 ( .A1(n8387), .A2(n8731), .ZN(n6635) );
  NAND2_X1 U8257 ( .A1(n6636), .A2(n6635), .ZN(n6895) );
  AND2_X1 U8258 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9874) );
  AOI21_X1 U8259 ( .B1(n8358), .B2(n6895), .A(n9874), .ZN(n6638) );
  AOI22_X1 U8260 ( .A1(n6886), .A2(n8374), .B1(n8345), .B2(n6883), .ZN(n6637)
         );
  OAI211_X1 U8261 ( .C1(n6639), .C2(n8376), .A(n6638), .B(n6637), .ZN(P2_U3215) );
  INV_X1 U8262 ( .A(n7288), .ZN(n6677) );
  OAI222_X1 U8263 ( .A1(n8237), .A2(n6640), .B1(n8236), .B2(n6677), .C1(n7860), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  NAND2_X1 U8264 ( .A1(n6645), .A2(n7449), .ZN(n6647) );
  AOI22_X1 U8265 ( .A1(n7450), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7382), .B2(
        n9599), .ZN(n6646) );
  NAND2_X1 U8266 ( .A1(n9649), .A2(n7995), .ZN(n6649) );
  NAND2_X1 U8267 ( .A1(n9047), .A2(n8004), .ZN(n6648) );
  NAND2_X1 U8268 ( .A1(n6649), .A2(n6648), .ZN(n6650) );
  XNOR2_X1 U8269 ( .A(n6650), .B(n7998), .ZN(n6741) );
  AND2_X1 U8270 ( .A1(n9047), .A2(n8007), .ZN(n6651) );
  AOI21_X1 U8271 ( .B1(n9649), .B2(n8004), .A(n6651), .ZN(n6740) );
  XNOR2_X1 U8272 ( .A(n6741), .B(n6740), .ZN(n6762) );
  XOR2_X1 U8273 ( .A(n6788), .B(n6762), .Z(n6664) );
  NAND2_X1 U8274 ( .A1(n7324), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6659) );
  NAND2_X1 U8275 ( .A1(n4417), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6658) );
  INV_X1 U8276 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6653) );
  NAND2_X1 U8277 ( .A1(n6654), .A2(n6653), .ZN(n6655) );
  AND2_X1 U8278 ( .A1(n6695), .A2(n6655), .ZN(n9468) );
  NAND2_X1 U8279 ( .A1(n7459), .A2(n9468), .ZN(n6657) );
  NAND2_X1 U8280 ( .A1(n4414), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6656) );
  NAND4_X1 U8281 ( .A1(n6659), .A2(n6658), .A3(n6657), .A4(n6656), .ZN(n9046)
         );
  AOI22_X1 U8282 ( .A1(n9030), .A2(n9046), .B1(n9653), .B2(n9029), .ZN(n6660)
         );
  NAND2_X1 U8283 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9592) );
  OAI211_X1 U8284 ( .C1(n9034), .C2(n6661), .A(n6660), .B(n9592), .ZN(n6662)
         );
  AOI21_X1 U8285 ( .B1(n9649), .B2(n9036), .A(n6662), .ZN(n6663) );
  OAI21_X1 U8286 ( .B1(n6664), .B2(n9038), .A(n6663), .ZN(P1_U3229) );
  INV_X1 U8287 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U8288 ( .A1(n9690), .A2(n9048), .ZN(n6665) );
  NOR2_X1 U8289 ( .A1(n9649), .A2(n9465), .ZN(n7542) );
  NAND2_X1 U8290 ( .A1(n9649), .A2(n9465), .ZN(n9456) );
  INV_X1 U8291 ( .A(n9456), .ZN(n6667) );
  OR2_X1 U8292 ( .A1(n7542), .A2(n6667), .ZN(n7484) );
  XNOR2_X1 U8293 ( .A(n6685), .B(n7484), .ZN(n9645) );
  INV_X1 U8294 ( .A(n7540), .ZN(n7545) );
  XNOR2_X1 U8295 ( .A(n6710), .B(n7484), .ZN(n6669) );
  AOI222_X1 U8296 ( .A1(n9296), .A2(n6669), .B1(n9048), .B2(n9291), .C1(n9046), 
        .C2(n9293), .ZN(n9646) );
  AOI21_X1 U8297 ( .B1(n9649), .B2(n6670), .A(n9473), .ZN(n9651) );
  AOI22_X1 U8298 ( .A1(n9651), .A2(n9471), .B1(n9392), .B2(n9649), .ZN(n6671)
         );
  OAI211_X1 U8299 ( .C1(n9645), .C2(n9396), .A(n9646), .B(n6671), .ZN(n6674)
         );
  NAND2_X1 U8300 ( .A1(n6674), .A2(n9671), .ZN(n6672) );
  OAI21_X1 U8301 ( .B1(n9671), .B2(n6673), .A(n6672), .ZN(P1_U3481) );
  INV_X1 U8302 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6676) );
  NAND2_X1 U8303 ( .A1(n6674), .A2(n9702), .ZN(n6675) );
  OAI21_X1 U8304 ( .B1(n9702), .B2(n6676), .A(n6675), .ZN(P1_U3532) );
  OAI222_X1 U8305 ( .A1(n8231), .A2(n6679), .B1(P1_U3084), .B2(n6678), .C1(
        n9424), .C2(n6677), .ZN(P1_U3333) );
  INV_X1 U8306 ( .A(n7277), .ZN(n6682) );
  OAI222_X1 U8307 ( .A1(n8237), .A2(n6681), .B1(n8236), .B2(n6682), .C1(n6680), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  OAI222_X1 U8308 ( .A1(n8231), .A2(n10056), .B1(P1_U3084), .B2(n7630), .C1(
        n9424), .C2(n6682), .ZN(P1_U3332) );
  AND2_X1 U8309 ( .A1(n9649), .A2(n9047), .ZN(n6684) );
  NAND2_X1 U8310 ( .A1(n6686), .A2(n7449), .ZN(n6689) );
  AOI22_X1 U8311 ( .A1(n7450), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7382), .B2(
        n6687), .ZN(n6688) );
  NAND2_X1 U8312 ( .A1(n6689), .A2(n6688), .ZN(n9470) );
  INV_X1 U8313 ( .A(n9046), .ZN(n6713) );
  OR2_X1 U8314 ( .A1(n9470), .A2(n6713), .ZN(n9460) );
  NAND2_X1 U8315 ( .A1(n9470), .A2(n6713), .ZN(n7551) );
  NAND2_X1 U8316 ( .A1(n9460), .A2(n7551), .ZN(n9454) );
  NAND2_X1 U8317 ( .A1(n9452), .A2(n9454), .ZN(n6690) );
  OR2_X1 U8318 ( .A1(n9470), .A2(n9046), .ZN(n6812) );
  NAND2_X1 U8319 ( .A1(n6690), .A2(n6812), .ZN(n6701) );
  NAND2_X1 U8320 ( .A1(n6691), .A2(n7449), .ZN(n6693) );
  AOI22_X1 U8321 ( .A1(n7450), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7382), .B2(
        n9603), .ZN(n6692) );
  NAND2_X1 U8322 ( .A1(n4414), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6700) );
  OR2_X1 U8323 ( .A1(n7456), .A2(n6170), .ZN(n6699) );
  NAND2_X1 U8324 ( .A1(n7324), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6698) );
  NAND2_X1 U8325 ( .A1(n6695), .A2(n6694), .ZN(n6696) );
  AND2_X1 U8326 ( .A1(n6704), .A2(n6696), .ZN(n6756) );
  NAND2_X1 U8327 ( .A1(n7459), .A2(n6756), .ZN(n6697) );
  NAND4_X1 U8328 ( .A1(n6700), .A2(n6699), .A3(n6698), .A4(n6697), .ZN(n9045)
         );
  XNOR2_X1 U8329 ( .A(n6859), .B(n9045), .ZN(n7552) );
  XNOR2_X1 U8330 ( .A(n6701), .B(n7552), .ZN(n6861) );
  NAND2_X1 U8331 ( .A1(n4414), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U8332 ( .A1(n7324), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U8333 ( .A1(n6704), .A2(n6703), .ZN(n6705) );
  AND2_X1 U8334 ( .A1(n6800), .A2(n6705), .ZN(n6848) );
  NAND2_X1 U8335 ( .A1(n7459), .A2(n6848), .ZN(n6707) );
  NAND2_X1 U8336 ( .A1(n4416), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6706) );
  NAND4_X1 U8337 ( .A1(n6709), .A2(n6708), .A3(n6707), .A4(n6706), .ZN(n9044)
         );
  INV_X1 U8338 ( .A(n9044), .ZN(n6816) );
  AND2_X1 U8339 ( .A1(n7551), .A2(n9456), .ZN(n7547) );
  XNOR2_X1 U8340 ( .A(n6818), .B(n7552), .ZN(n6712) );
  OAI222_X1 U8341 ( .A1(n9464), .A2(n6713), .B1(n9462), .B2(n6816), .C1(n6712), 
        .C2(n9459), .ZN(n6857) );
  INV_X1 U8342 ( .A(n6859), .ZN(n6761) );
  INV_X1 U8343 ( .A(n9470), .ZN(n9479) );
  INV_X1 U8344 ( .A(n6714), .ZN(n9472) );
  AOI211_X1 U8345 ( .C1(n6859), .C2(n9472), .A(n9692), .B(n6822), .ZN(n6858)
         );
  NAND2_X1 U8346 ( .A1(n6858), .A2(n9475), .ZN(n6716) );
  AOI22_X1 U8347 ( .A1(n4419), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n6756), .B2(
        n9652), .ZN(n6715) );
  OAI211_X1 U8348 ( .C1(n6761), .C2(n9656), .A(n6716), .B(n6715), .ZN(n6717)
         );
  AOI21_X1 U8349 ( .B1(n6857), .B2(n9281), .A(n6717), .ZN(n6718) );
  OAI21_X1 U8350 ( .B1(n6861), .B2(n9308), .A(n6718), .ZN(P1_U3280) );
  NAND2_X1 U8351 ( .A1(n6720), .A2(n6724), .ZN(n6721) );
  INV_X1 U8352 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9617) );
  NAND2_X1 U8353 ( .A1(n9618), .A2(n9617), .ZN(n9616) );
  NAND2_X1 U8354 ( .A1(n6721), .A2(n9616), .ZN(n6903) );
  XNOR2_X1 U8355 ( .A(n6903), .B(n7380), .ZN(n6723) );
  INV_X1 U8356 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6722) );
  NOR2_X1 U8357 ( .A1(n6722), .A2(n6723), .ZN(n6904) );
  AOI211_X1 U8358 ( .C1(n6723), .C2(n6722), .A(n6904), .B(n9629), .ZN(n6731)
         );
  INV_X1 U8359 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9523) );
  AOI22_X1 U8360 ( .A1(n9615), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n9523), .B2(
        n6724), .ZN(n9621) );
  NAND2_X1 U8361 ( .A1(n9621), .A2(n9620), .ZN(n9619) );
  OAI21_X1 U8362 ( .B1(n9615), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9619), .ZN(
        n6909) );
  XNOR2_X1 U8363 ( .A(n6909), .B(n7380), .ZN(n6727) );
  INV_X1 U8364 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6726) );
  AOI211_X1 U8365 ( .C1(n6727), .C2(n6726), .A(n6910), .B(n9060), .ZN(n6730)
         );
  NAND2_X1 U8366 ( .A1(n9640), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n6728) );
  NAND2_X1 U8367 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9031) );
  OAI211_X1 U8368 ( .C1(n9069), .C2(n7380), .A(n6728), .B(n9031), .ZN(n6729)
         );
  OR3_X1 U8369 ( .A1(n6731), .A2(n6730), .A3(n6729), .ZN(P1_U3256) );
  NAND2_X1 U8370 ( .A1(n9470), .A2(n7995), .ZN(n6733) );
  NAND2_X1 U8371 ( .A1(n9046), .A2(n8004), .ZN(n6732) );
  NAND2_X1 U8372 ( .A1(n6733), .A2(n6732), .ZN(n6734) );
  XNOR2_X1 U8373 ( .A(n6734), .B(n8005), .ZN(n6738) );
  INV_X1 U8374 ( .A(n6738), .ZN(n6736) );
  AND2_X1 U8375 ( .A1(n9046), .A2(n8007), .ZN(n6735) );
  AOI21_X1 U8376 ( .B1(n9470), .B2(n8004), .A(n6735), .ZN(n6737) );
  NAND2_X1 U8377 ( .A1(n6736), .A2(n6737), .ZN(n6742) );
  INV_X1 U8378 ( .A(n6742), .ZN(n6739) );
  XNOR2_X1 U8379 ( .A(n6738), .B(n6737), .ZN(n6766) );
  NOR2_X1 U8380 ( .A1(n6739), .A2(n6766), .ZN(n6744) );
  OR2_X1 U8381 ( .A1(n6762), .A2(n6744), .ZN(n6786) );
  OR2_X1 U8382 ( .A1(n6788), .A2(n6786), .ZN(n6753) );
  NAND2_X1 U8383 ( .A1(n6741), .A2(n6740), .ZN(n6763) );
  AND2_X1 U8384 ( .A1(n6763), .A2(n6742), .ZN(n6743) );
  OR2_X1 U8385 ( .A1(n6744), .A2(n6743), .ZN(n6752) );
  NAND2_X1 U8386 ( .A1(n6753), .A2(n6752), .ZN(n6749) );
  NAND2_X1 U8387 ( .A1(n6859), .A2(n7995), .ZN(n6746) );
  NAND2_X1 U8388 ( .A1(n9045), .A2(n8004), .ZN(n6745) );
  NAND2_X1 U8389 ( .A1(n6746), .A2(n6745), .ZN(n6747) );
  XNOR2_X1 U8390 ( .A(n6747), .B(n7998), .ZN(n6782) );
  AND2_X1 U8391 ( .A1(n9045), .A2(n8007), .ZN(n6748) );
  AOI21_X1 U8392 ( .B1(n6859), .B2(n8004), .A(n6748), .ZN(n6783) );
  XNOR2_X1 U8393 ( .A(n6782), .B(n6783), .ZN(n6750) );
  AOI21_X1 U8394 ( .B1(n6749), .B2(n6750), .A(n9038), .ZN(n6755) );
  INV_X1 U8395 ( .A(n6750), .ZN(n6751) );
  AND2_X1 U8396 ( .A1(n6752), .A2(n6751), .ZN(n6789) );
  NAND2_X1 U8397 ( .A1(n6753), .A2(n6789), .ZN(n6754) );
  NAND2_X1 U8398 ( .A1(n6755), .A2(n6754), .ZN(n6760) );
  AND2_X1 U8399 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9602) );
  INV_X1 U8400 ( .A(n6756), .ZN(n6757) );
  OAI22_X1 U8401 ( .A1(n9010), .A2(n6757), .B1(n9009), .B2(n6816), .ZN(n6758)
         );
  AOI211_X1 U8402 ( .C1(n8978), .C2(n9046), .A(n9602), .B(n6758), .ZN(n6759)
         );
  OAI211_X1 U8403 ( .C1(n6761), .C2(n9024), .A(n6760), .B(n6759), .ZN(P1_U3234) );
  OR2_X1 U8404 ( .A1(n6788), .A2(n6762), .ZN(n6764) );
  NAND2_X1 U8405 ( .A1(n6764), .A2(n6763), .ZN(n6765) );
  XOR2_X1 U8406 ( .A(n6766), .B(n6765), .Z(n6771) );
  AOI22_X1 U8407 ( .A1(n9030), .A2(n9045), .B1(n9468), .B2(n9029), .ZN(n6768)
         );
  OAI211_X1 U8408 ( .C1(n9034), .C2(n9465), .A(n6768), .B(n6767), .ZN(n6769)
         );
  AOI21_X1 U8409 ( .B1(n9470), .B2(n9036), .A(n6769), .ZN(n6770) );
  OAI21_X1 U8410 ( .B1(n6771), .B2(n9038), .A(n6770), .ZN(P1_U3215) );
  XNOR2_X1 U8411 ( .A(n6773), .B(n6772), .ZN(n6777) );
  INV_X1 U8412 ( .A(n8370), .ZN(n8316) );
  NAND2_X1 U8413 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8088) );
  OAI21_X1 U8414 ( .B1(n8368), .B2(n9742), .A(n8088), .ZN(n6775) );
  INV_X1 U8415 ( .A(n7062), .ZN(n9788) );
  OAI22_X1 U8416 ( .A1(n8348), .A2(n9788), .B1(n8369), .B2(n9733), .ZN(n6774)
         );
  AOI211_X1 U8417 ( .C1(n8316), .C2(n8732), .A(n6775), .B(n6774), .ZN(n6776)
         );
  OAI21_X1 U8418 ( .B1(n6777), .B2(n8376), .A(n6776), .ZN(P2_U3223) );
  NAND2_X1 U8419 ( .A1(n6778), .A2(n7449), .ZN(n6781) );
  AOI22_X1 U8420 ( .A1(n7450), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7382), .B2(
        n6779), .ZN(n6780) );
  INV_X1 U8421 ( .A(n7002), .ZN(n6850) );
  INV_X1 U8422 ( .A(n6782), .ZN(n6785) );
  INV_X1 U8423 ( .A(n6783), .ZN(n6784) );
  AND2_X1 U8424 ( .A1(n6785), .A2(n6784), .ZN(n6790) );
  OR2_X1 U8425 ( .A1(n6786), .A2(n6790), .ZN(n6787) );
  OR2_X1 U8426 ( .A1(n6790), .A2(n6789), .ZN(n6934) );
  AND2_X1 U8427 ( .A1(n6936), .A2(n6934), .ZN(n6796) );
  NAND2_X1 U8428 ( .A1(n7002), .A2(n7995), .ZN(n6792) );
  NAND2_X1 U8429 ( .A1(n9044), .A2(n8004), .ZN(n6791) );
  NAND2_X1 U8430 ( .A1(n6792), .A2(n6791), .ZN(n6793) );
  XNOR2_X1 U8431 ( .A(n6793), .B(n7998), .ZN(n6937) );
  AND2_X1 U8432 ( .A1(n9044), .A2(n8007), .ZN(n6794) );
  AOI21_X1 U8433 ( .B1(n7002), .B2(n8004), .A(n6794), .ZN(n6938) );
  XNOR2_X1 U8434 ( .A(n6937), .B(n6938), .ZN(n6795) );
  XNOR2_X1 U8435 ( .A(n6796), .B(n6795), .ZN(n6797) );
  NAND2_X1 U8436 ( .A1(n6797), .A2(n9015), .ZN(n6810) );
  INV_X1 U8437 ( .A(n6848), .ZN(n6806) );
  NAND2_X1 U8438 ( .A1(n7324), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6805) );
  INV_X1 U8439 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6798) );
  OR2_X1 U8440 ( .A1(n7456), .A2(n6798), .ZN(n6804) );
  NAND2_X1 U8441 ( .A1(n4414), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6803) );
  INV_X1 U8442 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6799) );
  NAND2_X1 U8443 ( .A1(n6800), .A2(n6799), .ZN(n6801) );
  AND2_X1 U8444 ( .A1(n6957), .A2(n6801), .ZN(n9300) );
  NAND2_X1 U8445 ( .A1(n7459), .A2(n9300), .ZN(n6802) );
  NAND4_X1 U8446 ( .A1(n6805), .A2(n6804), .A3(n6803), .A4(n6802), .ZN(n9043)
         );
  INV_X1 U8447 ( .A(n9043), .ZN(n7385) );
  OAI22_X1 U8448 ( .A1(n9010), .A2(n6806), .B1(n9009), .B2(n7385), .ZN(n6807)
         );
  AOI211_X1 U8449 ( .C1(n8978), .C2(n9045), .A(n6808), .B(n6807), .ZN(n6809)
         );
  OAI211_X1 U8450 ( .C1(n6850), .C2(n9024), .A(n6810), .B(n6809), .ZN(P1_U3222) );
  NAND2_X1 U8451 ( .A1(n6859), .A2(n9045), .ZN(n6811) );
  AND2_X1 U8452 ( .A1(n9454), .A2(n6811), .ZN(n7003) );
  NAND2_X1 U8453 ( .A1(n9452), .A2(n7003), .ZN(n6815) );
  INV_X1 U8454 ( .A(n6811), .ZN(n6814) );
  AND2_X1 U8455 ( .A1(n6812), .A2(n4994), .ZN(n6813) );
  OR2_X1 U8456 ( .A1(n6814), .A2(n6813), .ZN(n7006) );
  AND2_X1 U8457 ( .A1(n6815), .A2(n7006), .ZN(n6817) );
  NAND2_X1 U8458 ( .A1(n7002), .A2(n6816), .ZN(n7554) );
  NAND2_X1 U8459 ( .A1(n7557), .A2(n7554), .ZN(n7485) );
  XNOR2_X1 U8460 ( .A(n6817), .B(n7485), .ZN(n6856) );
  INV_X1 U8461 ( .A(n9045), .ZN(n9463) );
  NOR2_X1 U8462 ( .A1(n6859), .A2(n9463), .ZN(n7013) );
  NAND2_X1 U8463 ( .A1(n6859), .A2(n9463), .ZN(n7389) );
  AOI21_X1 U8464 ( .B1(n6819), .B2(n7485), .A(n9459), .ZN(n6821) );
  OAI22_X1 U8465 ( .A1(n9463), .A2(n9464), .B1(n7385), .B2(n9462), .ZN(n6820)
         );
  AOI21_X1 U8466 ( .B1(n6821), .B2(n7015), .A(n6820), .ZN(n6851) );
  INV_X1 U8467 ( .A(n6822), .ZN(n6824) );
  NAND2_X1 U8468 ( .A1(n6822), .A2(n6850), .ZN(n7040) );
  INV_X1 U8469 ( .A(n7040), .ZN(n6823) );
  AOI211_X1 U8470 ( .C1(n7002), .C2(n6824), .A(n9692), .B(n6823), .ZN(n6854)
         );
  AOI21_X1 U8471 ( .B1(n9392), .B2(n7002), .A(n6854), .ZN(n6825) );
  OAI211_X1 U8472 ( .C1(n6856), .C2(n9396), .A(n6851), .B(n6825), .ZN(n6827)
         );
  NAND2_X1 U8473 ( .A1(n6827), .A2(n9702), .ZN(n6826) );
  OAI21_X1 U8474 ( .B1(n9702), .B2(n6162), .A(n6826), .ZN(P1_U3535) );
  INV_X1 U8475 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n6829) );
  NAND2_X1 U8476 ( .A1(n6827), .A2(n9671), .ZN(n6828) );
  OAI21_X1 U8477 ( .B1(n9671), .B2(n6829), .A(n6828), .ZN(P1_U3490) );
  OR2_X1 U8478 ( .A1(n6834), .A2(n8546), .ZN(n7073) );
  NAND2_X1 U8479 ( .A1(n9740), .A2(n7073), .ZN(n6835) );
  OAI22_X1 U8480 ( .A1(n6837), .A2(n8727), .B1(n6836), .B2(n9745), .ZN(n6845)
         );
  NAND2_X1 U8481 ( .A1(n6838), .A2(n8546), .ZN(n7063) );
  INV_X1 U8482 ( .A(n7063), .ZN(n8756) );
  AOI22_X1 U8483 ( .A1(n8756), .A2(n6840), .B1(n6839), .B2(n8752), .ZN(n6843)
         );
  OR2_X1 U8484 ( .A1(n9747), .A2(n4677), .ZN(n6842) );
  OAI211_X1 U8485 ( .C1(n8394), .C2(n9749), .A(n6843), .B(n6842), .ZN(n6844)
         );
  OR2_X1 U8486 ( .A1(n6845), .A2(n6844), .ZN(P2_U3292) );
  INV_X1 U8487 ( .A(n7298), .ZN(n7886) );
  OAI222_X1 U8488 ( .A1(n8231), .A2(n6847), .B1(n9424), .B2(n7886), .C1(n6846), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  AOI22_X1 U8489 ( .A1(n4419), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n6848), .B2(
        n9652), .ZN(n6849) );
  OAI21_X1 U8490 ( .B1(n6850), .B2(n9656), .A(n6849), .ZN(n6853) );
  NOR2_X1 U8491 ( .A1(n6851), .A2(n4419), .ZN(n6852) );
  AOI211_X1 U8492 ( .C1(n6854), .C2(n9475), .A(n6853), .B(n6852), .ZN(n6855)
         );
  OAI21_X1 U8493 ( .B1(n9308), .B2(n6856), .A(n6855), .ZN(P1_U3279) );
  INV_X1 U8494 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n6863) );
  AOI211_X1 U8495 ( .C1(n9392), .C2(n6859), .A(n6858), .B(n6857), .ZN(n6860)
         );
  OAI21_X1 U8496 ( .B1(n9396), .B2(n6861), .A(n6860), .ZN(n6864) );
  NAND2_X1 U8497 ( .A1(n6864), .A2(n9671), .ZN(n6862) );
  OAI21_X1 U8498 ( .B1(n9671), .B2(n6863), .A(n6862), .ZN(P1_U3487) );
  NAND2_X1 U8499 ( .A1(n6864), .A2(n9702), .ZN(n6865) );
  OAI21_X1 U8500 ( .B1(n9702), .B2(n6866), .A(n6865), .ZN(P1_U3534) );
  NAND2_X1 U8501 ( .A1(n6322), .A2(n7729), .ZN(n7689) );
  INV_X1 U8502 ( .A(n7689), .ZN(n9765) );
  AOI22_X1 U8503 ( .A1(n7689), .A2(n9737), .B1(n8731), .B2(n6449), .ZN(n9761)
         );
  OAI21_X1 U8504 ( .B1(n6455), .B2(n9743), .A(n9761), .ZN(n6868) );
  INV_X1 U8505 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9712) );
  NOR2_X1 U8506 ( .A1(n9749), .A2(n9712), .ZN(n6867) );
  AOI21_X1 U8507 ( .B1(n9749), .B2(n6868), .A(n6867), .ZN(n6871) );
  OAI21_X1 U8508 ( .B1(n9727), .B2(n8749), .A(n6869), .ZN(n6870) );
  OAI211_X1 U8509 ( .C1(n9765), .C2(n8727), .A(n6871), .B(n6870), .ZN(P2_U3296) );
  NAND2_X1 U8510 ( .A1(n6872), .A2(n4677), .ZN(n6873) );
  NAND2_X1 U8511 ( .A1(n6875), .A2(n6987), .ZN(n7749) );
  INV_X1 U8512 ( .A(n6875), .ZN(n8730) );
  NAND2_X1 U8513 ( .A1(n8730), .A2(n9770), .ZN(n7721) );
  NAND2_X1 U8514 ( .A1(n7749), .A2(n7721), .ZN(n7690) );
  NAND2_X1 U8515 ( .A1(n6875), .A2(n9770), .ZN(n6876) );
  NAND2_X1 U8516 ( .A1(n6877), .A2(n6876), .ZN(n8736) );
  INV_X1 U8517 ( .A(n8736), .ZN(n6881) );
  NAND2_X1 U8518 ( .A1(n6878), .A2(n9773), .ZN(n7759) );
  INV_X1 U8519 ( .A(n6878), .ZN(n8388) );
  NAND2_X1 U8520 ( .A1(n8388), .A2(n6879), .ZN(n7753) );
  NAND2_X1 U8521 ( .A1(n8388), .A2(n9773), .ZN(n6882) );
  NAND2_X1 U8522 ( .A1(n9735), .A2(n6886), .ZN(n7760) );
  NAND2_X1 U8523 ( .A1(n8732), .A2(n9783), .ZN(n7761) );
  OAI21_X1 U8524 ( .B1(n5000), .B2(n6891), .A(n7050), .ZN(n9786) );
  INV_X1 U8525 ( .A(n9786), .ZN(n6902) );
  OAI211_X1 U8526 ( .C1(n8737), .C2(n9783), .A(n9774), .B(n9723), .ZN(n9782)
         );
  INV_X1 U8527 ( .A(n6883), .ZN(n6884) );
  OAI22_X1 U8528 ( .A1(n9782), .A2(n7063), .B1(n6884), .B2(n9743), .ZN(n6885)
         );
  AOI21_X1 U8529 ( .B1(n8749), .B2(n6886), .A(n6885), .ZN(n6901) );
  AND2_X1 U8530 ( .A1(n6977), .A2(n7721), .ZN(n7724) );
  NAND2_X1 U8531 ( .A1(n6887), .A2(n7724), .ZN(n6888) );
  NAND2_X1 U8532 ( .A1(n6888), .A2(n7749), .ZN(n8728) );
  NAND2_X1 U8533 ( .A1(n6893), .A2(n7759), .ZN(n6889) );
  NAND2_X1 U8534 ( .A1(n6889), .A2(n6891), .ZN(n6894) );
  INV_X1 U8535 ( .A(n7759), .ZN(n6890) );
  NOR2_X1 U8536 ( .A1(n6891), .A2(n6890), .ZN(n6892) );
  NAND2_X1 U8537 ( .A1(n6893), .A2(n6892), .ZN(n7045) );
  NAND3_X1 U8538 ( .A1(n6894), .A2(n9737), .A3(n7045), .ZN(n6897) );
  INV_X1 U8539 ( .A(n6895), .ZN(n6896) );
  NAND2_X1 U8540 ( .A1(n6897), .A2(n6896), .ZN(n9785) );
  INV_X1 U8541 ( .A(n9785), .ZN(n6899) );
  INV_X1 U8542 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6898) );
  MUX2_X1 U8543 ( .A(n6899), .B(n6898), .S(n9745), .Z(n6900) );
  OAI211_X1 U8544 ( .C1(n6902), .C2(n8727), .A(n6901), .B(n6900), .ZN(P2_U3289) );
  NOR2_X1 U8545 ( .A1(n7380), .A2(n6903), .ZN(n6905) );
  NAND2_X1 U8546 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n7655), .ZN(n6906) );
  OAI21_X1 U8547 ( .B1(n7655), .B2(P1_REG2_REG_16__SCAN_IN), .A(n6906), .ZN(
        n6907) );
  AOI211_X1 U8548 ( .C1(n6908), .C2(n6907), .A(n7650), .B(n9629), .ZN(n6919)
         );
  NOR2_X1 U8549 ( .A1(n7380), .A2(n6909), .ZN(n6911) );
  XNOR2_X1 U8550 ( .A(n7655), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n6912) );
  NOR2_X1 U8551 ( .A1(n6913), .A2(n6912), .ZN(n7654) );
  AOI211_X1 U8552 ( .C1(n6913), .C2(n6912), .A(n7654), .B(n9060), .ZN(n6918)
         );
  INV_X1 U8553 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n6916) );
  NAND2_X1 U8554 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n6915) );
  NAND2_X1 U8555 ( .A1(n9635), .A2(n7655), .ZN(n6914) );
  OAI211_X1 U8556 ( .C1(n9627), .C2(n6916), .A(n6915), .B(n6914), .ZN(n6917)
         );
  OR3_X1 U8557 ( .A1(n6919), .A2(n6918), .A3(n6917), .ZN(P1_U3257) );
  AOI22_X1 U8558 ( .A1(n6920), .A2(n8756), .B1(n8752), .B2(n10012), .ZN(n6921)
         );
  OAI21_X1 U8559 ( .B1(n6922), .B2(n9749), .A(n6921), .ZN(n6923) );
  INV_X1 U8560 ( .A(n6923), .ZN(n6927) );
  AOI22_X1 U8561 ( .A1(n6925), .A2(n8751), .B1(n8749), .B2(n4421), .ZN(n6926)
         );
  OAI211_X1 U8562 ( .C1(n9745), .C2(n6928), .A(n6927), .B(n6926), .ZN(P2_U3293) );
  NAND2_X1 U8563 ( .A1(n6929), .A2(n7449), .ZN(n6932) );
  AOI22_X1 U8564 ( .A1(n7450), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7382), .B2(
        n6930), .ZN(n6931) );
  INV_X1 U8565 ( .A(n7386), .ZN(n9302) );
  NAND2_X1 U8566 ( .A1(n6937), .A2(n6938), .ZN(n6933) );
  AND2_X1 U8567 ( .A1(n6934), .A2(n6933), .ZN(n6935) );
  NAND2_X1 U8568 ( .A1(n6936), .A2(n6935), .ZN(n6942) );
  INV_X1 U8569 ( .A(n6937), .ZN(n6940) );
  INV_X1 U8570 ( .A(n6938), .ZN(n6939) );
  NAND2_X1 U8571 ( .A1(n6940), .A2(n6939), .ZN(n6941) );
  NAND2_X1 U8572 ( .A1(n7386), .A2(n7995), .ZN(n6944) );
  NAND2_X1 U8573 ( .A1(n9043), .A2(n8004), .ZN(n6943) );
  NAND2_X1 U8574 ( .A1(n6944), .A2(n6943), .ZN(n6945) );
  XNOR2_X1 U8575 ( .A(n6945), .B(n8005), .ZN(n6948) );
  NAND2_X1 U8576 ( .A1(n7386), .A2(n8004), .ZN(n6947) );
  NAND2_X1 U8577 ( .A1(n9043), .A2(n8007), .ZN(n6946) );
  NAND2_X1 U8578 ( .A1(n6947), .A2(n6946), .ZN(n6949) );
  AND2_X1 U8579 ( .A1(n6948), .A2(n6949), .ZN(n6953) );
  INV_X1 U8580 ( .A(n6948), .ZN(n6951) );
  INV_X1 U8581 ( .A(n6949), .ZN(n6950) );
  NAND2_X1 U8582 ( .A1(n6951), .A2(n6950), .ZN(n7903) );
  INV_X1 U8583 ( .A(n7903), .ZN(n6955) );
  OAI21_X1 U8584 ( .B1(n6955), .B2(n6953), .A(n6952), .ZN(n6954) );
  OAI21_X1 U8585 ( .B1(n7904), .B2(n6955), .A(n6954), .ZN(n6956) );
  NAND2_X1 U8586 ( .A1(n6956), .A2(n9015), .ZN(n6967) );
  INV_X1 U8587 ( .A(n9300), .ZN(n6963) );
  NAND2_X1 U8588 ( .A1(n4414), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6962) );
  NAND2_X1 U8589 ( .A1(n7324), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6961) );
  INV_X1 U8590 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8910) );
  NAND2_X1 U8591 ( .A1(n6957), .A2(n8910), .ZN(n6958) );
  AND2_X1 U8592 ( .A1(n7020), .A2(n6958), .ZN(n8911) );
  NAND2_X1 U8593 ( .A1(n7459), .A2(n8911), .ZN(n6960) );
  NAND2_X1 U8594 ( .A1(n4417), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6959) );
  NAND4_X1 U8595 ( .A1(n6962), .A2(n6961), .A3(n6960), .A4(n6959), .ZN(n9292)
         );
  INV_X1 U8596 ( .A(n9292), .ZN(n9033) );
  OAI22_X1 U8597 ( .A1(n9010), .A2(n6963), .B1(n9009), .B2(n9033), .ZN(n6964)
         );
  AOI211_X1 U8598 ( .C1(n8978), .C2(n9044), .A(n6965), .B(n6964), .ZN(n6966)
         );
  OAI211_X1 U8599 ( .C1(n9302), .C2(n9024), .A(n6967), .B(n6966), .ZN(P1_U3232) );
  OAI21_X1 U8600 ( .B1(n6970), .B2(n6969), .A(n6968), .ZN(n6974) );
  INV_X1 U8601 ( .A(n7080), .ZN(n9795) );
  OAI22_X1 U8602 ( .A1(n8348), .A2(n9795), .B1(n8369), .B2(n7075), .ZN(n6973)
         );
  INV_X1 U8603 ( .A(n8387), .ZN(n7076) );
  NAND2_X1 U8604 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8076) );
  NAND2_X1 U8605 ( .A1(n8345), .A2(n7083), .ZN(n6971) );
  OAI211_X1 U8606 ( .C1(n8370), .C2(n7076), .A(n8076), .B(n6971), .ZN(n6972)
         );
  AOI211_X1 U8607 ( .C1(n6974), .C2(n8353), .A(n6973), .B(n6972), .ZN(n6975)
         );
  INV_X1 U8608 ( .A(n6975), .ZN(P2_U3233) );
  INV_X1 U8609 ( .A(n7351), .ZN(n7001) );
  AOI21_X1 U8610 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n7143), .A(n7867), .ZN(
        n6976) );
  OAI21_X1 U8611 ( .B1(n7001), .B2(n8236), .A(n6976), .ZN(P2_U3335) );
  NAND2_X1 U8612 ( .A1(n6887), .A2(n6977), .ZN(n6978) );
  XNOR2_X1 U8613 ( .A(n6978), .B(n7690), .ZN(n6980) );
  AOI21_X1 U8614 ( .B1(n6980), .B2(n9737), .A(n6979), .ZN(n9769) );
  INV_X1 U8615 ( .A(n6981), .ZN(n6982) );
  OAI22_X1 U8616 ( .A1(n9749), .A2(n9985), .B1(n6982), .B2(n9743), .ZN(n6986)
         );
  NOR2_X1 U8617 ( .A1(n8656), .A2(n7711), .ZN(n8672) );
  INV_X1 U8618 ( .A(n8672), .ZN(n6984) );
  OAI211_X1 U8619 ( .C1(n4676), .C2(n9770), .A(n9774), .B(n8738), .ZN(n9768)
         );
  NOR2_X1 U8620 ( .A1(n6984), .A2(n9768), .ZN(n6985) );
  AOI211_X1 U8621 ( .C1(n8749), .C2(n6987), .A(n6986), .B(n6985), .ZN(n6990)
         );
  XNOR2_X1 U8622 ( .A(n6988), .B(n7690), .ZN(n9772) );
  NAND2_X1 U8623 ( .A1(n9772), .A2(n8751), .ZN(n6989) );
  OAI211_X1 U8624 ( .C1(n9745), .C2(n9769), .A(n6990), .B(n6989), .ZN(P2_U3291) );
  XNOR2_X1 U8625 ( .A(n6992), .B(n6991), .ZN(n6997) );
  INV_X1 U8626 ( .A(n7137), .ZN(n6993) );
  NAND2_X1 U8627 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n8064) );
  OAI21_X1 U8628 ( .B1(n8368), .B2(n6993), .A(n8064), .ZN(n6995) );
  OAI22_X1 U8629 ( .A1(n9733), .A2(n8370), .B1(n8369), .B2(n7130), .ZN(n6994)
         );
  AOI211_X1 U8630 ( .C1(n7054), .C2(n8374), .A(n6995), .B(n6994), .ZN(n6996)
         );
  OAI21_X1 U8631 ( .B1(n6997), .B2(n8376), .A(n6996), .ZN(P2_U3219) );
  NAND2_X1 U8632 ( .A1(n9421), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7000) );
  INV_X1 U8633 ( .A(n6998), .ZN(n6999) );
  NAND2_X1 U8634 ( .A1(n6999), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7648) );
  OAI211_X1 U8635 ( .C1(n7001), .C2(n9424), .A(n7000), .B(n7648), .ZN(P1_U3330) );
  NAND2_X1 U8636 ( .A1(n7002), .A2(n9044), .ZN(n7005) );
  AND2_X1 U8637 ( .A1(n7003), .A2(n7005), .ZN(n7004) );
  INV_X1 U8638 ( .A(n7005), .ZN(n7008) );
  AND2_X1 U8639 ( .A1(n7006), .A2(n7485), .ZN(n7007) );
  AND2_X1 U8640 ( .A1(n7386), .A2(n9043), .ZN(n7009) );
  NAND2_X1 U8641 ( .A1(n7010), .A2(n7449), .ZN(n7012) );
  AOI22_X1 U8642 ( .A1(n7450), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7382), .B2(
        n9615), .ZN(n7011) );
  NAND2_X1 U8643 ( .A1(n8914), .A2(n9033), .ZN(n7563) );
  NAND2_X1 U8644 ( .A1(n8195), .A2(n7563), .ZN(n7471) );
  XNOR2_X1 U8645 ( .A(n8173), .B(n7471), .ZN(n9522) );
  INV_X1 U8646 ( .A(n9522), .ZN(n7034) );
  NAND2_X1 U8647 ( .A1(n7554), .A2(n7013), .ZN(n7014) );
  AND2_X1 U8648 ( .A1(n7014), .A2(n7557), .ZN(n7387) );
  XNOR2_X1 U8649 ( .A(n7386), .B(n9043), .ZN(n7486) );
  NAND2_X1 U8650 ( .A1(n7386), .A2(n7385), .ZN(n7392) );
  NAND2_X1 U8651 ( .A1(n7016), .A2(n7471), .ZN(n7017) );
  NAND3_X1 U8652 ( .A1(n8196), .A2(n9296), .A3(n7017), .ZN(n7027) );
  NAND2_X1 U8653 ( .A1(n4414), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7025) );
  NAND2_X1 U8654 ( .A1(n7324), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7024) );
  INV_X1 U8655 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7019) );
  NAND2_X1 U8656 ( .A1(n7020), .A2(n7019), .ZN(n7021) );
  AND2_X1 U8657 ( .A1(n7372), .A2(n7021), .ZN(n9286) );
  NAND2_X1 U8658 ( .A1(n7459), .A2(n9286), .ZN(n7023) );
  NAND2_X1 U8659 ( .A1(n4417), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7022) );
  NAND4_X1 U8660 ( .A1(n7025), .A2(n7024), .A3(n7023), .A4(n7022), .ZN(n9042)
         );
  AOI22_X1 U8661 ( .A1(n9293), .A2(n9042), .B1(n9043), .B2(n9291), .ZN(n7026)
         );
  NAND2_X1 U8662 ( .A1(n7027), .A2(n7026), .ZN(n9520) );
  INV_X1 U8663 ( .A(n8914), .ZN(n9518) );
  INV_X1 U8664 ( .A(n7028), .ZN(n7039) );
  NOR2_X1 U8665 ( .A1(n7028), .A2(n8914), .ZN(n7896) );
  INV_X1 U8666 ( .A(n7896), .ZN(n9285) );
  OAI211_X1 U8667 ( .C1(n9518), .C2(n7039), .A(n9285), .B(n9471), .ZN(n9517)
         );
  AOI22_X1 U8668 ( .A1(n4419), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8911), .B2(
        n9652), .ZN(n7030) );
  NAND2_X1 U8669 ( .A1(n8914), .A2(n9469), .ZN(n7029) );
  OAI211_X1 U8670 ( .C1(n9517), .C2(n7031), .A(n7030), .B(n7029), .ZN(n7032)
         );
  AOI21_X1 U8671 ( .B1(n9520), .B2(n9281), .A(n7032), .ZN(n7033) );
  OAI21_X1 U8672 ( .B1(n7034), .B2(n9308), .A(n7033), .ZN(P1_U3277) );
  XOR2_X1 U8673 ( .A(n7486), .B(n7035), .Z(n9309) );
  OAI21_X1 U8674 ( .B1(n7037), .B2(n7486), .A(n7036), .ZN(n7038) );
  AOI222_X1 U8675 ( .A1(n9296), .A2(n7038), .B1(n9292), .B2(n9293), .C1(n9044), 
        .C2(n9291), .ZN(n9303) );
  AOI21_X1 U8676 ( .B1(n7386), .B2(n7040), .A(n7039), .ZN(n9306) );
  AOI22_X1 U8677 ( .A1(n9306), .A2(n9471), .B1(n9392), .B2(n7386), .ZN(n7041)
         );
  OAI211_X1 U8678 ( .C1(n9309), .C2(n9396), .A(n9303), .B(n7041), .ZN(n7043)
         );
  NAND2_X1 U8679 ( .A1(n7043), .A2(n9702), .ZN(n7042) );
  OAI21_X1 U8680 ( .B1(n9702), .B2(n6257), .A(n7042), .ZN(P1_U3536) );
  INV_X1 U8681 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10045) );
  NAND2_X1 U8682 ( .A1(n7043), .A2(n9671), .ZN(n7044) );
  OAI21_X1 U8683 ( .B1(n9671), .B2(n10045), .A(n7044), .ZN(P1_U3493) );
  AND2_X2 U8684 ( .A1(n7045), .A2(n7761), .ZN(n9731) );
  NAND2_X1 U8685 ( .A1(n7076), .A2(n7062), .ZN(n7765) );
  NAND2_X1 U8686 ( .A1(n9733), .A2(n7080), .ZN(n7768) );
  INV_X1 U8687 ( .A(n9733), .ZN(n8386) );
  NAND2_X1 U8688 ( .A1(n8386), .A2(n9795), .ZN(n7771) );
  NAND2_X1 U8689 ( .A1(n7075), .A2(n7054), .ZN(n7773) );
  INV_X1 U8690 ( .A(n7075), .ZN(n8385) );
  NAND2_X1 U8691 ( .A1(n9802), .A2(n8385), .ZN(n7774) );
  NAND2_X1 U8692 ( .A1(n7773), .A2(n7774), .ZN(n7695) );
  INV_X1 U8693 ( .A(n7695), .ZN(n7046) );
  OR2_X1 U8694 ( .A1(n8334), .A2(n7130), .ZN(n7776) );
  NAND2_X1 U8695 ( .A1(n8334), .A2(n7130), .ZN(n7782) );
  NAND2_X1 U8696 ( .A1(n7776), .A2(n7782), .ZN(n7694) );
  XNOR2_X1 U8697 ( .A(n7089), .B(n7694), .ZN(n7049) );
  OR2_X1 U8698 ( .A1(n7163), .A2(n9732), .ZN(n7048) );
  OR2_X1 U8699 ( .A1(n7075), .A2(n9734), .ZN(n7047) );
  NAND2_X1 U8700 ( .A1(n7048), .A2(n7047), .ZN(n8333) );
  AOI21_X1 U8701 ( .B1(n7049), .B2(n9737), .A(n8333), .ZN(n9809) );
  INV_X1 U8702 ( .A(n9719), .ZN(n7052) );
  NAND2_X1 U8703 ( .A1(n8387), .A2(n7062), .ZN(n7053) );
  AND2_X1 U8704 ( .A1(n7054), .A2(n8385), .ZN(n7055) );
  OR2_X1 U8705 ( .A1(n7692), .A2(n7055), .ZN(n7093) );
  OR2_X1 U8706 ( .A1(n7113), .A2(n7093), .ZN(n7057) );
  NAND2_X1 U8707 ( .A1(n9733), .A2(n9795), .ZN(n7123) );
  OR2_X1 U8708 ( .A1(n7055), .A2(n7124), .ZN(n7056) );
  AND2_X1 U8709 ( .A1(n7057), .A2(n7056), .ZN(n7059) );
  NAND2_X1 U8710 ( .A1(n7057), .A2(n7094), .ZN(n7058) );
  OAI21_X1 U8711 ( .B1(n7059), .B2(n7694), .A(n7058), .ZN(n7060) );
  INV_X1 U8712 ( .A(n7060), .ZN(n9813) );
  NAND2_X1 U8713 ( .A1(n9813), .A2(n8751), .ZN(n7067) );
  INV_X1 U8714 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8055) );
  INV_X1 U8715 ( .A(n7061), .ZN(n8335) );
  OAI22_X1 U8716 ( .A1(n9749), .A2(n8055), .B1(n8335), .B2(n9743), .ZN(n7065)
         );
  INV_X1 U8717 ( .A(n8334), .ZN(n9811) );
  OAI211_X1 U8718 ( .C1(n7134), .C2(n9811), .A(n9774), .B(n4502), .ZN(n9808)
         );
  NOR2_X1 U8719 ( .A1(n9808), .A2(n7063), .ZN(n7064) );
  AOI211_X1 U8720 ( .C1(n8749), .C2(n8334), .A(n7065), .B(n7064), .ZN(n7066)
         );
  OAI211_X1 U8721 ( .C1(n9745), .C2(n9809), .A(n7067), .B(n7066), .ZN(P2_U3285) );
  INV_X1 U8722 ( .A(n7354), .ZN(n7070) );
  OAI222_X1 U8723 ( .A1(P2_U3152), .A2(n7069), .B1(n8236), .B2(n7070), .C1(
        n7068), .C2(n8881), .ZN(P2_U3334) );
  OAI222_X1 U8724 ( .A1(n8231), .A2(n10167), .B1(P1_U3084), .B2(n7071), .C1(
        n9424), .C2(n7070), .ZN(P1_U3329) );
  INV_X1 U8725 ( .A(n7125), .ZN(n7072) );
  AOI21_X1 U8726 ( .B1(n7692), .B2(n7113), .A(n7072), .ZN(n9794) );
  OR2_X1 U8727 ( .A1(n9745), .A2(n7073), .ZN(n9722) );
  XNOR2_X1 U8728 ( .A(n7074), .B(n7692), .ZN(n7078) );
  OAI22_X1 U8729 ( .A1(n7076), .A2(n9734), .B1(n7075), .B2(n9732), .ZN(n7077)
         );
  AOI21_X1 U8730 ( .B1(n7078), .B2(n9737), .A(n7077), .ZN(n7079) );
  OAI21_X1 U8731 ( .B1(n9794), .B2(n9740), .A(n7079), .ZN(n9797) );
  NAND2_X1 U8732 ( .A1(n9797), .A2(n9749), .ZN(n7088) );
  INV_X1 U8733 ( .A(n7136), .ZN(n7082) );
  NAND2_X1 U8734 ( .A1(n9724), .A2(n7080), .ZN(n7081) );
  NAND2_X1 U8735 ( .A1(n7082), .A2(n7081), .ZN(n9796) );
  INV_X1 U8736 ( .A(n9796), .ZN(n7086) );
  AOI22_X1 U8737 ( .A1(n8754), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7083), .B2(
        n8752), .ZN(n7084) );
  OAI21_X1 U8738 ( .B1(n9795), .B2(n9747), .A(n7084), .ZN(n7085) );
  AOI21_X1 U8739 ( .B1(n7086), .B2(n9727), .A(n7085), .ZN(n7087) );
  OAI211_X1 U8740 ( .C1(n9794), .C2(n9722), .A(n7088), .B(n7087), .ZN(P2_U3287) );
  NAND2_X1 U8741 ( .A1(n7110), .A2(n7776), .ZN(n7090) );
  OR2_X1 U8742 ( .A1(n9816), .A2(n7163), .ZN(n7786) );
  NAND2_X1 U8743 ( .A1(n9816), .A2(n7163), .ZN(n7787) );
  INV_X1 U8744 ( .A(n7698), .ZN(n7099) );
  XNOR2_X1 U8745 ( .A(n7090), .B(n7099), .ZN(n7092) );
  OAI22_X1 U8746 ( .A1(n7130), .A2(n9734), .B1(n7176), .B2(n9732), .ZN(n7091)
         );
  AOI21_X1 U8747 ( .B1(n7092), .B2(n9737), .A(n7091), .ZN(n9818) );
  INV_X1 U8748 ( .A(n7130), .ZN(n8384) );
  AND2_X1 U8749 ( .A1(n8334), .A2(n8384), .ZN(n7095) );
  OR2_X1 U8750 ( .A1(n7093), .A2(n7095), .ZN(n7112) );
  OR2_X1 U8751 ( .A1(n7113), .A2(n7112), .ZN(n7096) );
  OR2_X1 U8752 ( .A1(n7095), .A2(n7094), .ZN(n7114) );
  AND2_X1 U8753 ( .A1(n7096), .A2(n7114), .ZN(n7097) );
  INV_X1 U8754 ( .A(n7097), .ZN(n7100) );
  OR2_X1 U8755 ( .A1(n7097), .A2(n7698), .ZN(n7098) );
  OAI21_X1 U8756 ( .B1(n7100), .B2(n7099), .A(n7098), .ZN(n9823) );
  NAND2_X1 U8757 ( .A1(n9823), .A2(n8751), .ZN(n7108) );
  NAND2_X1 U8758 ( .A1(n4502), .A2(n9816), .ZN(n7101) );
  NAND2_X1 U8759 ( .A1(n7118), .A2(n7101), .ZN(n9819) );
  INV_X1 U8760 ( .A(n9819), .ZN(n7106) );
  INV_X1 U8761 ( .A(n7102), .ZN(n7152) );
  NOR2_X1 U8762 ( .A1(n9743), .A2(n7152), .ZN(n7103) );
  AOI21_X1 U8763 ( .B1(n9745), .B2(P2_REG2_REG_12__SCAN_IN), .A(n7103), .ZN(
        n7104) );
  OAI21_X1 U8764 ( .B1(n4688), .B2(n9747), .A(n7104), .ZN(n7105) );
  AOI21_X1 U8765 ( .B1(n7106), .B2(n9727), .A(n7105), .ZN(n7107) );
  OAI211_X1 U8766 ( .C1(n9745), .C2(n9818), .A(n7108), .B(n7107), .ZN(P2_U3284) );
  AND2_X1 U8767 ( .A1(n7786), .A2(n7776), .ZN(n7783) );
  INV_X1 U8768 ( .A(n7787), .ZN(n7109) );
  OR2_X1 U8769 ( .A1(n8855), .A2(n7176), .ZN(n7793) );
  NAND2_X1 U8770 ( .A1(n8855), .A2(n7176), .ZN(n7792) );
  NAND2_X1 U8771 ( .A1(n7793), .A2(n7792), .ZN(n7697) );
  XNOR2_X1 U8772 ( .A(n7202), .B(n7697), .ZN(n7111) );
  INV_X1 U8773 ( .A(n8371), .ZN(n8704) );
  INV_X1 U8774 ( .A(n7163), .ZN(n8383) );
  AOI222_X1 U8775 ( .A1(n9737), .A2(n7111), .B1(n8704), .B2(n8731), .C1(n8383), 
        .C2(n8729), .ZN(n8858) );
  OR2_X1 U8776 ( .A1(n9816), .A2(n8383), .ZN(n7115) );
  OR2_X1 U8777 ( .A1(n7117), .A2(n7697), .ZN(n8854) );
  NAND3_X1 U8778 ( .A1(n8854), .A2(n8751), .A3(n8853), .ZN(n7122) );
  AOI21_X1 U8779 ( .B1(n8855), .B2(n7118), .A(n8714), .ZN(n8856) );
  INV_X1 U8780 ( .A(n8855), .ZN(n7168) );
  AOI22_X1 U8781 ( .A1(n8754), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7165), .B2(
        n8752), .ZN(n7119) );
  OAI21_X1 U8782 ( .B1(n7168), .B2(n9747), .A(n7119), .ZN(n7120) );
  AOI21_X1 U8783 ( .B1(n8856), .B2(n9727), .A(n7120), .ZN(n7121) );
  OAI211_X1 U8784 ( .C1(n9745), .C2(n8858), .A(n7122), .B(n7121), .ZN(P2_U3283) );
  AND2_X1 U8785 ( .A1(n7125), .A2(n7123), .ZN(n7127) );
  NAND2_X1 U8786 ( .A1(n7125), .A2(n7124), .ZN(n7126) );
  OAI21_X1 U8787 ( .B1(n7127), .B2(n7695), .A(n7126), .ZN(n9801) );
  AOI21_X1 U8788 ( .B1(n7128), .B2(n7695), .A(n8620), .ZN(n7132) );
  OAI22_X1 U8789 ( .A1(n9733), .A2(n9734), .B1(n7130), .B2(n9732), .ZN(n7131)
         );
  AOI21_X1 U8790 ( .B1(n7132), .B2(n7129), .A(n7131), .ZN(n7133) );
  OAI21_X1 U8791 ( .B1(n9801), .B2(n9740), .A(n7133), .ZN(n9804) );
  NAND2_X1 U8792 ( .A1(n9804), .A2(n9749), .ZN(n7142) );
  INV_X1 U8793 ( .A(n7134), .ZN(n7135) );
  OAI21_X1 U8794 ( .B1(n9802), .B2(n7136), .A(n7135), .ZN(n9803) );
  INV_X1 U8795 ( .A(n9803), .ZN(n7140) );
  AOI22_X1 U8796 ( .A1(n8754), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7137), .B2(
        n8752), .ZN(n7138) );
  OAI21_X1 U8797 ( .B1(n9802), .B2(n9747), .A(n7138), .ZN(n7139) );
  AOI21_X1 U8798 ( .B1(n7140), .B2(n9727), .A(n7139), .ZN(n7141) );
  OAI211_X1 U8799 ( .C1(n9801), .C2(n9722), .A(n7142), .B(n7141), .ZN(P2_U3286) );
  INV_X1 U8800 ( .A(n7266), .ZN(n7170) );
  AOI22_X1 U8801 ( .A1(n7144), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n7143), .ZN(n7145) );
  OAI21_X1 U8802 ( .B1(n7170), .B2(n8236), .A(n7145), .ZN(P2_U3333) );
  NAND2_X1 U8803 ( .A1(n7158), .A2(n7156), .ZN(n7150) );
  NAND2_X1 U8804 ( .A1(n7147), .A2(n7146), .ZN(n8329) );
  NAND2_X1 U8805 ( .A1(n8329), .A2(n8330), .ZN(n7149) );
  NAND2_X1 U8806 ( .A1(n7149), .A2(n7148), .ZN(n7157) );
  XOR2_X1 U8807 ( .A(n7150), .B(n7157), .Z(n7155) );
  INV_X1 U8808 ( .A(n7176), .ZN(n8382) );
  AOI22_X1 U8809 ( .A1(n8316), .A2(n8384), .B1(n8315), .B2(n8382), .ZN(n7151)
         );
  NAND2_X1 U8810 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n8028) );
  OAI211_X1 U8811 ( .C1(n7152), .C2(n8368), .A(n7151), .B(n8028), .ZN(n7153)
         );
  AOI21_X1 U8812 ( .B1(n9816), .B2(n8374), .A(n7153), .ZN(n7154) );
  OAI21_X1 U8813 ( .B1(n7155), .B2(n8376), .A(n7154), .ZN(P2_U3226) );
  NAND2_X1 U8814 ( .A1(n7157), .A2(n7156), .ZN(n7159) );
  NAND2_X1 U8815 ( .A1(n7159), .A2(n7158), .ZN(n7162) );
  OAI211_X1 U8816 ( .C1(n7162), .C2(n7161), .A(n7160), .B(n8353), .ZN(n7167)
         );
  AND2_X1 U8817 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8152) );
  OAI22_X1 U8818 ( .A1(n7163), .A2(n8370), .B1(n8369), .B2(n8371), .ZN(n7164)
         );
  AOI211_X1 U8819 ( .C1(n8345), .C2(n7165), .A(n8152), .B(n7164), .ZN(n7166)
         );
  OAI211_X1 U8820 ( .C1(n7168), .C2(n8348), .A(n7167), .B(n7166), .ZN(P2_U3236) );
  OAI222_X1 U8821 ( .A1(n8231), .A2(n7171), .B1(n9424), .B2(n7170), .C1(n7169), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U8822 ( .A(n7172), .ZN(n7173) );
  AOI21_X1 U8823 ( .B1(n7175), .B2(n7174), .A(n7173), .ZN(n7184) );
  INV_X1 U8824 ( .A(n8717), .ZN(n7181) );
  OR2_X1 U8825 ( .A1(n8681), .A2(n9732), .ZN(n7178) );
  OR2_X1 U8826 ( .A1(n7176), .A2(n9734), .ZN(n7177) );
  NAND2_X1 U8827 ( .A1(n7178), .A2(n7177), .ZN(n8722) );
  NOR2_X1 U8828 ( .A1(n7179), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8143) );
  AOI21_X1 U8829 ( .B1(n8358), .B2(n8722), .A(n8143), .ZN(n7180) );
  OAI21_X1 U8830 ( .B1(n7181), .B2(n8368), .A(n7180), .ZN(n7182) );
  AOI21_X1 U8831 ( .B1(n8848), .B2(n8374), .A(n7182), .ZN(n7183) );
  OAI21_X1 U8832 ( .B1(n7184), .B2(n8376), .A(n7183), .ZN(P2_U3217) );
  INV_X1 U8833 ( .A(n7256), .ZN(n7188) );
  OAI222_X1 U8834 ( .A1(n8237), .A2(n7186), .B1(n8236), .B2(n7188), .C1(
        P2_U3152), .C2(n7185), .ZN(P2_U3332) );
  OAI222_X1 U8835 ( .A1(n8231), .A2(n9983), .B1(n9424), .B2(n7188), .C1(n7187), 
        .C2(P1_U3084), .ZN(P1_U3327) );
  INV_X1 U8836 ( .A(n7242), .ZN(n7215) );
  AOI21_X1 U8837 ( .B1(n9421), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7189), .ZN(
        n7190) );
  OAI21_X1 U8838 ( .B1(n7215), .B2(n9424), .A(n7190), .ZN(P1_U3326) );
  INV_X1 U8839 ( .A(n8680), .ZN(n8653) );
  NAND2_X1 U8840 ( .A1(n8855), .A2(n8382), .ZN(n7191) );
  OR2_X1 U8841 ( .A1(n8848), .A2(n8371), .ZN(n7796) );
  NAND2_X1 U8842 ( .A1(n8848), .A2(n8371), .ZN(n7797) );
  OR2_X1 U8843 ( .A1(n8848), .A2(n8704), .ZN(n7192) );
  OR2_X1 U8844 ( .A1(n8843), .A2(n8681), .ZN(n7801) );
  NAND2_X1 U8845 ( .A1(n8843), .A2(n8681), .ZN(n7800) );
  NAND2_X1 U8846 ( .A1(n7801), .A2(n7800), .ZN(n8702) );
  INV_X1 U8847 ( .A(n8681), .ZN(n8381) );
  NOR2_X1 U8848 ( .A1(n8843), .A2(n8381), .ZN(n7193) );
  OR2_X1 U8849 ( .A1(n8838), .A2(n8666), .ZN(n7804) );
  NAND2_X1 U8850 ( .A1(n8838), .A2(n8666), .ZN(n7717) );
  NAND2_X1 U8851 ( .A1(n7804), .A2(n7717), .ZN(n8682) );
  INV_X1 U8852 ( .A(n8666), .ZN(n8705) );
  NAND2_X1 U8853 ( .A1(n8835), .A2(n8680), .ZN(n7716) );
  NAND2_X1 U8854 ( .A1(n7715), .A2(n7716), .ZN(n8661) );
  NAND2_X1 U8855 ( .A1(n8828), .A2(n8669), .ZN(n7809) );
  INV_X1 U8856 ( .A(n8828), .ZN(n8649) );
  INV_X1 U8857 ( .A(n8824), .ZN(n8635) );
  NAND2_X1 U8858 ( .A1(n8818), .A2(n8257), .ZN(n7821) );
  NAND2_X1 U8859 ( .A1(n7816), .A2(n7821), .ZN(n8610) );
  INV_X1 U8860 ( .A(n8257), .ZN(n8604) );
  AOI21_X2 U8861 ( .B1(n8611), .B2(n8610), .A(n7194), .ZN(n8597) );
  NAND2_X1 U8862 ( .A1(n8597), .A2(n7195), .ZN(n7196) );
  NAND2_X1 U8863 ( .A1(n8808), .A2(n8248), .ZN(n7814) );
  NAND2_X1 U8864 ( .A1(n7824), .A2(n7814), .ZN(n8590) );
  AOI22_X1 U8865 ( .A1(n8581), .A2(n8590), .B1(n8587), .B2(n8248), .ZN(n8578)
         );
  OR2_X1 U8866 ( .A1(n8803), .A2(n8591), .ZN(n7829) );
  NAND2_X1 U8867 ( .A1(n8803), .A2(n8591), .ZN(n7713) );
  NAND2_X1 U8868 ( .A1(n7829), .A2(n7713), .ZN(n8577) );
  OAI21_X1 U8869 ( .B1(n4696), .B2(n8591), .A(n8801), .ZN(n8555) );
  NAND2_X1 U8870 ( .A1(n8796), .A2(n8570), .ZN(n7197) );
  NAND2_X1 U8871 ( .A1(n8792), .A2(n8561), .ZN(n7835) );
  NAND2_X1 U8872 ( .A1(n8787), .A2(n8275), .ZN(n7837) );
  INV_X1 U8873 ( .A(n8787), .ZN(n8527) );
  AOI22_X1 U8874 ( .A1(n8521), .A2(n8529), .B1(n8527), .B2(n8275), .ZN(n8508)
         );
  NAND2_X1 U8875 ( .A1(n8781), .A2(n8357), .ZN(n7844) );
  AND2_X2 U8876 ( .A1(n7843), .A2(n7844), .ZN(n8512) );
  NAND2_X1 U8877 ( .A1(n8776), .A2(n8494), .ZN(n7846) );
  XNOR2_X1 U8878 ( .A(n8487), .B(n7207), .ZN(n8780) );
  INV_X1 U8879 ( .A(n8848), .ZN(n8719) );
  INV_X1 U8880 ( .A(n8843), .ZN(n8701) );
  INV_X1 U8881 ( .A(n8818), .ZN(n8616) );
  INV_X1 U8882 ( .A(n8792), .ZN(n8549) );
  AOI21_X1 U8883 ( .B1(n8776), .B2(n4682), .A(n8498), .ZN(n8777) );
  INV_X1 U8884 ( .A(n7199), .ZN(n7200) );
  AOI22_X1 U8885 ( .A1(n8754), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n7200), .B2(
        n8752), .ZN(n7201) );
  OAI21_X1 U8886 ( .B1(n8485), .B2(n9747), .A(n7201), .ZN(n7212) );
  INV_X1 U8887 ( .A(n7717), .ZN(n7203) );
  NAND2_X1 U8888 ( .A1(n8665), .A2(n4645), .ZN(n8664) );
  NOR2_X1 U8889 ( .A1(n8824), .A2(n8624), .ZN(n7815) );
  NOR2_X1 U8890 ( .A1(n7815), .A2(n7818), .ZN(n8638) );
  INV_X1 U8891 ( .A(n8610), .ZN(n8618) );
  INV_X1 U8892 ( .A(n7816), .ZN(n7204) );
  XNOR2_X1 U8893 ( .A(n8813), .B(n8380), .ZN(n8602) );
  NAND2_X1 U8894 ( .A1(n8813), .A2(n8623), .ZN(n7820) );
  INV_X1 U8895 ( .A(n7824), .ZN(n7205) );
  INV_X1 U8896 ( .A(n8577), .ZN(n8569) );
  NAND2_X1 U8897 ( .A1(n8567), .A2(n7713), .ZN(n8560) );
  NOR2_X1 U8898 ( .A1(n8796), .A2(n8274), .ZN(n8537) );
  INV_X1 U8899 ( .A(n7208), .ZN(n7206) );
  AOI21_X1 U8900 ( .B1(n7206), .B2(n8486), .A(n8620), .ZN(n7210) );
  OAI22_X1 U8901 ( .A1(n7668), .A2(n9732), .B1(n8357), .B2(n9734), .ZN(n7209)
         );
  AOI21_X1 U8902 ( .B1(n7210), .B2(n7664), .A(n7209), .ZN(n8779) );
  NOR2_X1 U8903 ( .A1(n8779), .A2(n9745), .ZN(n7211) );
  AOI211_X1 U8904 ( .C1(n9727), .C2(n8777), .A(n7212), .B(n7211), .ZN(n7213)
         );
  OAI21_X1 U8905 ( .B1(n8780), .B2(n8727), .A(n7213), .ZN(P2_U3268) );
  OAI222_X1 U8906 ( .A1(n8237), .A2(n10091), .B1(n8236), .B2(n7215), .C1(n7214), .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U8907 ( .A(n7218), .ZN(n7219) );
  INV_X1 U8908 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8226) );
  INV_X1 U8909 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10079) );
  MUX2_X1 U8910 ( .A(n8226), .B(n10079), .S(n7220), .Z(n7446) );
  INV_X1 U8911 ( .A(SI_29_), .ZN(n9977) );
  AND2_X1 U8912 ( .A1(n7446), .A2(n9977), .ZN(n7223) );
  INV_X1 U8913 ( .A(n7446), .ZN(n7221) );
  NAND2_X1 U8914 ( .A1(n7221), .A2(SI_29_), .ZN(n7222) );
  MUX2_X1 U8915 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7229), .Z(n7225) );
  INV_X1 U8916 ( .A(n7235), .ZN(n7224) );
  NAND2_X1 U8917 ( .A1(n7224), .A2(SI_30_), .ZN(n7228) );
  NAND2_X1 U8918 ( .A1(n7226), .A2(n7225), .ZN(n7227) );
  NAND2_X1 U8919 ( .A1(n7228), .A2(n7227), .ZN(n7232) );
  MUX2_X1 U8920 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7229), .Z(n7230) );
  XNOR2_X1 U8921 ( .A(n7230), .B(SI_31_), .ZN(n7231) );
  XNOR2_X2 U8922 ( .A(n7232), .B(n7231), .ZN(n8879) );
  NAND2_X1 U8923 ( .A1(n8879), .A2(n7449), .ZN(n7234) );
  NAND2_X1 U8924 ( .A1(n6348), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7233) );
  INV_X1 U8925 ( .A(n7899), .ZN(n7522) );
  NAND2_X1 U8926 ( .A1(n7521), .A2(n7522), .ZN(n7628) );
  NAND2_X1 U8927 ( .A1(n8228), .A2(n7449), .ZN(n7237) );
  NAND2_X1 U8928 ( .A1(n6348), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7236) );
  NAND2_X1 U8929 ( .A1(n4414), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7240) );
  NAND2_X1 U8930 ( .A1(n4417), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7239) );
  NAND2_X1 U8931 ( .A1(n7324), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7238) );
  NAND3_X1 U8932 ( .A1(n7240), .A2(n7239), .A3(n7238), .ZN(n9040) );
  INV_X1 U8933 ( .A(n9040), .ZN(n7460) );
  NOR2_X1 U8934 ( .A1(n9075), .A2(n7460), .ZN(n7523) );
  INV_X1 U8935 ( .A(n7523), .ZN(n7241) );
  NAND2_X1 U8936 ( .A1(n7628), .A2(n7241), .ZN(n7496) );
  INV_X1 U8937 ( .A(n7496), .ZN(n7465) );
  NAND2_X1 U8938 ( .A1(n7242), .A2(n7449), .ZN(n7244) );
  NAND2_X1 U8939 ( .A1(n7450), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7243) );
  NAND2_X2 U8940 ( .A1(n7244), .A2(n7243), .ZN(n9328) );
  INV_X1 U8941 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8972) );
  INV_X1 U8942 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7330) );
  INV_X1 U8943 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n7280) );
  INV_X1 U8944 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n7357) );
  INV_X1 U8945 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8955) );
  XNOR2_X1 U8946 ( .A(n7432), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U8947 ( .A1(n9101), .A2(n7459), .ZN(n7255) );
  INV_X1 U8948 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10171) );
  NAND2_X1 U8949 ( .A1(n4414), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7252) );
  NAND2_X1 U8950 ( .A1(n4416), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7251) );
  OAI211_X1 U8951 ( .C1(n7314), .C2(n10171), .A(n7252), .B(n7251), .ZN(n7253)
         );
  INV_X1 U8952 ( .A(n7253), .ZN(n7254) );
  INV_X1 U8953 ( .A(n9117), .ZN(n7427) );
  INV_X1 U8954 ( .A(n7615), .ZN(n8216) );
  NAND2_X1 U8955 ( .A1(n7256), .A2(n7449), .ZN(n7258) );
  NAND2_X1 U8956 ( .A1(n7450), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7257) );
  INV_X1 U8957 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n7259) );
  NAND2_X1 U8958 ( .A1(n7270), .A2(n7259), .ZN(n7260) );
  NAND2_X1 U8959 ( .A1(n7432), .A2(n7260), .ZN(n9019) );
  INV_X1 U8960 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10146) );
  NAND2_X1 U8961 ( .A1(n4417), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7262) );
  NAND2_X1 U8962 ( .A1(n7324), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7261) );
  OAI211_X1 U8963 ( .C1(n6097), .C2(n10146), .A(n7262), .B(n7261), .ZN(n7263)
         );
  INV_X1 U8964 ( .A(n7263), .ZN(n7264) );
  OR2_X1 U8965 ( .A1(n9332), .A2(n9096), .ZN(n7612) );
  NAND2_X1 U8966 ( .A1(n7266), .A2(n7449), .ZN(n7268) );
  NAND2_X1 U8967 ( .A1(n7450), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7267) );
  NAND2_X1 U8968 ( .A1(n7360), .A2(n8955), .ZN(n7269) );
  NAND2_X1 U8969 ( .A1(n9125), .A2(n7459), .ZN(n7276) );
  INV_X1 U8970 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n7273) );
  NAND2_X1 U8971 ( .A1(n4414), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n7272) );
  NAND2_X1 U8972 ( .A1(n7324), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7271) );
  OAI211_X1 U8973 ( .C1(n7273), .C2(n7456), .A(n7272), .B(n7271), .ZN(n7274)
         );
  INV_X1 U8974 ( .A(n7274), .ZN(n7275) );
  NAND2_X1 U8975 ( .A1(n7612), .A2(n9113), .ZN(n8215) );
  OR2_X1 U8976 ( .A1(n8216), .A2(n8215), .ZN(n7516) );
  INV_X1 U8977 ( .A(n7516), .ZN(n7445) );
  NAND2_X1 U8978 ( .A1(n7277), .A2(n7449), .ZN(n7279) );
  NAND2_X1 U8979 ( .A1(n7450), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7278) );
  NAND2_X1 U8980 ( .A1(n7292), .A2(n7280), .ZN(n7281) );
  AND2_X1 U8981 ( .A1(n7301), .A2(n7281), .ZN(n9185) );
  NAND2_X1 U8982 ( .A1(n9185), .A2(n7459), .ZN(n7287) );
  INV_X1 U8983 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n7284) );
  NAND2_X1 U8984 ( .A1(n7324), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7283) );
  NAND2_X1 U8985 ( .A1(n4414), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n7282) );
  OAI211_X1 U8986 ( .C1(n7456), .C2(n7284), .A(n7283), .B(n7282), .ZN(n7285)
         );
  INV_X1 U8987 ( .A(n7285), .ZN(n7286) );
  NAND2_X1 U8988 ( .A1(n7287), .A2(n7286), .ZN(n9177) );
  INV_X1 U8989 ( .A(n7596), .ZN(n7309) );
  NAND2_X1 U8990 ( .A1(n7288), .A2(n7449), .ZN(n7290) );
  NAND2_X1 U8991 ( .A1(n7450), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7289) );
  INV_X1 U8992 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U8993 ( .A1(n7333), .A2(n8989), .ZN(n7291) );
  NAND2_X1 U8994 ( .A1(n7292), .A2(n7291), .ZN(n9209) );
  OR2_X1 U8995 ( .A1(n9209), .A2(n7434), .ZN(n7297) );
  INV_X1 U8996 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10062) );
  NAND2_X1 U8997 ( .A1(n7324), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7294) );
  NAND2_X1 U8998 ( .A1(n4414), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n7293) );
  OAI211_X1 U8999 ( .C1(n7456), .C2(n10062), .A(n7294), .B(n7293), .ZN(n7295)
         );
  INV_X1 U9000 ( .A(n7295), .ZN(n7296) );
  NAND2_X1 U9001 ( .A1(n7297), .A2(n7296), .ZN(n9228) );
  INV_X1 U9002 ( .A(n9228), .ZN(n9192) );
  AND2_X1 U9003 ( .A1(n9368), .A2(n9192), .ZN(n7585) );
  INV_X1 U9004 ( .A(n7585), .ZN(n7308) );
  NAND2_X1 U9005 ( .A1(n7298), .A2(n7449), .ZN(n7300) );
  NAND2_X1 U9006 ( .A1(n7450), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7299) );
  INV_X1 U9007 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9000) );
  NAND2_X1 U9008 ( .A1(n7301), .A2(n9000), .ZN(n7302) );
  NAND2_X1 U9009 ( .A1(n7343), .A2(n7302), .ZN(n9170) );
  OR2_X1 U9010 ( .A1(n9170), .A2(n7434), .ZN(n7307) );
  INV_X1 U9011 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10096) );
  NAND2_X1 U9012 ( .A1(n4414), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n7304) );
  NAND2_X1 U9013 ( .A1(n4416), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n7303) );
  OAI211_X1 U9014 ( .C1(n7314), .C2(n10096), .A(n7304), .B(n7303), .ZN(n7305)
         );
  INV_X1 U9015 ( .A(n7305), .ZN(n7306) );
  NAND2_X1 U9016 ( .A1(n7307), .A2(n7306), .ZN(n9162) );
  INV_X1 U9017 ( .A(n8209), .ZN(n9156) );
  NAND2_X1 U9018 ( .A1(n9362), .A2(n9207), .ZN(n8206) );
  OAI211_X1 U9019 ( .C1(n7309), .C2(n7308), .A(n9156), .B(n8206), .ZN(n7419)
         );
  INV_X1 U9020 ( .A(n7419), .ZN(n7595) );
  NAND2_X1 U9021 ( .A1(n7310), .A2(n7449), .ZN(n7312) );
  AOI22_X1 U9022 ( .A1(n7450), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7382), .B2(
        n9059), .ZN(n7311) );
  NAND2_X1 U9023 ( .A1(n7374), .A2(n8972), .ZN(n7313) );
  NAND2_X1 U9024 ( .A1(n7322), .A2(n7313), .ZN(n9259) );
  INV_X1 U9025 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9260) );
  OAI22_X1 U9026 ( .A1(n9259), .A2(n7434), .B1(n7456), .B2(n9260), .ZN(n7317)
         );
  INV_X1 U9027 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7315) );
  INV_X1 U9028 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10106) );
  OAI22_X1 U9029 ( .A1(n6097), .A2(n7315), .B1(n7314), .B2(n10106), .ZN(n7316)
         );
  NOR2_X1 U9030 ( .A1(n9383), .A2(n9271), .ZN(n8200) );
  NAND2_X1 U9031 ( .A1(n7318), .A2(n7449), .ZN(n7320) );
  AOI22_X1 U9032 ( .A1(n7450), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7382), .B2(
        n9636), .ZN(n7319) );
  INV_X1 U9033 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10158) );
  INV_X1 U9034 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7321) );
  NAND2_X1 U9035 ( .A1(n7322), .A2(n7321), .ZN(n7323) );
  NAND2_X1 U9036 ( .A1(n7331), .A2(n7323), .ZN(n9245) );
  OR2_X1 U9037 ( .A1(n9245), .A2(n7434), .ZN(n7326) );
  AOI22_X1 U9038 ( .A1(n4416), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n7324), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n7325) );
  OAI211_X1 U9039 ( .C1(n6097), .C2(n10158), .A(n7326), .B(n7325), .ZN(n9227)
         );
  INV_X1 U9040 ( .A(n9227), .ZN(n9254) );
  OR2_X1 U9041 ( .A1(n9377), .A2(n9254), .ZN(n7582) );
  NAND2_X1 U9042 ( .A1(n4592), .A2(n7582), .ZN(n7579) );
  INV_X1 U9043 ( .A(n7579), .ZN(n7340) );
  NAND2_X1 U9044 ( .A1(n7327), .A2(n7449), .ZN(n7329) );
  AOI22_X1 U9045 ( .A1(n7450), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7661), .B2(
        n7382), .ZN(n7328) );
  NAND2_X1 U9046 ( .A1(n7331), .A2(n7330), .ZN(n7332) );
  NAND2_X1 U9047 ( .A1(n7333), .A2(n7332), .ZN(n9220) );
  AOI22_X1 U9048 ( .A1(n4414), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n7324), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n7336) );
  INV_X1 U9049 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n7334) );
  OR2_X1 U9050 ( .A1(n7456), .A2(n7334), .ZN(n7335) );
  OAI211_X1 U9051 ( .C1(n9220), .C2(n7434), .A(n7336), .B(n7335), .ZN(n9240)
         );
  INV_X1 U9052 ( .A(n9240), .ZN(n9206) );
  NAND2_X1 U9053 ( .A1(n9377), .A2(n9254), .ZN(n8202) );
  NOR2_X1 U9054 ( .A1(n8203), .A2(n4589), .ZN(n7587) );
  INV_X1 U9055 ( .A(n7587), .ZN(n7339) );
  NOR2_X1 U9056 ( .A1(n9368), .A2(n9192), .ZN(n7468) );
  INV_X1 U9057 ( .A(n7468), .ZN(n8204) );
  NOR2_X1 U9058 ( .A1(n9372), .A2(n9206), .ZN(n7583) );
  INV_X1 U9059 ( .A(n7583), .ZN(n7337) );
  NAND2_X1 U9060 ( .A1(n8204), .A2(n7337), .ZN(n7589) );
  INV_X1 U9061 ( .A(n7589), .ZN(n7338) );
  OAI21_X1 U9062 ( .B1(n7340), .B2(n7339), .A(n7338), .ZN(n7366) );
  OR2_X1 U9063 ( .A1(n7419), .A2(n7596), .ZN(n7342) );
  NOR2_X1 U9064 ( .A1(n9354), .A2(n9191), .ZN(n8208) );
  INV_X1 U9065 ( .A(n8208), .ZN(n7341) );
  NAND2_X1 U9066 ( .A1(n7342), .A2(n7341), .ZN(n7594) );
  INV_X1 U9067 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8921) );
  NAND2_X1 U9068 ( .A1(n7343), .A2(n8921), .ZN(n7344) );
  NAND2_X1 U9069 ( .A1(n7358), .A2(n7344), .ZN(n9152) );
  OR2_X1 U9070 ( .A1(n9152), .A2(n7434), .ZN(n7350) );
  INV_X1 U9071 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n7347) );
  NAND2_X1 U9072 ( .A1(n7324), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n7346) );
  NAND2_X1 U9073 ( .A1(n4414), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n7345) );
  OAI211_X1 U9074 ( .C1(n7347), .C2(n7456), .A(n7346), .B(n7345), .ZN(n7348)
         );
  INV_X1 U9075 ( .A(n7348), .ZN(n7349) );
  NAND2_X1 U9076 ( .A1(n7350), .A2(n7349), .ZN(n9176) );
  INV_X1 U9077 ( .A(n9176), .ZN(n9142) );
  NAND2_X1 U9078 ( .A1(n7351), .A2(n7449), .ZN(n7353) );
  NAND2_X1 U9079 ( .A1(n7450), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7352) );
  NAND2_X1 U9080 ( .A1(n7354), .A2(n7449), .ZN(n7356) );
  NAND2_X1 U9081 ( .A1(n7450), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7355) );
  NAND2_X1 U9082 ( .A1(n7358), .A2(n7357), .ZN(n7359) );
  NAND2_X1 U9083 ( .A1(n7360), .A2(n7359), .ZN(n9137) );
  INV_X1 U9084 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n10188) );
  NAND2_X1 U9085 ( .A1(n7324), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7362) );
  NAND2_X1 U9086 ( .A1(n4414), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n7361) );
  OAI211_X1 U9087 ( .C1(n7456), .C2(n10188), .A(n7362), .B(n7361), .ZN(n7363)
         );
  INV_X1 U9088 ( .A(n7363), .ZN(n7364) );
  NAND2_X1 U9089 ( .A1(n7365), .A2(n7364), .ZN(n9161) );
  INV_X1 U9090 ( .A(n9161), .ZN(n8956) );
  OAI21_X1 U9091 ( .B1(n9142), .B2(n9349), .A(n4799), .ZN(n7604) );
  AOI211_X1 U9092 ( .C1(n7595), .C2(n7366), .A(n7594), .B(n7604), .ZN(n7514)
         );
  INV_X1 U9093 ( .A(n7514), .ZN(n7426) );
  NAND2_X1 U9094 ( .A1(n7367), .A2(n7449), .ZN(n7369) );
  AOI22_X1 U9095 ( .A1(n7450), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7382), .B2(
        n7655), .ZN(n7368) );
  NAND2_X1 U9096 ( .A1(n7324), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7378) );
  NAND2_X1 U9097 ( .A1(n4417), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7377) );
  INV_X1 U9098 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7371) );
  NAND2_X1 U9099 ( .A1(n7372), .A2(n7371), .ZN(n7373) );
  AND2_X1 U9100 ( .A1(n7374), .A2(n7373), .ZN(n9276) );
  NAND2_X1 U9101 ( .A1(n7459), .A2(n9276), .ZN(n7376) );
  NAND2_X1 U9102 ( .A1(n4414), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7375) );
  NAND4_X1 U9103 ( .A1(n7378), .A2(n7377), .A3(n7376), .A4(n7375), .ZN(n9294)
         );
  INV_X1 U9104 ( .A(n9294), .ZN(n9253) );
  OR2_X1 U9105 ( .A1(n9388), .A2(n9253), .ZN(n7574) );
  NAND2_X1 U9106 ( .A1(n7379), .A2(n7449), .ZN(n7384) );
  INV_X1 U9107 ( .A(n7380), .ZN(n7381) );
  AOI22_X1 U9108 ( .A1(n7450), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7382), .B2(
        n7381), .ZN(n7383) );
  INV_X1 U9109 ( .A(n9042), .ZN(n9272) );
  OR2_X1 U9110 ( .A1(n9391), .A2(n9272), .ZN(n9266) );
  AND2_X1 U9111 ( .A1(n7574), .A2(n9266), .ZN(n8199) );
  OR2_X1 U9112 ( .A1(n7386), .A2(n7385), .ZN(n7565) );
  NAND2_X1 U9113 ( .A1(n7387), .A2(n7565), .ZN(n7555) );
  INV_X1 U9114 ( .A(n7555), .ZN(n7394) );
  INV_X1 U9115 ( .A(n7388), .ZN(n7541) );
  NOR2_X1 U9116 ( .A1(n7542), .A2(n7541), .ZN(n7544) );
  INV_X1 U9117 ( .A(n7544), .ZN(n7391) );
  NAND2_X1 U9118 ( .A1(n7554), .A2(n7389), .ZN(n7558) );
  NOR2_X1 U9119 ( .A1(n7547), .A2(n4788), .ZN(n7390) );
  NOR2_X1 U9120 ( .A1(n7558), .A2(n7390), .ZN(n7414) );
  OAI21_X1 U9121 ( .B1(n4788), .B2(n7391), .A(n7414), .ZN(n7393) );
  NAND2_X1 U9122 ( .A1(n7563), .A2(n7392), .ZN(n7556) );
  AOI21_X1 U9123 ( .B1(n7394), .B2(n7393), .A(n7556), .ZN(n7395) );
  INV_X1 U9124 ( .A(n8195), .ZN(n7561) );
  NAND2_X1 U9125 ( .A1(n9391), .A2(n9272), .ZN(n8197) );
  OAI21_X1 U9126 ( .B1(n7395), .B2(n7561), .A(n8197), .ZN(n7397) );
  NAND2_X1 U9127 ( .A1(n9383), .A2(n9271), .ZN(n8201) );
  INV_X1 U9128 ( .A(n8201), .ZN(n7469) );
  NAND2_X1 U9129 ( .A1(n9388), .A2(n9253), .ZN(n7470) );
  INV_X1 U9130 ( .A(n7470), .ZN(n8198) );
  NOR3_X1 U9131 ( .A1(n4589), .A2(n7469), .A3(n8198), .ZN(n7415) );
  INV_X1 U9132 ( .A(n7415), .ZN(n7396) );
  AOI21_X1 U9133 ( .B1(n8199), .B2(n7397), .A(n7396), .ZN(n7512) );
  INV_X1 U9134 ( .A(n7512), .ZN(n7422) );
  INV_X1 U9135 ( .A(n7398), .ZN(n7399) );
  OAI211_X1 U9136 ( .C1(n7401), .C2(n7400), .A(n5807), .B(n7399), .ZN(n7403)
         );
  NAND2_X1 U9137 ( .A1(n7403), .A2(n7402), .ZN(n7406) );
  OAI22_X1 U9138 ( .A1(n7407), .A2(n7406), .B1(n7405), .B2(n7404), .ZN(n7410)
         );
  AND2_X1 U9139 ( .A1(n7499), .A2(n7408), .ZN(n7504) );
  INV_X1 U9140 ( .A(n7504), .ZN(n7409) );
  AOI21_X1 U9141 ( .B1(n7410), .B2(n7498), .A(n7409), .ZN(n7412) );
  OAI21_X1 U9142 ( .B1(n7412), .B2(n4584), .A(n7503), .ZN(n7418) );
  NAND2_X1 U9143 ( .A1(n7537), .A2(n7413), .ZN(n7539) );
  INV_X1 U9144 ( .A(n7556), .ZN(n7562) );
  NAND4_X1 U9145 ( .A1(n7415), .A2(n7562), .A3(n7414), .A4(n7538), .ZN(n7509)
         );
  INV_X1 U9146 ( .A(n7509), .ZN(n7417) );
  NAND2_X1 U9147 ( .A1(n8197), .A2(n7540), .ZN(n7507) );
  INV_X1 U9148 ( .A(n7507), .ZN(n7416) );
  OAI211_X1 U9149 ( .C1(n7418), .C2(n7539), .A(n7417), .B(n7416), .ZN(n7421)
         );
  NOR2_X1 U9150 ( .A1(n7419), .A2(n8203), .ZN(n7510) );
  INV_X1 U9151 ( .A(n7510), .ZN(n7420) );
  AOI21_X1 U9152 ( .B1(n7422), .B2(n7421), .A(n7420), .ZN(n7425) );
  INV_X1 U9153 ( .A(n7605), .ZN(n7423) );
  NAND2_X1 U9154 ( .A1(n9349), .A2(n9142), .ZN(n9138) );
  NAND2_X1 U9155 ( .A1(n9337), .A2(n9141), .ZN(n8212) );
  OAI21_X1 U9156 ( .B1(n8210), .B2(n8211), .A(n8212), .ZN(n7607) );
  INV_X1 U9157 ( .A(n7607), .ZN(n7424) );
  OAI21_X1 U9158 ( .B1(n7426), .B2(n7425), .A(n7424), .ZN(n7444) );
  NAND2_X1 U9159 ( .A1(n9332), .A2(n9096), .ZN(n8214) );
  NAND2_X1 U9160 ( .A1(n9328), .A2(n7427), .ZN(n7616) );
  INV_X1 U9161 ( .A(n7616), .ZN(n7442) );
  NAND2_X1 U9162 ( .A1(n8235), .A2(n7449), .ZN(n7429) );
  NAND2_X1 U9163 ( .A1(n6348), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n7428) );
  NAND2_X2 U9164 ( .A1(n7429), .A2(n7428), .ZN(n9322) );
  INV_X1 U9165 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7431) );
  INV_X1 U9166 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7430) );
  OAI21_X1 U9167 ( .B1(n7432), .B2(n7431), .A(n7430), .ZN(n7433) );
  NAND2_X1 U9168 ( .A1(n7433), .A2(n7453), .ZN(n8011) );
  INV_X1 U9169 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n7437) );
  NAND2_X1 U9170 ( .A1(n4414), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n7436) );
  NAND2_X1 U9171 ( .A1(n7324), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7435) );
  OAI211_X1 U9172 ( .C1(n7437), .C2(n7456), .A(n7436), .B(n7435), .ZN(n7438)
         );
  INV_X1 U9173 ( .A(n7438), .ZN(n7439) );
  NAND2_X1 U9174 ( .A1(n9322), .A2(n9097), .ZN(n8217) );
  INV_X1 U9175 ( .A(n8217), .ZN(n7441) );
  AOI211_X1 U9176 ( .C1(n4791), .C2(n7615), .A(n7442), .B(n7441), .ZN(n7515)
         );
  INV_X1 U9177 ( .A(n7515), .ZN(n7443) );
  AOI21_X1 U9178 ( .B1(n7445), .B2(n7444), .A(n7443), .ZN(n7462) );
  XNOR2_X1 U9179 ( .A(n7446), .B(SI_29_), .ZN(n7447) );
  NAND2_X1 U9180 ( .A1(n8225), .A2(n7449), .ZN(n7452) );
  NAND2_X1 U9181 ( .A1(n7450), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7451) );
  INV_X1 U9182 ( .A(n7453), .ZN(n8190) );
  INV_X1 U9183 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n7457) );
  NAND2_X1 U9184 ( .A1(n7324), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7455) );
  NAND2_X1 U9185 ( .A1(n4414), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7454) );
  OAI211_X1 U9186 ( .C1(n7457), .C2(n7456), .A(n7455), .B(n7454), .ZN(n7458)
         );
  AOI21_X1 U9187 ( .B1(n8190), .B2(n7459), .A(n7458), .ZN(n8014) );
  NAND2_X1 U9188 ( .A1(n9075), .A2(n7460), .ZN(n7494) );
  INV_X1 U9189 ( .A(n8014), .ZN(n9089) );
  INV_X1 U9190 ( .A(n7622), .ZN(n7461) );
  OAI211_X1 U9191 ( .C1(n7462), .C2(n7619), .A(n7494), .B(n7461), .ZN(n7464)
         );
  NAND2_X2 U9192 ( .A1(n9311), .A2(n7899), .ZN(n7632) );
  INV_X1 U9193 ( .A(n7632), .ZN(n7463) );
  AOI21_X1 U9194 ( .B1(n7465), .B2(n7464), .A(n7463), .ZN(n7466) );
  XNOR2_X1 U9195 ( .A(n7466), .B(n9243), .ZN(n7640) );
  INV_X1 U9196 ( .A(n9088), .ZN(n7493) );
  NAND2_X1 U9197 ( .A1(n9113), .A2(n8212), .ZN(n9129) );
  NOR2_X1 U9198 ( .A1(n7468), .A2(n7585), .ZN(n9204) );
  NAND2_X1 U9199 ( .A1(n9266), .A2(n8197), .ZN(n9289) );
  NAND2_X1 U9200 ( .A1(n7574), .A2(n7470), .ZN(n9269) );
  NAND4_X1 U9201 ( .A1(n7475), .A2(n7474), .A3(n7473), .A4(n7472), .ZN(n7478)
         );
  NOR4_X1 U9202 ( .A1(n7478), .A2(n6345), .A3(n7535), .A4(n7477), .ZN(n7482)
         );
  INV_X1 U9203 ( .A(n7479), .ZN(n7480) );
  NAND3_X1 U9204 ( .A1(n7482), .A2(n7481), .A3(n7480), .ZN(n7483) );
  NOR4_X1 U9205 ( .A1(n7485), .A2(n9454), .A3(n7484), .A4(n7483), .ZN(n7487)
         );
  NAND4_X1 U9206 ( .A1(n4525), .A2(n7487), .A3(n7552), .A4(n7486), .ZN(n7488)
         );
  NOR4_X1 U9207 ( .A1(n9251), .A2(n9289), .A3(n9269), .A4(n7488), .ZN(n7489)
         );
  NAND4_X1 U9208 ( .A1(n9204), .A2(n9226), .A3(n9238), .A4(n7489), .ZN(n7490)
         );
  NOR3_X1 U9209 ( .A1(n9174), .A2(n9189), .A3(n7490), .ZN(n7491) );
  XNOR2_X1 U9210 ( .A(n9349), .B(n9176), .ZN(n9155) );
  NAND4_X1 U9211 ( .A1(n9115), .A2(n9144), .A3(n7491), .A4(n9155), .ZN(n7492)
         );
  NAND4_X1 U9212 ( .A1(n7632), .A2(n8218), .A3(n7495), .A4(n7494), .ZN(n7497)
         );
  OAI21_X1 U9213 ( .B1(n7497), .B2(n7496), .A(n7630), .ZN(n7528) );
  INV_X1 U9214 ( .A(n7619), .ZN(n7520) );
  INV_X1 U9215 ( .A(n7498), .ZN(n7502) );
  NAND3_X1 U9216 ( .A1(n7536), .A2(n4583), .A3(n7500), .ZN(n7501) );
  OAI211_X1 U9217 ( .C1(n4584), .C2(n7502), .A(n7503), .B(n7501), .ZN(n7506)
         );
  NAND3_X1 U9218 ( .A1(n6232), .A2(n7504), .A3(n7503), .ZN(n7505) );
  AOI21_X1 U9219 ( .B1(n7506), .B2(n7505), .A(n7539), .ZN(n7508) );
  NOR3_X1 U9220 ( .A1(n7509), .A2(n7508), .A3(n7507), .ZN(n7511) );
  OAI21_X1 U9221 ( .B1(n7512), .B2(n7511), .A(n7510), .ZN(n7513) );
  AOI21_X1 U9222 ( .B1(n7514), .B2(n7513), .A(n7607), .ZN(n7517) );
  OAI21_X1 U9223 ( .B1(n7517), .B2(n7516), .A(n7515), .ZN(n7519) );
  NAND2_X1 U9224 ( .A1(n7899), .A2(n9040), .ZN(n7518) );
  AND2_X1 U9225 ( .A1(n9075), .A2(n7518), .ZN(n7624) );
  AOI211_X1 U9226 ( .C1(n7520), .C2(n7519), .A(n7622), .B(n7624), .ZN(n7525)
         );
  OAI21_X1 U9227 ( .B1(n7523), .B2(n7522), .A(n7521), .ZN(n7626) );
  INV_X1 U9228 ( .A(n7626), .ZN(n7524) );
  OAI211_X1 U9229 ( .C1(n7525), .C2(n7524), .A(n5807), .B(n7632), .ZN(n7526)
         );
  NAND2_X1 U9230 ( .A1(n7526), .A2(n7528), .ZN(n7527) );
  MUX2_X1 U9231 ( .A(n7528), .B(n7527), .S(n9243), .Z(n7637) );
  INV_X1 U9232 ( .A(n7624), .ZN(n7529) );
  NOR2_X1 U9233 ( .A1(n7529), .A2(n7627), .ZN(n7629) );
  INV_X1 U9234 ( .A(n7533), .ZN(n7534) );
  OAI211_X1 U9235 ( .C1(n7546), .C2(n7541), .A(n7540), .B(n9456), .ZN(n7543)
         );
  OAI21_X1 U9236 ( .B1(n7546), .B2(n7545), .A(n7544), .ZN(n7548) );
  INV_X1 U9237 ( .A(n7557), .ZN(n7549) );
  NOR2_X1 U9238 ( .A1(n7549), .A2(n4788), .ZN(n7550) );
  MUX2_X1 U9239 ( .A(n7551), .B(n7550), .S(n7627), .Z(n7553) );
  NOR2_X1 U9240 ( .A1(n7561), .A2(n7555), .ZN(n7560) );
  AOI21_X1 U9241 ( .B1(n7558), .B2(n7557), .A(n7556), .ZN(n7559) );
  MUX2_X1 U9242 ( .A(n7560), .B(n7559), .S(n7627), .Z(n7569) );
  NOR2_X1 U9243 ( .A1(n7562), .A2(n7561), .ZN(n7567) );
  INV_X1 U9244 ( .A(n7563), .ZN(n7564) );
  AOI21_X1 U9245 ( .B1(n8195), .B2(n7565), .A(n7564), .ZN(n7566) );
  MUX2_X1 U9246 ( .A(n7567), .B(n7566), .S(n7627), .Z(n7568) );
  INV_X1 U9247 ( .A(n9266), .ZN(n7571) );
  INV_X1 U9248 ( .A(n8197), .ZN(n7570) );
  MUX2_X1 U9249 ( .A(n7571), .B(n7570), .S(n7627), .Z(n7572) );
  INV_X1 U9250 ( .A(n7574), .ZN(n7575) );
  MUX2_X1 U9251 ( .A(n8198), .B(n7575), .S(n7627), .Z(n7576) );
  NOR3_X1 U9252 ( .A1(n7577), .A2(n7576), .A3(n9251), .ZN(n7581) );
  NAND2_X1 U9253 ( .A1(n8202), .A2(n8201), .ZN(n7578) );
  MUX2_X1 U9254 ( .A(n7579), .B(n7578), .S(n7627), .Z(n7580) );
  INV_X1 U9255 ( .A(n7582), .ZN(n7584) );
  INV_X1 U9256 ( .A(n7586), .ZN(n7588) );
  NAND2_X1 U9257 ( .A1(n7588), .A2(n7587), .ZN(n7592) );
  OAI22_X1 U9258 ( .A1(n7590), .A2(n8203), .B1(n7627), .B2(n7589), .ZN(n7591)
         );
  OAI21_X1 U9259 ( .B1(n7593), .B2(n7592), .A(n7591), .ZN(n7597) );
  AOI21_X1 U9260 ( .B1(n7597), .B2(n7595), .A(n7594), .ZN(n7601) );
  NAND3_X1 U9261 ( .A1(n7597), .A2(n7596), .A3(n8204), .ZN(n7598) );
  AOI21_X1 U9262 ( .B1(n7598), .B2(n8206), .A(n8208), .ZN(n7599) );
  NOR2_X1 U9263 ( .A1(n7599), .A2(n8209), .ZN(n7600) );
  MUX2_X1 U9264 ( .A(n7601), .B(n7600), .S(n7627), .Z(n7603) );
  INV_X1 U9265 ( .A(n8211), .ZN(n7602) );
  NOR3_X1 U9266 ( .A1(n7603), .A2(n7602), .A3(n7604), .ZN(n7611) );
  INV_X1 U9267 ( .A(n7604), .ZN(n7606) );
  OAI21_X1 U9268 ( .B1(n7606), .B2(n7605), .A(n9113), .ZN(n7608) );
  MUX2_X1 U9269 ( .A(n7608), .B(n7607), .S(n7627), .Z(n7610) );
  MUX2_X1 U9270 ( .A(n8212), .B(n9113), .S(n7627), .Z(n7609) );
  OAI211_X1 U9271 ( .C1(n7611), .C2(n7610), .A(n9115), .B(n7609), .ZN(n7614)
         );
  MUX2_X1 U9272 ( .A(n7612), .B(n8214), .S(n7627), .Z(n7613) );
  NAND3_X1 U9273 ( .A1(n7614), .A2(n8188), .A3(n7613), .ZN(n7618) );
  MUX2_X1 U9274 ( .A(n7616), .B(n7615), .S(n7627), .Z(n7617) );
  NAND3_X1 U9275 ( .A1(n7618), .A2(n9088), .A3(n7617), .ZN(n7621) );
  NAND2_X1 U9276 ( .A1(n7619), .A2(n4706), .ZN(n7620) );
  NAND2_X1 U9277 ( .A1(n7623), .A2(n7627), .ZN(n7625) );
  NOR2_X1 U9278 ( .A1(n7646), .A2(n7630), .ZN(n7634) );
  OAI21_X1 U9279 ( .B1(n9243), .B2(n7631), .A(n7635), .ZN(n7633) );
  OAI211_X1 U9280 ( .C1(n7635), .C2(n7634), .A(n7633), .B(n7632), .ZN(n7636)
         );
  AND2_X1 U9281 ( .A1(n7637), .A2(n7636), .ZN(n7639) );
  NAND4_X1 U9282 ( .A1(n7644), .A2(n7643), .A3(n7642), .A4(n7641), .ZN(n7645)
         );
  OAI211_X1 U9283 ( .C1(n7646), .C2(n7648), .A(n7645), .B(P1_B_REG_SCAN_IN), 
        .ZN(n7647) );
  OAI21_X1 U9284 ( .B1(n7649), .B2(n7648), .A(n7647), .ZN(P1_U3240) );
  NAND2_X1 U9285 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9059), .ZN(n7651) );
  OAI21_X1 U9286 ( .B1(n9059), .B2(P1_REG2_REG_17__SCAN_IN), .A(n7651), .ZN(
        n9057) );
  AOI21_X1 U9287 ( .B1(n9059), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9056), .ZN(
        n9632) );
  XNOR2_X1 U9288 ( .A(n9636), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n9631) );
  NOR2_X1 U9289 ( .A1(n9632), .A2(n9631), .ZN(n9630) );
  AOI21_X1 U9290 ( .B1(n9636), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9630), .ZN(
        n7652) );
  XNOR2_X1 U9291 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n7652), .ZN(n7660) );
  INV_X1 U9292 ( .A(n7660), .ZN(n7656) );
  AOI22_X1 U9293 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n9636), .B1(n7653), .B2(
        n10158), .ZN(n9639) );
  AOI21_X1 U9294 ( .B1(n7655), .B2(P1_REG1_REG_16__SCAN_IN), .A(n7654), .ZN(
        n9063) );
  XNOR2_X1 U9295 ( .A(n9059), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9062) );
  NOR2_X1 U9296 ( .A1(n9063), .A2(n9062), .ZN(n9061) );
  AOI21_X1 U9297 ( .B1(n9059), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9061), .ZN(
        n9638) );
  NAND2_X1 U9298 ( .A1(n9639), .A2(n9638), .ZN(n9637) );
  OAI22_X1 U9299 ( .A1(n7656), .A2(n9629), .B1(n7657), .B2(n9060), .ZN(n7663)
         );
  AOI21_X1 U9300 ( .B1(n7657), .B2(n9641), .A(n9635), .ZN(n7658) );
  OAI21_X1 U9301 ( .B1(n7660), .B2(n7659), .A(n7658), .ZN(n7662) );
  NAND2_X1 U9302 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8939) );
  NAND2_X1 U9303 ( .A1(n7664), .A2(n7847), .ZN(n8490) );
  NAND2_X1 U9304 ( .A1(n8225), .A2(n7673), .ZN(n7667) );
  NAND2_X1 U9305 ( .A1(n7665), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7666) );
  INV_X1 U9306 ( .A(n7849), .ZN(n7669) );
  NAND2_X1 U9307 ( .A1(n7873), .A2(n7668), .ZN(n7850) );
  NAND2_X1 U9308 ( .A1(n8228), .A2(n7673), .ZN(n7671) );
  INV_X1 U9309 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8233) );
  OR2_X1 U9310 ( .A1(n7674), .A2(n8233), .ZN(n7670) );
  OAI211_X1 U9311 ( .C1(n7672), .C2(n8481), .A(n7728), .B(n7876), .ZN(n7679)
         );
  NAND2_X1 U9312 ( .A1(n8879), .A2(n7673), .ZN(n7676) );
  OR2_X1 U9313 ( .A1(n7674), .A2(n5948), .ZN(n7675) );
  OR2_X1 U9314 ( .A1(n8761), .A2(n7876), .ZN(n7854) );
  NAND2_X1 U9315 ( .A1(n8481), .A2(n8492), .ZN(n7852) );
  NAND2_X1 U9316 ( .A1(n7854), .A2(n7852), .ZN(n7857) );
  NAND3_X1 U9317 ( .A1(n7679), .A2(n7678), .A3(n7677), .ZN(n7680) );
  NAND2_X1 U9318 ( .A1(n8761), .A2(n7876), .ZN(n7856) );
  NAND2_X1 U9319 ( .A1(n7680), .A2(n7856), .ZN(n7681) );
  XNOR2_X1 U9320 ( .A(n7681), .B(n7711), .ZN(n7684) );
  NAND2_X1 U9321 ( .A1(n7856), .A2(n4436), .ZN(n7855) );
  INV_X1 U9322 ( .A(n7855), .ZN(n7707) );
  NAND4_X1 U9323 ( .A1(n6495), .A2(n7687), .A3(n7686), .A4(n7709), .ZN(n7691)
         );
  NOR4_X1 U9324 ( .A1(n7691), .A2(n7690), .A3(n7689), .A4(n7688), .ZN(n7693)
         );
  NAND4_X1 U9325 ( .A1(n7693), .A2(n7692), .A3(n7757), .A4(n8735), .ZN(n7696)
         );
  NOR4_X1 U9326 ( .A1(n7696), .A2(n7051), .A3(n7695), .A4(n7694), .ZN(n7699)
         );
  INV_X1 U9327 ( .A(n7697), .ZN(n7789) );
  NAND3_X1 U9328 ( .A1(n7699), .A2(n7789), .A3(n7698), .ZN(n7700) );
  NOR4_X1 U9329 ( .A1(n8682), .A2(n7700), .A3(n8702), .A4(n8711), .ZN(n7701)
         );
  NAND4_X1 U9330 ( .A1(n8638), .A2(n4468), .A3(n4645), .A4(n7701), .ZN(n7702)
         );
  NOR4_X1 U9331 ( .A1(n8577), .A2(n8590), .A3(n8610), .A4(n7702), .ZN(n7703)
         );
  NAND4_X1 U9332 ( .A1(n8520), .A2(n7703), .A3(n8602), .A4(n8556), .ZN(n7704)
         );
  NOR4_X1 U9333 ( .A1(n8486), .A2(n8507), .A3(n7705), .A4(n7704), .ZN(n7706)
         );
  NAND4_X1 U9334 ( .A1(n7677), .A2(n7707), .A3(n8488), .A4(n7706), .ZN(n7708)
         );
  XNOR2_X1 U9335 ( .A(n7708), .B(n8546), .ZN(n7710) );
  OAI22_X1 U9336 ( .A1(n7710), .A2(n7728), .B1(n7709), .B2(n7863), .ZN(n7862)
         );
  NAND2_X1 U9337 ( .A1(n7728), .A2(n7711), .ZN(n7712) );
  OR2_X1 U9338 ( .A1(n5140), .A2(n7712), .ZN(n7842) );
  INV_X1 U9339 ( .A(n7713), .ZN(n7714) );
  AOI22_X1 U9340 ( .A1(n8556), .A2(n7714), .B1(n8274), .B2(n8796), .ZN(n7828)
         );
  INV_X1 U9341 ( .A(n7842), .ZN(n7859) );
  INV_X1 U9342 ( .A(n7715), .ZN(n7719) );
  OAI211_X1 U9343 ( .C1(n8661), .C2(n7717), .A(n7809), .B(n7716), .ZN(n7718)
         );
  MUX2_X1 U9344 ( .A(n7719), .B(n7718), .S(n7859), .Z(n7808) );
  AND2_X1 U9345 ( .A1(n7749), .A2(n7746), .ZN(n7720) );
  MUX2_X1 U9346 ( .A(n7720), .B(n7724), .S(n7842), .Z(n7748) );
  INV_X1 U9347 ( .A(n7748), .ZN(n7722) );
  NAND2_X1 U9348 ( .A1(n7722), .A2(n7721), .ZN(n7727) );
  NAND2_X1 U9349 ( .A1(n7724), .A2(n7723), .ZN(n7726) );
  INV_X1 U9350 ( .A(n7753), .ZN(n7725) );
  AOI21_X1 U9351 ( .B1(n7727), .B2(n7726), .A(n7725), .ZN(n7756) );
  AND2_X1 U9352 ( .A1(n7729), .A2(n7728), .ZN(n7732) );
  AND2_X1 U9353 ( .A1(n7731), .A2(n7730), .ZN(n7740) );
  OAI21_X1 U9354 ( .B1(n7733), .B2(n7732), .A(n7740), .ZN(n7736) );
  AND2_X1 U9355 ( .A1(n7742), .A2(n7842), .ZN(n7735) );
  AOI21_X1 U9356 ( .B1(n7736), .B2(n7735), .A(n7734), .ZN(n7737) );
  NAND2_X1 U9357 ( .A1(n7737), .A2(n7748), .ZN(n7751) );
  NAND2_X1 U9358 ( .A1(n7739), .A2(n7738), .ZN(n7741) );
  NAND2_X1 U9359 ( .A1(n7741), .A2(n7740), .ZN(n7743) );
  NAND2_X1 U9360 ( .A1(n7743), .A2(n7742), .ZN(n7744) );
  OAI21_X1 U9361 ( .B1(n7751), .B2(n7744), .A(n7859), .ZN(n7754) );
  NAND2_X1 U9362 ( .A1(n7746), .A2(n7745), .ZN(n7747) );
  NAND2_X1 U9363 ( .A1(n7748), .A2(n7747), .ZN(n7750) );
  NAND4_X1 U9364 ( .A1(n7751), .A2(n7750), .A3(n7759), .A4(n7749), .ZN(n7752)
         );
  NAND3_X1 U9365 ( .A1(n7754), .A2(n7753), .A3(n7752), .ZN(n7755) );
  OAI21_X1 U9366 ( .B1(n7756), .B2(n7842), .A(n7755), .ZN(n7758) );
  OAI211_X1 U9367 ( .C1(n7759), .C2(n7842), .A(n7758), .B(n7757), .ZN(n7763)
         );
  MUX2_X1 U9368 ( .A(n7761), .B(n7760), .S(n7842), .Z(n7762) );
  NAND3_X1 U9369 ( .A1(n7763), .A2(n9730), .A3(n7762), .ZN(n7767) );
  NAND2_X1 U9370 ( .A1(n8387), .A2(n9788), .ZN(n7764) );
  MUX2_X1 U9371 ( .A(n7765), .B(n7764), .S(n7842), .Z(n7766) );
  NAND3_X1 U9372 ( .A1(n7767), .A2(n7768), .A3(n7766), .ZN(n7781) );
  NAND2_X1 U9373 ( .A1(n7773), .A2(n7768), .ZN(n7770) );
  NAND2_X1 U9374 ( .A1(n7774), .A2(n7771), .ZN(n7769) );
  AOI21_X1 U9375 ( .B1(n7770), .B2(n7842), .A(n7769), .ZN(n7780) );
  NAND2_X1 U9376 ( .A1(n7782), .A2(n7773), .ZN(n7778) );
  INV_X1 U9377 ( .A(n7771), .ZN(n7772) );
  NAND2_X1 U9378 ( .A1(n7773), .A2(n7772), .ZN(n7775) );
  NAND3_X1 U9379 ( .A1(n7776), .A2(n7775), .A3(n7774), .ZN(n7777) );
  MUX2_X1 U9380 ( .A(n7778), .B(n7777), .S(n7842), .Z(n7779) );
  AOI21_X1 U9381 ( .B1(n7781), .B2(n7780), .A(n7779), .ZN(n7791) );
  NAND2_X1 U9382 ( .A1(n7787), .A2(n7782), .ZN(n7785) );
  INV_X1 U9383 ( .A(n7783), .ZN(n7784) );
  MUX2_X1 U9384 ( .A(n7785), .B(n7784), .S(n7859), .Z(n7790) );
  MUX2_X1 U9385 ( .A(n7787), .B(n7786), .S(n7842), .Z(n7788) );
  OAI211_X1 U9386 ( .C1(n7791), .C2(n7790), .A(n7789), .B(n7788), .ZN(n7795)
         );
  INV_X1 U9387 ( .A(n8711), .ZN(n8720) );
  MUX2_X1 U9388 ( .A(n7793), .B(n7792), .S(n7842), .Z(n7794) );
  NAND3_X1 U9389 ( .A1(n7795), .A2(n8720), .A3(n7794), .ZN(n7799) );
  INV_X1 U9390 ( .A(n8702), .ZN(n8694) );
  MUX2_X1 U9391 ( .A(n7797), .B(n7796), .S(n7842), .Z(n7798) );
  NAND3_X1 U9392 ( .A1(n7799), .A2(n8694), .A3(n7798), .ZN(n7803) );
  INV_X1 U9393 ( .A(n8682), .ZN(n8678) );
  MUX2_X1 U9394 ( .A(n7801), .B(n7800), .S(n7842), .Z(n7802) );
  NAND3_X1 U9395 ( .A1(n7803), .A2(n8678), .A3(n7802), .ZN(n7806) );
  OR2_X1 U9396 ( .A1(n7804), .A2(n7859), .ZN(n7805) );
  INV_X1 U9397 ( .A(n7807), .ZN(n8636) );
  AOI21_X1 U9398 ( .B1(n7819), .B2(n7809), .A(n7815), .ZN(n7811) );
  NAND2_X1 U9399 ( .A1(n7821), .A2(n8619), .ZN(n7810) );
  NAND2_X1 U9400 ( .A1(n8600), .A2(n8380), .ZN(n7822) );
  OAI211_X1 U9401 ( .C1(n7811), .C2(n7810), .A(n7816), .B(n7822), .ZN(n7812)
         );
  NAND3_X1 U9402 ( .A1(n7812), .A2(n7814), .A3(n7820), .ZN(n7813) );
  MUX2_X1 U9403 ( .A(n7814), .B(n7813), .S(n7842), .Z(n7827) );
  AOI21_X1 U9404 ( .B1(n8636), .B2(n8619), .A(n7815), .ZN(n7817) );
  NAND3_X1 U9405 ( .A1(n7823), .A2(n7824), .A3(n7822), .ZN(n7825) );
  MUX2_X1 U9406 ( .A(n7825), .B(n7824), .S(n7842), .Z(n7826) );
  INV_X1 U9407 ( .A(n8537), .ZN(n7832) );
  INV_X1 U9408 ( .A(n7829), .ZN(n7830) );
  NAND2_X1 U9409 ( .A1(n8556), .A2(n7830), .ZN(n7831) );
  NAND3_X1 U9410 ( .A1(n8528), .A2(n7832), .A3(n7831), .ZN(n7833) );
  INV_X1 U9411 ( .A(n7835), .ZN(n7834) );
  AOI21_X1 U9412 ( .B1(n7837), .B2(n7835), .A(n7859), .ZN(n7836) );
  AOI21_X1 U9413 ( .B1(n7838), .B2(n7837), .A(n7836), .ZN(n7841) );
  OAI21_X1 U9414 ( .B1(n7859), .B2(n7839), .A(n8512), .ZN(n7840) );
  AOI21_X1 U9415 ( .B1(n7846), .B2(n7844), .A(n7859), .ZN(n7845) );
  OAI21_X1 U9416 ( .B1(n7859), .B2(n7847), .A(n8488), .ZN(n7848) );
  MUX2_X1 U9417 ( .A(n7850), .B(n7849), .S(n7859), .Z(n7851) );
  NAND2_X1 U9418 ( .A1(n7862), .A2(n7861), .ZN(n7866) );
  NAND3_X1 U9419 ( .A1(n7864), .A2(n7863), .A3(n9763), .ZN(n7865) );
  NAND4_X1 U9420 ( .A1(n7869), .A2(n7874), .A3(n8729), .A4(n7868), .ZN(n7870)
         );
  OAI211_X1 U9421 ( .C1(n5140), .C2(n7871), .A(n7870), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7872) );
  XOR2_X1 U9422 ( .A(n8761), .B(n8480), .Z(n8763) );
  NAND2_X1 U9423 ( .A1(n7874), .A2(P2_B_REG_SCAN_IN), .ZN(n7875) );
  NAND2_X1 U9424 ( .A1(n8731), .A2(n7875), .ZN(n8493) );
  NOR2_X1 U9425 ( .A1(n7876), .A2(n8493), .ZN(n8760) );
  INV_X1 U9426 ( .A(n8760), .ZN(n8766) );
  NOR2_X1 U9427 ( .A1(n8656), .A2(n8766), .ZN(n8482) );
  AOI21_X1 U9428 ( .B1(n9745), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8482), .ZN(
        n7878) );
  NAND2_X1 U9429 ( .A1(n8761), .A2(n8749), .ZN(n7877) );
  OAI211_X1 U9430 ( .C1(n8763), .C2(n8499), .A(n7878), .B(n7877), .ZN(P2_U3265) );
  AOI22_X1 U9431 ( .A1(n8358), .A2(n7879), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n7893), .ZN(n7884) );
  XOR2_X1 U9432 ( .A(n7881), .B(n7880), .Z(n7882) );
  NAND2_X1 U9433 ( .A1(n7882), .A2(n8353), .ZN(n7883) );
  OAI211_X1 U9434 ( .C1(n7885), .C2(n8348), .A(n7884), .B(n7883), .ZN(P2_U3239) );
  OAI222_X1 U9435 ( .A1(n8237), .A2(n7887), .B1(n8236), .B2(n7886), .C1(
        P2_U3152), .C2(n5702), .ZN(P2_U3336) );
  OAI21_X1 U9436 ( .B1(n7890), .B2(n7889), .A(n7888), .ZN(n7892) );
  AOI22_X1 U9437 ( .A1(n8353), .A2(n7892), .B1(n8358), .B2(n7891), .ZN(n7895)
         );
  AOI22_X1 U9438 ( .A1(n8374), .A2(n6270), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n7893), .ZN(n7894) );
  NAND2_X1 U9439 ( .A1(n7895), .A2(n7894), .ZN(P2_U3224) );
  INV_X1 U9440 ( .A(n9322), .ZN(n9085) );
  INV_X1 U9441 ( .A(n9362), .ZN(n8949) );
  INV_X1 U9442 ( .A(n9372), .ZN(n9223) );
  INV_X1 U9443 ( .A(n9388), .ZN(n9279) );
  INV_X1 U9444 ( .A(n9391), .ZN(n9288) );
  NOR2_X2 U9445 ( .A1(n9337), .A2(n9135), .ZN(n9124) );
  NAND2_X1 U9446 ( .A1(n9112), .A2(n9124), .ZN(n9107) );
  NAND2_X1 U9447 ( .A1(n9085), .A2(n9100), .ZN(n9080) );
  NAND2_X1 U9448 ( .A1(n9316), .A2(n9073), .ZN(n9313) );
  NAND2_X1 U9449 ( .A1(n9310), .A2(n9650), .ZN(n7901) );
  INV_X1 U9450 ( .A(P1_B_REG_SCAN_IN), .ZN(n7897) );
  NOR2_X1 U9451 ( .A1(n9532), .A2(n7897), .ZN(n7898) );
  NOR2_X1 U9452 ( .A1(n9462), .A2(n7898), .ZN(n8193) );
  NAND2_X1 U9453 ( .A1(n7899), .A2(n8193), .ZN(n9314) );
  NOR2_X1 U9454 ( .A1(n4419), .A2(n9314), .ZN(n9076) );
  AOI21_X1 U9455 ( .B1(n4419), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9076), .ZN(
        n7900) );
  OAI211_X1 U9456 ( .C1(n9311), .C2(n9656), .A(n7901), .B(n7900), .ZN(P1_U3261) );
  AND2_X1 U9457 ( .A1(n9176), .A2(n8007), .ZN(n7902) );
  AOI21_X1 U9458 ( .B1(n9349), .B2(n8004), .A(n7902), .ZN(n8919) );
  NAND2_X1 U9459 ( .A1(n8914), .A2(n7995), .ZN(n7906) );
  NAND2_X1 U9460 ( .A1(n9292), .A2(n8004), .ZN(n7905) );
  NAND2_X1 U9461 ( .A1(n7906), .A2(n7905), .ZN(n7907) );
  XNOR2_X1 U9462 ( .A(n7907), .B(n7998), .ZN(n7914) );
  NAND2_X1 U9463 ( .A1(n7913), .A2(n7914), .ZN(n8906) );
  NAND2_X1 U9464 ( .A1(n8914), .A2(n6394), .ZN(n7909) );
  NAND2_X1 U9465 ( .A1(n9292), .A2(n8007), .ZN(n7908) );
  NAND2_X1 U9466 ( .A1(n7909), .A2(n7908), .ZN(n8909) );
  NAND2_X1 U9467 ( .A1(n8906), .A2(n8909), .ZN(n7919) );
  NAND2_X1 U9468 ( .A1(n9391), .A2(n7995), .ZN(n7911) );
  NAND2_X1 U9469 ( .A1(n9042), .A2(n8004), .ZN(n7910) );
  NAND2_X1 U9470 ( .A1(n7911), .A2(n7910), .ZN(n7912) );
  XNOR2_X1 U9471 ( .A(n7912), .B(n7998), .ZN(n7920) );
  INV_X1 U9472 ( .A(n7914), .ZN(n7915) );
  NAND2_X1 U9473 ( .A1(n7916), .A2(n7915), .ZN(n8907) );
  NAND2_X1 U9474 ( .A1(n9391), .A2(n6394), .ZN(n7918) );
  NAND2_X1 U9475 ( .A1(n9042), .A2(n8007), .ZN(n7917) );
  NAND2_X1 U9476 ( .A1(n7918), .A2(n7917), .ZN(n9028) );
  INV_X1 U9477 ( .A(n7920), .ZN(n7921) );
  NAND2_X1 U9478 ( .A1(n9388), .A2(n7995), .ZN(n7923) );
  NAND2_X1 U9479 ( .A1(n9294), .A2(n8004), .ZN(n7922) );
  NAND2_X1 U9480 ( .A1(n7923), .A2(n7922), .ZN(n7924) );
  XNOR2_X1 U9481 ( .A(n7924), .B(n8005), .ZN(n7926) );
  AND2_X1 U9482 ( .A1(n9294), .A2(n8007), .ZN(n7925) );
  AOI21_X1 U9483 ( .B1(n9388), .B2(n8004), .A(n7925), .ZN(n7927) );
  XNOR2_X1 U9484 ( .A(n7926), .B(n7927), .ZN(n8963) );
  INV_X1 U9485 ( .A(n7926), .ZN(n7928) );
  NAND2_X1 U9486 ( .A1(n7928), .A2(n7927), .ZN(n7929) );
  NAND2_X1 U9487 ( .A1(n9383), .A2(n7995), .ZN(n7931) );
  NAND2_X1 U9488 ( .A1(n9239), .A2(n8004), .ZN(n7930) );
  NAND2_X1 U9489 ( .A1(n7931), .A2(n7930), .ZN(n7932) );
  XNOR2_X1 U9490 ( .A(n7932), .B(n8005), .ZN(n7934) );
  AND2_X1 U9491 ( .A1(n9239), .A2(n8007), .ZN(n7933) );
  AOI21_X1 U9492 ( .B1(n9383), .B2(n8004), .A(n7933), .ZN(n7935) );
  XNOR2_X1 U9493 ( .A(n7934), .B(n7935), .ZN(n8971) );
  INV_X1 U9494 ( .A(n7934), .ZN(n7936) );
  NAND2_X1 U9495 ( .A1(n9377), .A2(n7995), .ZN(n7938) );
  NAND2_X1 U9496 ( .A1(n9227), .A2(n8004), .ZN(n7937) );
  NAND2_X1 U9497 ( .A1(n7938), .A2(n7937), .ZN(n7939) );
  XNOR2_X1 U9498 ( .A(n7939), .B(n7998), .ZN(n9006) );
  AND2_X1 U9499 ( .A1(n9227), .A2(n8007), .ZN(n7940) );
  AOI21_X1 U9500 ( .B1(n9377), .B2(n8004), .A(n7940), .ZN(n9005) );
  NAND2_X1 U9501 ( .A1(n9372), .A2(n7995), .ZN(n7942) );
  NAND2_X1 U9502 ( .A1(n9240), .A2(n8004), .ZN(n7941) );
  NAND2_X1 U9503 ( .A1(n7942), .A2(n7941), .ZN(n7943) );
  XNOR2_X1 U9504 ( .A(n7943), .B(n7998), .ZN(n8937) );
  AND2_X1 U9505 ( .A1(n9240), .A2(n8007), .ZN(n7944) );
  AOI21_X1 U9506 ( .B1(n9372), .B2(n8004), .A(n7944), .ZN(n8936) );
  AND2_X1 U9507 ( .A1(n8937), .A2(n8936), .ZN(n7945) );
  INV_X1 U9508 ( .A(n8937), .ZN(n7947) );
  INV_X1 U9509 ( .A(n8936), .ZN(n7946) );
  NAND2_X1 U9510 ( .A1(n9368), .A2(n7995), .ZN(n7949) );
  NAND2_X1 U9511 ( .A1(n9228), .A2(n8004), .ZN(n7948) );
  NAND2_X1 U9512 ( .A1(n7949), .A2(n7948), .ZN(n7950) );
  XNOR2_X1 U9513 ( .A(n7950), .B(n8005), .ZN(n7953) );
  NAND2_X1 U9514 ( .A1(n9368), .A2(n8004), .ZN(n7952) );
  NAND2_X1 U9515 ( .A1(n9228), .A2(n8007), .ZN(n7951) );
  NAND2_X1 U9516 ( .A1(n7952), .A2(n7951), .ZN(n7954) );
  INV_X1 U9517 ( .A(n7953), .ZN(n7956) );
  INV_X1 U9518 ( .A(n7954), .ZN(n7955) );
  NAND2_X1 U9519 ( .A1(n7956), .A2(n7955), .ZN(n8987) );
  NAND2_X1 U9520 ( .A1(n9362), .A2(n7995), .ZN(n7958) );
  NAND2_X1 U9521 ( .A1(n9177), .A2(n8004), .ZN(n7957) );
  NAND2_X1 U9522 ( .A1(n7958), .A2(n7957), .ZN(n7959) );
  XNOR2_X1 U9523 ( .A(n7959), .B(n8005), .ZN(n7961) );
  AND2_X1 U9524 ( .A1(n9177), .A2(n8007), .ZN(n7960) );
  AOI21_X1 U9525 ( .B1(n9362), .B2(n6394), .A(n7960), .ZN(n7962) );
  XNOR2_X1 U9526 ( .A(n7961), .B(n7962), .ZN(n8946) );
  NAND2_X1 U9527 ( .A1(n8945), .A2(n8946), .ZN(n8944) );
  INV_X1 U9528 ( .A(n7961), .ZN(n7963) );
  NAND2_X1 U9529 ( .A1(n7963), .A2(n7962), .ZN(n7964) );
  AND2_X1 U9530 ( .A1(n9162), .A2(n8007), .ZN(n7965) );
  AOI21_X1 U9531 ( .B1(n9354), .B2(n6394), .A(n7965), .ZN(n7969) );
  NAND2_X1 U9532 ( .A1(n7970), .A2(n7969), .ZN(n8994) );
  NAND2_X1 U9533 ( .A1(n9354), .A2(n7995), .ZN(n7967) );
  NAND2_X1 U9534 ( .A1(n9162), .A2(n8004), .ZN(n7966) );
  NAND2_X1 U9535 ( .A1(n7967), .A2(n7966), .ZN(n7968) );
  XNOR2_X1 U9536 ( .A(n7968), .B(n8005), .ZN(n8997) );
  NAND2_X1 U9537 ( .A1(n9349), .A2(n7995), .ZN(n7972) );
  NAND2_X1 U9538 ( .A1(n9176), .A2(n6394), .ZN(n7971) );
  NAND2_X1 U9539 ( .A1(n7972), .A2(n7971), .ZN(n7973) );
  XNOR2_X1 U9540 ( .A(n7973), .B(n8005), .ZN(n7974) );
  AOI22_X1 U9541 ( .A1(n9345), .A2(n6394), .B1(n8007), .B2(n9161), .ZN(n7978)
         );
  NAND2_X1 U9542 ( .A1(n9345), .A2(n7995), .ZN(n7976) );
  NAND2_X1 U9543 ( .A1(n9161), .A2(n6394), .ZN(n7975) );
  NAND2_X1 U9544 ( .A1(n7976), .A2(n7975), .ZN(n7977) );
  XNOR2_X1 U9545 ( .A(n7977), .B(n8005), .ZN(n7980) );
  XOR2_X1 U9546 ( .A(n7978), .B(n7980), .Z(n8977) );
  INV_X1 U9547 ( .A(n7978), .ZN(n7979) );
  NAND2_X1 U9548 ( .A1(n9337), .A2(n7995), .ZN(n7983) );
  NAND2_X1 U9549 ( .A1(n9118), .A2(n6394), .ZN(n7982) );
  NAND2_X1 U9550 ( .A1(n7983), .A2(n7982), .ZN(n7984) );
  XNOR2_X1 U9551 ( .A(n7984), .B(n8005), .ZN(n7985) );
  AOI22_X1 U9552 ( .A1(n9337), .A2(n6394), .B1(n8007), .B2(n9118), .ZN(n7986)
         );
  XNOR2_X1 U9553 ( .A(n7985), .B(n7986), .ZN(n8954) );
  INV_X1 U9554 ( .A(n7985), .ZN(n7987) );
  NAND2_X1 U9555 ( .A1(n9332), .A2(n7995), .ZN(n7989) );
  NAND2_X1 U9556 ( .A1(n9130), .A2(n8004), .ZN(n7988) );
  NAND2_X1 U9557 ( .A1(n7989), .A2(n7988), .ZN(n7990) );
  XNOR2_X1 U9558 ( .A(n7990), .B(n8005), .ZN(n7992) );
  AND2_X1 U9559 ( .A1(n9130), .A2(n8007), .ZN(n7991) );
  AOI21_X1 U9560 ( .B1(n9332), .B2(n8004), .A(n7991), .ZN(n7993) );
  XNOR2_X1 U9561 ( .A(n7992), .B(n7993), .ZN(n9017) );
  NAND2_X1 U9562 ( .A1(n9328), .A2(n7995), .ZN(n7997) );
  NAND2_X1 U9563 ( .A1(n9117), .A2(n6394), .ZN(n7996) );
  NAND2_X1 U9564 ( .A1(n7997), .A2(n7996), .ZN(n7999) );
  XNOR2_X1 U9565 ( .A(n7999), .B(n7998), .ZN(n8898) );
  AND2_X1 U9566 ( .A1(n9117), .A2(n8007), .ZN(n8000) );
  AOI21_X1 U9567 ( .B1(n9328), .B2(n8004), .A(n8000), .ZN(n8001) );
  NAND2_X1 U9568 ( .A1(n8898), .A2(n8001), .ZN(n8003) );
  INV_X1 U9569 ( .A(n8898), .ZN(n8002) );
  INV_X1 U9570 ( .A(n8001), .ZN(n8897) );
  AOI22_X1 U9571 ( .A1(n9322), .A2(n6077), .B1(n8004), .B2(n9041), .ZN(n8006)
         );
  XNOR2_X1 U9572 ( .A(n8006), .B(n8005), .ZN(n8009) );
  AOI22_X1 U9573 ( .A1(n9322), .A2(n6394), .B1(n8007), .B2(n9041), .ZN(n8008)
         );
  XNOR2_X1 U9574 ( .A(n8009), .B(n8008), .ZN(n8010) );
  INV_X1 U9575 ( .A(n8011), .ZN(n9083) );
  AOI22_X1 U9576 ( .A1(n9083), .A2(n9029), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8013) );
  NAND2_X1 U9577 ( .A1(n9117), .A2(n8978), .ZN(n8012) );
  OAI211_X1 U9578 ( .C1(n8014), .C2(n9009), .A(n8013), .B(n8012), .ZN(n8015)
         );
  AOI21_X1 U9579 ( .B1(n9322), .B2(n9036), .A(n8015), .ZN(n8016) );
  INV_X1 U9580 ( .A(n8099), .ZN(n8021) );
  NAND2_X1 U9581 ( .A1(n8041), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8018) );
  OAI21_X1 U9582 ( .B1(n8041), .B2(P2_REG1_REG_6__SCAN_IN), .A(n8018), .ZN(
        n8102) );
  NOR2_X1 U9583 ( .A1(n8103), .A2(n8102), .ZN(n8101) );
  AOI21_X1 U9584 ( .B1(n8041), .B2(P2_REG1_REG_6__SCAN_IN), .A(n8101), .ZN(
        n9872) );
  NAND2_X1 U9585 ( .A1(n8039), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8019) );
  OAI21_X1 U9586 ( .B1(n8039), .B2(P2_REG1_REG_7__SCAN_IN), .A(n8019), .ZN(
        n9871) );
  NOR2_X1 U9587 ( .A1(n9872), .A2(n9871), .ZN(n9870) );
  INV_X1 U9588 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8020) );
  MUX2_X1 U9589 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n8020), .S(n8099), .Z(n8090)
         );
  NOR2_X1 U9590 ( .A1(n8091), .A2(n8090), .ZN(n8089) );
  AOI21_X1 U9591 ( .B1(n8021), .B2(P2_REG1_REG_8__SCAN_IN), .A(n8089), .ZN(
        n8079) );
  NAND2_X1 U9592 ( .A1(n8036), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8022) );
  OAI21_X1 U9593 ( .B1(n8036), .B2(P2_REG1_REG_9__SCAN_IN), .A(n8022), .ZN(
        n8078) );
  NOR2_X1 U9594 ( .A1(n8079), .A2(n8078), .ZN(n8077) );
  INV_X1 U9595 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8023) );
  MUX2_X1 U9596 ( .A(n8023), .B(P2_REG1_REG_10__SCAN_IN), .S(n8033), .Z(n8066)
         );
  NOR2_X1 U9597 ( .A1(n8067), .A2(n8066), .ZN(n8065) );
  AOI21_X1 U9598 ( .B1(n8033), .B2(P2_REG1_REG_10__SCAN_IN), .A(n8065), .ZN(
        n8165) );
  INV_X1 U9599 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8024) );
  MUX2_X1 U9600 ( .A(n8024), .B(P2_REG1_REG_11__SCAN_IN), .S(n8167), .Z(n8164)
         );
  NOR2_X1 U9601 ( .A1(n8165), .A2(n8164), .ZN(n8163) );
  INV_X1 U9602 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8025) );
  MUX2_X1 U9603 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8025), .S(n8122), .Z(n8026)
         );
  NAND2_X1 U9604 ( .A1(n8027), .A2(n8026), .ZN(n8121) );
  OAI21_X1 U9605 ( .B1(n8027), .B2(n8026), .A(n8121), .ZN(n8032) );
  INV_X1 U9606 ( .A(n8028), .ZN(n8031) );
  INV_X1 U9607 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8029) );
  NOR2_X1 U9608 ( .A1(n8479), .A2(n8029), .ZN(n8030) );
  AOI211_X1 U9609 ( .C1(n9714), .C2(n8032), .A(n8031), .B(n8030), .ZN(n8062)
         );
  NAND2_X1 U9610 ( .A1(n8033), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8054) );
  INV_X1 U9611 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8034) );
  MUX2_X1 U9612 ( .A(n8034), .B(P2_REG2_REG_10__SCAN_IN), .S(n8033), .Z(n8035)
         );
  INV_X1 U9613 ( .A(n8035), .ZN(n8071) );
  NAND2_X1 U9614 ( .A1(n8036), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8053) );
  INV_X1 U9615 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8037) );
  MUX2_X1 U9616 ( .A(n8037), .B(P2_REG2_REG_9__SCAN_IN), .S(n8036), .Z(n8038)
         );
  INV_X1 U9617 ( .A(n8038), .ZN(n8084) );
  INV_X1 U9618 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8052) );
  MUX2_X1 U9619 ( .A(n8052), .B(P2_REG2_REG_8__SCAN_IN), .S(n8099), .Z(n8095)
         );
  NAND2_X1 U9620 ( .A1(n8039), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8051) );
  MUX2_X1 U9621 ( .A(n6898), .B(P2_REG2_REG_7__SCAN_IN), .S(n8039), .Z(n8040)
         );
  INV_X1 U9622 ( .A(n8040), .ZN(n9878) );
  NAND2_X1 U9623 ( .A1(n8041), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8050) );
  INV_X1 U9624 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n8042) );
  MUX2_X1 U9625 ( .A(n8042), .B(P2_REG2_REG_6__SCAN_IN), .S(n8041), .Z(n8043)
         );
  INV_X1 U9626 ( .A(n8043), .ZN(n8107) );
  NAND2_X1 U9627 ( .A1(n8044), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8049) );
  INV_X1 U9628 ( .A(n8045), .ZN(n8046) );
  NAND2_X1 U9629 ( .A1(n8047), .A2(n8046), .ZN(n8048) );
  NAND2_X1 U9630 ( .A1(n8049), .A2(n8048), .ZN(n8108) );
  NAND2_X1 U9631 ( .A1(n8107), .A2(n8108), .ZN(n8106) );
  NAND2_X1 U9632 ( .A1(n8050), .A2(n8106), .ZN(n9879) );
  NAND2_X1 U9633 ( .A1(n9878), .A2(n9879), .ZN(n9876) );
  NAND2_X1 U9634 ( .A1(n8051), .A2(n9876), .ZN(n8096) );
  NAND2_X1 U9635 ( .A1(n8095), .A2(n8096), .ZN(n8094) );
  OAI21_X1 U9636 ( .B1(n8099), .B2(n8052), .A(n8094), .ZN(n8083) );
  NAND2_X1 U9637 ( .A1(n8084), .A2(n8083), .ZN(n8082) );
  NAND2_X1 U9638 ( .A1(n8053), .A2(n8082), .ZN(n8072) );
  NAND2_X1 U9639 ( .A1(n8071), .A2(n8072), .ZN(n8070) );
  NAND2_X1 U9640 ( .A1(n8054), .A2(n8070), .ZN(n8162) );
  MUX2_X1 U9641 ( .A(n8055), .B(P2_REG2_REG_11__SCAN_IN), .S(n8167), .Z(n8161)
         );
  NOR2_X1 U9642 ( .A1(n8162), .A2(n8161), .ZN(n8160) );
  AOI21_X1 U9643 ( .B1(n8056), .B2(n8055), .A(n8160), .ZN(n8060) );
  INV_X1 U9644 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8057) );
  MUX2_X1 U9645 ( .A(n8057), .B(P2_REG2_REG_12__SCAN_IN), .S(n8122), .Z(n8058)
         );
  INV_X1 U9646 ( .A(n8058), .ZN(n8059) );
  NAND2_X1 U9647 ( .A1(n8059), .A2(n8060), .ZN(n8112) );
  OAI211_X1 U9648 ( .C1(n8060), .C2(n8059), .A(n9877), .B(n8112), .ZN(n8061)
         );
  OAI211_X1 U9649 ( .C1(n9883), .C2(n8063), .A(n8062), .B(n8061), .ZN(P2_U3257) );
  INV_X1 U9650 ( .A(n8064), .ZN(n8069) );
  AOI211_X1 U9651 ( .C1(n8067), .C2(n8066), .A(n8065), .B(n9869), .ZN(n8068)
         );
  AOI211_X1 U9652 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n9875), .A(n8069), .B(
        n8068), .ZN(n8074) );
  OAI211_X1 U9653 ( .C1(n8072), .C2(n8071), .A(n9877), .B(n8070), .ZN(n8073)
         );
  OAI211_X1 U9654 ( .C1(n9883), .C2(n8075), .A(n8074), .B(n8073), .ZN(P2_U3255) );
  INV_X1 U9655 ( .A(n8076), .ZN(n8081) );
  AOI211_X1 U9656 ( .C1(n8079), .C2(n8078), .A(n8077), .B(n9869), .ZN(n8080)
         );
  AOI211_X1 U9657 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n9875), .A(n8081), .B(
        n8080), .ZN(n8086) );
  OAI211_X1 U9658 ( .C1(n8084), .C2(n8083), .A(n9877), .B(n8082), .ZN(n8085)
         );
  OAI211_X1 U9659 ( .C1(n9883), .C2(n8087), .A(n8086), .B(n8085), .ZN(P2_U3254) );
  INV_X1 U9660 ( .A(n8088), .ZN(n8093) );
  AOI211_X1 U9661 ( .C1(n8091), .C2(n8090), .A(n8089), .B(n9869), .ZN(n8092)
         );
  AOI211_X1 U9662 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n9875), .A(n8093), .B(
        n8092), .ZN(n8098) );
  OAI211_X1 U9663 ( .C1(n8096), .C2(n8095), .A(n9877), .B(n8094), .ZN(n8097)
         );
  OAI211_X1 U9664 ( .C1(n9883), .C2(n8099), .A(n8098), .B(n8097), .ZN(P2_U3253) );
  INV_X1 U9665 ( .A(n8100), .ZN(n8105) );
  AOI211_X1 U9666 ( .C1(n8103), .C2(n8102), .A(n8101), .B(n9869), .ZN(n8104)
         );
  AOI211_X1 U9667 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n9875), .A(n8105), .B(
        n8104), .ZN(n8110) );
  OAI211_X1 U9668 ( .C1(n8108), .C2(n8107), .A(n9877), .B(n8106), .ZN(n8109)
         );
  OAI211_X1 U9669 ( .C1(n9883), .C2(n8111), .A(n8110), .B(n8109), .ZN(P2_U3251) );
  NOR2_X1 U9670 ( .A1(n8124), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8117) );
  NOR2_X1 U9671 ( .A1(n8123), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8115) );
  NAND2_X1 U9672 ( .A1(n8122), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8113) );
  NAND2_X1 U9673 ( .A1(n8113), .A2(n8112), .ZN(n8149) );
  INV_X1 U9674 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8114) );
  AOI22_X1 U9675 ( .A1(n8123), .A2(n8114), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n8150), .ZN(n8148) );
  NOR2_X1 U9676 ( .A1(n8149), .A2(n8148), .ZN(n8147) );
  NOR2_X1 U9677 ( .A1(n8115), .A2(n8147), .ZN(n8136) );
  INV_X1 U9678 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8116) );
  AOI22_X1 U9679 ( .A1(n8124), .A2(n8116), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n8141), .ZN(n8135) );
  NOR2_X1 U9680 ( .A1(n8136), .A2(n8135), .ZN(n8134) );
  NOR2_X1 U9681 ( .A1(n8117), .A2(n8134), .ZN(n8421) );
  XNOR2_X1 U9682 ( .A(n8421), .B(n8422), .ZN(n8118) );
  NOR2_X1 U9683 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n8118), .ZN(n8423) );
  AOI21_X1 U9684 ( .B1(n8118), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8423), .ZN(
        n8133) );
  INV_X1 U9685 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8119) );
  AOI22_X1 U9686 ( .A1(n8124), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n8119), .B2(
        n8141), .ZN(n8139) );
  INV_X1 U9687 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8120) );
  AOI22_X1 U9688 ( .A1(n8123), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n8120), .B2(
        n8150), .ZN(n8155) );
  OAI21_X1 U9689 ( .B1(n8122), .B2(P2_REG1_REG_12__SCAN_IN), .A(n8121), .ZN(
        n8154) );
  NAND2_X1 U9690 ( .A1(n8155), .A2(n8154), .ZN(n8153) );
  OAI21_X1 U9691 ( .B1(n8123), .B2(P2_REG1_REG_13__SCAN_IN), .A(n8153), .ZN(
        n8138) );
  NAND2_X1 U9692 ( .A1(n8139), .A2(n8138), .ZN(n8137) );
  OAI21_X1 U9693 ( .B1(n8124), .B2(P2_REG1_REG_14__SCAN_IN), .A(n8137), .ZN(
        n8412) );
  XNOR2_X1 U9694 ( .A(n8412), .B(n8413), .ZN(n8125) );
  INV_X1 U9695 ( .A(n8125), .ZN(n8128) );
  INV_X1 U9696 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8126) );
  NOR2_X1 U9697 ( .A1(n8126), .A2(n8125), .ZN(n8414) );
  INV_X1 U9698 ( .A(n8414), .ZN(n8127) );
  OAI211_X1 U9699 ( .C1(n8128), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9714), .B(
        n8127), .ZN(n8132) );
  AND2_X1 U9700 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8130) );
  NOR2_X1 U9701 ( .A1(n9883), .A2(n8413), .ZN(n8129) );
  AOI211_X1 U9702 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n9875), .A(n8130), .B(
        n8129), .ZN(n8131) );
  OAI211_X1 U9703 ( .C1(n8133), .C2(n8474), .A(n8132), .B(n8131), .ZN(P2_U3260) );
  AOI21_X1 U9704 ( .B1(n8136), .B2(n8135), .A(n8134), .ZN(n8146) );
  OAI21_X1 U9705 ( .B1(n8139), .B2(n8138), .A(n8137), .ZN(n8140) );
  NAND2_X1 U9706 ( .A1(n8140), .A2(n9714), .ZN(n8145) );
  NOR2_X1 U9707 ( .A1(n9883), .A2(n8141), .ZN(n8142) );
  AOI211_X1 U9708 ( .C1(P2_ADDR_REG_14__SCAN_IN), .C2(n9875), .A(n8143), .B(
        n8142), .ZN(n8144) );
  OAI211_X1 U9709 ( .C1(n8146), .C2(n8474), .A(n8145), .B(n8144), .ZN(P2_U3259) );
  AOI21_X1 U9710 ( .B1(n8149), .B2(n8148), .A(n8147), .ZN(n8159) );
  NOR2_X1 U9711 ( .A1(n9883), .A2(n8150), .ZN(n8151) );
  AOI211_X1 U9712 ( .C1(P2_ADDR_REG_13__SCAN_IN), .C2(n9875), .A(n8152), .B(
        n8151), .ZN(n8158) );
  OAI21_X1 U9713 ( .B1(n8155), .B2(n8154), .A(n8153), .ZN(n8156) );
  NAND2_X1 U9714 ( .A1(n8156), .A2(n9714), .ZN(n8157) );
  OAI211_X1 U9715 ( .C1(n8159), .C2(n8474), .A(n8158), .B(n8157), .ZN(P2_U3258) );
  AOI21_X1 U9716 ( .B1(n8162), .B2(n8161), .A(n8160), .ZN(n8170) );
  NOR2_X1 U9717 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9953), .ZN(n8332) );
  AOI211_X1 U9718 ( .C1(n8165), .C2(n8164), .A(n8163), .B(n9869), .ZN(n8166)
         );
  AOI211_X1 U9719 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n9875), .A(n8332), .B(
        n8166), .ZN(n8169) );
  NAND2_X1 U9720 ( .A1(n9433), .A2(n8167), .ZN(n8168) );
  OAI211_X1 U9721 ( .C1(n8170), .C2(n8474), .A(n8169), .B(n8168), .ZN(P2_U3256) );
  INV_X1 U9722 ( .A(n9354), .ZN(n9173) );
  NOR2_X1 U9723 ( .A1(n8914), .A2(n9292), .ZN(n8172) );
  NAND2_X1 U9724 ( .A1(n8914), .A2(n9292), .ZN(n8171) );
  OAI21_X2 U9725 ( .B1(n8173), .B2(n8172), .A(n8171), .ZN(n9283) );
  OR2_X1 U9726 ( .A1(n9391), .A2(n9042), .ZN(n8174) );
  NAND2_X1 U9727 ( .A1(n9283), .A2(n8174), .ZN(n8176) );
  NAND2_X1 U9728 ( .A1(n9391), .A2(n9042), .ZN(n8175) );
  NAND2_X1 U9729 ( .A1(n8176), .A2(n8175), .ZN(n9265) );
  NAND2_X1 U9730 ( .A1(n9388), .A2(n9294), .ZN(n8177) );
  OR2_X1 U9731 ( .A1(n9383), .A2(n9239), .ZN(n8178) );
  NOR2_X1 U9732 ( .A1(n9372), .A2(n9240), .ZN(n8181) );
  NAND2_X1 U9733 ( .A1(n9377), .A2(n9227), .ZN(n9216) );
  NAND2_X1 U9734 ( .A1(n9372), .A2(n9240), .ZN(n8179) );
  AND2_X1 U9735 ( .A1(n9216), .A2(n8179), .ZN(n8180) );
  OR2_X1 U9736 ( .A1(n8181), .A2(n8180), .ZN(n8182) );
  AND2_X1 U9737 ( .A1(n9368), .A2(n9228), .ZN(n8184) );
  OAI21_X1 U9738 ( .B1(n4734), .B2(n9142), .A(n9150), .ZN(n8185) );
  OAI21_X1 U9739 ( .B1(n9176), .B2(n9349), .A(n8185), .ZN(n9145) );
  NOR2_X1 U9740 ( .A1(n9145), .A2(n9144), .ZN(n9348) );
  NOR2_X1 U9741 ( .A1(n9332), .A2(n9130), .ZN(n8187) );
  XNOR2_X1 U9742 ( .A(n8189), .B(n8218), .ZN(n9321) );
  AOI21_X1 U9743 ( .B1(n9317), .B2(n9080), .A(n9073), .ZN(n9318) );
  AOI22_X1 U9744 ( .A1(n8190), .A2(n9652), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n4419), .ZN(n8191) );
  OAI21_X1 U9745 ( .B1(n8192), .B2(n9656), .A(n8191), .ZN(n8223) );
  AND2_X1 U9746 ( .A1(n9040), .A2(n8193), .ZN(n8194) );
  AOI21_X1 U9747 ( .B1(n9041), .B2(n9291), .A(n8194), .ZN(n8221) );
  NAND2_X1 U9748 ( .A1(n8196), .A2(n8195), .ZN(n9290) );
  NAND2_X1 U9749 ( .A1(n9290), .A2(n8197), .ZN(n9267) );
  AOI21_X2 U9750 ( .B1(n9267), .B2(n8199), .A(n8198), .ZN(n9250) );
  INV_X1 U9751 ( .A(n8203), .ZN(n9202) );
  NAND3_X1 U9752 ( .A1(n9224), .A2(n9204), .A3(n9202), .ZN(n8205) );
  NAND2_X1 U9753 ( .A1(n8205), .A2(n8204), .ZN(n9188) );
  NOR2_X1 U9754 ( .A1(n9188), .A2(n9189), .ZN(n9187) );
  INV_X1 U9755 ( .A(n8206), .ZN(n8207) );
  NOR2_X1 U9756 ( .A1(n9187), .A2(n8207), .ZN(n9175) );
  INV_X1 U9757 ( .A(n8212), .ZN(n8213) );
  NOR2_X1 U9758 ( .A1(n9093), .A2(n8216), .ZN(n9087) );
  NAND2_X1 U9759 ( .A1(n9087), .A2(n9088), .ZN(n9086) );
  NAND2_X1 U9760 ( .A1(n9086), .A2(n8217), .ZN(n8219) );
  XNOR2_X1 U9761 ( .A(n8219), .B(n8218), .ZN(n8220) );
  OAI21_X1 U9762 ( .B1(n9321), .B2(n9308), .A(n8224), .ZN(P1_U3355) );
  INV_X1 U9763 ( .A(n8225), .ZN(n9420) );
  OAI222_X1 U9764 ( .A1(P2_U3152), .A2(n8227), .B1(n8236), .B2(n9420), .C1(
        n8226), .C2(n8881), .ZN(P2_U3329) );
  INV_X1 U9765 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8230) );
  INV_X1 U9766 ( .A(n8228), .ZN(n8234) );
  OAI222_X1 U9767 ( .A1(n8231), .A2(n8230), .B1(n9424), .B2(n8234), .C1(n8229), 
        .C2(P1_U3084), .ZN(P1_U3323) );
  INV_X1 U9768 ( .A(n8235), .ZN(n9425) );
  OAI222_X1 U9769 ( .A1(n8237), .A2(n10185), .B1(n8236), .B2(n9425), .C1(n5721), .C2(P2_U3152), .ZN(P2_U3330) );
  OAI211_X1 U9770 ( .C1(n8240), .C2(n8239), .A(n8238), .B(n8353), .ZN(n8244)
         );
  NOR2_X1 U9771 ( .A1(n10144), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8242) );
  OAI22_X1 U9772 ( .A1(n8275), .A2(n8370), .B1(n8369), .B2(n8494), .ZN(n8241)
         );
  AOI211_X1 U9773 ( .C1(n8345), .C2(n8510), .A(n8242), .B(n8241), .ZN(n8243)
         );
  OAI211_X1 U9774 ( .C1(n4679), .C2(n8348), .A(n8244), .B(n8243), .ZN(P2_U3216) );
  INV_X1 U9775 ( .A(n8301), .ZN(n8245) );
  OAI211_X1 U9776 ( .C1(n8247), .C2(n8246), .A(n8245), .B(n8353), .ZN(n8252)
         );
  AOI22_X1 U9777 ( .A1(n8345), .A2(n8574), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8251) );
  INV_X1 U9778 ( .A(n8248), .ZN(n8605) );
  AOI22_X1 U9779 ( .A1(n8316), .A2(n8605), .B1(n8315), .B2(n8570), .ZN(n8250)
         );
  NAND2_X1 U9780 ( .A1(n8803), .A2(n8374), .ZN(n8249) );
  NAND4_X1 U9781 ( .A1(n8252), .A2(n8251), .A3(n8250), .A4(n8249), .ZN(
        P2_U3218) );
  INV_X1 U9782 ( .A(n8253), .ZN(n8254) );
  AOI21_X1 U9783 ( .B1(n8256), .B2(n8255), .A(n8254), .ZN(n8264) );
  INV_X1 U9784 ( .A(n8633), .ZN(n8261) );
  OR2_X1 U9785 ( .A1(n8669), .A2(n9734), .ZN(n8259) );
  OR2_X1 U9786 ( .A1(n8257), .A2(n9732), .ZN(n8258) );
  NAND2_X1 U9787 ( .A1(n8259), .A2(n8258), .ZN(n8640) );
  AOI22_X1 U9788 ( .A1(n8358), .A2(n8640), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8260) );
  OAI21_X1 U9789 ( .B1(n8261), .B2(n8368), .A(n8260), .ZN(n8262) );
  AOI21_X1 U9790 ( .B1(n8824), .B2(n8374), .A(n8262), .ZN(n8263) );
  OAI21_X1 U9791 ( .B1(n8264), .B2(n8376), .A(n8263), .ZN(P2_U3221) );
  OAI211_X1 U9792 ( .C1(n8267), .C2(n8266), .A(n8265), .B(n8353), .ZN(n8271)
         );
  AOI22_X1 U9793 ( .A1(n8345), .A2(n8598), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8270) );
  AOI22_X1 U9794 ( .A1(n8316), .A2(n8604), .B1(n8315), .B2(n8605), .ZN(n8269)
         );
  NAND2_X1 U9795 ( .A1(n8813), .A2(n8374), .ZN(n8268) );
  NAND4_X1 U9796 ( .A1(n8271), .A2(n8270), .A3(n8269), .A4(n8268), .ZN(
        P2_U3225) );
  INV_X1 U9797 ( .A(n8273), .ZN(n8545) );
  OAI22_X1 U9798 ( .A1(n8275), .A2(n9732), .B1(n8274), .B2(n9734), .ZN(n8540)
         );
  INV_X1 U9799 ( .A(n8540), .ZN(n8277) );
  OAI22_X1 U9800 ( .A1(n8278), .A2(n8277), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8276), .ZN(n8279) );
  AOI21_X1 U9801 ( .B1(n8545), .B2(n8345), .A(n8279), .ZN(n8280) );
  OAI211_X1 U9802 ( .C1(n8549), .C2(n8348), .A(n8281), .B(n8280), .ZN(P2_U3227) );
  XNOR2_X1 U9803 ( .A(n8282), .B(n8283), .ZN(n8365) );
  NOR2_X1 U9804 ( .A1(n8365), .A2(n8364), .ZN(n8363) );
  AOI21_X1 U9805 ( .B1(n8283), .B2(n8282), .A(n8363), .ZN(n8287) );
  XNOR2_X1 U9806 ( .A(n8285), .B(n8284), .ZN(n8286) );
  XNOR2_X1 U9807 ( .A(n8287), .B(n8286), .ZN(n8292) );
  INV_X1 U9808 ( .A(n8689), .ZN(n8289) );
  AOI22_X1 U9809 ( .A1(n8316), .A2(n8381), .B1(n8315), .B2(n8653), .ZN(n8288)
         );
  NAND2_X1 U9810 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8419) );
  OAI211_X1 U9811 ( .C1(n8289), .C2(n8368), .A(n8288), .B(n8419), .ZN(n8290)
         );
  AOI21_X1 U9812 ( .B1(n8838), .B2(n8374), .A(n8290), .ZN(n8291) );
  OAI21_X1 U9813 ( .B1(n8292), .B2(n8376), .A(n8291), .ZN(P2_U3228) );
  AOI21_X1 U9814 ( .B1(n8294), .B2(n8293), .A(n8376), .ZN(n8296) );
  NAND2_X1 U9815 ( .A1(n8296), .A2(n8295), .ZN(n8299) );
  NOR2_X1 U9816 ( .A1(n9951), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8437) );
  OAI22_X1 U9817 ( .A1(n8666), .A2(n8370), .B1(n8369), .B2(n8669), .ZN(n8297)
         );
  AOI211_X1 U9818 ( .C1(n8345), .C2(n8673), .A(n8437), .B(n8297), .ZN(n8298)
         );
  OAI211_X1 U9819 ( .C1(n4814), .C2(n8348), .A(n8299), .B(n8298), .ZN(P2_U3230) );
  NOR2_X1 U9820 ( .A1(n8301), .A2(n8300), .ZN(n8303) );
  XNOR2_X1 U9821 ( .A(n8303), .B(n8302), .ZN(n8305) );
  AOI21_X1 U9822 ( .B1(n8305), .B2(n8306), .A(n8376), .ZN(n8304) );
  OAI21_X1 U9823 ( .B1(n8306), .B2(n8305), .A(n8304), .ZN(n8311) );
  INV_X1 U9824 ( .A(n8557), .ZN(n8307) );
  NOR2_X1 U9825 ( .A1(n8368), .A2(n8307), .ZN(n8309) );
  OAI22_X1 U9826 ( .A1(n8591), .A2(n8370), .B1(n8369), .B2(n8561), .ZN(n8308)
         );
  AOI211_X1 U9827 ( .C1(P2_REG3_REG_24__SCAN_IN), .C2(P2_U3152), .A(n8309), 
        .B(n8308), .ZN(n8310) );
  OAI211_X1 U9828 ( .C1(n4695), .C2(n8348), .A(n8311), .B(n8310), .ZN(P2_U3231) );
  OAI211_X1 U9829 ( .C1(n8314), .C2(n8313), .A(n8312), .B(n8353), .ZN(n8320)
         );
  AOI22_X1 U9830 ( .A1(n8345), .A2(n8614), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8319) );
  AOI22_X1 U9831 ( .A1(n8316), .A2(n8652), .B1(n8315), .B2(n8380), .ZN(n8318)
         );
  NAND2_X1 U9832 ( .A1(n8818), .A2(n8374), .ZN(n8317) );
  NAND4_X1 U9833 ( .A1(n8320), .A2(n8319), .A3(n8318), .A4(n8317), .ZN(
        P2_U3235) );
  XOR2_X1 U9834 ( .A(n8322), .B(n8321), .Z(n8328) );
  INV_X1 U9835 ( .A(n8585), .ZN(n8324) );
  OAI22_X1 U9836 ( .A1(n8368), .A2(n8324), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8323), .ZN(n8326) );
  OAI22_X1 U9837 ( .A1(n8623), .A2(n8370), .B1(n8369), .B2(n8591), .ZN(n8325)
         );
  AOI211_X1 U9838 ( .C1(n8808), .C2(n8374), .A(n8326), .B(n8325), .ZN(n8327)
         );
  OAI21_X1 U9839 ( .B1(n8328), .B2(n8376), .A(n8327), .ZN(P2_U3237) );
  XOR2_X1 U9840 ( .A(n8330), .B(n8329), .Z(n8331) );
  NAND2_X1 U9841 ( .A1(n8331), .A2(n8353), .ZN(n8339) );
  AOI21_X1 U9842 ( .B1(n8358), .B2(n8333), .A(n8332), .ZN(n8338) );
  NAND2_X1 U9843 ( .A1(n8374), .A2(n8334), .ZN(n8337) );
  OR2_X1 U9844 ( .A1(n8368), .A2(n8335), .ZN(n8336) );
  NAND4_X1 U9845 ( .A1(n8339), .A2(n8338), .A3(n8337), .A4(n8336), .ZN(
        P2_U3238) );
  OAI211_X1 U9846 ( .C1(n8342), .C2(n8341), .A(n8340), .B(n8353), .ZN(n8347)
         );
  NOR2_X1 U9847 ( .A1(n8343), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8452) );
  OAI22_X1 U9848 ( .A1(n8680), .A2(n8370), .B1(n8369), .B2(n8624), .ZN(n8344)
         );
  AOI211_X1 U9849 ( .C1(n8345), .C2(n8647), .A(n8452), .B(n8344), .ZN(n8346)
         );
  OAI211_X1 U9850 ( .C1(n8649), .C2(n8348), .A(n8347), .B(n8346), .ZN(P2_U3240) );
  NAND2_X1 U9851 ( .A1(n8350), .A2(n8349), .ZN(n8356) );
  AND2_X1 U9852 ( .A1(n8352), .A2(n8351), .ZN(n8354) );
  OAI211_X1 U9853 ( .C1(n8356), .C2(n8355), .A(n8354), .B(n8353), .ZN(n8362)
         );
  OAI22_X1 U9854 ( .A1(n8357), .A2(n9732), .B1(n8561), .B2(n9734), .ZN(n8531)
         );
  AOI22_X1 U9855 ( .A1(n8358), .A2(n8531), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8359) );
  OAI21_X1 U9856 ( .B1(n8524), .B2(n8368), .A(n8359), .ZN(n8360) );
  AOI21_X1 U9857 ( .B1(n8787), .B2(n8374), .A(n8360), .ZN(n8361) );
  NAND2_X1 U9858 ( .A1(n8362), .A2(n8361), .ZN(P2_U3242) );
  AOI21_X1 U9859 ( .B1(n8365), .B2(n8364), .A(n8363), .ZN(n8377) );
  INV_X1 U9860 ( .A(n8699), .ZN(n8367) );
  OAI22_X1 U9861 ( .A1(n8368), .A2(n8367), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8366), .ZN(n8373) );
  OAI22_X1 U9862 ( .A1(n8371), .A2(n8370), .B1(n8369), .B2(n8666), .ZN(n8372)
         );
  AOI211_X1 U9863 ( .C1(n8843), .C2(n8374), .A(n8373), .B(n8372), .ZN(n8375)
         );
  OAI21_X1 U9864 ( .B1(n8377), .B2(n8376), .A(n8375), .ZN(P2_U3243) );
  INV_X1 U9865 ( .A(n8494), .ZN(n8515) );
  MUX2_X1 U9866 ( .A(n8515), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8392), .Z(
        P2_U3580) );
  MUX2_X1 U9867 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8378), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9868 ( .A(n8514), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8392), .Z(
        P2_U3578) );
  MUX2_X1 U9869 ( .A(n8379), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8392), .Z(
        P2_U3577) );
  MUX2_X1 U9870 ( .A(n8570), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8392), .Z(
        P2_U3576) );
  MUX2_X1 U9871 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8605), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9872 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8380), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9873 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8604), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9874 ( .A(n8652), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8392), .Z(
        P2_U3571) );
  MUX2_X1 U9875 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8653), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9876 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8705), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9877 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8381), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9878 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8704), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9879 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8382), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9880 ( .A(n8383), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8392), .Z(
        P2_U3564) );
  MUX2_X1 U9881 ( .A(n8384), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8392), .Z(
        P2_U3563) );
  MUX2_X1 U9882 ( .A(n8385), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8392), .Z(
        P2_U3562) );
  MUX2_X1 U9883 ( .A(n8386), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8392), .Z(
        P2_U3561) );
  MUX2_X1 U9884 ( .A(n8387), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8392), .Z(
        P2_U3560) );
  MUX2_X1 U9885 ( .A(n8732), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8392), .Z(
        P2_U3559) );
  MUX2_X1 U9886 ( .A(n8388), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8392), .Z(
        P2_U3558) );
  MUX2_X1 U9887 ( .A(n8730), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8392), .Z(
        P2_U3557) );
  MUX2_X1 U9888 ( .A(n8389), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8392), .Z(
        P2_U3556) );
  MUX2_X1 U9889 ( .A(n8390), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8392), .Z(
        P2_U3555) );
  MUX2_X1 U9890 ( .A(n8391), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8392), .Z(
        P2_U3554) );
  MUX2_X1 U9891 ( .A(n6449), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8392), .Z(
        P2_U3553) );
  INV_X1 U9892 ( .A(n8393), .ZN(n8396) );
  MUX2_X1 U9893 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n8394), .S(n8402), .Z(n8395)
         );
  NAND2_X1 U9894 ( .A1(n8396), .A2(n8395), .ZN(n8398) );
  OAI211_X1 U9895 ( .C1(n8399), .C2(n8398), .A(n9877), .B(n8397), .ZN(n8411)
         );
  NOR2_X1 U9896 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8400), .ZN(n8401) );
  AOI21_X1 U9897 ( .B1(n9875), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n8401), .ZN(
        n8410) );
  INV_X1 U9898 ( .A(n8402), .ZN(n8403) );
  NAND2_X1 U9899 ( .A1(n9433), .A2(n8403), .ZN(n8409) );
  OAI21_X1 U9900 ( .B1(n8406), .B2(n8405), .A(n8404), .ZN(n8407) );
  OR2_X1 U9901 ( .A1(n9869), .A2(n8407), .ZN(n8408) );
  NAND4_X1 U9902 ( .A1(n8411), .A2(n8410), .A3(n8409), .A4(n8408), .ZN(
        P2_U3249) );
  NOR2_X1 U9903 ( .A1(n8413), .A2(n8412), .ZN(n8415) );
  XOR2_X1 U9904 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8439), .Z(n8416) );
  NAND2_X1 U9905 ( .A1(n8416), .A2(n8417), .ZN(n8440) );
  OAI21_X1 U9906 ( .B1(n8417), .B2(n8416), .A(n8440), .ZN(n8418) );
  NAND2_X1 U9907 ( .A1(n8418), .A2(n9714), .ZN(n8431) );
  INV_X1 U9908 ( .A(n8419), .ZN(n8420) );
  AOI21_X1 U9909 ( .B1(n9875), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8420), .ZN(
        n8430) );
  NOR2_X1 U9910 ( .A1(n8422), .A2(n8421), .ZN(n8424) );
  NOR2_X1 U9911 ( .A1(n8424), .A2(n8423), .ZN(n8427) );
  OR2_X1 U9912 ( .A1(n8439), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U9913 ( .A1(n8439), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8433) );
  AND2_X1 U9914 ( .A1(n8425), .A2(n8433), .ZN(n8426) );
  NAND2_X1 U9915 ( .A1(n8426), .A2(n8427), .ZN(n8432) );
  OAI211_X1 U9916 ( .C1(n8427), .C2(n8426), .A(n9877), .B(n8432), .ZN(n8429)
         );
  NAND2_X1 U9917 ( .A1(n9433), .A2(n8439), .ZN(n8428) );
  NAND4_X1 U9918 ( .A1(n8431), .A2(n8430), .A3(n8429), .A4(n8428), .ZN(
        P2_U3261) );
  NAND2_X1 U9919 ( .A1(n8433), .A2(n8432), .ZN(n8436) );
  INV_X1 U9920 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8434) );
  MUX2_X1 U9921 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n8434), .S(n8455), .Z(n8435)
         );
  NAND2_X1 U9922 ( .A1(n8435), .A2(n8436), .ZN(n8449) );
  OAI211_X1 U9923 ( .C1(n8436), .C2(n8435), .A(n9877), .B(n8449), .ZN(n8448)
         );
  AOI21_X1 U9924 ( .B1(n9875), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8437), .ZN(
        n8447) );
  OR2_X1 U9925 ( .A1(n9883), .A2(n8438), .ZN(n8446) );
  XNOR2_X1 U9926 ( .A(n8455), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8443) );
  OR2_X1 U9927 ( .A1(n8439), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8441) );
  NAND2_X1 U9928 ( .A1(n8441), .A2(n8440), .ZN(n8442) );
  NOR2_X1 U9929 ( .A1(n8443), .A2(n8442), .ZN(n8454) );
  AOI21_X1 U9930 ( .B1(n8443), .B2(n8442), .A(n8454), .ZN(n8444) );
  NAND2_X1 U9931 ( .A1(n9714), .A2(n8444), .ZN(n8445) );
  NAND4_X1 U9932 ( .A1(n8448), .A2(n8447), .A3(n8446), .A4(n8445), .ZN(
        P2_U3262) );
  NAND2_X1 U9933 ( .A1(n8455), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8450) );
  NAND2_X1 U9934 ( .A1(n8450), .A2(n8449), .ZN(n8463) );
  XOR2_X1 U9935 ( .A(n8468), .B(n8463), .Z(n8451) );
  NAND2_X1 U9936 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8451), .ZN(n8465) );
  OAI211_X1 U9937 ( .C1(n8451), .C2(P2_REG2_REG_18__SCAN_IN), .A(n9877), .B(
        n8465), .ZN(n8462) );
  AOI21_X1 U9938 ( .B1(n9875), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8452), .ZN(
        n8461) );
  OR2_X1 U9939 ( .A1(n9883), .A2(n8453), .ZN(n8460) );
  INV_X1 U9940 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n10042) );
  XNOR2_X1 U9941 ( .A(n8468), .B(n10042), .ZN(n8457) );
  NAND2_X1 U9942 ( .A1(n8456), .A2(n8457), .ZN(n8467) );
  OAI21_X1 U9943 ( .B1(n8457), .B2(n8456), .A(n8467), .ZN(n8458) );
  NAND2_X1 U9944 ( .A1(n9714), .A2(n8458), .ZN(n8459) );
  NAND4_X1 U9945 ( .A1(n8462), .A2(n8461), .A3(n8460), .A4(n8459), .ZN(
        P2_U3263) );
  NAND2_X1 U9946 ( .A1(n8468), .A2(n8463), .ZN(n8464) );
  NAND2_X1 U9947 ( .A1(n8465), .A2(n8464), .ZN(n8466) );
  XNOR2_X1 U9948 ( .A(n8466), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U9949 ( .A1(n8475), .A2(n9877), .ZN(n8472) );
  OAI21_X1 U9950 ( .B1(n8468), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8467), .ZN(
        n8470) );
  INV_X1 U9951 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8469) );
  XNOR2_X1 U9952 ( .A(n8470), .B(n8469), .ZN(n8473) );
  NAND2_X1 U9953 ( .A1(n8473), .A2(n9714), .ZN(n8471) );
  NAND3_X1 U9954 ( .A1(n8472), .A2(n8471), .A3(n9883), .ZN(n8477) );
  OAI22_X1 U9955 ( .A1(n8475), .A2(n8474), .B1(n8473), .B2(n9869), .ZN(n8476)
         );
  NAND2_X1 U9956 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8478) );
  INV_X1 U9957 ( .A(n8481), .ZN(n8768) );
  INV_X1 U9958 ( .A(n8480), .ZN(n8765) );
  NAND2_X1 U9959 ( .A1(n8481), .A2(n4455), .ZN(n8764) );
  NAND3_X1 U9960 ( .A1(n8765), .A2(n9727), .A3(n8764), .ZN(n8484) );
  AOI21_X1 U9961 ( .B1(n9745), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8482), .ZN(
        n8483) );
  OAI211_X1 U9962 ( .C1(n8768), .C2(n9747), .A(n8484), .B(n8483), .ZN(P2_U3266) );
  INV_X1 U9963 ( .A(n8769), .ZN(n8506) );
  INV_X1 U9964 ( .A(n8488), .ZN(n8489) );
  XNOR2_X1 U9965 ( .A(n8490), .B(n8489), .ZN(n8491) );
  NAND2_X1 U9966 ( .A1(n8491), .A2(n9737), .ZN(n8497) );
  OAI22_X1 U9967 ( .A1(n8494), .A2(n9734), .B1(n8493), .B2(n8492), .ZN(n8495)
         );
  INV_X1 U9968 ( .A(n8495), .ZN(n8496) );
  NAND2_X1 U9969 ( .A1(n8497), .A2(n8496), .ZN(n8773) );
  OAI21_X1 U9970 ( .B1(n8498), .B2(n8770), .A(n4455), .ZN(n8771) );
  NOR2_X1 U9971 ( .A1(n8771), .A2(n8499), .ZN(n8504) );
  INV_X1 U9972 ( .A(n8500), .ZN(n8501) );
  AOI22_X1 U9973 ( .A1(n9745), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8501), .B2(
        n8752), .ZN(n8502) );
  OAI21_X1 U9974 ( .B1(n8770), .B2(n9747), .A(n8502), .ZN(n8503) );
  AOI211_X1 U9975 ( .C1(n8773), .C2(n9749), .A(n8504), .B(n8503), .ZN(n8505)
         );
  OAI21_X1 U9976 ( .B1(n8506), .B2(n8727), .A(n8505), .ZN(P2_U3267) );
  XNOR2_X1 U9977 ( .A(n8508), .B(n8507), .ZN(n8785) );
  AOI21_X1 U9978 ( .B1(n8781), .B2(n8522), .A(n8509), .ZN(n8782) );
  AOI22_X1 U9979 ( .A1(n8754), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8510), .B2(
        n8752), .ZN(n8511) );
  OAI21_X1 U9980 ( .B1(n4679), .B2(n9747), .A(n8511), .ZN(n8518) );
  XNOR2_X1 U9981 ( .A(n8513), .B(n8512), .ZN(n8516) );
  AOI222_X1 U9982 ( .A1(n9737), .A2(n8516), .B1(n8515), .B2(n8731), .C1(n8514), 
        .C2(n8729), .ZN(n8784) );
  NOR2_X1 U9983 ( .A1(n8784), .A2(n8754), .ZN(n8517) );
  OAI21_X1 U9984 ( .B1(n8785), .B2(n8727), .A(n8519), .ZN(P2_U3269) );
  XNOR2_X1 U9985 ( .A(n8521), .B(n8520), .ZN(n8790) );
  INV_X1 U9986 ( .A(n8522), .ZN(n8523) );
  AOI211_X1 U9987 ( .C1(n8787), .C2(n8543), .A(n9820), .B(n8523), .ZN(n8786)
         );
  INV_X1 U9988 ( .A(n8524), .ZN(n8525) );
  AOI22_X1 U9989 ( .A1(n8754), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8525), .B2(
        n8752), .ZN(n8526) );
  OAI21_X1 U9990 ( .B1(n8527), .B2(n9747), .A(n8526), .ZN(n8534) );
  NAND2_X1 U9991 ( .A1(n8541), .A2(n8528), .ZN(n8530) );
  XNOR2_X1 U9992 ( .A(n8530), .B(n8529), .ZN(n8532) );
  AOI21_X1 U9993 ( .B1(n8532), .B2(n9737), .A(n8531), .ZN(n8789) );
  NOR2_X1 U9994 ( .A1(n8789), .A2(n8754), .ZN(n8533) );
  AOI211_X1 U9995 ( .C1(n8786), .C2(n8672), .A(n8534), .B(n8533), .ZN(n8535)
         );
  OAI21_X1 U9996 ( .B1(n8790), .B2(n8727), .A(n8535), .ZN(P2_U3270) );
  XNOR2_X1 U9997 ( .A(n8536), .B(n8538), .ZN(n8795) );
  NOR3_X1 U9998 ( .A1(n8559), .A2(n8538), .A3(n8537), .ZN(n8539) );
  NOR2_X1 U9999 ( .A1(n8539), .A2(n8620), .ZN(n8542) );
  AOI21_X1 U10000 ( .B1(n8542), .B2(n8541), .A(n8540), .ZN(n8794) );
  INV_X1 U10001 ( .A(n8543), .ZN(n8544) );
  AOI211_X1 U10002 ( .C1(n8792), .C2(n4495), .A(n9820), .B(n8544), .ZN(n8791)
         );
  AOI22_X1 U10003 ( .A1(n8791), .A2(n8546), .B1(n8752), .B2(n8545), .ZN(n8547)
         );
  AOI21_X1 U10004 ( .B1(n8794), .B2(n8547), .A(n8656), .ZN(n8551) );
  OAI22_X1 U10005 ( .A1(n8549), .A2(n9747), .B1(n9749), .B2(n8548), .ZN(n8550)
         );
  NOR2_X1 U10006 ( .A1(n8551), .A2(n8550), .ZN(n8552) );
  OAI21_X1 U10007 ( .B1(n8795), .B2(n8727), .A(n8552), .ZN(P2_U3271) );
  INV_X1 U10008 ( .A(n8553), .ZN(n8554) );
  AOI21_X1 U10009 ( .B1(n8556), .B2(n8555), .A(n8554), .ZN(n8800) );
  XNOR2_X1 U10010 ( .A(n8572), .B(n4695), .ZN(n8797) );
  AOI22_X1 U10011 ( .A1(n8754), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8557), .B2(
        n8752), .ZN(n8558) );
  OAI21_X1 U10012 ( .B1(n4695), .B2(n9747), .A(n8558), .ZN(n8565) );
  AOI211_X1 U10013 ( .C1(n4661), .C2(n8560), .A(n8620), .B(n8559), .ZN(n8563)
         );
  OAI22_X1 U10014 ( .A1(n8561), .A2(n9732), .B1(n8591), .B2(n9734), .ZN(n8562)
         );
  NOR2_X1 U10015 ( .A1(n8563), .A2(n8562), .ZN(n8799) );
  NOR2_X1 U10016 ( .A1(n8799), .A2(n9745), .ZN(n8564) );
  AOI211_X1 U10017 ( .C1(n8797), .C2(n9727), .A(n8565), .B(n8564), .ZN(n8566)
         );
  OAI21_X1 U10018 ( .B1(n8800), .B2(n8727), .A(n8566), .ZN(P2_U3272) );
  OAI21_X1 U10019 ( .B1(n8569), .B2(n8568), .A(n8567), .ZN(n8571) );
  AOI222_X1 U10020 ( .A1(n9737), .A2(n8571), .B1(n8570), .B2(n8731), .C1(n8605), .C2(n8729), .ZN(n8806) );
  INV_X1 U10021 ( .A(n8572), .ZN(n8573) );
  AOI21_X1 U10022 ( .B1(n8803), .B2(n8582), .A(n8573), .ZN(n8804) );
  AOI22_X1 U10023 ( .A1(n9745), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8574), .B2(
        n8752), .ZN(n8575) );
  OAI21_X1 U10024 ( .B1(n4696), .B2(n9747), .A(n8575), .ZN(n8576) );
  AOI21_X1 U10025 ( .B1(n8804), .B2(n9727), .A(n8576), .ZN(n8580) );
  OR2_X1 U10026 ( .A1(n8578), .A2(n8577), .ZN(n8802) );
  NAND3_X1 U10027 ( .A1(n8802), .A2(n8801), .A3(n8751), .ZN(n8579) );
  OAI211_X1 U10028 ( .C1(n8806), .C2(n8656), .A(n8580), .B(n8579), .ZN(
        P2_U3273) );
  XOR2_X1 U10029 ( .A(n8590), .B(n8581), .Z(n8812) );
  INV_X1 U10030 ( .A(n8582), .ZN(n8584) );
  AOI21_X1 U10031 ( .B1(n8612), .B2(n8600), .A(n8587), .ZN(n8583) );
  NOR2_X1 U10032 ( .A1(n8584), .A2(n8583), .ZN(n8809) );
  AOI22_X1 U10033 ( .A1(n8656), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8585), .B2(
        n8752), .ZN(n8586) );
  OAI21_X1 U10034 ( .B1(n8587), .B2(n9747), .A(n8586), .ZN(n8595) );
  AOI211_X1 U10035 ( .C1(n8590), .C2(n8589), .A(n8620), .B(n8588), .ZN(n8593)
         );
  OAI22_X1 U10036 ( .A1(n8623), .A2(n9734), .B1(n8591), .B2(n9732), .ZN(n8592)
         );
  NOR2_X1 U10037 ( .A1(n8593), .A2(n8592), .ZN(n8811) );
  NOR2_X1 U10038 ( .A1(n8811), .A2(n8656), .ZN(n8594) );
  AOI211_X1 U10039 ( .C1(n8809), .C2(n9727), .A(n8595), .B(n8594), .ZN(n8596)
         );
  OAI21_X1 U10040 ( .B1(n8812), .B2(n8727), .A(n8596), .ZN(P2_U3274) );
  XNOR2_X1 U10041 ( .A(n8597), .B(n8602), .ZN(n8817) );
  XNOR2_X1 U10042 ( .A(n8612), .B(n8813), .ZN(n8814) );
  AOI22_X1 U10043 ( .A1(n9745), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8598), .B2(
        n8752), .ZN(n8599) );
  OAI21_X1 U10044 ( .B1(n8600), .B2(n9747), .A(n8599), .ZN(n8608) );
  OAI21_X1 U10045 ( .B1(n8603), .B2(n8602), .A(n8601), .ZN(n8606) );
  AOI222_X1 U10046 ( .A1(n9737), .A2(n8606), .B1(n8605), .B2(n8731), .C1(n8604), .C2(n8729), .ZN(n8816) );
  NOR2_X1 U10047 ( .A1(n8816), .A2(n8656), .ZN(n8607) );
  AOI211_X1 U10048 ( .C1(n8814), .C2(n9727), .A(n8608), .B(n8607), .ZN(n8609)
         );
  OAI21_X1 U10049 ( .B1(n8817), .B2(n8727), .A(n8609), .ZN(P2_U3275) );
  XNOR2_X1 U10050 ( .A(n8611), .B(n8610), .ZN(n8822) );
  INV_X1 U10051 ( .A(n8631), .ZN(n8613) );
  AOI21_X1 U10052 ( .B1(n8818), .B2(n8613), .A(n8612), .ZN(n8819) );
  AOI22_X1 U10053 ( .A1(n8754), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8614), .B2(
        n8752), .ZN(n8615) );
  OAI21_X1 U10054 ( .B1(n8616), .B2(n9747), .A(n8615), .ZN(n8628) );
  AOI21_X1 U10055 ( .B1(n8617), .B2(n8619), .A(n8618), .ZN(n8621) );
  NOR3_X1 U10056 ( .A1(n8622), .A2(n8621), .A3(n8620), .ZN(n8626) );
  OAI22_X1 U10057 ( .A1(n8624), .A2(n9734), .B1(n8623), .B2(n9732), .ZN(n8625)
         );
  NOR2_X1 U10058 ( .A1(n8626), .A2(n8625), .ZN(n8821) );
  NOR2_X1 U10059 ( .A1(n8821), .A2(n8656), .ZN(n8627) );
  AOI211_X1 U10060 ( .C1(n8819), .C2(n9727), .A(n8628), .B(n8627), .ZN(n8629)
         );
  OAI21_X1 U10061 ( .B1(n8727), .B2(n8822), .A(n8629), .ZN(P2_U3276) );
  XOR2_X1 U10062 ( .A(n8638), .B(n8630), .Z(n8827) );
  INV_X1 U10063 ( .A(n8646), .ZN(n8632) );
  AOI211_X1 U10064 ( .C1(n8824), .C2(n8632), .A(n9820), .B(n8631), .ZN(n8823)
         );
  AOI22_X1 U10065 ( .A1(n8754), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8633), .B2(
        n8752), .ZN(n8634) );
  OAI21_X1 U10066 ( .B1(n8635), .B2(n9747), .A(n8634), .ZN(n8643) );
  INV_X1 U10067 ( .A(n8650), .ZN(n8637) );
  NOR2_X1 U10068 ( .A1(n8637), .A2(n8636), .ZN(n8639) );
  OAI21_X1 U10069 ( .B1(n8639), .B2(n8638), .A(n8617), .ZN(n8641) );
  AOI21_X1 U10070 ( .B1(n8641), .B2(n9737), .A(n8640), .ZN(n8826) );
  NOR2_X1 U10071 ( .A1(n8826), .A2(n8656), .ZN(n8642) );
  AOI211_X1 U10072 ( .C1(n8823), .C2(n8672), .A(n8643), .B(n8642), .ZN(n8644)
         );
  OAI21_X1 U10073 ( .B1(n8827), .B2(n8727), .A(n8644), .ZN(P2_U3277) );
  XNOR2_X1 U10074 ( .A(n8645), .B(n4468), .ZN(n8832) );
  AOI21_X1 U10075 ( .B1(n8828), .B2(n8670), .A(n8646), .ZN(n8829) );
  AOI22_X1 U10076 ( .A1(n8754), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8647), .B2(
        n8752), .ZN(n8648) );
  OAI21_X1 U10077 ( .B1(n8649), .B2(n9747), .A(n8648), .ZN(n8658) );
  OAI211_X1 U10078 ( .C1(n4468), .C2(n8651), .A(n8650), .B(n9737), .ZN(n8655)
         );
  AOI22_X1 U10079 ( .A1(n8653), .A2(n8729), .B1(n8731), .B2(n8652), .ZN(n8654)
         );
  NOR2_X1 U10080 ( .A1(n8831), .A2(n8656), .ZN(n8657) );
  AOI211_X1 U10081 ( .C1(n8829), .C2(n9727), .A(n8658), .B(n8657), .ZN(n8659)
         );
  OAI21_X1 U10082 ( .B1(n8832), .B2(n8727), .A(n8659), .ZN(P2_U3278) );
  OAI21_X1 U10083 ( .B1(n8662), .B2(n8661), .A(n8660), .ZN(n8663) );
  INV_X1 U10084 ( .A(n8663), .ZN(n8837) );
  OAI211_X1 U10085 ( .C1(n8665), .C2(n4645), .A(n8664), .B(n9737), .ZN(n8668)
         );
  OR2_X1 U10086 ( .A1(n8666), .A2(n9734), .ZN(n8667) );
  OAI211_X1 U10087 ( .C1(n8669), .C2(n9732), .A(n8668), .B(n8667), .ZN(n8833)
         );
  INV_X1 U10088 ( .A(n8670), .ZN(n8671) );
  AOI211_X1 U10089 ( .C1(n8835), .C2(n8687), .A(n9820), .B(n8671), .ZN(n8834)
         );
  NAND2_X1 U10090 ( .A1(n8834), .A2(n8672), .ZN(n8675) );
  AOI22_X1 U10091 ( .A1(n8754), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8673), .B2(
        n8752), .ZN(n8674) );
  OAI211_X1 U10092 ( .C1(n4814), .C2(n9747), .A(n8675), .B(n8674), .ZN(n8676)
         );
  AOI21_X1 U10093 ( .B1(n8833), .B2(n9749), .A(n8676), .ZN(n8677) );
  OAI21_X1 U10094 ( .B1(n8837), .B2(n8727), .A(n8677), .ZN(P2_U3279) );
  XNOR2_X1 U10095 ( .A(n8679), .B(n8678), .ZN(n8686) );
  OAI22_X1 U10096 ( .A1(n8681), .A2(n9734), .B1(n8680), .B2(n9732), .ZN(n8685)
         );
  XNOR2_X1 U10097 ( .A(n8683), .B(n8682), .ZN(n8842) );
  NOR2_X1 U10098 ( .A1(n8842), .A2(n9740), .ZN(n8684) );
  AOI211_X1 U10099 ( .C1(n8686), .C2(n9737), .A(n8685), .B(n8684), .ZN(n8841)
         );
  INV_X1 U10100 ( .A(n8687), .ZN(n8688) );
  AOI21_X1 U10101 ( .B1(n8838), .B2(n8696), .A(n8688), .ZN(n8839) );
  AOI22_X1 U10102 ( .A1(n8754), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8689), .B2(
        n8752), .ZN(n8690) );
  OAI21_X1 U10103 ( .B1(n4684), .B2(n9747), .A(n8690), .ZN(n8692) );
  NOR2_X1 U10104 ( .A1(n8842), .A2(n9722), .ZN(n8691) );
  AOI211_X1 U10105 ( .C1(n8839), .C2(n9727), .A(n8692), .B(n8691), .ZN(n8693)
         );
  OAI21_X1 U10106 ( .B1(n8841), .B2(n8754), .A(n8693), .ZN(P2_U3280) );
  XNOR2_X1 U10107 ( .A(n8695), .B(n8694), .ZN(n8847) );
  INV_X1 U10108 ( .A(n8715), .ZN(n8698) );
  INV_X1 U10109 ( .A(n8696), .ZN(n8697) );
  AOI21_X1 U10110 ( .B1(n8843), .B2(n8698), .A(n8697), .ZN(n8844) );
  AOI22_X1 U10111 ( .A1(n8754), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8699), .B2(
        n8752), .ZN(n8700) );
  OAI21_X1 U10112 ( .B1(n8701), .B2(n9747), .A(n8700), .ZN(n8708) );
  XNOR2_X1 U10113 ( .A(n8703), .B(n8702), .ZN(n8706) );
  AOI222_X1 U10114 ( .A1(n9737), .A2(n8706), .B1(n8705), .B2(n8731), .C1(n8704), .C2(n8729), .ZN(n8846) );
  NOR2_X1 U10115 ( .A1(n8846), .A2(n9745), .ZN(n8707) );
  AOI211_X1 U10116 ( .C1(n8844), .C2(n9727), .A(n8708), .B(n8707), .ZN(n8709)
         );
  OAI21_X1 U10117 ( .B1(n8847), .B2(n8727), .A(n8709), .ZN(P2_U3281) );
  OAI21_X1 U10118 ( .B1(n8712), .B2(n8711), .A(n8710), .ZN(n8713) );
  INV_X1 U10119 ( .A(n8713), .ZN(n8852) );
  INV_X1 U10120 ( .A(n8714), .ZN(n8716) );
  AOI21_X1 U10121 ( .B1(n8848), .B2(n8716), .A(n8715), .ZN(n8849) );
  AOI22_X1 U10122 ( .A1(n8754), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8717), .B2(
        n8752), .ZN(n8718) );
  OAI21_X1 U10123 ( .B1(n8719), .B2(n9747), .A(n8718), .ZN(n8725) );
  XNOR2_X1 U10124 ( .A(n8721), .B(n8720), .ZN(n8723) );
  AOI21_X1 U10125 ( .B1(n8723), .B2(n9737), .A(n8722), .ZN(n8851) );
  NOR2_X1 U10126 ( .A1(n8851), .A2(n8754), .ZN(n8724) );
  AOI211_X1 U10127 ( .C1(n8849), .C2(n9727), .A(n8725), .B(n8724), .ZN(n8726)
         );
  OAI21_X1 U10128 ( .B1(n8852), .B2(n8727), .A(n8726), .ZN(P2_U3282) );
  XNOR2_X1 U10129 ( .A(n8728), .B(n8735), .ZN(n8733) );
  AOI222_X1 U10130 ( .A1(n9737), .A2(n8733), .B1(n8732), .B2(n8731), .C1(n8730), .C2(n8729), .ZN(n9780) );
  MUX2_X1 U10131 ( .A(n8042), .B(n9780), .S(n9749), .Z(n8742) );
  AOI22_X1 U10132 ( .A1(n8749), .A2(n9773), .B1(n8752), .B2(n8734), .ZN(n8741)
         );
  NAND2_X1 U10133 ( .A1(n8736), .A2(n8735), .ZN(n9776) );
  NAND3_X1 U10134 ( .A1(n9777), .A2(n9776), .A3(n8751), .ZN(n8740) );
  AOI21_X1 U10135 ( .B1(n9773), .B2(n8738), .A(n8737), .ZN(n9775) );
  NAND2_X1 U10136 ( .A1(n9775), .A2(n9727), .ZN(n8739) );
  NAND4_X1 U10137 ( .A1(n8742), .A2(n8741), .A3(n8740), .A4(n8739), .ZN(
        P2_U3290) );
  AOI22_X1 U10138 ( .A1(n8751), .A2(n8743), .B1(n8749), .B2(n4411), .ZN(n8748)
         );
  AOI22_X1 U10139 ( .A1(n8756), .A2(n8744), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n8752), .ZN(n8747) );
  MUX2_X1 U10140 ( .A(n8745), .B(n5194), .S(n9745), .Z(n8746) );
  NAND3_X1 U10141 ( .A1(n8748), .A2(n8747), .A3(n8746), .ZN(P2_U3294) );
  AOI22_X1 U10142 ( .A1(n8751), .A2(n8750), .B1(n8749), .B2(n6270), .ZN(n8759)
         );
  AOI22_X1 U10143 ( .A1(n9749), .A2(n8753), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8752), .ZN(n8758) );
  AOI22_X1 U10144 ( .A1(n8756), .A2(n8755), .B1(P2_REG2_REG_1__SCAN_IN), .B2(
        n8754), .ZN(n8757) );
  NAND3_X1 U10145 ( .A1(n8759), .A2(n8758), .A3(n8757), .ZN(P2_U3295) );
  AOI21_X1 U10146 ( .B1(n8761), .B2(n9815), .A(n8760), .ZN(n8762) );
  OAI21_X1 U10147 ( .B1(n8763), .B2(n9820), .A(n8762), .ZN(n8860) );
  MUX2_X1 U10148 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8860), .S(n9839), .Z(
        P2_U3551) );
  NAND3_X1 U10149 ( .A1(n8765), .A2(n9774), .A3(n8764), .ZN(n8767) );
  OAI211_X1 U10150 ( .C1(n8768), .C2(n9810), .A(n8767), .B(n8766), .ZN(n8861)
         );
  MUX2_X1 U10151 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8861), .S(n9839), .Z(
        P2_U3550) );
  NAND2_X1 U10152 ( .A1(n8769), .A2(n9822), .ZN(n8775) );
  OAI22_X1 U10153 ( .A1(n8771), .A2(n9820), .B1(n8770), .B2(n9810), .ZN(n8772)
         );
  NOR2_X1 U10154 ( .A1(n8773), .A2(n8772), .ZN(n8774) );
  NAND2_X1 U10155 ( .A1(n8775), .A2(n8774), .ZN(n8862) );
  MUX2_X1 U10156 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8862), .S(n9839), .Z(
        P2_U3549) );
  AOI22_X1 U10157 ( .A1(n8777), .A2(n9774), .B1(n9815), .B2(n8776), .ZN(n8778)
         );
  OAI211_X1 U10158 ( .C1(n8780), .C2(n9764), .A(n8779), .B(n8778), .ZN(n8863)
         );
  MUX2_X1 U10159 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8863), .S(n9839), .Z(
        P2_U3548) );
  AOI22_X1 U10160 ( .A1(n8782), .A2(n9774), .B1(n9815), .B2(n8781), .ZN(n8783)
         );
  OAI211_X1 U10161 ( .C1(n8785), .C2(n9764), .A(n8784), .B(n8783), .ZN(n8864)
         );
  MUX2_X1 U10162 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8864), .S(n9839), .Z(
        P2_U3547) );
  AOI21_X1 U10163 ( .B1(n9815), .B2(n8787), .A(n8786), .ZN(n8788) );
  OAI211_X1 U10164 ( .C1(n8790), .C2(n9764), .A(n8789), .B(n8788), .ZN(n8865)
         );
  MUX2_X1 U10165 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8865), .S(n9839), .Z(
        P2_U3546) );
  AOI21_X1 U10166 ( .B1(n9815), .B2(n8792), .A(n8791), .ZN(n8793) );
  OAI211_X1 U10167 ( .C1(n8795), .C2(n9764), .A(n8794), .B(n8793), .ZN(n8866)
         );
  MUX2_X1 U10168 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8866), .S(n9839), .Z(
        P2_U3545) );
  AOI22_X1 U10169 ( .A1(n8797), .A2(n9774), .B1(n9815), .B2(n8796), .ZN(n8798)
         );
  OAI211_X1 U10170 ( .C1(n8800), .C2(n9764), .A(n8799), .B(n8798), .ZN(n8867)
         );
  MUX2_X1 U10171 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8867), .S(n9839), .Z(
        P2_U3544) );
  NAND3_X1 U10172 ( .A1(n8802), .A2(n8801), .A3(n9822), .ZN(n8807) );
  AOI22_X1 U10173 ( .A1(n8804), .A2(n9774), .B1(n9815), .B2(n8803), .ZN(n8805)
         );
  NAND3_X1 U10174 ( .A1(n8807), .A2(n8806), .A3(n8805), .ZN(n8868) );
  MUX2_X1 U10175 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8868), .S(n9839), .Z(
        P2_U3543) );
  AOI22_X1 U10176 ( .A1(n8809), .A2(n9774), .B1(n9815), .B2(n8808), .ZN(n8810)
         );
  OAI211_X1 U10177 ( .C1(n8812), .C2(n9764), .A(n8811), .B(n8810), .ZN(n8869)
         );
  MUX2_X1 U10178 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8869), .S(n9839), .Z(
        P2_U3542) );
  AOI22_X1 U10179 ( .A1(n8814), .A2(n9774), .B1(n9815), .B2(n8813), .ZN(n8815)
         );
  OAI211_X1 U10180 ( .C1(n8817), .C2(n9764), .A(n8816), .B(n8815), .ZN(n8870)
         );
  MUX2_X1 U10181 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8870), .S(n9839), .Z(
        P2_U3541) );
  AOI22_X1 U10182 ( .A1(n8819), .A2(n9774), .B1(n9815), .B2(n8818), .ZN(n8820)
         );
  OAI211_X1 U10183 ( .C1(n8822), .C2(n9764), .A(n8821), .B(n8820), .ZN(n8871)
         );
  MUX2_X1 U10184 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8871), .S(n9839), .Z(
        P2_U3540) );
  AOI21_X1 U10185 ( .B1(n9815), .B2(n8824), .A(n8823), .ZN(n8825) );
  OAI211_X1 U10186 ( .C1(n8827), .C2(n9764), .A(n8826), .B(n8825), .ZN(n8872)
         );
  MUX2_X1 U10187 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8872), .S(n9839), .Z(
        P2_U3539) );
  AOI22_X1 U10188 ( .A1(n8829), .A2(n9774), .B1(n9815), .B2(n8828), .ZN(n8830)
         );
  OAI211_X1 U10189 ( .C1(n8832), .C2(n9764), .A(n8831), .B(n8830), .ZN(n8873)
         );
  MUX2_X1 U10190 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8873), .S(n9839), .Z(
        P2_U3538) );
  AOI211_X1 U10191 ( .C1(n9815), .C2(n8835), .A(n8834), .B(n8833), .ZN(n8836)
         );
  OAI21_X1 U10192 ( .B1(n8837), .B2(n9764), .A(n8836), .ZN(n8874) );
  MUX2_X1 U10193 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8874), .S(n9839), .Z(
        P2_U3537) );
  AOI22_X1 U10194 ( .A1(n8839), .A2(n9774), .B1(n9815), .B2(n8838), .ZN(n8840)
         );
  OAI211_X1 U10195 ( .C1(n8842), .C2(n9787), .A(n8841), .B(n8840), .ZN(n8875)
         );
  MUX2_X1 U10196 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8875), .S(n9839), .Z(
        P2_U3536) );
  AOI22_X1 U10197 ( .A1(n8844), .A2(n9774), .B1(n9815), .B2(n8843), .ZN(n8845)
         );
  OAI211_X1 U10198 ( .C1(n8847), .C2(n9764), .A(n8846), .B(n8845), .ZN(n8876)
         );
  MUX2_X1 U10199 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8876), .S(n9839), .Z(
        P2_U3535) );
  AOI22_X1 U10200 ( .A1(n8849), .A2(n9774), .B1(n9815), .B2(n8848), .ZN(n8850)
         );
  OAI211_X1 U10201 ( .C1(n8852), .C2(n9764), .A(n8851), .B(n8850), .ZN(n8877)
         );
  MUX2_X1 U10202 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8877), .S(n9839), .Z(
        P2_U3534) );
  NAND3_X1 U10203 ( .A1(n8854), .A2(n9822), .A3(n8853), .ZN(n8859) );
  AOI22_X1 U10204 ( .A1(n8856), .A2(n9774), .B1(n9815), .B2(n8855), .ZN(n8857)
         );
  NAND3_X1 U10205 ( .A1(n8859), .A2(n8858), .A3(n8857), .ZN(n8878) );
  MUX2_X1 U10206 ( .A(n8878), .B(P2_REG1_REG_13__SCAN_IN), .S(n9837), .Z(
        P2_U3533) );
  MUX2_X1 U10207 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8860), .S(n9826), .Z(
        P2_U3519) );
  MUX2_X1 U10208 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8861), .S(n9826), .Z(
        P2_U3518) );
  MUX2_X1 U10209 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8862), .S(n9826), .Z(
        P2_U3517) );
  MUX2_X1 U10210 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8863), .S(n9826), .Z(
        P2_U3516) );
  MUX2_X1 U10211 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8864), .S(n9826), .Z(
        P2_U3515) );
  MUX2_X1 U10212 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8865), .S(n9826), .Z(
        P2_U3514) );
  MUX2_X1 U10213 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8866), .S(n9826), .Z(
        P2_U3513) );
  MUX2_X1 U10214 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8867), .S(n9826), .Z(
        P2_U3512) );
  MUX2_X1 U10215 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8868), .S(n9826), .Z(
        P2_U3511) );
  MUX2_X1 U10216 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8869), .S(n9826), .Z(
        P2_U3510) );
  MUX2_X1 U10217 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8870), .S(n9826), .Z(
        P2_U3509) );
  MUX2_X1 U10218 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8871), .S(n9826), .Z(
        P2_U3508) );
  MUX2_X1 U10219 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8872), .S(n9826), .Z(
        P2_U3507) );
  MUX2_X1 U10220 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8873), .S(n9826), .Z(
        P2_U3505) );
  MUX2_X1 U10221 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8874), .S(n9826), .Z(
        P2_U3502) );
  MUX2_X1 U10222 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8875), .S(n9826), .Z(
        P2_U3499) );
  MUX2_X1 U10223 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8876), .S(n9826), .Z(
        P2_U3496) );
  MUX2_X1 U10224 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8877), .S(n9826), .Z(
        P2_U3493) );
  MUX2_X1 U10225 ( .A(n8878), .B(P2_REG0_REG_13__SCAN_IN), .S(n9824), .Z(
        P2_U3490) );
  INV_X1 U10226 ( .A(n8879), .ZN(n9418) );
  NAND3_X1 U10227 ( .A1(n8880), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8882) );
  OAI22_X1 U10228 ( .A1(n8883), .A2(n8882), .B1(n5948), .B2(n8881), .ZN(n8884)
         );
  INV_X1 U10229 ( .A(n8884), .ZN(n8885) );
  OAI21_X1 U10230 ( .B1(n9418), .B2(n8236), .A(n8885), .ZN(P2_U3327) );
  MUX2_X1 U10231 ( .A(n8886), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  OAI21_X1 U10232 ( .B1(n8889), .B2(n8888), .A(n8887), .ZN(n8890) );
  NAND2_X1 U10233 ( .A1(n8890), .A2(n9015), .ZN(n8896) );
  AOI22_X1 U10234 ( .A1(n8978), .A2(n9050), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3084), .ZN(n8895) );
  AOI22_X1 U10235 ( .A1(n9030), .A2(n9048), .B1(n8891), .B2(n9029), .ZN(n8894)
         );
  NAND2_X1 U10236 ( .A1(n9036), .A2(n8892), .ZN(n8893) );
  NAND4_X1 U10237 ( .A1(n8896), .A2(n8895), .A3(n8894), .A4(n8893), .ZN(
        P1_U3211) );
  XNOR2_X1 U10238 ( .A(n8898), .B(n8897), .ZN(n8899) );
  XNOR2_X1 U10239 ( .A(n8900), .B(n8899), .ZN(n8905) );
  AOI22_X1 U10240 ( .A1(n9130), .A2(n8978), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8902) );
  NAND2_X1 U10241 ( .A1(n9101), .A2(n9029), .ZN(n8901) );
  OAI211_X1 U10242 ( .C1(n9097), .C2(n9009), .A(n8902), .B(n8901), .ZN(n8903)
         );
  AOI21_X1 U10243 ( .B1(n9328), .B2(n9036), .A(n8903), .ZN(n8904) );
  OAI21_X1 U10244 ( .B1(n8905), .B2(n9038), .A(n8904), .ZN(P1_U3212) );
  NAND2_X1 U10245 ( .A1(n8907), .A2(n8906), .ZN(n8908) );
  XOR2_X1 U10246 ( .A(n8909), .B(n8908), .Z(n8917) );
  NOR2_X1 U10247 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8910), .ZN(n9614) );
  INV_X1 U10248 ( .A(n8911), .ZN(n8912) );
  OAI22_X1 U10249 ( .A1(n9010), .A2(n8912), .B1(n9009), .B2(n9272), .ZN(n8913)
         );
  AOI211_X1 U10250 ( .C1(n8978), .C2(n9043), .A(n9614), .B(n8913), .ZN(n8916)
         );
  NAND2_X1 U10251 ( .A1(n8914), .A2(n9036), .ZN(n8915) );
  OAI211_X1 U10252 ( .C1(n8917), .C2(n9038), .A(n8916), .B(n8915), .ZN(
        P1_U3213) );
  NAND2_X1 U10253 ( .A1(n4477), .A2(n8918), .ZN(n8920) );
  XNOR2_X1 U10254 ( .A(n8920), .B(n8919), .ZN(n8925) );
  OAI22_X1 U10255 ( .A1(n8956), .A2(n9009), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8921), .ZN(n8923) );
  OAI22_X1 U10256 ( .A1(n9191), .A2(n9034), .B1(n9010), .B2(n9152), .ZN(n8922)
         );
  AOI211_X1 U10257 ( .C1(n9349), .C2(n9036), .A(n8923), .B(n8922), .ZN(n8924)
         );
  OAI21_X1 U10258 ( .B1(n8925), .B2(n9038), .A(n8924), .ZN(P1_U3214) );
  OAI21_X1 U10259 ( .B1(n8928), .B2(n8927), .A(n8926), .ZN(n8929) );
  NAND2_X1 U10260 ( .A1(n8929), .A2(n9015), .ZN(n8934) );
  AOI22_X1 U10261 ( .A1(n8978), .A2(n9054), .B1(n9030), .B2(n9052), .ZN(n8933)
         );
  AOI22_X1 U10262 ( .A1(n9036), .A2(n8930), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3084), .ZN(n8932) );
  NAND2_X1 U10263 ( .A1(n9029), .A2(n5810), .ZN(n8931) );
  NAND4_X1 U10264 ( .A1(n8934), .A2(n8933), .A3(n8932), .A4(n8931), .ZN(
        P1_U3216) );
  XNOR2_X1 U10265 ( .A(n8937), .B(n8936), .ZN(n8938) );
  XNOR2_X1 U10266 ( .A(n8935), .B(n8938), .ZN(n8943) );
  OAI21_X1 U10267 ( .B1(n9192), .B2(n9009), .A(n8939), .ZN(n8941) );
  OAI22_X1 U10268 ( .A1(n9034), .A2(n9254), .B1(n9010), .B2(n9220), .ZN(n8940)
         );
  AOI211_X1 U10269 ( .C1(n9372), .C2(n9036), .A(n8941), .B(n8940), .ZN(n8942)
         );
  OAI21_X1 U10270 ( .B1(n8943), .B2(n9038), .A(n8942), .ZN(P1_U3217) );
  OAI21_X1 U10271 ( .B1(n8946), .B2(n8945), .A(n8944), .ZN(n8951) );
  AOI22_X1 U10272 ( .A1(n9162), .A2(n9030), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8948) );
  AOI22_X1 U10273 ( .A1(n8978), .A2(n9228), .B1(n9185), .B2(n9029), .ZN(n8947)
         );
  OAI211_X1 U10274 ( .C1(n8949), .C2(n9024), .A(n8948), .B(n8947), .ZN(n8950)
         );
  AOI21_X1 U10275 ( .B1(n8951), .B2(n9015), .A(n8950), .ZN(n8952) );
  INV_X1 U10276 ( .A(n8952), .ZN(P1_U3221) );
  XOR2_X1 U10277 ( .A(n8954), .B(n8953), .Z(n8961) );
  OAI22_X1 U10278 ( .A1(n8956), .A2(n9034), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8955), .ZN(n8957) );
  AOI21_X1 U10279 ( .B1(n9125), .B2(n9029), .A(n8957), .ZN(n8958) );
  OAI21_X1 U10280 ( .B1(n9096), .B2(n9009), .A(n8958), .ZN(n8959) );
  AOI21_X1 U10281 ( .B1(n9337), .B2(n9036), .A(n8959), .ZN(n8960) );
  OAI21_X1 U10282 ( .B1(n8961), .B2(n9038), .A(n8960), .ZN(P1_U3223) );
  OAI21_X1 U10283 ( .B1(n8963), .B2(n4491), .A(n8962), .ZN(n8964) );
  NAND2_X1 U10284 ( .A1(n8964), .A2(n9015), .ZN(n8969) );
  NOR2_X1 U10285 ( .A1(n9009), .A2(n9271), .ZN(n8967) );
  INV_X1 U10286 ( .A(n9276), .ZN(n8965) );
  OAI22_X1 U10287 ( .A1(n9034), .A2(n9272), .B1(n9010), .B2(n8965), .ZN(n8966)
         );
  AOI211_X1 U10288 ( .C1(P1_REG3_REG_16__SCAN_IN), .C2(P1_U3084), .A(n8967), 
        .B(n8966), .ZN(n8968) );
  OAI211_X1 U10289 ( .C1(n9279), .C2(n9024), .A(n8969), .B(n8968), .ZN(
        P1_U3224) );
  XOR2_X1 U10290 ( .A(n8971), .B(n8970), .Z(n8976) );
  OAI22_X1 U10291 ( .A1(n9009), .A2(n9254), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8972), .ZN(n8974) );
  OAI22_X1 U10292 ( .A1(n9034), .A2(n9253), .B1(n9010), .B2(n9259), .ZN(n8973)
         );
  AOI211_X1 U10293 ( .C1(n9383), .C2(n9036), .A(n8974), .B(n8973), .ZN(n8975)
         );
  OAI21_X1 U10294 ( .B1(n8976), .B2(n9038), .A(n8975), .ZN(P1_U3226) );
  XOR2_X1 U10295 ( .A(n8977), .B(n4446), .Z(n8983) );
  NAND2_X1 U10296 ( .A1(n9118), .A2(n9030), .ZN(n8980) );
  AOI22_X1 U10297 ( .A1(n9176), .A2(n8978), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8979) );
  OAI211_X1 U10298 ( .C1(n9010), .C2(n9137), .A(n8980), .B(n8979), .ZN(n8981)
         );
  AOI21_X1 U10299 ( .B1(n9345), .B2(n9036), .A(n8981), .ZN(n8982) );
  OAI21_X1 U10300 ( .B1(n8983), .B2(n9038), .A(n8982), .ZN(P1_U3227) );
  INV_X1 U10301 ( .A(n8984), .ZN(n8988) );
  NAND2_X1 U10302 ( .A1(n4496), .A2(n8987), .ZN(n8985) );
  AOI22_X1 U10303 ( .A1(n8988), .A2(n8987), .B1(n8986), .B2(n8985), .ZN(n8993)
         );
  OAI22_X1 U10304 ( .A1(n9207), .A2(n9009), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8989), .ZN(n8991) );
  OAI22_X1 U10305 ( .A1(n9034), .A2(n9206), .B1(n9010), .B2(n9209), .ZN(n8990)
         );
  AOI211_X1 U10306 ( .C1(n9368), .C2(n9036), .A(n8991), .B(n8990), .ZN(n8992)
         );
  OAI21_X1 U10307 ( .B1(n8993), .B2(n9038), .A(n8992), .ZN(P1_U3231) );
  INV_X1 U10308 ( .A(n8994), .ZN(n8996) );
  INV_X1 U10309 ( .A(n8997), .ZN(n8995) );
  OAI21_X1 U10310 ( .B1(n8998), .B2(n8996), .A(n8995), .ZN(n8999) );
  AOI22_X1 U10311 ( .A1(n8999), .A2(n4919), .B1(n8998), .B2(n8997), .ZN(n9004)
         );
  OAI22_X1 U10312 ( .A1(n9142), .A2(n9009), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9000), .ZN(n9002) );
  OAI22_X1 U10313 ( .A1(n9207), .A2(n9034), .B1(n9010), .B2(n9170), .ZN(n9001)
         );
  AOI211_X1 U10314 ( .C1(n9354), .C2(n9036), .A(n9002), .B(n9001), .ZN(n9003)
         );
  OAI21_X1 U10315 ( .B1(n9004), .B2(n9038), .A(n9003), .ZN(P1_U3233) );
  XNOR2_X1 U10316 ( .A(n9006), .B(n9005), .ZN(n9007) );
  XNOR2_X1 U10317 ( .A(n9008), .B(n9007), .ZN(n9014) );
  NAND2_X1 U10318 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9628) );
  OAI21_X1 U10319 ( .B1(n9206), .B2(n9009), .A(n9628), .ZN(n9012) );
  OAI22_X1 U10320 ( .A1(n9034), .A2(n9271), .B1(n9010), .B2(n9245), .ZN(n9011)
         );
  AOI211_X1 U10321 ( .C1(n9377), .C2(n9036), .A(n9012), .B(n9011), .ZN(n9013)
         );
  OAI21_X1 U10322 ( .B1(n9014), .B2(n9038), .A(n9013), .ZN(P1_U3236) );
  OAI211_X1 U10323 ( .C1(n9018), .C2(n9017), .A(n9016), .B(n9015), .ZN(n9023)
         );
  INV_X1 U10324 ( .A(n9019), .ZN(n9110) );
  AOI22_X1 U10325 ( .A1(n9110), .A2(n9029), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9020) );
  OAI21_X1 U10326 ( .B1(n9141), .B2(n9034), .A(n9020), .ZN(n9021) );
  AOI21_X1 U10327 ( .B1(n9030), .B2(n9117), .A(n9021), .ZN(n9022) );
  OAI211_X1 U10328 ( .C1(n9112), .C2(n9024), .A(n9023), .B(n9022), .ZN(
        P1_U3238) );
  NAND2_X1 U10329 ( .A1(n9026), .A2(n9025), .ZN(n9027) );
  XOR2_X1 U10330 ( .A(n9028), .B(n9027), .Z(n9039) );
  AOI22_X1 U10331 ( .A1(n9030), .A2(n9294), .B1(n9286), .B2(n9029), .ZN(n9032)
         );
  OAI211_X1 U10332 ( .C1(n9034), .C2(n9033), .A(n9032), .B(n9031), .ZN(n9035)
         );
  AOI21_X1 U10333 ( .B1(n9391), .B2(n9036), .A(n9035), .ZN(n9037) );
  OAI21_X1 U10334 ( .B1(n9039), .B2(n9038), .A(n9037), .ZN(P1_U3239) );
  MUX2_X1 U10335 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9040), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10336 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9089), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10337 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9041), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10338 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9117), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10339 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9130), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10340 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9118), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10341 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9161), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10342 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9176), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10343 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9162), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10344 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9177), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10345 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9228), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10346 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9240), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10347 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9227), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10348 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9239), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10349 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9294), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10350 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9042), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10351 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9292), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10352 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9043), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10353 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9044), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10354 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9045), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10355 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9046), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10356 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9047), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10357 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9048), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10358 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9049), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10359 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9050), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10360 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9051), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10361 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9052), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10362 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9053), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10363 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9054), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10364 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9055), .S(P1_U4006), .Z(
        P1_U3556) );
  AOI211_X1 U10365 ( .C1(n9058), .C2(n9057), .A(n9056), .B(n9629), .ZN(n9071)
         );
  INV_X1 U10366 ( .A(n9059), .ZN(n9068) );
  AOI211_X1 U10367 ( .C1(n9063), .C2(n9062), .A(n9061), .B(n9060), .ZN(n9064)
         );
  INV_X1 U10368 ( .A(n9064), .ZN(n9067) );
  NAND2_X1 U10369 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9066) );
  OAI211_X1 U10370 ( .C1(n9069), .C2(n9068), .A(n9067), .B(n9066), .ZN(n9070)
         );
  AOI211_X1 U10371 ( .C1(P1_ADDR_REG_17__SCAN_IN), .C2(n9640), .A(n9071), .B(
        n9070), .ZN(n9072) );
  INV_X1 U10372 ( .A(n9072), .ZN(P1_U3258) );
  INV_X1 U10373 ( .A(n9073), .ZN(n9074) );
  NAND2_X1 U10374 ( .A1(n9075), .A2(n9074), .ZN(n9312) );
  NAND3_X1 U10375 ( .A1(n9313), .A2(n9650), .A3(n9312), .ZN(n9078) );
  AOI21_X1 U10376 ( .B1(n4419), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9076), .ZN(
        n9077) );
  OAI211_X1 U10377 ( .C1(n9316), .C2(n9656), .A(n9078), .B(n9077), .ZN(
        P1_U3262) );
  INV_X1 U10378 ( .A(n9100), .ZN(n9082) );
  INV_X1 U10379 ( .A(n9080), .ZN(n9081) );
  AOI21_X1 U10380 ( .B1(n9322), .B2(n9082), .A(n9081), .ZN(n9323) );
  AOI22_X1 U10381 ( .A1(n9083), .A2(n9652), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n4419), .ZN(n9084) );
  OAI21_X1 U10382 ( .B1(n9085), .B2(n9656), .A(n9084), .ZN(n9091) );
  OAI21_X1 U10383 ( .B1(n9088), .B2(n9087), .A(n9086), .ZN(n9090) );
  XNOR2_X1 U10384 ( .A(n9092), .B(n9095), .ZN(n9331) );
  AOI22_X1 U10385 ( .A1(n9328), .A2(n9469), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n4419), .ZN(n9105) );
  AOI211_X1 U10386 ( .C1(n9095), .C2(n9094), .A(n9459), .B(n9093), .ZN(n9099)
         );
  OAI22_X1 U10387 ( .A1(n9097), .A2(n9462), .B1(n9096), .B2(n9464), .ZN(n9098)
         );
  NOR2_X1 U10388 ( .A1(n9099), .A2(n9098), .ZN(n9330) );
  AOI211_X1 U10389 ( .C1(n9328), .C2(n9107), .A(n9692), .B(n9100), .ZN(n9327)
         );
  AOI22_X1 U10390 ( .A1(n9327), .A2(n9243), .B1(n9652), .B2(n9101), .ZN(n9102)
         );
  AOI21_X1 U10391 ( .B1(n9330), .B2(n9102), .A(n4419), .ZN(n9103) );
  INV_X1 U10392 ( .A(n9103), .ZN(n9104) );
  OAI211_X1 U10393 ( .C1(n9331), .C2(n9308), .A(n9105), .B(n9104), .ZN(
        P1_U3264) );
  XNOR2_X1 U10394 ( .A(n9106), .B(n9115), .ZN(n9336) );
  INV_X1 U10395 ( .A(n9124), .ZN(n9109) );
  INV_X1 U10396 ( .A(n9107), .ZN(n9108) );
  AOI21_X1 U10397 ( .B1(n9332), .B2(n9109), .A(n9108), .ZN(n9333) );
  AOI22_X1 U10398 ( .A1(n9110), .A2(n9652), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n4419), .ZN(n9111) );
  OAI21_X1 U10399 ( .B1(n9112), .B2(n9656), .A(n9111), .ZN(n9120) );
  INV_X1 U10400 ( .A(n9113), .ZN(n9114) );
  NOR2_X1 U10401 ( .A1(n4483), .A2(n9114), .ZN(n9116) );
  XNOR2_X1 U10402 ( .A(n9116), .B(n9115), .ZN(n9119) );
  OAI21_X1 U10403 ( .B1(n9122), .B2(n9129), .A(n9121), .ZN(n9123) );
  INV_X1 U10404 ( .A(n9123), .ZN(n9341) );
  AOI21_X1 U10405 ( .B1(n9337), .B2(n9135), .A(n9124), .ZN(n9338) );
  INV_X1 U10406 ( .A(n9337), .ZN(n9127) );
  AOI22_X1 U10407 ( .A1(n9125), .A2(n9652), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n4419), .ZN(n9126) );
  OAI21_X1 U10408 ( .B1(n9127), .B2(n9656), .A(n9126), .ZN(n9133) );
  XOR2_X1 U10409 ( .A(n9129), .B(n9128), .Z(n9131) );
  AOI222_X1 U10410 ( .A1(n9296), .A2(n9131), .B1(n9130), .B2(n9293), .C1(n9161), .C2(n9291), .ZN(n9340) );
  NOR2_X1 U10411 ( .A1(n9340), .A2(n4419), .ZN(n9132) );
  AOI211_X1 U10412 ( .C1(n9338), .C2(n9650), .A(n9133), .B(n9132), .ZN(n9134)
         );
  OAI21_X1 U10413 ( .B1(n9341), .B2(n9308), .A(n9134), .ZN(P1_U3266) );
  INV_X1 U10414 ( .A(n9135), .ZN(n9136) );
  AOI211_X1 U10415 ( .C1(n9345), .C2(n4736), .A(n9692), .B(n9136), .ZN(n9344)
         );
  NOR2_X1 U10416 ( .A1(n9137), .A2(n9258), .ZN(n9143) );
  NAND2_X1 U10417 ( .A1(n9158), .A2(n9138), .ZN(n9139) );
  XOR2_X1 U10418 ( .A(n9144), .B(n9139), .Z(n9140) );
  OAI222_X1 U10419 ( .A1(n9464), .A2(n9142), .B1(n9462), .B2(n9141), .C1(n9140), .C2(n9459), .ZN(n9343) );
  AOI211_X1 U10420 ( .C1(n9344), .C2(n9243), .A(n9143), .B(n9343), .ZN(n9149)
         );
  INV_X1 U10421 ( .A(n9348), .ZN(n9146) );
  NAND2_X1 U10422 ( .A1(n9145), .A2(n9144), .ZN(n9342) );
  NAND3_X1 U10423 ( .A1(n9146), .A2(n9196), .A3(n9342), .ZN(n9148) );
  AOI22_X1 U10424 ( .A1(n9345), .A2(n9469), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n4419), .ZN(n9147) );
  OAI211_X1 U10425 ( .C1(n4419), .C2(n9149), .A(n9148), .B(n9147), .ZN(
        P1_U3267) );
  XNOR2_X1 U10426 ( .A(n9150), .B(n9155), .ZN(n9353) );
  AOI21_X1 U10427 ( .B1(n9349), .B2(n9168), .A(n9151), .ZN(n9350) );
  INV_X1 U10428 ( .A(n9152), .ZN(n9153) );
  AOI22_X1 U10429 ( .A1(n9153), .A2(n9652), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n4419), .ZN(n9154) );
  OAI21_X1 U10430 ( .B1(n4734), .B2(n9656), .A(n9154), .ZN(n9165) );
  INV_X1 U10431 ( .A(n9155), .ZN(n9157) );
  NAND2_X1 U10432 ( .A1(n9157), .A2(n9156), .ZN(n9159) );
  OAI21_X1 U10433 ( .B1(n9160), .B2(n9159), .A(n9158), .ZN(n9163) );
  AOI222_X1 U10434 ( .A1(n9296), .A2(n9163), .B1(n9162), .B2(n9291), .C1(n9161), .C2(n9293), .ZN(n9352) );
  NOR2_X1 U10435 ( .A1(n9352), .A2(n4419), .ZN(n9164) );
  AOI211_X1 U10436 ( .C1(n9350), .C2(n9650), .A(n9165), .B(n9164), .ZN(n9166)
         );
  OAI21_X1 U10437 ( .B1(n9353), .B2(n9308), .A(n9166), .ZN(P1_U3268) );
  XOR2_X1 U10438 ( .A(n9174), .B(n9167), .Z(n9358) );
  INV_X1 U10439 ( .A(n9168), .ZN(n9169) );
  AOI21_X1 U10440 ( .B1(n9354), .B2(n9182), .A(n9169), .ZN(n9355) );
  INV_X1 U10441 ( .A(n9170), .ZN(n9171) );
  AOI22_X1 U10442 ( .A1(n9171), .A2(n9652), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n4419), .ZN(n9172) );
  OAI21_X1 U10443 ( .B1(n9173), .B2(n9656), .A(n9172), .ZN(n9180) );
  XNOR2_X1 U10444 ( .A(n9175), .B(n9174), .ZN(n9178) );
  AOI222_X1 U10445 ( .A1(n9296), .A2(n9178), .B1(n9177), .B2(n9291), .C1(n9176), .C2(n9293), .ZN(n9357) );
  NOR2_X1 U10446 ( .A1(n9357), .A2(n4419), .ZN(n9179) );
  AOI211_X1 U10447 ( .C1(n9355), .C2(n9650), .A(n9180), .B(n9179), .ZN(n9181)
         );
  OAI21_X1 U10448 ( .B1(n9308), .B2(n9358), .A(n9181), .ZN(P1_U3269) );
  INV_X1 U10449 ( .A(n9182), .ZN(n9183) );
  AOI211_X1 U10450 ( .C1(n9362), .C2(n9184), .A(n9692), .B(n9183), .ZN(n9361)
         );
  INV_X1 U10451 ( .A(n9185), .ZN(n9186) );
  NOR2_X1 U10452 ( .A1(n9186), .A2(n9258), .ZN(n9193) );
  AOI21_X1 U10453 ( .B1(n9189), .B2(n9188), .A(n9187), .ZN(n9190) );
  OAI222_X1 U10454 ( .A1(n9464), .A2(n9192), .B1(n9462), .B2(n9191), .C1(n9459), .C2(n9190), .ZN(n9360) );
  AOI211_X1 U10455 ( .C1(n9361), .C2(n9243), .A(n9193), .B(n9360), .ZN(n9200)
         );
  AOI22_X1 U10456 ( .A1(n9362), .A2(n9469), .B1(n4419), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9199) );
  INV_X1 U10457 ( .A(n9365), .ZN(n9197) );
  NAND2_X1 U10458 ( .A1(n9195), .A2(n9194), .ZN(n9359) );
  NAND3_X1 U10459 ( .A1(n9197), .A2(n9196), .A3(n9359), .ZN(n9198) );
  OAI211_X1 U10460 ( .C1(n9200), .C2(n4419), .A(n9199), .B(n9198), .ZN(
        P1_U3270) );
  XOR2_X1 U10461 ( .A(n9204), .B(n9201), .Z(n9370) );
  NAND2_X1 U10462 ( .A1(n9224), .A2(n9202), .ZN(n9203) );
  XOR2_X1 U10463 ( .A(n9204), .B(n9203), .Z(n9205) );
  OAI222_X1 U10464 ( .A1(n9462), .A2(n9207), .B1(n9464), .B2(n9206), .C1(n9205), .C2(n9459), .ZN(n9366) );
  INV_X1 U10465 ( .A(n9368), .ZN(n9213) );
  AOI211_X1 U10466 ( .C1(n9368), .C2(n9218), .A(n9692), .B(n9208), .ZN(n9367)
         );
  NAND2_X1 U10467 ( .A1(n9367), .A2(n9475), .ZN(n9212) );
  INV_X1 U10468 ( .A(n9209), .ZN(n9210) );
  AOI22_X1 U10469 ( .A1(n9210), .A2(n9652), .B1(n4419), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9211) );
  OAI211_X1 U10470 ( .C1(n9213), .C2(n9656), .A(n9212), .B(n9211), .ZN(n9214)
         );
  AOI21_X1 U10471 ( .B1(n9366), .B2(n9281), .A(n9214), .ZN(n9215) );
  OAI21_X1 U10472 ( .B1(n9370), .B2(n9308), .A(n9215), .ZN(P1_U3271) );
  NAND2_X1 U10473 ( .A1(n9234), .A2(n9216), .ZN(n9217) );
  XOR2_X1 U10474 ( .A(n9226), .B(n9217), .Z(n9375) );
  INV_X1 U10475 ( .A(n9218), .ZN(n9219) );
  AOI211_X1 U10476 ( .C1(n9372), .C2(n4742), .A(n9692), .B(n9219), .ZN(n9371)
         );
  INV_X1 U10477 ( .A(n9220), .ZN(n9221) );
  AOI22_X1 U10478 ( .A1(n4419), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9221), .B2(
        n9652), .ZN(n9222) );
  OAI21_X1 U10479 ( .B1(n9223), .B2(n9656), .A(n9222), .ZN(n9231) );
  OAI21_X1 U10480 ( .B1(n9226), .B2(n9225), .A(n9224), .ZN(n9229) );
  AOI222_X1 U10481 ( .A1(n9296), .A2(n9229), .B1(n9228), .B2(n9293), .C1(n9227), .C2(n9291), .ZN(n9374) );
  NOR2_X1 U10482 ( .A1(n9374), .A2(n4419), .ZN(n9230) );
  AOI211_X1 U10483 ( .C1(n9371), .C2(n9475), .A(n9231), .B(n9230), .ZN(n9232)
         );
  OAI21_X1 U10484 ( .B1(n9308), .B2(n9375), .A(n9232), .ZN(P1_U3272) );
  INV_X1 U10485 ( .A(n9233), .ZN(n9236) );
  INV_X1 U10486 ( .A(n9238), .ZN(n9235) );
  OAI21_X1 U10487 ( .B1(n9236), .B2(n9235), .A(n9234), .ZN(n9380) );
  OAI21_X1 U10488 ( .B1(n9238), .B2(n4500), .A(n9237), .ZN(n9241) );
  AOI222_X1 U10489 ( .A1(n9296), .A2(n9241), .B1(n9240), .B2(n9293), .C1(n9239), .C2(n9291), .ZN(n9379) );
  AOI211_X1 U10490 ( .C1(n9377), .C2(n9255), .A(n9692), .B(n9242), .ZN(n9376)
         );
  NAND2_X1 U10491 ( .A1(n9376), .A2(n9243), .ZN(n9244) );
  OAI211_X1 U10492 ( .C1(n9258), .C2(n9245), .A(n9379), .B(n9244), .ZN(n9246)
         );
  NAND2_X1 U10493 ( .A1(n9246), .A2(n9281), .ZN(n9248) );
  AOI22_X1 U10494 ( .A1(n9377), .A2(n9469), .B1(n4419), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n9247) );
  OAI211_X1 U10495 ( .C1(n9380), .C2(n9308), .A(n9248), .B(n9247), .ZN(
        P1_U3273) );
  XNOR2_X1 U10496 ( .A(n9249), .B(n9251), .ZN(n9385) );
  XOR2_X1 U10497 ( .A(n9251), .B(n9250), .Z(n9252) );
  OAI222_X1 U10498 ( .A1(n9462), .A2(n9254), .B1(n9464), .B2(n9253), .C1(n9252), .C2(n9459), .ZN(n9381) );
  NAND2_X1 U10499 ( .A1(n9381), .A2(n9281), .ZN(n9264) );
  INV_X1 U10500 ( .A(n9255), .ZN(n9256) );
  AOI211_X1 U10501 ( .C1(n9383), .C2(n9273), .A(n9692), .B(n9256), .ZN(n9382)
         );
  INV_X1 U10502 ( .A(n9383), .ZN(n9257) );
  NOR2_X1 U10503 ( .A1(n9257), .A2(n9656), .ZN(n9262) );
  OAI22_X1 U10504 ( .A1(n9281), .A2(n9260), .B1(n9259), .B2(n9258), .ZN(n9261)
         );
  AOI211_X1 U10505 ( .C1(n9382), .C2(n9475), .A(n9262), .B(n9261), .ZN(n9263)
         );
  OAI211_X1 U10506 ( .C1(n9385), .C2(n9308), .A(n9264), .B(n9263), .ZN(
        P1_U3274) );
  XNOR2_X1 U10507 ( .A(n9265), .B(n9269), .ZN(n9390) );
  NAND2_X1 U10508 ( .A1(n9267), .A2(n9266), .ZN(n9268) );
  XOR2_X1 U10509 ( .A(n9269), .B(n9268), .Z(n9270) );
  OAI222_X1 U10510 ( .A1(n9464), .A2(n9272), .B1(n9462), .B2(n9271), .C1(n9459), .C2(n9270), .ZN(n9386) );
  INV_X1 U10511 ( .A(n9284), .ZN(n9275) );
  INV_X1 U10512 ( .A(n9273), .ZN(n9274) );
  AOI211_X1 U10513 ( .C1(n9388), .C2(n9275), .A(n9692), .B(n9274), .ZN(n9387)
         );
  NAND2_X1 U10514 ( .A1(n9387), .A2(n9475), .ZN(n9278) );
  AOI22_X1 U10515 ( .A1(n4419), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9276), .B2(
        n9652), .ZN(n9277) );
  OAI211_X1 U10516 ( .C1(n9279), .C2(n9656), .A(n9278), .B(n9277), .ZN(n9280)
         );
  AOI21_X1 U10517 ( .B1(n9386), .B2(n9281), .A(n9280), .ZN(n9282) );
  OAI21_X1 U10518 ( .B1(n9308), .B2(n9390), .A(n9282), .ZN(P1_U3275) );
  XNOR2_X1 U10519 ( .A(n9283), .B(n9289), .ZN(n9397) );
  AOI21_X1 U10520 ( .B1(n9391), .B2(n9285), .A(n9284), .ZN(n9393) );
  AOI22_X1 U10521 ( .A1(n4419), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9286), .B2(
        n9652), .ZN(n9287) );
  OAI21_X1 U10522 ( .B1(n9288), .B2(n9656), .A(n9287), .ZN(n9298) );
  XNOR2_X1 U10523 ( .A(n9290), .B(n9289), .ZN(n9295) );
  AOI222_X1 U10524 ( .A1(n9296), .A2(n9295), .B1(n9294), .B2(n9293), .C1(n9292), .C2(n9291), .ZN(n9395) );
  NOR2_X1 U10525 ( .A1(n9395), .A2(n4419), .ZN(n9297) );
  AOI211_X1 U10526 ( .C1(n9393), .C2(n9650), .A(n9298), .B(n9297), .ZN(n9299)
         );
  OAI21_X1 U10527 ( .B1(n9308), .B2(n9397), .A(n9299), .ZN(P1_U3276) );
  AOI22_X1 U10528 ( .A1(n4419), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9300), .B2(
        n9652), .ZN(n9301) );
  OAI21_X1 U10529 ( .B1(n9302), .B2(n9656), .A(n9301), .ZN(n9305) );
  NOR2_X1 U10530 ( .A1(n9303), .A2(n4419), .ZN(n9304) );
  AOI211_X1 U10531 ( .C1(n9306), .C2(n9650), .A(n9305), .B(n9304), .ZN(n9307)
         );
  OAI21_X1 U10532 ( .B1(n9309), .B2(n9308), .A(n9307), .ZN(P1_U3278) );
  MUX2_X1 U10533 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9398), .S(n9702), .Z(
        P1_U3554) );
  NAND3_X1 U10534 ( .A1(n9313), .A2(n9471), .A3(n9312), .ZN(n9315) );
  OAI211_X1 U10535 ( .C1(n9316), .C2(n9691), .A(n9315), .B(n9314), .ZN(n9399)
         );
  MUX2_X1 U10536 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9399), .S(n9702), .Z(
        P1_U3553) );
  AOI22_X1 U10537 ( .A1(n9318), .A2(n9471), .B1(n9392), .B2(n9317), .ZN(n9319)
         );
  OAI211_X1 U10538 ( .C1(n9321), .C2(n9396), .A(n9320), .B(n9319), .ZN(n9400)
         );
  MUX2_X1 U10539 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9400), .S(n9702), .Z(
        P1_U3552) );
  AOI22_X1 U10540 ( .A1(n9323), .A2(n9471), .B1(n9392), .B2(n9322), .ZN(n9324)
         );
  OAI211_X1 U10541 ( .C1(n9326), .C2(n9396), .A(n9325), .B(n9324), .ZN(n9401)
         );
  MUX2_X1 U10542 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9401), .S(n9702), .Z(
        P1_U3551) );
  AOI21_X1 U10543 ( .B1(n9392), .B2(n9328), .A(n9327), .ZN(n9329) );
  OAI211_X1 U10544 ( .C1(n9331), .C2(n9396), .A(n9330), .B(n9329), .ZN(n9402)
         );
  MUX2_X1 U10545 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9402), .S(n9702), .Z(
        P1_U3550) );
  AOI22_X1 U10546 ( .A1(n9333), .A2(n9471), .B1(n9392), .B2(n9332), .ZN(n9334)
         );
  OAI211_X1 U10547 ( .C1(n9336), .C2(n9396), .A(n9335), .B(n9334), .ZN(n9403)
         );
  MUX2_X1 U10548 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9403), .S(n9702), .Z(
        P1_U3549) );
  AOI22_X1 U10549 ( .A1(n9338), .A2(n9471), .B1(n9392), .B2(n9337), .ZN(n9339)
         );
  OAI211_X1 U10550 ( .C1(n9341), .C2(n9396), .A(n9340), .B(n9339), .ZN(n9404)
         );
  MUX2_X1 U10551 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9404), .S(n9702), .Z(
        P1_U3548) );
  NAND2_X1 U10552 ( .A1(n9342), .A2(n9521), .ZN(n9347) );
  AOI211_X1 U10553 ( .C1(n9392), .C2(n9345), .A(n9344), .B(n9343), .ZN(n9346)
         );
  OAI21_X1 U10554 ( .B1(n9348), .B2(n9347), .A(n9346), .ZN(n9405) );
  MUX2_X1 U10555 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9405), .S(n9702), .Z(
        P1_U3547) );
  AOI22_X1 U10556 ( .A1(n9350), .A2(n9471), .B1(n9392), .B2(n9349), .ZN(n9351)
         );
  OAI211_X1 U10557 ( .C1(n9353), .C2(n9396), .A(n9352), .B(n9351), .ZN(n9406)
         );
  MUX2_X1 U10558 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9406), .S(n9702), .Z(
        P1_U3546) );
  AOI22_X1 U10559 ( .A1(n9355), .A2(n9471), .B1(n9392), .B2(n9354), .ZN(n9356)
         );
  OAI211_X1 U10560 ( .C1(n9358), .C2(n9396), .A(n9357), .B(n9356), .ZN(n9407)
         );
  MUX2_X1 U10561 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9407), .S(n9702), .Z(
        P1_U3545) );
  NAND2_X1 U10562 ( .A1(n9359), .A2(n9521), .ZN(n9364) );
  AOI211_X1 U10563 ( .C1(n9392), .C2(n9362), .A(n9361), .B(n9360), .ZN(n9363)
         );
  OAI21_X1 U10564 ( .B1(n9365), .B2(n9364), .A(n9363), .ZN(n9408) );
  MUX2_X1 U10565 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9408), .S(n9702), .Z(
        P1_U3544) );
  AOI211_X1 U10566 ( .C1(n9392), .C2(n9368), .A(n9367), .B(n9366), .ZN(n9369)
         );
  OAI21_X1 U10567 ( .B1(n9396), .B2(n9370), .A(n9369), .ZN(n9409) );
  MUX2_X1 U10568 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9409), .S(n9702), .Z(
        P1_U3543) );
  AOI21_X1 U10569 ( .B1(n9392), .B2(n9372), .A(n9371), .ZN(n9373) );
  OAI211_X1 U10570 ( .C1(n9375), .C2(n9396), .A(n9374), .B(n9373), .ZN(n9410)
         );
  MUX2_X1 U10571 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9410), .S(n9702), .Z(
        P1_U3542) );
  AOI21_X1 U10572 ( .B1(n9392), .B2(n9377), .A(n9376), .ZN(n9378) );
  OAI211_X1 U10573 ( .C1(n9380), .C2(n9396), .A(n9379), .B(n9378), .ZN(n9411)
         );
  MUX2_X1 U10574 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9411), .S(n9702), .Z(
        P1_U3541) );
  AOI211_X1 U10575 ( .C1(n9392), .C2(n9383), .A(n9382), .B(n9381), .ZN(n9384)
         );
  OAI21_X1 U10576 ( .B1(n9396), .B2(n9385), .A(n9384), .ZN(n9412) );
  MUX2_X1 U10577 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9412), .S(n9702), .Z(
        P1_U3540) );
  AOI211_X1 U10578 ( .C1(n9392), .C2(n9388), .A(n9387), .B(n9386), .ZN(n9389)
         );
  OAI21_X1 U10579 ( .B1(n9396), .B2(n9390), .A(n9389), .ZN(n9413) );
  MUX2_X1 U10580 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9413), .S(n9702), .Z(
        P1_U3539) );
  AOI22_X1 U10581 ( .A1(n9393), .A2(n9471), .B1(n9392), .B2(n9391), .ZN(n9394)
         );
  OAI211_X1 U10582 ( .C1(n9397), .C2(n9396), .A(n9395), .B(n9394), .ZN(n9414)
         );
  MUX2_X1 U10583 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9414), .S(n9702), .Z(
        P1_U3538) );
  MUX2_X1 U10584 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9399), .S(n9671), .Z(
        P1_U3521) );
  MUX2_X1 U10585 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9400), .S(n9671), .Z(
        P1_U3520) );
  MUX2_X1 U10586 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9401), .S(n9671), .Z(
        P1_U3519) );
  MUX2_X1 U10587 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9402), .S(n9671), .Z(
        P1_U3518) );
  MUX2_X1 U10588 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9403), .S(n9671), .Z(
        P1_U3517) );
  MUX2_X1 U10589 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9404), .S(n9671), .Z(
        P1_U3516) );
  MUX2_X1 U10590 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9405), .S(n9671), .Z(
        P1_U3515) );
  MUX2_X1 U10591 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9406), .S(n9671), .Z(
        P1_U3514) );
  MUX2_X1 U10592 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9407), .S(n9671), .Z(
        P1_U3513) );
  MUX2_X1 U10593 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9408), .S(n9671), .Z(
        P1_U3512) );
  MUX2_X1 U10594 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9409), .S(n9671), .Z(
        P1_U3511) );
  MUX2_X1 U10595 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9410), .S(n9671), .Z(
        P1_U3510) );
  MUX2_X1 U10596 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9411), .S(n9671), .Z(
        P1_U3508) );
  MUX2_X1 U10597 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9412), .S(n9671), .Z(
        P1_U3505) );
  MUX2_X1 U10598 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9413), .S(n9671), .Z(
        P1_U3502) );
  MUX2_X1 U10599 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9414), .S(n9671), .Z(
        P1_U3499) );
  NOR4_X1 U10600 ( .A1(n4961), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9415), .A4(
        P1_U3084), .ZN(n9416) );
  AOI21_X1 U10601 ( .B1(n9421), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9416), .ZN(
        n9417) );
  OAI21_X1 U10602 ( .B1(n9418), .B2(n9424), .A(n9417), .ZN(P1_U3322) );
  OAI222_X1 U10603 ( .A1(n9424), .A2(n9420), .B1(P1_U3084), .B2(n9419), .C1(
        n10079), .C2(n8231), .ZN(P1_U3324) );
  NAND2_X1 U10604 ( .A1(n9421), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9423) );
  OAI211_X1 U10605 ( .C1(n9425), .C2(n9424), .A(n9423), .B(n9422), .ZN(
        P1_U3325) );
  MUX2_X1 U10606 ( .A(n9426), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10607 ( .A1(n9875), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9439) );
  INV_X1 U10608 ( .A(n9427), .ZN(n9432) );
  AOI211_X1 U10609 ( .C1(n9430), .C2(n9429), .A(n9428), .B(n9869), .ZN(n9431)
         );
  AOI21_X1 U10610 ( .B1(n9433), .B2(n9432), .A(n9431), .ZN(n9438) );
  INV_X1 U10611 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9716) );
  NOR2_X1 U10612 ( .A1(n9716), .A2(n9712), .ZN(n9436) );
  OAI211_X1 U10613 ( .C1(n9436), .C2(n9435), .A(n9877), .B(n9434), .ZN(n9437)
         );
  NAND3_X1 U10614 ( .A1(n9439), .A2(n9438), .A3(n9437), .ZN(P2_U3246) );
  AOI22_X1 U10615 ( .A1(n9875), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9451) );
  OAI21_X1 U10616 ( .B1(n9442), .B2(n9441), .A(n9440), .ZN(n9443) );
  OAI22_X1 U10617 ( .A1(n9883), .A2(n9444), .B1(n9869), .B2(n9443), .ZN(n9445)
         );
  INV_X1 U10618 ( .A(n9445), .ZN(n9450) );
  OAI211_X1 U10619 ( .C1(n9448), .C2(n9447), .A(n9877), .B(n9446), .ZN(n9449)
         );
  NAND3_X1 U10620 ( .A1(n9451), .A2(n9450), .A3(n9449), .ZN(P2_U3247) );
  XNOR2_X1 U10621 ( .A(n9452), .B(n9454), .ZN(n9483) );
  INV_X1 U10622 ( .A(n9453), .ZN(n9461) );
  INV_X1 U10623 ( .A(n9454), .ZN(n9455) );
  AOI21_X1 U10624 ( .B1(n9457), .B2(n9456), .A(n9455), .ZN(n9458) );
  AOI211_X1 U10625 ( .C1(n9461), .C2(n9460), .A(n9459), .B(n9458), .ZN(n9467)
         );
  OAI22_X1 U10626 ( .A1(n9465), .A2(n9464), .B1(n9463), .B2(n9462), .ZN(n9466)
         );
  AOI211_X1 U10627 ( .C1(n9483), .C2(n9648), .A(n9467), .B(n9466), .ZN(n9480)
         );
  AOI222_X1 U10628 ( .A1(n9470), .A2(n9469), .B1(n9468), .B2(n9652), .C1(
        P1_REG2_REG_10__SCAN_IN), .C2(n4419), .ZN(n9477) );
  OAI211_X1 U10629 ( .C1(n9479), .C2(n9473), .A(n9472), .B(n9471), .ZN(n9478)
         );
  INV_X1 U10630 ( .A(n9478), .ZN(n9474) );
  AOI22_X1 U10631 ( .A1(n9483), .A2(n9659), .B1(n9475), .B2(n9474), .ZN(n9476)
         );
  OAI211_X1 U10632 ( .C1(n4419), .C2(n9480), .A(n9477), .B(n9476), .ZN(
        P1_U3281) );
  OAI21_X1 U10633 ( .B1(n9479), .B2(n9691), .A(n9478), .ZN(n9482) );
  INV_X1 U10634 ( .A(n9480), .ZN(n9481) );
  AOI211_X1 U10635 ( .C1(n9697), .C2(n9483), .A(n9482), .B(n9481), .ZN(n9485)
         );
  INV_X1 U10636 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9484) );
  AOI22_X1 U10637 ( .A1(n9671), .A2(n9485), .B1(n9484), .B2(n9698), .ZN(
        P1_U3484) );
  AOI22_X1 U10638 ( .A1(n9702), .A2(n9485), .B1(n5992), .B2(n9707), .ZN(
        P1_U3533) );
  INV_X1 U10639 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10219) );
  NOR2_X1 U10640 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9486) );
  AOI21_X1 U10641 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9486), .ZN(n9847) );
  NOR2_X1 U10642 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9487) );
  AOI21_X1 U10643 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9487), .ZN(n9850) );
  NOR2_X1 U10644 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9488) );
  AOI21_X1 U10645 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9488), .ZN(n9853) );
  NOR2_X1 U10646 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9489) );
  AOI21_X1 U10647 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9489), .ZN(n9856) );
  NOR2_X1 U10648 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9490) );
  AOI21_X1 U10649 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9490), .ZN(n9859) );
  NOR2_X1 U10650 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9497) );
  XNOR2_X1 U10651 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10227) );
  NAND2_X1 U10652 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9495) );
  XOR2_X1 U10653 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10225) );
  NAND2_X1 U10654 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9493) );
  XOR2_X1 U10655 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10222) );
  AOI21_X1 U10656 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9840) );
  INV_X1 U10657 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9491) );
  NAND3_X1 U10658 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9842) );
  OAI21_X1 U10659 ( .B1(n9840), .B2(n9491), .A(n9842), .ZN(n10221) );
  NAND2_X1 U10660 ( .A1(n10222), .A2(n10221), .ZN(n9492) );
  NAND2_X1 U10661 ( .A1(n9493), .A2(n9492), .ZN(n10224) );
  NAND2_X1 U10662 ( .A1(n10225), .A2(n10224), .ZN(n9494) );
  NAND2_X1 U10663 ( .A1(n9495), .A2(n9494), .ZN(n10226) );
  NOR2_X1 U10664 ( .A1(n10227), .A2(n10226), .ZN(n9496) );
  NOR2_X1 U10665 ( .A1(n9497), .A2(n9496), .ZN(n9498) );
  NOR2_X1 U10666 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9498), .ZN(n10215) );
  AND2_X1 U10667 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9498), .ZN(n10214) );
  NOR2_X1 U10668 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10214), .ZN(n9499) );
  NOR2_X1 U10669 ( .A1(n10215), .A2(n9499), .ZN(n9500) );
  NAND2_X1 U10670 ( .A1(n9500), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9502) );
  XOR2_X1 U10671 ( .A(n9500), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10213) );
  NAND2_X1 U10672 ( .A1(n10213), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9501) );
  NAND2_X1 U10673 ( .A1(n9502), .A2(n9501), .ZN(n9503) );
  NAND2_X1 U10674 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9503), .ZN(n9505) );
  XOR2_X1 U10675 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9503), .Z(n10208) );
  NAND2_X1 U10676 ( .A1(n10208), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9504) );
  NAND2_X1 U10677 ( .A1(n9505), .A2(n9504), .ZN(n9506) );
  NAND2_X1 U10678 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9506), .ZN(n9508) );
  XOR2_X1 U10679 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9506), .Z(n10223) );
  NAND2_X1 U10680 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10223), .ZN(n9507) );
  NAND2_X1 U10681 ( .A1(n9508), .A2(n9507), .ZN(n9509) );
  AND2_X1 U10682 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9509), .ZN(n9510) );
  XNOR2_X1 U10683 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9509), .ZN(n10211) );
  INV_X1 U10684 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10210) );
  NAND2_X1 U10685 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9511) );
  OAI21_X1 U10686 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9511), .ZN(n9867) );
  NAND2_X1 U10687 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9512) );
  OAI21_X1 U10688 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9512), .ZN(n9864) );
  AOI21_X1 U10689 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9863), .ZN(n9862) );
  NOR2_X1 U10690 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9513) );
  AOI21_X1 U10691 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9513), .ZN(n9861) );
  NAND2_X1 U10692 ( .A1(n9862), .A2(n9861), .ZN(n9860) );
  OAI21_X1 U10693 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9860), .ZN(n9858) );
  NAND2_X1 U10694 ( .A1(n9859), .A2(n9858), .ZN(n9857) );
  OAI21_X1 U10695 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9857), .ZN(n9855) );
  NAND2_X1 U10696 ( .A1(n9856), .A2(n9855), .ZN(n9854) );
  OAI21_X1 U10697 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9854), .ZN(n9852) );
  NAND2_X1 U10698 ( .A1(n9853), .A2(n9852), .ZN(n9851) );
  OAI21_X1 U10699 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9851), .ZN(n9849) );
  NAND2_X1 U10700 ( .A1(n9850), .A2(n9849), .ZN(n9848) );
  OAI21_X1 U10701 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9848), .ZN(n9846) );
  NAND2_X1 U10702 ( .A1(n9847), .A2(n9846), .ZN(n9845) );
  OAI21_X1 U10703 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9845), .ZN(n10218) );
  NOR2_X1 U10704 ( .A1(n10219), .A2(n10218), .ZN(n9514) );
  NAND2_X1 U10705 ( .A1(n10219), .A2(n10218), .ZN(n10217) );
  OAI21_X1 U10706 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9514), .A(n10217), .ZN(
        n9516) );
  XOR2_X1 U10707 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n9515) );
  XNOR2_X1 U10708 ( .A(n9516), .B(n9515), .ZN(ADD_1071_U4) );
  OAI21_X1 U10709 ( .B1(n9518), .B2(n9691), .A(n9517), .ZN(n9519) );
  AOI211_X1 U10710 ( .C1(n9522), .C2(n9521), .A(n9520), .B(n9519), .ZN(n9525)
         );
  AOI22_X1 U10711 ( .A1(n9702), .A2(n9525), .B1(n9523), .B2(n9707), .ZN(
        P1_U3537) );
  INV_X1 U10712 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9524) );
  AOI22_X1 U10713 ( .A1(n9671), .A2(n9525), .B1(n9524), .B2(n9698), .ZN(
        P1_U3496) );
  XNOR2_X1 U10714 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10715 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U10716 ( .B1(n9528), .B2(n9527), .A(n9526), .ZN(n9531) );
  NAND2_X1 U10717 ( .A1(n9635), .A2(n9529), .ZN(n9530) );
  OAI21_X1 U10718 ( .B1(n9629), .B2(n9531), .A(n9530), .ZN(n9539) );
  MUX2_X1 U10719 ( .A(n9534), .B(n9533), .S(n9532), .Z(n9537) );
  OAI211_X1 U10720 ( .C1(n9537), .C2(n9536), .A(P1_U4006), .B(n9535), .ZN(
        n9559) );
  INV_X1 U10721 ( .A(n9559), .ZN(n9538) );
  AOI211_X1 U10722 ( .C1(n9640), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n9539), .B(
        n9538), .ZN(n9544) );
  OAI211_X1 U10723 ( .C1(n9542), .C2(n9541), .A(n9641), .B(n9540), .ZN(n9543)
         );
  OAI211_X1 U10724 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n6150), .A(n9544), .B(
        n9543), .ZN(P1_U3243) );
  INV_X1 U10725 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9552) );
  MUX2_X1 U10726 ( .A(n5931), .B(P1_REG2_REG_4__SCAN_IN), .S(n9545), .Z(n9547)
         );
  OAI21_X1 U10727 ( .B1(n4510), .B2(n9547), .A(n9546), .ZN(n9548) );
  NAND2_X1 U10728 ( .A1(n9623), .A2(n9548), .ZN(n9551) );
  NAND2_X1 U10729 ( .A1(n9635), .A2(n9549), .ZN(n9550) );
  OAI211_X1 U10730 ( .C1(n9627), .C2(n9552), .A(n9551), .B(n9550), .ZN(n9553)
         );
  INV_X1 U10731 ( .A(n9553), .ZN(n9561) );
  OAI21_X1 U10732 ( .B1(n9556), .B2(n9555), .A(n9554), .ZN(n9557) );
  NAND2_X1 U10733 ( .A1(n9641), .A2(n9557), .ZN(n9558) );
  NAND4_X1 U10734 ( .A1(n9561), .A2(n9560), .A3(n9559), .A4(n9558), .ZN(
        P1_U3245) );
  AOI22_X1 U10735 ( .A1(n9640), .A2(P1_ADDR_REG_7__SCAN_IN), .B1(n9635), .B2(
        n9562), .ZN(n9574) );
  NAND2_X1 U10736 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3084), .ZN(n9573) );
  NOR2_X1 U10737 ( .A1(n9564), .A2(n9563), .ZN(n9565) );
  OAI21_X1 U10738 ( .B1(n9566), .B2(n9565), .A(n9623), .ZN(n9572) );
  NOR2_X1 U10739 ( .A1(n9568), .A2(n9567), .ZN(n9569) );
  OAI21_X1 U10740 ( .B1(n9570), .B2(n9569), .A(n9641), .ZN(n9571) );
  NAND4_X1 U10741 ( .A1(n9574), .A2(n9573), .A3(n9572), .A4(n9571), .ZN(
        P1_U3248) );
  OAI21_X1 U10742 ( .B1(n6576), .B2(n9582), .A(n9575), .ZN(n9576) );
  XNOR2_X1 U10743 ( .A(n9577), .B(n9576), .ZN(n9578) );
  AOI22_X1 U10744 ( .A1(n9578), .A2(n9623), .B1(n9640), .B2(
        P1_ADDR_REG_8__SCAN_IN), .ZN(n9588) );
  INV_X1 U10745 ( .A(n9579), .ZN(n9587) );
  AND3_X1 U10746 ( .A1(n9584), .A2(P1_REG1_REG_8__SCAN_IN), .A3(n9641), .ZN(
        n9581) );
  OAI21_X1 U10747 ( .B1(n9581), .B2(n9635), .A(n9580), .ZN(n9586) );
  NAND2_X1 U10748 ( .A1(n9582), .A2(n9708), .ZN(n9583) );
  OAI211_X1 U10749 ( .C1(n9584), .C2(n9583), .A(n9590), .B(n9641), .ZN(n9585)
         );
  NAND4_X1 U10750 ( .A1(n9588), .A2(n9587), .A3(n9586), .A4(n9585), .ZN(
        P1_U3249) );
  OAI21_X1 U10751 ( .B1(n9591), .B2(n9590), .A(n9589), .ZN(n9594) );
  INV_X1 U10752 ( .A(n9592), .ZN(n9593) );
  AOI21_X1 U10753 ( .B1(n9594), .B2(n9641), .A(n9593), .ZN(n9601) );
  AOI211_X1 U10754 ( .C1(n9597), .C2(n9596), .A(n9595), .B(n9629), .ZN(n9598)
         );
  AOI21_X1 U10755 ( .B1(n9635), .B2(n9599), .A(n9598), .ZN(n9600) );
  OAI211_X1 U10756 ( .C1(n9627), .C2(n10210), .A(n9601), .B(n9600), .ZN(
        P1_U3250) );
  INV_X1 U10757 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9613) );
  AOI21_X1 U10758 ( .B1(n9635), .B2(n9603), .A(n9602), .ZN(n9612) );
  OAI21_X1 U10759 ( .B1(n9606), .B2(n9605), .A(n9604), .ZN(n9610) );
  OAI21_X1 U10760 ( .B1(n4504), .B2(n9608), .A(n9607), .ZN(n9609) );
  AOI22_X1 U10761 ( .A1(n9610), .A2(n9641), .B1(n9623), .B2(n9609), .ZN(n9611)
         );
  OAI211_X1 U10762 ( .C1(n9627), .C2(n9613), .A(n9612), .B(n9611), .ZN(
        P1_U3252) );
  INV_X1 U10763 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10138) );
  AOI21_X1 U10764 ( .B1(n9635), .B2(n9615), .A(n9614), .ZN(n9626) );
  OAI21_X1 U10765 ( .B1(n9618), .B2(n9617), .A(n9616), .ZN(n9624) );
  OAI21_X1 U10766 ( .B1(n9621), .B2(n9620), .A(n9619), .ZN(n9622) );
  AOI22_X1 U10767 ( .A1(n9624), .A2(n9623), .B1(n9641), .B2(n9622), .ZN(n9625)
         );
  OAI211_X1 U10768 ( .C1(n9627), .C2(n10138), .A(n9626), .B(n9625), .ZN(
        P1_U3255) );
  INV_X1 U10769 ( .A(n9628), .ZN(n9634) );
  AOI211_X1 U10770 ( .C1(n9632), .C2(n9631), .A(n9630), .B(n9629), .ZN(n9633)
         );
  AOI211_X1 U10771 ( .C1(n9636), .C2(n9635), .A(n9634), .B(n9633), .ZN(n9644)
         );
  OAI21_X1 U10772 ( .B1(n9639), .B2(n9638), .A(n9637), .ZN(n9642) );
  AOI22_X1 U10773 ( .A1(n9642), .A2(n9641), .B1(n9640), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n9643) );
  NAND2_X1 U10774 ( .A1(n9644), .A2(n9643), .ZN(P1_U3259) );
  INV_X1 U10775 ( .A(n9645), .ZN(n9660) );
  INV_X1 U10776 ( .A(n9646), .ZN(n9647) );
  AOI21_X1 U10777 ( .B1(n9648), .B2(n9660), .A(n9647), .ZN(n9662) );
  INV_X1 U10778 ( .A(n9649), .ZN(n9657) );
  NAND2_X1 U10779 ( .A1(n9651), .A2(n9650), .ZN(n9655) );
  AOI22_X1 U10780 ( .A1(n4419), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n9653), .B2(
        n9652), .ZN(n9654) );
  OAI211_X1 U10781 ( .C1(n9657), .C2(n9656), .A(n9655), .B(n9654), .ZN(n9658)
         );
  AOI21_X1 U10782 ( .B1(n9660), .B2(n9659), .A(n9658), .ZN(n9661) );
  OAI21_X1 U10783 ( .B1(n4419), .B2(n9662), .A(n9661), .ZN(P1_U3282) );
  AND2_X1 U10784 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9664), .ZN(P1_U3292) );
  AND2_X1 U10785 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9664), .ZN(P1_U3293) );
  AND2_X1 U10786 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9664), .ZN(P1_U3294) );
  AND2_X1 U10787 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9664), .ZN(P1_U3295) );
  AND2_X1 U10788 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9664), .ZN(P1_U3296) );
  NOR2_X1 U10789 ( .A1(n9663), .A2(n10123), .ZN(P1_U3297) );
  AND2_X1 U10790 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9664), .ZN(P1_U3298) );
  AND2_X1 U10791 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9664), .ZN(P1_U3299) );
  INV_X1 U10792 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10029) );
  NOR2_X1 U10793 ( .A1(n9663), .A2(n10029), .ZN(P1_U3300) );
  INV_X1 U10794 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9965) );
  NOR2_X1 U10795 ( .A1(n9663), .A2(n9965), .ZN(P1_U3301) );
  AND2_X1 U10796 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9664), .ZN(P1_U3302) );
  AND2_X1 U10797 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9664), .ZN(P1_U3303) );
  INV_X1 U10798 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10018) );
  NOR2_X1 U10799 ( .A1(n9663), .A2(n10018), .ZN(P1_U3304) );
  NOR2_X1 U10800 ( .A1(n9663), .A2(n10137), .ZN(P1_U3305) );
  AND2_X1 U10801 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9664), .ZN(P1_U3306) );
  NOR2_X1 U10802 ( .A1(n9663), .A2(n10181), .ZN(P1_U3307) );
  AND2_X1 U10803 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9664), .ZN(P1_U3308) );
  AND2_X1 U10804 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9664), .ZN(P1_U3309) );
  AND2_X1 U10805 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9664), .ZN(P1_U3310) );
  NOR2_X1 U10806 ( .A1(n9663), .A2(n10094), .ZN(P1_U3311) );
  AND2_X1 U10807 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9664), .ZN(P1_U3312) );
  INV_X1 U10808 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10105) );
  NOR2_X1 U10809 ( .A1(n9663), .A2(n10105), .ZN(P1_U3313) );
  AND2_X1 U10810 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9664), .ZN(P1_U3314) );
  AND2_X1 U10811 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9664), .ZN(P1_U3315) );
  AND2_X1 U10812 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9664), .ZN(P1_U3316) );
  AND2_X1 U10813 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9664), .ZN(P1_U3317) );
  AND2_X1 U10814 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9664), .ZN(P1_U3318) );
  AND2_X1 U10815 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9664), .ZN(P1_U3319) );
  AND2_X1 U10816 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9664), .ZN(P1_U3320) );
  AND2_X1 U10817 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9664), .ZN(P1_U3321) );
  INV_X1 U10818 ( .A(n9665), .ZN(n9669) );
  OAI21_X1 U10819 ( .B1(n4636), .B2(n9691), .A(n9666), .ZN(n9668) );
  AOI211_X1 U10820 ( .C1(n9697), .C2(n9669), .A(n9668), .B(n9667), .ZN(n9701)
         );
  INV_X1 U10821 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9670) );
  AOI22_X1 U10822 ( .A1(n9671), .A2(n9701), .B1(n9670), .B2(n9698), .ZN(
        P1_U3457) );
  OR3_X1 U10823 ( .A1(n9672), .A2(n4508), .A3(n9692), .ZN(n9673) );
  OAI21_X1 U10824 ( .B1(n9674), .B2(n9691), .A(n9673), .ZN(n9676) );
  AOI211_X1 U10825 ( .C1(n9697), .C2(n9677), .A(n9676), .B(n9675), .ZN(n9703)
         );
  INV_X1 U10826 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10189) );
  AOI22_X1 U10827 ( .A1(n9671), .A2(n9703), .B1(n10189), .B2(n9698), .ZN(
        P1_U3460) );
  INV_X1 U10828 ( .A(n9678), .ZN(n9680) );
  OAI22_X1 U10829 ( .A1(n9680), .A2(n9692), .B1(n9679), .B2(n9691), .ZN(n9682)
         );
  AOI211_X1 U10830 ( .C1(n9697), .C2(n9683), .A(n9682), .B(n9681), .ZN(n9704)
         );
  INV_X1 U10831 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10141) );
  AOI22_X1 U10832 ( .A1(n9671), .A2(n9704), .B1(n10141), .B2(n9698), .ZN(
        P1_U3466) );
  OAI22_X1 U10833 ( .A1(n9685), .A2(n9692), .B1(n9684), .B2(n9691), .ZN(n9687)
         );
  AOI211_X1 U10834 ( .C1(n9697), .C2(n9688), .A(n9687), .B(n9686), .ZN(n9706)
         );
  INV_X1 U10835 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9954) );
  AOI22_X1 U10836 ( .A1(n9671), .A2(n9706), .B1(n9954), .B2(n9698), .ZN(
        P1_U3472) );
  INV_X1 U10837 ( .A(n9689), .ZN(n9696) );
  OAI22_X1 U10838 ( .A1(n9693), .A2(n9692), .B1(n4729), .B2(n9691), .ZN(n9695)
         );
  AOI211_X1 U10839 ( .C1(n9697), .C2(n9696), .A(n9695), .B(n9694), .ZN(n9709)
         );
  INV_X1 U10840 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9699) );
  AOI22_X1 U10841 ( .A1(n9671), .A2(n9709), .B1(n9699), .B2(n9698), .ZN(
        P1_U3478) );
  AOI22_X1 U10842 ( .A1(n9702), .A2(n9701), .B1(n9700), .B2(n9707), .ZN(
        P1_U3524) );
  AOI22_X1 U10843 ( .A1(n9702), .A2(n9703), .B1(n5906), .B2(n9707), .ZN(
        P1_U3525) );
  AOI22_X1 U10844 ( .A1(n9702), .A2(n9704), .B1(n10032), .B2(n9707), .ZN(
        P1_U3527) );
  AOI22_X1 U10845 ( .A1(n9702), .A2(n9706), .B1(n9705), .B2(n9707), .ZN(
        P1_U3529) );
  AOI22_X1 U10846 ( .A1(n9702), .A2(n9709), .B1(n9708), .B2(n9707), .ZN(
        P1_U3531) );
  INV_X1 U10847 ( .A(n9710), .ZN(n9713) );
  OAI211_X1 U10848 ( .C1(n9869), .C2(P2_REG1_REG_0__SCAN_IN), .A(
        P2_IR_REG_0__SCAN_IN), .B(n9883), .ZN(n9711) );
  AOI21_X1 U10849 ( .B1(n9713), .B2(n9712), .A(n9711), .ZN(n9718) );
  AOI22_X1 U10850 ( .A1(n9877), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9714), .ZN(n9717) );
  AOI22_X1 U10851 ( .A1(n9875), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9715) );
  OAI221_X1 U10852 ( .B1(n9718), .B2(n9717), .C1(n9718), .C2(n9716), .A(n9715), 
        .ZN(P2_U3245) );
  NAND2_X1 U10853 ( .A1(n9719), .A2(n9730), .ZN(n9720) );
  NAND2_X1 U10854 ( .A1(n9721), .A2(n9720), .ZN(n9741) );
  INV_X1 U10855 ( .A(n9741), .ZN(n9792) );
  INV_X1 U10856 ( .A(n9722), .ZN(n9728) );
  INV_X1 U10857 ( .A(n9723), .ZN(n9725) );
  OAI21_X1 U10858 ( .B1(n9725), .B2(n9788), .A(n9724), .ZN(n9789) );
  INV_X1 U10859 ( .A(n9789), .ZN(n9726) );
  AOI22_X1 U10860 ( .A1(n9792), .A2(n9728), .B1(n9727), .B2(n9726), .ZN(n9751)
         );
  OAI21_X1 U10861 ( .B1(n9731), .B2(n9730), .A(n9729), .ZN(n9738) );
  OAI22_X1 U10862 ( .A1(n9735), .A2(n9734), .B1(n9733), .B2(n9732), .ZN(n9736)
         );
  AOI21_X1 U10863 ( .B1(n9738), .B2(n9737), .A(n9736), .ZN(n9739) );
  OAI21_X1 U10864 ( .B1(n9741), .B2(n9740), .A(n9739), .ZN(n9790) );
  NOR2_X1 U10865 ( .A1(n9743), .A2(n9742), .ZN(n9744) );
  AOI21_X1 U10866 ( .B1(n9745), .B2(P2_REG2_REG_8__SCAN_IN), .A(n9744), .ZN(
        n9746) );
  OAI21_X1 U10867 ( .B1(n9788), .B2(n9747), .A(n9746), .ZN(n9748) );
  AOI21_X1 U10868 ( .B1(n9790), .B2(n9749), .A(n9748), .ZN(n9750) );
  NAND2_X1 U10869 ( .A1(n9751), .A2(n9750), .ZN(P2_U3288) );
  AND2_X1 U10870 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9757), .ZN(P2_U3297) );
  INV_X1 U10871 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n10043) );
  NOR2_X1 U10872 ( .A1(n9754), .A2(n10043), .ZN(P2_U3298) );
  AND2_X1 U10873 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9757), .ZN(P2_U3299) );
  AND2_X1 U10874 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9757), .ZN(P2_U3300) );
  AND2_X1 U10875 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9757), .ZN(P2_U3301) );
  AND2_X1 U10876 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9757), .ZN(P2_U3302) );
  AND2_X1 U10877 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9757), .ZN(P2_U3303) );
  INV_X1 U10878 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10060) );
  NOR2_X1 U10879 ( .A1(n9754), .A2(n10060), .ZN(P2_U3304) );
  AND2_X1 U10880 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9757), .ZN(P2_U3305) );
  AND2_X1 U10881 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9757), .ZN(P2_U3306) );
  INV_X1 U10882 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10082) );
  NOR2_X1 U10883 ( .A1(n9754), .A2(n10082), .ZN(P2_U3307) );
  AND2_X1 U10884 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9757), .ZN(P2_U3308) );
  AND2_X1 U10885 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9757), .ZN(P2_U3309) );
  AND2_X1 U10886 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9757), .ZN(P2_U3310) );
  INV_X1 U10887 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10035) );
  NOR2_X1 U10888 ( .A1(n9754), .A2(n10035), .ZN(P2_U3311) );
  INV_X1 U10889 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9978) );
  NOR2_X1 U10890 ( .A1(n9754), .A2(n9978), .ZN(P2_U3312) );
  AND2_X1 U10891 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9757), .ZN(P2_U3313) );
  INV_X1 U10892 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10030) );
  NOR2_X1 U10893 ( .A1(n9754), .A2(n10030), .ZN(P2_U3314) );
  AND2_X1 U10894 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9757), .ZN(P2_U3315) );
  AND2_X1 U10895 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9757), .ZN(P2_U3316) );
  AND2_X1 U10896 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9757), .ZN(P2_U3317) );
  AND2_X1 U10897 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9757), .ZN(P2_U3318) );
  AND2_X1 U10898 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9757), .ZN(P2_U3319) );
  INV_X1 U10899 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10093) );
  NOR2_X1 U10900 ( .A1(n9754), .A2(n10093), .ZN(P2_U3320) );
  AND2_X1 U10901 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9757), .ZN(P2_U3321) );
  AND2_X1 U10902 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9757), .ZN(P2_U3322) );
  AND2_X1 U10903 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9757), .ZN(P2_U3323) );
  INV_X1 U10904 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n9964) );
  NOR2_X1 U10905 ( .A1(n9754), .A2(n9964), .ZN(P2_U3324) );
  INV_X1 U10906 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10090) );
  NOR2_X1 U10907 ( .A1(n9754), .A2(n10090), .ZN(P2_U3325) );
  INV_X1 U10908 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10000) );
  NOR2_X1 U10909 ( .A1(n9754), .A2(n10000), .ZN(P2_U3326) );
  AOI22_X1 U10910 ( .A1(n9760), .A2(n9756), .B1(n9755), .B2(n9757), .ZN(
        P2_U3437) );
  AOI22_X1 U10911 ( .A1(n9760), .A2(n9759), .B1(n9758), .B2(n9757), .ZN(
        P2_U3438) );
  INV_X1 U10912 ( .A(n9761), .ZN(n9767) );
  OAI22_X1 U10913 ( .A1(n9765), .A2(n9764), .B1(n9763), .B2(n9762), .ZN(n9766)
         );
  NOR2_X1 U10914 ( .A1(n9767), .A2(n9766), .ZN(n9827) );
  INV_X1 U10915 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10183) );
  AOI22_X1 U10916 ( .A1(n9826), .A2(n9827), .B1(n10183), .B2(n9824), .ZN(
        P2_U3451) );
  OAI211_X1 U10917 ( .C1(n9770), .C2(n9810), .A(n9769), .B(n9768), .ZN(n9771)
         );
  AOI21_X1 U10918 ( .B1(n9822), .B2(n9772), .A(n9771), .ZN(n9828) );
  INV_X1 U10919 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U10920 ( .A1(n9826), .A2(n9828), .B1(n10175), .B2(n9824), .ZN(
        P2_U3466) );
  AOI22_X1 U10921 ( .A1(n9775), .A2(n9774), .B1(n9815), .B2(n9773), .ZN(n9779)
         );
  NAND3_X1 U10922 ( .A1(n9777), .A2(n9776), .A3(n9822), .ZN(n9778) );
  AND3_X1 U10923 ( .A1(n9780), .A2(n9779), .A3(n9778), .ZN(n9830) );
  INV_X1 U10924 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9781) );
  AOI22_X1 U10925 ( .A1(n9826), .A2(n9830), .B1(n9781), .B2(n9824), .ZN(
        P2_U3469) );
  OAI21_X1 U10926 ( .B1(n9783), .B2(n9810), .A(n9782), .ZN(n9784) );
  AOI211_X1 U10927 ( .C1(n9786), .C2(n9822), .A(n9785), .B(n9784), .ZN(n9831)
         );
  INV_X1 U10928 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9967) );
  AOI22_X1 U10929 ( .A1(n9826), .A2(n9831), .B1(n9967), .B2(n9824), .ZN(
        P2_U3472) );
  INV_X1 U10930 ( .A(n9787), .ZN(n9807) );
  OAI22_X1 U10931 ( .A1(n9789), .A2(n9820), .B1(n9788), .B2(n9810), .ZN(n9791)
         );
  AOI211_X1 U10932 ( .C1(n9807), .C2(n9792), .A(n9791), .B(n9790), .ZN(n9832)
         );
  INV_X1 U10933 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9793) );
  AOI22_X1 U10934 ( .A1(n9826), .A2(n9832), .B1(n9793), .B2(n9824), .ZN(
        P2_U3475) );
  INV_X1 U10935 ( .A(n9794), .ZN(n9799) );
  OAI22_X1 U10936 ( .A1(n9796), .A2(n9820), .B1(n9795), .B2(n9810), .ZN(n9798)
         );
  AOI211_X1 U10937 ( .C1(n9807), .C2(n9799), .A(n9798), .B(n9797), .ZN(n9834)
         );
  INV_X1 U10938 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9800) );
  AOI22_X1 U10939 ( .A1(n9826), .A2(n9834), .B1(n9800), .B2(n9824), .ZN(
        P2_U3478) );
  INV_X1 U10940 ( .A(n9801), .ZN(n9806) );
  OAI22_X1 U10941 ( .A1(n9803), .A2(n9820), .B1(n9802), .B2(n9810), .ZN(n9805)
         );
  AOI211_X1 U10942 ( .C1(n9807), .C2(n9806), .A(n9805), .B(n9804), .ZN(n9835)
         );
  INV_X1 U10943 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10036) );
  AOI22_X1 U10944 ( .A1(n9826), .A2(n9835), .B1(n10036), .B2(n9824), .ZN(
        P2_U3481) );
  OAI211_X1 U10945 ( .C1(n9811), .C2(n9810), .A(n9809), .B(n9808), .ZN(n9812)
         );
  AOI21_X1 U10946 ( .B1(n9813), .B2(n9822), .A(n9812), .ZN(n9836) );
  INV_X1 U10947 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9814) );
  AOI22_X1 U10948 ( .A1(n9826), .A2(n9836), .B1(n9814), .B2(n9824), .ZN(
        P2_U3484) );
  NAND2_X1 U10949 ( .A1(n9816), .A2(n9815), .ZN(n9817) );
  OAI211_X1 U10950 ( .C1(n9820), .C2(n9819), .A(n9818), .B(n9817), .ZN(n9821)
         );
  AOI21_X1 U10951 ( .B1(n9823), .B2(n9822), .A(n9821), .ZN(n9838) );
  INV_X1 U10952 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9825) );
  AOI22_X1 U10953 ( .A1(n9826), .A2(n9838), .B1(n9825), .B2(n9824), .ZN(
        P2_U3487) );
  INV_X1 U10954 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10143) );
  AOI22_X1 U10955 ( .A1(n9839), .A2(n9827), .B1(n10143), .B2(n9837), .ZN(
        P2_U3520) );
  INV_X1 U10956 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10046) );
  AOI22_X1 U10957 ( .A1(n9839), .A2(n9828), .B1(n10046), .B2(n9837), .ZN(
        P2_U3525) );
  INV_X1 U10958 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9829) );
  AOI22_X1 U10959 ( .A1(n9839), .A2(n9830), .B1(n9829), .B2(n9837), .ZN(
        P2_U3526) );
  INV_X1 U10960 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10113) );
  AOI22_X1 U10961 ( .A1(n9839), .A2(n9831), .B1(n10113), .B2(n9837), .ZN(
        P2_U3527) );
  AOI22_X1 U10962 ( .A1(n9839), .A2(n9832), .B1(n8020), .B2(n9837), .ZN(
        P2_U3528) );
  INV_X1 U10963 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9833) );
  AOI22_X1 U10964 ( .A1(n9839), .A2(n9834), .B1(n9833), .B2(n9837), .ZN(
        P2_U3529) );
  AOI22_X1 U10965 ( .A1(n9839), .A2(n9835), .B1(n8023), .B2(n9837), .ZN(
        P2_U3530) );
  AOI22_X1 U10966 ( .A1(n9839), .A2(n9836), .B1(n8024), .B2(n9837), .ZN(
        P2_U3531) );
  AOI22_X1 U10967 ( .A1(n9839), .A2(n9838), .B1(n8025), .B2(n9837), .ZN(
        P2_U3532) );
  INV_X1 U10968 ( .A(n9840), .ZN(n9841) );
  NAND2_X1 U10969 ( .A1(n9842), .A2(n9841), .ZN(n9843) );
  XNOR2_X1 U10970 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9843), .ZN(ADD_1071_U5) );
  INV_X1 U10971 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10076) );
  INV_X1 U10972 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9844) );
  AOI22_X1 U10973 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n10076), .B2(n9844), .ZN(ADD_1071_U46) );
  OAI21_X1 U10974 ( .B1(n9847), .B2(n9846), .A(n9845), .ZN(ADD_1071_U56) );
  OAI21_X1 U10975 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(ADD_1071_U57) );
  OAI21_X1 U10976 ( .B1(n9853), .B2(n9852), .A(n9851), .ZN(ADD_1071_U58) );
  OAI21_X1 U10977 ( .B1(n9856), .B2(n9855), .A(n9854), .ZN(ADD_1071_U59) );
  OAI21_X1 U10978 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(ADD_1071_U60) );
  OAI21_X1 U10979 ( .B1(n9862), .B2(n9861), .A(n9860), .ZN(ADD_1071_U61) );
  AOI21_X1 U10980 ( .B1(n9865), .B2(n9864), .A(n9863), .ZN(ADD_1071_U62) );
  AOI21_X1 U10981 ( .B1(n9868), .B2(n9867), .A(n9866), .ZN(ADD_1071_U63) );
  AOI211_X1 U10982 ( .C1(n9872), .C2(n9871), .A(n9870), .B(n9869), .ZN(n9873)
         );
  AOI211_X1 U10983 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n9875), .A(n9874), .B(
        n9873), .ZN(n9881) );
  OAI211_X1 U10984 ( .C1(n9879), .C2(n9878), .A(n9877), .B(n9876), .ZN(n9880)
         );
  OAI211_X1 U10985 ( .C1(n9883), .C2(n9882), .A(n9881), .B(n9880), .ZN(n10206)
         );
  INV_X1 U10986 ( .A(keyinput50), .ZN(n9884) );
  NOR4_X1 U10987 ( .A1(keyinput89), .A2(keyinput64), .A3(keyinput101), .A4(
        n9884), .ZN(n9947) );
  NAND2_X1 U10988 ( .A1(keyinput2), .A2(keyinput9), .ZN(n9885) );
  NOR3_X1 U10989 ( .A1(keyinput29), .A2(keyinput33), .A3(n9885), .ZN(n9946) );
  NAND2_X1 U10990 ( .A1(keyinput66), .A2(keyinput87), .ZN(n9886) );
  NOR3_X1 U10991 ( .A1(keyinput56), .A2(keyinput121), .A3(n9886), .ZN(n9887)
         );
  NAND3_X1 U10992 ( .A1(keyinput21), .A2(keyinput47), .A3(n9887), .ZN(n9896)
         );
  NAND2_X1 U10993 ( .A1(keyinput22), .A2(keyinput11), .ZN(n9888) );
  NOR3_X1 U10994 ( .A1(keyinput83), .A2(keyinput71), .A3(n9888), .ZN(n9894) );
  NAND3_X1 U10995 ( .A1(keyinput67), .A2(keyinput73), .A3(keyinput16), .ZN(
        n9889) );
  NOR2_X1 U10996 ( .A1(keyinput30), .A2(n9889), .ZN(n9893) );
  NAND3_X1 U10997 ( .A1(keyinput107), .A2(keyinput118), .A3(keyinput112), .ZN(
        n9890) );
  NOR2_X1 U10998 ( .A1(keyinput84), .A2(n9890), .ZN(n9892) );
  NOR4_X1 U10999 ( .A1(keyinput34), .A2(keyinput114), .A3(keyinput62), .A4(
        keyinput15), .ZN(n9891) );
  NAND4_X1 U11000 ( .A1(n9894), .A2(n9893), .A3(n9892), .A4(n9891), .ZN(n9895)
         );
  NOR4_X1 U11001 ( .A1(keyinput0), .A2(keyinput105), .A3(n9896), .A4(n9895), 
        .ZN(n9945) );
  NAND2_X1 U11002 ( .A1(keyinput104), .A2(keyinput4), .ZN(n9897) );
  NOR3_X1 U11003 ( .A1(keyinput28), .A2(keyinput39), .A3(n9897), .ZN(n9899) );
  INV_X1 U11004 ( .A(keyinput120), .ZN(n9898) );
  NAND4_X1 U11005 ( .A1(keyinput113), .A2(keyinput116), .A3(n9899), .A4(n9898), 
        .ZN(n9943) );
  NOR2_X1 U11006 ( .A1(keyinput99), .A2(keyinput38), .ZN(n9900) );
  NAND3_X1 U11007 ( .A1(keyinput17), .A2(keyinput123), .A3(n9900), .ZN(n9901)
         );
  NOR3_X1 U11008 ( .A1(keyinput81), .A2(keyinput7), .A3(n9901), .ZN(n9910) );
  NOR2_X1 U11009 ( .A1(keyinput127), .A2(keyinput40), .ZN(n9902) );
  NAND3_X1 U11010 ( .A1(keyinput60), .A2(keyinput98), .A3(n9902), .ZN(n9908)
         );
  INV_X1 U11011 ( .A(keyinput61), .ZN(n9903) );
  NAND4_X1 U11012 ( .A1(keyinput35), .A2(keyinput55), .A3(keyinput37), .A4(
        n9903), .ZN(n9907) );
  OR4_X1 U11013 ( .A1(keyinput77), .A2(keyinput54), .A3(keyinput70), .A4(
        keyinput80), .ZN(n9906) );
  INV_X1 U11014 ( .A(keyinput85), .ZN(n9904) );
  NAND4_X1 U11015 ( .A1(keyinput44), .A2(keyinput6), .A3(keyinput12), .A4(
        n9904), .ZN(n9905) );
  NOR4_X1 U11016 ( .A1(n9908), .A2(n9907), .A3(n9906), .A4(n9905), .ZN(n9909)
         );
  NAND4_X1 U11017 ( .A1(keyinput58), .A2(keyinput19), .A3(n9910), .A4(n9909), 
        .ZN(n9942) );
  NOR2_X1 U11018 ( .A1(keyinput27), .A2(keyinput5), .ZN(n9911) );
  NAND3_X1 U11019 ( .A1(keyinput102), .A2(keyinput24), .A3(n9911), .ZN(n9912)
         );
  NOR3_X1 U11020 ( .A1(keyinput82), .A2(keyinput51), .A3(n9912), .ZN(n9924) );
  NAND2_X1 U11021 ( .A1(keyinput45), .A2(keyinput126), .ZN(n9913) );
  NOR3_X1 U11022 ( .A1(keyinput72), .A2(keyinput25), .A3(n9913), .ZN(n9914) );
  NAND3_X1 U11023 ( .A1(keyinput13), .A2(keyinput97), .A3(n9914), .ZN(n9922)
         );
  AND4_X1 U11024 ( .A1(keyinput92), .A2(keyinput23), .A3(keyinput18), .A4(
        keyinput76), .ZN(n9920) );
  NOR4_X1 U11025 ( .A1(keyinput42), .A2(keyinput103), .A3(keyinput57), .A4(
        keyinput65), .ZN(n9919) );
  NAND2_X1 U11026 ( .A1(keyinput48), .A2(keyinput124), .ZN(n9915) );
  NOR3_X1 U11027 ( .A1(keyinput46), .A2(keyinput41), .A3(n9915), .ZN(n9918) );
  INV_X1 U11028 ( .A(keyinput3), .ZN(n9916) );
  NOR4_X1 U11029 ( .A1(keyinput100), .A2(keyinput91), .A3(keyinput88), .A4(
        n9916), .ZN(n9917) );
  NAND4_X1 U11030 ( .A1(n9920), .A2(n9919), .A3(n9918), .A4(n9917), .ZN(n9921)
         );
  NOR4_X1 U11031 ( .A1(keyinput110), .A2(keyinput74), .A3(n9922), .A4(n9921), 
        .ZN(n9923) );
  NAND4_X1 U11032 ( .A1(keyinput90), .A2(keyinput1), .A3(n9924), .A4(n9923), 
        .ZN(n9941) );
  NOR4_X1 U11033 ( .A1(keyinput26), .A2(keyinput10), .A3(keyinput68), .A4(
        keyinput79), .ZN(n9939) );
  NAND2_X1 U11034 ( .A1(keyinput75), .A2(keyinput115), .ZN(n9925) );
  NOR3_X1 U11035 ( .A1(keyinput43), .A2(keyinput86), .A3(n9925), .ZN(n9938) );
  INV_X1 U11036 ( .A(keyinput96), .ZN(n9926) );
  NOR4_X1 U11037 ( .A1(keyinput69), .A2(keyinput49), .A3(keyinput36), .A4(
        n9926), .ZN(n9927) );
  NAND3_X1 U11038 ( .A1(keyinput109), .A2(keyinput14), .A3(n9927), .ZN(n9928)
         );
  NOR3_X1 U11039 ( .A1(keyinput94), .A2(keyinput53), .A3(n9928), .ZN(n9937) );
  INV_X1 U11040 ( .A(keyinput8), .ZN(n9929) );
  NAND4_X1 U11041 ( .A1(keyinput111), .A2(keyinput31), .A3(keyinput122), .A4(
        n9929), .ZN(n9935) );
  NOR2_X1 U11042 ( .A1(keyinput117), .A2(keyinput108), .ZN(n9930) );
  NAND3_X1 U11043 ( .A1(keyinput78), .A2(keyinput52), .A3(n9930), .ZN(n9934)
         );
  NAND4_X1 U11044 ( .A1(keyinput106), .A2(keyinput20), .A3(keyinput119), .A4(
        keyinput59), .ZN(n9933) );
  NOR2_X1 U11045 ( .A1(keyinput125), .A2(keyinput95), .ZN(n9931) );
  NAND3_X1 U11046 ( .A1(keyinput63), .A2(keyinput32), .A3(n9931), .ZN(n9932)
         );
  NOR4_X1 U11047 ( .A1(n9935), .A2(n9934), .A3(n9933), .A4(n9932), .ZN(n9936)
         );
  NAND4_X1 U11048 ( .A1(n9939), .A2(n9938), .A3(n9937), .A4(n9936), .ZN(n9940)
         );
  NOR4_X1 U11049 ( .A1(n9943), .A2(n9942), .A3(n9941), .A4(n9940), .ZN(n9944)
         );
  NAND4_X1 U11050 ( .A1(n9947), .A2(n9946), .A3(n9945), .A4(n9944), .ZN(n10203) );
  AOI22_X1 U11051 ( .A1(n5810), .A2(keyinput122), .B1(n9949), .B2(keyinput43), 
        .ZN(n9948) );
  OAI221_X1 U11052 ( .B1(n5810), .B2(keyinput122), .C1(n9949), .C2(keyinput43), 
        .A(n9948), .ZN(n9960) );
  AOI22_X1 U11053 ( .A1(n9951), .A2(keyinput111), .B1(n5449), .B2(keyinput8), 
        .ZN(n9950) );
  OAI221_X1 U11054 ( .B1(n9951), .B2(keyinput111), .C1(n5449), .C2(keyinput8), 
        .A(n9950), .ZN(n9959) );
  AOI22_X1 U11055 ( .A1(n9954), .A2(keyinput117), .B1(keyinput52), .B2(n9953), 
        .ZN(n9952) );
  OAI221_X1 U11056 ( .B1(n9954), .B2(keyinput117), .C1(n9953), .C2(keyinput52), 
        .A(n9952), .ZN(n9958) );
  XNOR2_X1 U11057 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput108), .ZN(n9956) );
  XNOR2_X1 U11058 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(keyinput31), .ZN(n9955)
         );
  NAND2_X1 U11059 ( .A1(n9956), .A2(n9955), .ZN(n9957) );
  NOR4_X1 U11060 ( .A1(n9960), .A2(n9959), .A3(n9958), .A4(n9957), .ZN(n10009)
         );
  INV_X1 U11061 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9962) );
  AOI22_X1 U11062 ( .A1(n9962), .A2(keyinput115), .B1(n8055), .B2(keyinput86), 
        .ZN(n9961) );
  OAI221_X1 U11063 ( .B1(n9962), .B2(keyinput115), .C1(n8055), .C2(keyinput86), 
        .A(n9961), .ZN(n9975) );
  AOI22_X1 U11064 ( .A1(n9965), .A2(keyinput75), .B1(keyinput26), .B2(n9964), 
        .ZN(n9963) );
  OAI221_X1 U11065 ( .B1(n9965), .B2(keyinput75), .C1(n9964), .C2(keyinput26), 
        .A(n9963), .ZN(n9974) );
  INV_X1 U11066 ( .A(SI_4_), .ZN(n9968) );
  AOI22_X1 U11067 ( .A1(n9968), .A2(keyinput10), .B1(keyinput68), .B2(n9967), 
        .ZN(n9966) );
  OAI221_X1 U11068 ( .B1(n9968), .B2(keyinput10), .C1(n9967), .C2(keyinput68), 
        .A(n9966), .ZN(n9973) );
  INV_X1 U11069 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9970) );
  AOI22_X1 U11070 ( .A1(n9971), .A2(keyinput79), .B1(keyinput125), .B2(n9970), 
        .ZN(n9969) );
  OAI221_X1 U11071 ( .B1(n9971), .B2(keyinput79), .C1(n9970), .C2(keyinput125), 
        .A(n9969), .ZN(n9972) );
  NOR4_X1 U11072 ( .A1(n9975), .A2(n9974), .A3(n9973), .A4(n9972), .ZN(n10008)
         );
  AOI22_X1 U11073 ( .A1(n9978), .A2(keyinput59), .B1(keyinput94), .B2(n9977), 
        .ZN(n9976) );
  OAI221_X1 U11074 ( .B1(n9978), .B2(keyinput59), .C1(n9977), .C2(keyinput94), 
        .A(n9976), .ZN(n9991) );
  INV_X1 U11075 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9980) );
  AOI22_X1 U11076 ( .A1(n9981), .A2(keyinput20), .B1(keyinput95), .B2(n9980), 
        .ZN(n9979) );
  OAI221_X1 U11077 ( .B1(n9981), .B2(keyinput20), .C1(n9980), .C2(keyinput95), 
        .A(n9979), .ZN(n9990) );
  INV_X1 U11078 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9984) );
  AOI22_X1 U11079 ( .A1(n9984), .A2(keyinput63), .B1(n9983), .B2(keyinput106), 
        .ZN(n9982) );
  OAI221_X1 U11080 ( .B1(n9984), .B2(keyinput63), .C1(n9983), .C2(keyinput106), 
        .A(n9982), .ZN(n9989) );
  XOR2_X1 U11081 ( .A(n9985), .B(keyinput32), .Z(n9987) );
  XNOR2_X1 U11082 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput119), .ZN(n9986) );
  NAND2_X1 U11083 ( .A1(n9987), .A2(n9986), .ZN(n9988) );
  NOR4_X1 U11084 ( .A1(n9991), .A2(n9990), .A3(n9989), .A4(n9988), .ZN(n10007)
         );
  INV_X1 U11085 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9993) );
  AOI22_X1 U11086 ( .A1(n9993), .A2(keyinput53), .B1(keyinput109), .B2(n6455), 
        .ZN(n9992) );
  OAI221_X1 U11087 ( .B1(n9993), .B2(keyinput53), .C1(n6455), .C2(keyinput109), 
        .A(n9992), .ZN(n10005) );
  INV_X1 U11088 ( .A(keyinput69), .ZN(n9995) );
  AOI22_X1 U11089 ( .A1(n9996), .A2(keyinput14), .B1(P2_WR_REG_SCAN_IN), .B2(
        n9995), .ZN(n9994) );
  OAI221_X1 U11090 ( .B1(n9996), .B2(keyinput14), .C1(n9995), .C2(
        P2_WR_REG_SCAN_IN), .A(n9994), .ZN(n10004) );
  AOI22_X1 U11091 ( .A1(n9998), .A2(keyinput49), .B1(keyinput36), .B2(n7334), 
        .ZN(n9997) );
  OAI221_X1 U11092 ( .B1(n9998), .B2(keyinput49), .C1(n7334), .C2(keyinput36), 
        .A(n9997), .ZN(n10003) );
  AOI22_X1 U11093 ( .A1(n10001), .A2(keyinput96), .B1(keyinput87), .B2(n10000), 
        .ZN(n9999) );
  OAI221_X1 U11094 ( .B1(n10001), .B2(keyinput96), .C1(n10000), .C2(keyinput87), .A(n9999), .ZN(n10002) );
  NOR4_X1 U11095 ( .A1(n10005), .A2(n10004), .A3(n10003), .A4(n10002), .ZN(
        n10006) );
  NAND4_X1 U11096 ( .A1(n10009), .A2(n10008), .A3(n10007), .A4(n10006), .ZN(
        n10201) );
  AOI22_X1 U11097 ( .A1(n10012), .A2(keyinput56), .B1(n10011), .B2(keyinput66), 
        .ZN(n10010) );
  OAI221_X1 U11098 ( .B1(n10012), .B2(keyinput56), .C1(n10011), .C2(keyinput66), .A(n10010), .ZN(n10013) );
  INV_X1 U11099 ( .A(n10013), .ZN(n10024) );
  XNOR2_X1 U11100 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput121), .ZN(n10016)
         );
  XNOR2_X1 U11101 ( .A(P1_REG1_REG_16__SCAN_IN), .B(keyinput0), .ZN(n10015) );
  XNOR2_X1 U11102 ( .A(keyinput21), .B(P2_REG2_REG_24__SCAN_IN), .ZN(n10014)
         );
  AND3_X1 U11103 ( .A1(n10016), .A2(n10015), .A3(n10014), .ZN(n10023) );
  INV_X1 U11104 ( .A(keyinput47), .ZN(n10017) );
  XNOR2_X1 U11105 ( .A(n10018), .B(n10017), .ZN(n10022) );
  XNOR2_X1 U11106 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput9), .ZN(n10020) );
  XNOR2_X1 U11107 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput105), .ZN(n10019) );
  AND2_X1 U11108 ( .A1(n10020), .A2(n10019), .ZN(n10021) );
  AND4_X1 U11109 ( .A1(n10024), .A2(n10023), .A3(n10022), .A4(n10021), .ZN(
        n10073) );
  AOI22_X1 U11110 ( .A1(n10027), .A2(keyinput33), .B1(n10026), .B2(keyinput29), 
        .ZN(n10025) );
  OAI221_X1 U11111 ( .B1(n10027), .B2(keyinput33), .C1(n10026), .C2(keyinput29), .A(n10025), .ZN(n10040) );
  AOI22_X1 U11112 ( .A1(n10030), .A2(keyinput2), .B1(n10029), .B2(keyinput89), 
        .ZN(n10028) );
  OAI221_X1 U11113 ( .B1(n10030), .B2(keyinput2), .C1(n10029), .C2(keyinput89), 
        .A(n10028), .ZN(n10039) );
  AOI22_X1 U11114 ( .A1(n10033), .A2(keyinput64), .B1(n10032), .B2(keyinput101), .ZN(n10031) );
  OAI221_X1 U11115 ( .B1(n10033), .B2(keyinput64), .C1(n10032), .C2(
        keyinput101), .A(n10031), .ZN(n10038) );
  AOI22_X1 U11116 ( .A1(n10036), .A2(keyinput50), .B1(n10035), .B2(keyinput30), 
        .ZN(n10034) );
  OAI221_X1 U11117 ( .B1(n10036), .B2(keyinput50), .C1(n10035), .C2(keyinput30), .A(n10034), .ZN(n10037) );
  NOR4_X1 U11118 ( .A1(n10040), .A2(n10039), .A3(n10038), .A4(n10037), .ZN(
        n10072) );
  AOI22_X1 U11119 ( .A1(n10043), .A2(keyinput67), .B1(keyinput11), .B2(n10042), 
        .ZN(n10041) );
  OAI221_X1 U11120 ( .B1(n10043), .B2(keyinput67), .C1(n10042), .C2(keyinput11), .A(n10041), .ZN(n10054) );
  AOI22_X1 U11121 ( .A1(n10046), .A2(keyinput16), .B1(n10045), .B2(keyinput73), 
        .ZN(n10044) );
  OAI221_X1 U11122 ( .B1(n10046), .B2(keyinput16), .C1(n10045), .C2(keyinput73), .A(n10044), .ZN(n10053) );
  INV_X1 U11123 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n10048) );
  AOI22_X1 U11124 ( .A1(n4655), .A2(keyinput71), .B1(keyinput83), .B2(n10048), 
        .ZN(n10047) );
  OAI221_X1 U11125 ( .B1(n4655), .B2(keyinput71), .C1(n10048), .C2(keyinput83), 
        .A(n10047), .ZN(n10052) );
  XNOR2_X1 U11126 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput34), .ZN(n10050) );
  XNOR2_X1 U11127 ( .A(keyinput22), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n10049)
         );
  NAND2_X1 U11128 ( .A1(n10050), .A2(n10049), .ZN(n10051) );
  NOR4_X1 U11129 ( .A1(n10054), .A2(n10053), .A3(n10052), .A4(n10051), .ZN(
        n10071) );
  INV_X1 U11130 ( .A(SI_11_), .ZN(n10057) );
  AOI22_X1 U11131 ( .A1(n10057), .A2(keyinput116), .B1(n10056), .B2(keyinput15), .ZN(n10055) );
  OAI221_X1 U11132 ( .B1(n10057), .B2(keyinput116), .C1(n10056), .C2(
        keyinput15), .A(n10055), .ZN(n10069) );
  AOI22_X1 U11133 ( .A1(n10060), .A2(keyinput107), .B1(keyinput62), .B2(n10059), .ZN(n10058) );
  OAI221_X1 U11134 ( .B1(n10060), .B2(keyinput107), .C1(n10059), .C2(
        keyinput62), .A(n10058), .ZN(n10068) );
  AOI22_X1 U11135 ( .A1(n10063), .A2(keyinput114), .B1(n10062), .B2(
        keyinput118), .ZN(n10061) );
  OAI221_X1 U11136 ( .B1(n10063), .B2(keyinput114), .C1(n10062), .C2(
        keyinput118), .A(n10061), .ZN(n10067) );
  XNOR2_X1 U11137 ( .A(P2_REG0_REG_31__SCAN_IN), .B(keyinput84), .ZN(n10065)
         );
  XNOR2_X1 U11138 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput112), .ZN(n10064) );
  NAND2_X1 U11139 ( .A1(n10065), .A2(n10064), .ZN(n10066) );
  NOR4_X1 U11140 ( .A1(n10069), .A2(n10068), .A3(n10067), .A4(n10066), .ZN(
        n10070) );
  NAND4_X1 U11141 ( .A1(n10073), .A2(n10072), .A3(n10071), .A4(n10070), .ZN(
        n10200) );
  AOI22_X1 U11142 ( .A1(n10076), .A2(keyinput65), .B1(n10075), .B2(keyinput92), 
        .ZN(n10074) );
  OAI221_X1 U11143 ( .B1(n10076), .B2(keyinput65), .C1(n10075), .C2(keyinput92), .A(n10074), .ZN(n10088) );
  INV_X1 U11144 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10078) );
  AOI22_X1 U11145 ( .A1(n10079), .A2(keyinput103), .B1(n10078), .B2(keyinput57), .ZN(n10077) );
  OAI221_X1 U11146 ( .B1(n10079), .B2(keyinput103), .C1(n10078), .C2(
        keyinput57), .A(n10077), .ZN(n10087) );
  AOI22_X1 U11147 ( .A1(n10082), .A2(keyinput76), .B1(n10081), .B2(keyinput13), 
        .ZN(n10080) );
  OAI221_X1 U11148 ( .B1(n10082), .B2(keyinput76), .C1(n10081), .C2(keyinput13), .A(n10080), .ZN(n10086) );
  AOI22_X1 U11149 ( .A1(n10084), .A2(keyinput23), .B1(keyinput18), .B2(n6150), 
        .ZN(n10083) );
  OAI221_X1 U11150 ( .B1(n10084), .B2(keyinput23), .C1(n6150), .C2(keyinput18), 
        .A(n10083), .ZN(n10085) );
  NOR4_X1 U11151 ( .A1(n10088), .A2(n10087), .A3(n10086), .A4(n10085), .ZN(
        n10135) );
  AOI22_X1 U11152 ( .A1(n10091), .A2(keyinput24), .B1(keyinput90), .B2(n10090), 
        .ZN(n10089) );
  OAI221_X1 U11153 ( .B1(n10091), .B2(keyinput24), .C1(n10090), .C2(keyinput90), .A(n10089), .ZN(n10103) );
  AOI22_X1 U11154 ( .A1(n10094), .A2(keyinput102), .B1(keyinput5), .B2(n10093), 
        .ZN(n10092) );
  OAI221_X1 U11155 ( .B1(n10094), .B2(keyinput102), .C1(n10093), .C2(keyinput5), .A(n10092), .ZN(n10102) );
  AOI22_X1 U11156 ( .A1(n5698), .A2(keyinput51), .B1(n10096), .B2(keyinput27), 
        .ZN(n10095) );
  OAI221_X1 U11157 ( .B1(n5698), .B2(keyinput51), .C1(n10096), .C2(keyinput27), 
        .A(n10095), .ZN(n10101) );
  INV_X1 U11158 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n10097) );
  XOR2_X1 U11159 ( .A(n10097), .B(keyinput1), .Z(n10099) );
  XNOR2_X1 U11160 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput42), .ZN(n10098)
         );
  NAND2_X1 U11161 ( .A1(n10099), .A2(n10098), .ZN(n10100) );
  NOR4_X1 U11162 ( .A1(n10103), .A2(n10102), .A3(n10101), .A4(n10100), .ZN(
        n10134) );
  AOI22_X1 U11163 ( .A1(n10106), .A2(keyinput3), .B1(n10105), .B2(keyinput91), 
        .ZN(n10104) );
  OAI221_X1 U11164 ( .B1(n10106), .B2(keyinput3), .C1(n10105), .C2(keyinput91), 
        .A(n10104), .ZN(n10119) );
  AOI22_X1 U11165 ( .A1(n10109), .A2(keyinput124), .B1(keyinput41), .B2(n10108), .ZN(n10107) );
  OAI221_X1 U11166 ( .B1(n10109), .B2(keyinput124), .C1(n10108), .C2(
        keyinput41), .A(n10107), .ZN(n10118) );
  AOI22_X1 U11167 ( .A1(n10112), .A2(keyinput88), .B1(n10111), .B2(keyinput46), 
        .ZN(n10110) );
  OAI221_X1 U11168 ( .B1(n10112), .B2(keyinput88), .C1(n10111), .C2(keyinput46), .A(n10110), .ZN(n10117) );
  XOR2_X1 U11169 ( .A(n10113), .B(keyinput78), .Z(n10115) );
  XNOR2_X1 U11170 ( .A(SI_2_), .B(keyinput48), .ZN(n10114) );
  NAND2_X1 U11171 ( .A1(n10115), .A2(n10114), .ZN(n10116) );
  NOR4_X1 U11172 ( .A1(n10119), .A2(n10118), .A3(n10117), .A4(n10116), .ZN(
        n10133) );
  INV_X1 U11173 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n10121) );
  AOI22_X1 U11174 ( .A1(n10121), .A2(keyinput74), .B1(n5750), .B2(keyinput72), 
        .ZN(n10120) );
  OAI221_X1 U11175 ( .B1(n10121), .B2(keyinput74), .C1(n5750), .C2(keyinput72), 
        .A(n10120), .ZN(n10126) );
  XNOR2_X1 U11176 ( .A(n10122), .B(keyinput110), .ZN(n10125) );
  XNOR2_X1 U11177 ( .A(n10123), .B(keyinput97), .ZN(n10124) );
  OR3_X1 U11178 ( .A1(n10126), .A2(n10125), .A3(n10124), .ZN(n10131) );
  INV_X1 U11179 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10207) );
  AOI22_X1 U11180 ( .A1(n5729), .A2(keyinput45), .B1(keyinput100), .B2(n10207), 
        .ZN(n10127) );
  OAI221_X1 U11181 ( .B1(n5729), .B2(keyinput45), .C1(n10207), .C2(keyinput100), .A(n10127), .ZN(n10130) );
  AOI22_X1 U11182 ( .A1(n7457), .A2(keyinput126), .B1(keyinput25), .B2(n5674), 
        .ZN(n10128) );
  OAI221_X1 U11183 ( .B1(n7457), .B2(keyinput126), .C1(n5674), .C2(keyinput25), 
        .A(n10128), .ZN(n10129) );
  NOR3_X1 U11184 ( .A1(n10131), .A2(n10130), .A3(n10129), .ZN(n10132) );
  NAND4_X1 U11185 ( .A1(n10135), .A2(n10134), .A3(n10133), .A4(n10132), .ZN(
        n10199) );
  AOI22_X1 U11186 ( .A1(n10138), .A2(keyinput37), .B1(n10137), .B2(keyinput60), 
        .ZN(n10136) );
  OAI221_X1 U11187 ( .B1(n10138), .B2(keyinput37), .C1(n10137), .C2(keyinput60), .A(n10136), .ZN(n10151) );
  AOI22_X1 U11188 ( .A1(n10141), .A2(keyinput35), .B1(n10140), .B2(keyinput61), 
        .ZN(n10139) );
  OAI221_X1 U11189 ( .B1(n10141), .B2(keyinput35), .C1(n10140), .C2(keyinput61), .A(n10139), .ZN(n10150) );
  AOI22_X1 U11190 ( .A1(n10144), .A2(keyinput98), .B1(keyinput58), .B2(n10143), 
        .ZN(n10142) );
  OAI221_X1 U11191 ( .B1(n10144), .B2(keyinput98), .C1(n10143), .C2(keyinput58), .A(n10142), .ZN(n10149) );
  INV_X1 U11192 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n10147) );
  AOI22_X1 U11193 ( .A1(n10147), .A2(keyinput40), .B1(n10146), .B2(keyinput127), .ZN(n10145) );
  OAI221_X1 U11194 ( .B1(n10147), .B2(keyinput40), .C1(n10146), .C2(
        keyinput127), .A(n10145), .ZN(n10148) );
  NOR4_X1 U11195 ( .A1(n10151), .A2(n10150), .A3(n10149), .A4(n10148), .ZN(
        n10197) );
  INV_X1 U11196 ( .A(SI_1_), .ZN(n10153) );
  AOI22_X1 U11197 ( .A1(n10154), .A2(keyinput39), .B1(keyinput55), .B2(n10153), 
        .ZN(n10152) );
  OAI221_X1 U11198 ( .B1(n10154), .B2(keyinput39), .C1(n10153), .C2(keyinput55), .A(n10152), .ZN(n10165) );
  INV_X1 U11199 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10156) );
  AOI22_X1 U11200 ( .A1(n5992), .A2(keyinput113), .B1(n10156), .B2(keyinput120), .ZN(n10155) );
  OAI221_X1 U11201 ( .B1(n5992), .B2(keyinput113), .C1(n10156), .C2(
        keyinput120), .A(n10155), .ZN(n10164) );
  AOI22_X1 U11202 ( .A1(keyinput28), .A2(n10158), .B1(keyinput93), .B2(n10204), 
        .ZN(n10157) );
  OAI21_X1 U11203 ( .B1(n10158), .B2(keyinput28), .A(n10157), .ZN(n10163) );
  INV_X1 U11204 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n10159) );
  XOR2_X1 U11205 ( .A(n10159), .B(keyinput104), .Z(n10161) );
  XNOR2_X1 U11206 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput4), .ZN(n10160) );
  NAND2_X1 U11207 ( .A1(n10161), .A2(n10160), .ZN(n10162) );
  NOR4_X1 U11208 ( .A1(n10165), .A2(n10164), .A3(n10163), .A4(n10162), .ZN(
        n10196) );
  AOI22_X1 U11209 ( .A1(n10168), .A2(keyinput54), .B1(n10167), .B2(keyinput12), 
        .ZN(n10166) );
  OAI221_X1 U11210 ( .B1(n10168), .B2(keyinput54), .C1(n10167), .C2(keyinput12), .A(n10166), .ZN(n10179) );
  INV_X1 U11211 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U11212 ( .A1(n10171), .A2(keyinput44), .B1(keyinput77), .B2(n10170), 
        .ZN(n10169) );
  OAI221_X1 U11213 ( .B1(n10171), .B2(keyinput44), .C1(n10170), .C2(keyinput77), .A(n10169), .ZN(n10178) );
  AOI22_X1 U11214 ( .A1(n6221), .A2(keyinput80), .B1(keyinput82), .B2(n5855), 
        .ZN(n10172) );
  OAI221_X1 U11215 ( .B1(n6221), .B2(keyinput80), .C1(n5855), .C2(keyinput82), 
        .A(n10172), .ZN(n10177) );
  AOI22_X1 U11216 ( .A1(n10175), .A2(keyinput85), .B1(n10174), .B2(keyinput70), 
        .ZN(n10173) );
  OAI221_X1 U11217 ( .B1(n10175), .B2(keyinput85), .C1(n10174), .C2(keyinput70), .A(n10173), .ZN(n10176) );
  NOR4_X1 U11218 ( .A1(n10179), .A2(n10178), .A3(n10177), .A4(n10176), .ZN(
        n10195) );
  INV_X1 U11219 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U11220 ( .A1(n10212), .A2(keyinput38), .B1(n10181), .B2(keyinput81), 
        .ZN(n10180) );
  OAI221_X1 U11221 ( .B1(n10212), .B2(keyinput38), .C1(n10181), .C2(keyinput81), .A(n10180), .ZN(n10193) );
  AOI22_X1 U11222 ( .A1(n10183), .A2(keyinput19), .B1(n5745), .B2(keyinput17), 
        .ZN(n10182) );
  OAI221_X1 U11223 ( .B1(n10183), .B2(keyinput19), .C1(n5745), .C2(keyinput17), 
        .A(n10182), .ZN(n10192) );
  INV_X1 U11224 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10186) );
  AOI22_X1 U11225 ( .A1(n10186), .A2(keyinput123), .B1(n10185), .B2(keyinput6), 
        .ZN(n10184) );
  OAI221_X1 U11226 ( .B1(n10186), .B2(keyinput123), .C1(n10185), .C2(keyinput6), .A(n10184), .ZN(n10191) );
  AOI22_X1 U11227 ( .A1(n10189), .A2(keyinput7), .B1(n10188), .B2(keyinput99), 
        .ZN(n10187) );
  OAI221_X1 U11228 ( .B1(n10189), .B2(keyinput7), .C1(n10188), .C2(keyinput99), 
        .A(n10187), .ZN(n10190) );
  NOR4_X1 U11229 ( .A1(n10193), .A2(n10192), .A3(n10191), .A4(n10190), .ZN(
        n10194) );
  NAND4_X1 U11230 ( .A1(n10197), .A2(n10196), .A3(n10195), .A4(n10194), .ZN(
        n10198) );
  NOR4_X1 U11231 ( .A1(n10201), .A2(n10200), .A3(n10199), .A4(n10198), .ZN(
        n10202) );
  OAI221_X1 U11232 ( .B1(keyinput93), .B2(n10204), .C1(keyinput93), .C2(n10203), .A(n10202), .ZN(n10205) );
  XNOR2_X1 U11233 ( .A(n10206), .B(n10205), .ZN(P2_U3252) );
  XNOR2_X1 U11234 ( .A(n10208), .B(n10207), .ZN(ADD_1071_U49) );
  AOI21_X1 U11235 ( .B1(n10211), .B2(n10210), .A(n10209), .ZN(ADD_1071_U47) );
  XNOR2_X1 U11236 ( .A(n10213), .B(n10212), .ZN(ADD_1071_U50) );
  NOR2_X1 U11237 ( .A1(n10215), .A2(n10214), .ZN(n10216) );
  XOR2_X1 U11238 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10216), .Z(ADD_1071_U51) );
  OAI21_X1 U11239 ( .B1(n10219), .B2(n10218), .A(n10217), .ZN(n10220) );
  XNOR2_X1 U11240 ( .A(n10220), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11241 ( .A(n10222), .B(n10221), .Z(ADD_1071_U54) );
  XOR2_X1 U11242 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10223), .Z(ADD_1071_U48) );
  XOR2_X1 U11243 ( .A(n10225), .B(n10224), .Z(ADD_1071_U53) );
  XNOR2_X1 U11244 ( .A(n10227), .B(n10226), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4924 ( .A(n7370), .Z(n4417) );
  CLKBUF_X1 U4925 ( .A(n6077), .Z(n7995) );
  CLKBUF_X1 U4928 ( .A(n5200), .Z(n5569) );
  CLKBUF_X1 U4929 ( .A(n5212), .Z(n4422) );
  CLKBUF_X1 U4930 ( .A(n5222), .Z(n5314) );
  CLKBUF_X1 U4935 ( .A(n5212), .Z(n4423) );
  INV_X2 U4968 ( .A(n10230), .ZN(n4414) );
  NAND2_X1 U4969 ( .A1(n8229), .A2(n5773), .ZN(n10230) );
endmodule

