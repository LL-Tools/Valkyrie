

module b20_C_SARLock_k_128_9 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297;

  OAI21_X1 U4922 ( .B1(n8157), .B2(n4991), .A(n4989), .ZN(n4992) );
  INV_X4 U4923 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OR2_X1 U4924 ( .A1(n5526), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U4925 ( .A1(n6196), .A2(n6195), .ZN(n8711) );
  CLKBUF_X2 U4926 ( .A(n6035), .Z(n4418) );
  CLKBUF_X2 U4927 ( .A(n5278), .Z(n5620) );
  INV_X2 U4928 ( .A(n6070), .ZN(n6516) );
  BUF_X1 U4929 ( .A(n4674), .Z(n4673) );
  XNOR2_X1 U4930 ( .A(n5986), .B(n5985), .ZN(n7768) );
  INV_X1 U4931 ( .A(n5666), .ZN(n5941) );
  NOR2_X1 U4932 ( .A1(n7147), .A2(n7241), .ZN(n7244) );
  OR2_X1 U4933 ( .A1(n5501), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U4934 ( .A1(n4641), .A2(n4640), .ZN(n5657) );
  OR2_X1 U4935 ( .A1(n5223), .A2(n5190), .ZN(n4672) );
  INV_X1 U4936 ( .A(n6476), .ZN(n7931) );
  INV_X1 U4937 ( .A(n6035), .ZN(n7927) );
  OR2_X1 U4938 ( .A1(n5589), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5600) );
  INV_X1 U4939 ( .A(n5291), .ZN(n5616) );
  NAND2_X1 U4940 ( .A1(n5900), .A2(n8439), .ZN(n8426) );
  INV_X1 U4941 ( .A(n8011), .ZN(n9888) );
  INV_X1 U4942 ( .A(n9062), .ZN(n4420) );
  NOR2_X1 U4943 ( .A1(n7232), .A2(n7480), .ZN(n7606) );
  INV_X1 U4944 ( .A(n6982), .ZN(n9756) );
  AOI21_X1 U4945 ( .B1(n9920), .B2(n8569), .A(n8568), .ZN(n8632) );
  AND4_X1 U4946 ( .A1(n6046), .A2(n6045), .A3(n6044), .A4(n6043), .ZN(n6979)
         );
  INV_X1 U4947 ( .A(n7973), .ZN(n8369) );
  NAND2_X1 U4948 ( .A1(n6479), .A2(n6478), .ZN(n7946) );
  AOI211_X1 U4949 ( .C1(n9482), .C2(n9724), .A(n7922), .B(n7921), .ZN(n7923)
         );
  AOI21_X2 U4950 ( .B1(n4894), .B2(n9715), .A(n4891), .ZN(n9485) );
  NAND2_X1 U4952 ( .A1(n7140), .A2(n5855), .ZN(n4415) );
  NAND2_X2 U4953 ( .A1(n7140), .A2(n5855), .ZN(n5261) );
  NAND2_X1 U4954 ( .A1(n5229), .A2(n5228), .ZN(n4416) );
  NAND2_X2 U4955 ( .A1(n5229), .A2(n5228), .ZN(n5291) );
  OR2_X1 U4956 ( .A1(n4430), .A2(n6578), .ZN(n5290) );
  NAND2_X2 U4957 ( .A1(n8426), .A2(n5901), .ZN(n8415) );
  AOI21_X2 U4958 ( .B1(n9333), .B2(n9339), .A(n7886), .ZN(n9317) );
  AOI21_X2 U4959 ( .B1(n7877), .B2(n9033), .A(n7876), .ZN(n9456) );
  NAND2_X2 U4960 ( .A1(n7748), .A2(n7747), .ZN(n7877) );
  BUF_X2 U4961 ( .A(n7202), .Z(n4417) );
  XNOR2_X1 U4962 ( .A(n5272), .B(n5271), .ZN(n7202) );
  INV_X2 U4963 ( .A(n6041), .ZN(n6275) );
  OAI21_X2 U4964 ( .B1(n6531), .B2(n9922), .A(n6530), .ZN(n6553) );
  OR2_X1 U4965 ( .A1(n8204), .A2(n9882), .ZN(n5664) );
  AND3_X2 U4966 ( .A1(n5275), .A2(n5274), .A3(n5273), .ZN(n9882) );
  OAI21_X2 U4967 ( .B1(n7819), .B2(n4998), .A(n4994), .ZN(n8111) );
  AOI22_X4 U4968 ( .A1(n7703), .A2(n7702), .B1(n8198), .B2(n7701), .ZN(n7819)
         );
  AOI21_X2 U4969 ( .B1(n5919), .B2(n8494), .A(n5918), .ZN(n6530) );
  XNOR2_X2 U4970 ( .A(n6101), .B(n6100), .ZN(n7310) );
  NAND2_X2 U4971 ( .A1(n6939), .A2(n6087), .ZN(n6101) );
  NAND2_X2 U4972 ( .A1(n4545), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5971) );
  NAND3_X1 U4973 ( .A1(n7494), .A2(n6572), .A3(n6001), .ZN(n6035) );
  OAI21_X2 U4974 ( .B1(n7650), .B2(n7651), .A(n5698), .ZN(n7677) );
  OAI21_X2 U4975 ( .B1(n7585), .B2(n7586), .A(n5684), .ZN(n7650) );
  NAND2_X2 U4976 ( .A1(n6221), .A2(n6220), .ZN(n8738) );
  AOI21_X2 U4977 ( .B1(n6880), .B2(n6917), .A(n6878), .ZN(n6885) );
  AND2_X1 U4978 ( .A1(n8419), .A2(n5800), .ZN(n8410) );
  CLKBUF_X1 U4979 ( .A(n8444), .Z(n8458) );
  NAND2_X1 U4980 ( .A1(n5886), .A2(n5885), .ZN(n8542) );
  AOI21_X1 U4981 ( .B1(n4789), .B2(n4791), .A(n4421), .ZN(n4786) );
  INV_X1 U4982 ( .A(n7820), .ZN(n4421) );
  NAND2_X1 U4983 ( .A1(n5704), .A2(n5705), .ZN(n7820) );
  NAND2_X1 U4984 ( .A1(n9073), .A2(n9552), .ZN(n9028) );
  INV_X1 U4985 ( .A(n7692), .ZN(n9905) );
  NAND2_X1 U4986 ( .A1(n5867), .A2(n5866), .ZN(n7301) );
  OR2_X1 U4987 ( .A1(n5442), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5456) );
  INV_X2 U4988 ( .A(n9471), .ZN(n4419) );
  NAND2_X1 U4989 ( .A1(n6978), .A2(n9061), .ZN(n9720) );
  OAI22_X1 U4990 ( .A1(n6979), .A2(n6320), .B1(n9756), .B2(n4521), .ZN(n6050)
         );
  AND4_X1 U4991 ( .A1(n6056), .A2(n6055), .A3(n6054), .A4(n6053), .ZN(n6997)
         );
  AND2_X1 U4992 ( .A1(n5242), .A2(n5241), .ZN(n5245) );
  CLKBUF_X2 U4993 ( .A(n9147), .Z(P1_U3973) );
  INV_X1 U4994 ( .A(n6987), .ZN(n9800) );
  OR2_X1 U4995 ( .A1(n4416), .A2(n9817), .ZN(n5243) );
  INV_X1 U4996 ( .A(n6572), .ZN(n6022) );
  CLKBUF_X2 U4997 ( .A(n5252), .Z(n5486) );
  AND2_X1 U4998 ( .A1(n7963), .A2(n5229), .ZN(n5253) );
  INV_X4 U4999 ( .A(n7135), .ZN(n8334) );
  MUX2_X1 U5000 ( .A(n6563), .B(n6566), .S(n9941), .Z(n6565) );
  AOI21_X1 U5001 ( .B1(n8370), .B2(n8494), .A(n4512), .ZN(n8564) );
  NOR2_X1 U5002 ( .A1(n4519), .A2(n4470), .ZN(n4518) );
  NAND2_X1 U5003 ( .A1(n4553), .A2(n4552), .ZN(n4551) );
  OAI22_X1 U5004 ( .A1(n6558), .A2(n5908), .B1(n7873), .B2(n8369), .ZN(n5909)
         );
  OAI21_X1 U5005 ( .B1(n4510), .B2(n9869), .A(n4508), .ZN(n8565) );
  NOR3_X1 U5006 ( .A1(n5955), .A2(n5954), .A3(n5036), .ZN(n5956) );
  NAND2_X1 U5007 ( .A1(n6440), .A2(n6439), .ZN(n8741) );
  XNOR2_X1 U5008 ( .A(n8691), .B(n8693), .ZN(n8811) );
  NAND2_X1 U5009 ( .A1(n4900), .A2(n6387), .ZN(n8691) );
  OR2_X1 U5010 ( .A1(n7891), .A2(n4972), .ZN(n4971) );
  INV_X1 U5011 ( .A(n9224), .ZN(n9565) );
  OAI21_X1 U5012 ( .B1(n8410), .B2(n4664), .A(n4662), .ZN(n8372) );
  OAI21_X1 U5013 ( .B1(n8410), .B2(n5766), .A(n5825), .ZN(n8395) );
  XNOR2_X1 U5014 ( .A(n5175), .B(n5174), .ZN(n9609) );
  NAND2_X1 U5015 ( .A1(n4649), .A2(n4648), .ZN(n8440) );
  INV_X1 U5016 ( .A(n5828), .ZN(n8379) );
  OR2_X1 U5017 ( .A1(n9389), .A2(n9390), .ZN(n9387) );
  NAND2_X1 U5018 ( .A1(n8527), .A2(n8532), .ZN(n4801) );
  NOR2_X1 U5019 ( .A1(n4493), .A2(n7884), .ZN(n4976) );
  NAND2_X1 U5020 ( .A1(n4878), .A2(n4877), .ZN(n7909) );
  AND2_X1 U5021 ( .A1(n8912), .A2(n8910), .ZN(n9551) );
  NAND2_X1 U5022 ( .A1(n5412), .A2(n5411), .ZN(n9926) );
  INV_X2 U5023 ( .A(n9696), .ZN(n4422) );
  XNOR2_X1 U5024 ( .A(n5408), .B(n5407), .ZN(n6618) );
  NAND2_X1 U5025 ( .A1(n6164), .A2(n6163), .ZN(n7627) );
  AND2_X1 U5026 ( .A1(n5693), .A2(n7464), .ZN(n7434) );
  NAND2_X1 U5027 ( .A1(n4844), .A2(n4458), .ZN(n9842) );
  OR2_X1 U5028 ( .A1(n7271), .A2(n4845), .ZN(n4844) );
  AND3_X1 U5029 ( .A1(n4826), .A2(n4487), .A3(n4825), .ZN(n7356) );
  NOR2_X1 U5030 ( .A1(n5953), .A2(n9858), .ZN(n8524) );
  XNOR2_X1 U5031 ( .A(n6034), .B(n4428), .ZN(n6036) );
  OR2_X1 U5032 ( .A1(n7167), .A2(n7136), .ZN(n7253) );
  NAND2_X2 U5033 ( .A1(n6926), .A2(n9701), .ZN(n9471) );
  INV_X1 U5034 ( .A(n7244), .ZN(n4423) );
  CLKBUF_X2 U5035 ( .A(n6476), .Z(n4521) );
  NAND2_X1 U5036 ( .A1(n9756), .A2(n9146), .ZN(n9061) );
  AND3_X2 U5037 ( .A1(n6808), .A2(n6925), .A3(n6923), .ZN(n9788) );
  INV_X2 U5038 ( .A(n6207), .ZN(n6136) );
  NAND2_X1 U5039 ( .A1(n7166), .A2(n7165), .ZN(n7251) );
  NAND3_X1 U5040 ( .A1(n5258), .A2(n5257), .A3(n5256), .ZN(n7012) );
  NAND4_X1 U5041 ( .A1(n5298), .A2(n5297), .A3(n5295), .A4(n5296), .ZN(n8202)
         );
  NAND2_X1 U5042 ( .A1(n5924), .A2(n4452), .ZN(n5008) );
  NAND2_X1 U5043 ( .A1(n4679), .A2(n4444), .ZN(n6964) );
  NAND4_X1 U5044 ( .A1(n5312), .A2(n5311), .A3(n5310), .A4(n5309), .ZN(n8201)
         );
  NAND2_X1 U5045 ( .A1(n5999), .A2(n9125), .ZN(n6207) );
  NAND3_X2 U5046 ( .A1(n5245), .A2(n5244), .A3(n5243), .ZN(n5860) );
  NOR2_X1 U5047 ( .A1(n6022), .A2(n9121), .ZN(n5999) );
  NAND4_X2 U5048 ( .A1(n5268), .A2(n5267), .A3(n5266), .A4(n5265), .ZN(n8204)
         );
  NAND2_X1 U5049 ( .A1(n4682), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4592) );
  XNOR2_X1 U5050 ( .A(n5643), .B(n5642), .ZN(n7334) );
  CLKBUF_X2 U5051 ( .A(n5253), .Z(n4426) );
  AND2_X1 U5052 ( .A1(n7035), .A2(n4550), .ZN(n9121) );
  OR2_X1 U5053 ( .A1(n9843), .A2(n5337), .ZN(n4845) );
  CLKBUF_X2 U5054 ( .A(n6008), .Z(n7924) );
  NOR2_X1 U5055 ( .A1(n7768), .A2(n7684), .ZN(n5991) );
  INV_X1 U5056 ( .A(n9054), .ZN(n7035) );
  CLKBUF_X1 U5057 ( .A(n9054), .Z(n4539) );
  XNOR2_X1 U5058 ( .A(n5977), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9054) );
  NAND2_X1 U5059 ( .A1(n5998), .A2(n5997), .ZN(n7279) );
  XNOR2_X1 U5060 ( .A(n6004), .B(n9603), .ZN(n6008) );
  INV_X1 U5061 ( .A(n6011), .ZN(n6012) );
  XNOR2_X1 U5062 ( .A(n5224), .B(n8670), .ZN(n7963) );
  NAND2_X1 U5063 ( .A1(n5990), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U5064 ( .A1(n8669), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U5065 ( .A1(n9606), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6004) );
  XNOR2_X1 U5066 ( .A(n5193), .B(n5192), .ZN(n7140) );
  INV_X1 U5067 ( .A(n9050), .ZN(n4550) );
  NAND2_X1 U5068 ( .A1(n5976), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5977) );
  INV_X2 U5069 ( .A(n9608), .ZN(n7925) );
  INV_X2 U5070 ( .A(n4503), .ZN(n7962) );
  OAI21_X1 U5071 ( .B1(n5247), .B2(n5246), .A(n5042), .ZN(n5270) );
  NOR2_X1 U5072 ( .A1(n5191), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5223) );
  AND2_X1 U5073 ( .A1(n4676), .A2(n5018), .ZN(n5189) );
  BUF_X2 U5074 ( .A(n5259), .Z(n4632) );
  AND4_X1 U5075 ( .A1(n5002), .A2(n5188), .A3(n4677), .A4(n5313), .ZN(n4675)
         );
  OAI21_X1 U5076 ( .B1(n5194), .B2(n5039), .A(n5038), .ZN(n5041) );
  AND2_X1 U5077 ( .A1(n5021), .A2(n5178), .ZN(n5018) );
  AND2_X1 U5078 ( .A1(n4939), .A2(n4938), .ZN(n4937) );
  AND2_X1 U5079 ( .A1(n5031), .A2(n5979), .ZN(n4983) );
  NOR2_X1 U5080 ( .A1(n5183), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5021) );
  AND2_X1 U5081 ( .A1(n5187), .A2(n5373), .ZN(n4677) );
  NAND2_X1 U5082 ( .A1(n5010), .A2(n4674), .ZN(n5299) );
  AND2_X1 U5083 ( .A1(n4448), .A2(n5177), .ZN(n5004) );
  AND2_X1 U5084 ( .A1(n4941), .A2(n4940), .ZN(n4939) );
  NAND2_X2 U5085 ( .A1(n4761), .A2(n4759), .ZN(n5194) );
  AND2_X1 U5086 ( .A1(n5271), .A2(n5176), .ZN(n5010) );
  AND4_X1 U5087 ( .A1(n5992), .A2(n5965), .A3(n5964), .A4(n5963), .ZN(n5031)
         );
  AND2_X1 U5088 ( .A1(n5973), .A2(n10189), .ZN(n4941) );
  NAND3_X1 U5089 ( .A1(n4760), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4759) );
  AND2_X1 U5090 ( .A1(n4785), .A2(n4784), .ZN(n4674) );
  NAND3_X1 U5091 ( .A1(n4764), .A2(n4763), .A3(n4762), .ZN(n4761) );
  INV_X1 U5092 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4762) );
  INV_X1 U5093 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4760) );
  NOR2_X1 U5094 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5958) );
  INV_X2 U5095 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5271) );
  NOR2_X1 U5096 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5992) );
  NOR2_X1 U5097 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4946) );
  INV_X4 U5098 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5099 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6179) );
  INV_X1 U5100 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4763) );
  NAND2_X1 U5101 ( .A1(n4805), .A2(n4804), .ZN(n5886) );
  AND2_X4 U5102 ( .A1(n6115), .A2(n5962), .ZN(n5972) );
  AND2_X2 U5103 ( .A1(n6207), .A2(n4427), .ZN(n6476) );
  AOI22_X1 U5104 ( .A1(n9317), .A2(n7887), .B1(n8947), .B2(n9330), .ZN(n9302)
         );
  OAI222_X1 U5105 ( .A1(n9616), .A2(n9615), .B1(P1_U3086), .B2(n9651), .C1(
        n7925), .C2(n9613), .ZN(P1_U3328) );
  OR2_X4 U5106 ( .A1(n9125), .A2(n6022), .ZN(n6062) );
  INV_X1 U5107 ( .A(n5252), .ZN(n4425) );
  INV_X1 U5108 ( .A(n5252), .ZN(n4511) );
  OR2_X4 U5109 ( .A1(n5229), .A2(n7963), .ZN(n5252) );
  INV_X2 U5110 ( .A(n5860), .ZN(n4640) );
  NOR2_X2 U5111 ( .A1(n6907), .A2(n6906), .ZN(n8009) );
  NOR2_X2 U5112 ( .A1(n6905), .A2(n6904), .ZN(n6907) );
  BUF_X4 U5113 ( .A(n6062), .Z(n6320) );
  NOR3_X2 U5114 ( .A1(n5786), .A2(n5785), .A3(n5944), .ZN(n5791) );
  AOI21_X2 U5115 ( .B1(n5782), .B2(n5781), .A(n5780), .ZN(n5786) );
  INV_X4 U5117 ( .A(n6275), .ZN(n8870) );
  NOR2_X4 U5118 ( .A1(n7547), .A2(n8711), .ZN(n7669) );
  NAND2_X2 U5119 ( .A1(n8387), .A2(n8394), .ZN(n8386) );
  AOI22_X2 U5120 ( .A1(n8400), .A2(n5904), .B1(n8638), .B2(n8388), .ZN(n8387)
         );
  OAI21_X4 U5121 ( .B1(n7467), .B2(n5877), .A(n5876), .ZN(n7583) );
  OAI21_X2 U5122 ( .B1(n7433), .B2(n5874), .A(n5875), .ZN(n7467) );
  NAND3_X1 U5123 ( .A1(n7494), .A2(n6572), .A3(n6001), .ZN(n4427) );
  NAND2_X1 U5124 ( .A1(n6724), .A2(n6723), .ZN(n6722) );
  INV_X1 U5125 ( .A(n6136), .ZN(n4428) );
  INV_X2 U5126 ( .A(n6136), .ZN(n4429) );
  CLKBUF_X1 U5127 ( .A(n5285), .Z(n4430) );
  CLKBUF_X3 U5128 ( .A(n5285), .Z(n4431) );
  NAND2_X1 U5129 ( .A1(n4415), .A2(n4633), .ZN(n5285) );
  OAI22_X2 U5130 ( .A1(n7301), .A2(n5868), .B1(n9864), .B2(n9888), .ZN(n7053)
         );
  AOI21_X2 U5131 ( .B1(n8704), .B2(n6216), .A(n6215), .ZN(n8732) );
  OAI21_X2 U5132 ( .B1(n8780), .B2(n8776), .A(n8777), .ZN(n8704) );
  XNOR2_X2 U5133 ( .A(n4672), .B(n5222), .ZN(n5855) );
  NAND2_X1 U5134 ( .A1(n5084), .A2(n5083), .ZN(n5087) );
  AOI21_X1 U5135 ( .B1(n5535), .B2(n4752), .A(n4749), .ZN(n4748) );
  NAND2_X1 U5136 ( .A1(n4750), .A2(n5136), .ZN(n4749) );
  NAND2_X1 U5137 ( .A1(n4752), .A2(n4754), .ZN(n4750) );
  NAND2_X1 U5138 ( .A1(n5120), .A2(n5119), .ZN(n5523) );
  NAND2_X1 U5139 ( .A1(n7201), .A2(n7200), .ZN(n7199) );
  NAND2_X1 U5140 ( .A1(n5683), .A2(n5682), .ZN(n4611) );
  NAND2_X1 U5141 ( .A1(n4634), .A2(n5750), .ZN(n5759) );
  OR2_X1 U5142 ( .A1(n9279), .A2(n9256), .ZN(n8987) );
  NAND2_X1 U5143 ( .A1(n9279), .A2(n9256), .ZN(n9000) );
  AND2_X1 U5144 ( .A1(n4737), .A2(n5492), .ZN(n4736) );
  INV_X1 U5145 ( .A(n5448), .ZN(n5099) );
  NOR2_X1 U5146 ( .A1(n7816), .A2(n7817), .ZN(n4996) );
  NAND2_X1 U5147 ( .A1(n4840), .A2(n4447), .ZN(n4841) );
  INV_X1 U5148 ( .A(n7361), .ZN(n4840) );
  NAND2_X1 U5149 ( .A1(n4437), .A2(n4461), .ZN(n4798) );
  OR2_X1 U5150 ( .A1(n8051), .A2(n8402), .ZN(n5771) );
  NAND2_X1 U5151 ( .A1(n8051), .A2(n8402), .ZN(n5772) );
  OR2_X1 U5152 ( .A1(n8094), .A2(n8450), .ZN(n5804) );
  OR2_X1 U5153 ( .A1(n8660), .A2(n8514), .ZN(n5737) );
  OR2_X1 U5154 ( .A1(n8197), .A2(n7618), .ZN(n5697) );
  NOR2_X1 U5155 ( .A1(n7334), .A2(n7484), .ZN(n5666) );
  NAND2_X1 U5156 ( .A1(n5191), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U5157 ( .A1(n4562), .A2(n8970), .ZN(n4561) );
  AND2_X1 U5158 ( .A1(n9223), .A2(n8976), .ZN(n8972) );
  INV_X1 U5159 ( .A(n4549), .ZN(n4548) );
  OAI21_X1 U5160 ( .B1(n4551), .B2(n4554), .A(n4550), .ZN(n4549) );
  AOI21_X1 U5161 ( .B1(n4548), .B2(n4551), .A(n9062), .ZN(n4546) );
  NAND2_X1 U5162 ( .A1(n9068), .A2(n9027), .ZN(n9072) );
  NAND2_X1 U5163 ( .A1(n4577), .A2(n9063), .ZN(n4576) );
  NAND3_X1 U5164 ( .A1(n5627), .A2(n4778), .A3(n8877), .ZN(n4776) );
  AND2_X1 U5165 ( .A1(n5141), .A2(n5140), .ZN(n5566) );
  INV_X1 U5166 ( .A(n5476), .ZN(n4742) );
  NOR2_X1 U5167 ( .A1(n4747), .A2(n5103), .ZN(n4746) );
  NOR2_X1 U5168 ( .A1(n5102), .A2(SI_16_), .ZN(n5103) );
  INV_X1 U5169 ( .A(n5100), .ZN(n4747) );
  NAND2_X1 U5170 ( .A1(n5097), .A2(n5096), .ZN(n5450) );
  INV_X1 U5171 ( .A(n5435), .ZN(n5094) );
  INV_X1 U5172 ( .A(n5081), .ZN(n4723) );
  XNOR2_X1 U5173 ( .A(n5079), .B(SI_10_), .ZN(n5391) );
  NAND2_X1 U5174 ( .A1(n5066), .A2(n4630), .ZN(n4629) );
  NOR2_X1 U5175 ( .A1(n5357), .A2(n4631), .ZN(n4630) );
  INV_X1 U5176 ( .A(n5065), .ZN(n4631) );
  NAND2_X1 U5177 ( .A1(n5068), .A2(n5067), .ZN(n5071) );
  NAND2_X1 U5178 ( .A1(n7688), .A2(n7687), .ZN(n4986) );
  NAND2_X1 U5179 ( .A1(n8056), .A2(n7862), .ZN(n8157) );
  OR2_X1 U5180 ( .A1(n6554), .A2(n7871), .ZN(n5784) );
  BUF_X1 U5181 ( .A(n4426), .Z(n5617) );
  INV_X1 U5182 ( .A(n4426), .ZN(n5602) );
  NAND2_X1 U5183 ( .A1(n7199), .A2(n4859), .ZN(n4858) );
  NOR2_X1 U5184 ( .A1(n4860), .A2(n7287), .ZN(n4859) );
  NAND2_X1 U5185 ( .A1(n4832), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4829) );
  INV_X1 U5186 ( .A(n8214), .ZN(n4832) );
  OAI21_X1 U5187 ( .B1(n8244), .B2(n4871), .A(n4870), .ZN(n8279) );
  NAND2_X1 U5188 ( .A1(n4875), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4871) );
  NAND2_X1 U5189 ( .A1(n4876), .A2(n4875), .ZN(n4870) );
  INV_X1 U5190 ( .A(n8262), .ZN(n4875) );
  OR2_X1 U5191 ( .A1(n8244), .A2(n8615), .ZN(n4873) );
  OR2_X1 U5192 ( .A1(n5778), .A2(n5779), .ZN(n8371) );
  OR2_X1 U5193 ( .A1(n8477), .A2(n8463), .ZN(n5743) );
  NAND2_X1 U5194 ( .A1(n5878), .A2(n4460), .ZN(n4791) );
  INV_X1 U5195 ( .A(n4431), .ZN(n5511) );
  NAND2_X1 U5197 ( .A1(n6546), .A2(n5911), .ZN(n8494) );
  NAND2_X1 U5198 ( .A1(n6125), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6149) );
  INV_X1 U5199 ( .A(n6126), .ZN(n6125) );
  OR2_X1 U5200 ( .A1(n6443), .A2(n8743), .ZN(n6459) );
  INV_X1 U5201 ( .A(n8873), .ZN(n7915) );
  AND4_X1 U5202 ( .A1(n6131), .A2(n6130), .A3(n6129), .A4(n6128), .ZN(n7491)
         );
  AND4_X1 U5203 ( .A1(n6094), .A2(n6093), .A3(n6092), .A4(n6091), .ZN(n7229)
         );
  NAND2_X1 U5204 ( .A1(n8980), .A2(n9008), .ZN(n9046) );
  NAND2_X1 U5205 ( .A1(n4967), .A2(n4964), .ZN(n7950) );
  INV_X1 U5206 ( .A(n4965), .ZN(n4964) );
  OAI22_X1 U5207 ( .A1(n9238), .A2(n4966), .B1(n9245), .B2(n9134), .ZN(n4965)
         );
  NAND2_X1 U5208 ( .A1(n4975), .A2(n7892), .ZN(n4972) );
  AOI21_X2 U5209 ( .B1(n9510), .B2(n9312), .A(n9288), .ZN(n7891) );
  NOR2_X1 U5210 ( .A1(n4981), .A2(n4979), .ZN(n4978) );
  AND2_X1 U5211 ( .A1(n9370), .A2(n9135), .ZN(n4981) );
  INV_X1 U5212 ( .A(n5029), .ZN(n4979) );
  AND2_X1 U5213 ( .A1(n9429), .A2(n9136), .ZN(n4942) );
  NOR2_X1 U5214 ( .A1(n6992), .A2(n4584), .ZN(n4583) );
  INV_X1 U5215 ( .A(n9061), .ZN(n4584) );
  NAND2_X1 U5216 ( .A1(n9730), .A2(n9728), .ZN(n6977) );
  NAND2_X1 U5217 ( .A1(n5523), .A2(n5520), .ZN(n5122) );
  AND4_X1 U5218 ( .A1(n5961), .A2(n5960), .A3(n5959), .A4(n6179), .ZN(n5962)
         );
  NAND2_X1 U5219 ( .A1(n6326), .A2(n4934), .ZN(n5998) );
  AND2_X1 U5220 ( .A1(n5994), .A2(n4935), .ZN(n4934) );
  INV_X1 U5221 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4935) );
  INV_X1 U5222 ( .A(n5259), .ZN(n4633) );
  NAND2_X1 U5223 ( .A1(n4623), .A2(n7197), .ZN(n4520) );
  XNOR2_X1 U5224 ( .A(n4624), .B(n8338), .ZN(n4623) );
  NOR2_X1 U5225 ( .A1(n5842), .A2(n5025), .ZN(n4519) );
  NAND2_X1 U5226 ( .A1(n7896), .A2(n7895), .ZN(n9489) );
  NAND2_X1 U5227 ( .A1(n5720), .A2(n4620), .ZN(n4619) );
  INV_X1 U5228 ( .A(n8551), .ZN(n4620) );
  INV_X1 U5229 ( .A(n4618), .ZN(n4617) );
  NAND2_X1 U5230 ( .A1(n8886), .A2(n8885), .ZN(n4543) );
  NOR2_X1 U5231 ( .A1(n8884), .A2(n8976), .ZN(n4542) );
  NAND2_X1 U5232 ( .A1(n4566), .A2(n4490), .ZN(n4565) );
  INV_X1 U5233 ( .A(n4569), .ZN(n4566) );
  AOI21_X1 U5234 ( .B1(n4571), .B2(n8913), .A(n4690), .ZN(n4569) );
  NOR2_X1 U5235 ( .A1(n4570), .A2(n4568), .ZN(n4567) );
  INV_X1 U5236 ( .A(n8913), .ZN(n4570) );
  INV_X1 U5237 ( .A(n8950), .ZN(n4587) );
  OAI21_X1 U5238 ( .B1(n4591), .B2(n4590), .A(n4589), .ZN(n4588) );
  INV_X1 U5239 ( .A(n8951), .ZN(n4589) );
  OAI21_X1 U5240 ( .B1(n8944), .B2(n8976), .A(n9319), .ZN(n4590) );
  NOR2_X1 U5241 ( .A1(n8945), .A2(n8970), .ZN(n4591) );
  AND2_X1 U5242 ( .A1(n7813), .A2(n7863), .ZN(n5776) );
  NAND3_X1 U5243 ( .A1(n4454), .A2(n5861), .A3(n5862), .ZN(n4641) );
  NAND2_X1 U5244 ( .A1(n4917), .A2(n4918), .ZN(n4916) );
  OR2_X1 U5245 ( .A1(n4912), .A2(n4914), .ZN(n4911) );
  INV_X1 U5246 ( .A(n8981), .ZN(n4886) );
  INV_X1 U5247 ( .A(n4770), .ZN(n4769) );
  OAI21_X1 U5248 ( .B1(n5596), .B2(n4771), .A(n5609), .ZN(n4770) );
  INV_X1 U5249 ( .A(n5158), .ZN(n4771) );
  NOR2_X1 U5250 ( .A1(n7144), .A2(n4861), .ZN(n7146) );
  INV_X1 U5251 ( .A(n7245), .ZN(n4827) );
  AOI21_X1 U5252 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7638), .A(n7634), .ZN(
        n7711) );
  NOR2_X1 U5253 ( .A1(n8279), .A2(n4874), .ZN(n8300) );
  NOR2_X1 U5254 ( .A1(n8266), .A2(n8261), .ZN(n4874) );
  INV_X1 U5255 ( .A(n5778), .ZN(n4661) );
  NOR2_X1 U5256 ( .A1(n4668), .A2(n5776), .ZN(n4666) );
  OR2_X1 U5257 ( .A1(n4472), .A2(n5776), .ZN(n5828) );
  OR2_X1 U5258 ( .A1(n8420), .A2(n8401), .ZN(n5800) );
  OR2_X1 U5259 ( .A1(n8024), .A2(n8190), .ZN(n8428) );
  OR2_X1 U5260 ( .A1(n8646), .A2(n8451), .ZN(n5751) );
  INV_X1 U5261 ( .A(n4653), .ZN(n4651) );
  NOR2_X1 U5262 ( .A1(n5532), .A2(n4657), .ZN(n4656) );
  INV_X1 U5263 ( .A(n5743), .ZN(n4657) );
  INV_X1 U5264 ( .A(n8461), .ZN(n5898) );
  OR2_X1 U5265 ( .A1(n8599), .A2(n8078), .ZN(n5738) );
  OR2_X1 U5266 ( .A1(n8609), .A2(n8530), .ZN(n5735) );
  OR2_X1 U5267 ( .A1(n9622), .A2(n8529), .ZN(n5718) );
  OR2_X1 U5268 ( .A1(n9926), .A2(n8137), .ZN(n5710) );
  NAND2_X1 U5269 ( .A1(n7997), .A2(n8036), .ZN(n5698) );
  OR2_X1 U5270 ( .A1(n8198), .A2(n9905), .ZN(n5811) );
  NAND2_X1 U5271 ( .A1(n5922), .A2(n5921), .ZN(n5924) );
  AND2_X1 U5272 ( .A1(n5021), .A2(n5020), .ZN(n5019) );
  NOR2_X1 U5273 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5020) );
  INV_X1 U5274 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5177) );
  INV_X1 U5275 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4784) );
  INV_X1 U5276 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4785) );
  INV_X1 U5277 ( .A(n4916), .ZN(n4914) );
  OAI22_X1 U5278 ( .A1(n8801), .A2(n4915), .B1(n4916), .B2(n4913), .ZN(n4912)
         );
  INV_X1 U5279 ( .A(n4917), .ZN(n4915) );
  INV_X1 U5280 ( .A(n8731), .ZN(n4913) );
  INV_X1 U5281 ( .A(n6387), .ZN(n4904) );
  INV_X1 U5282 ( .A(n6455), .ZN(n4924) );
  AND2_X1 U5283 ( .A1(n4485), .A2(n4560), .ZN(n4559) );
  NAND2_X1 U5284 ( .A1(n4731), .A2(n9223), .ZN(n4560) );
  NAND2_X1 U5285 ( .A1(n9131), .A2(n9132), .ZN(n4727) );
  AOI21_X1 U5286 ( .B1(n4561), .B2(n4441), .A(n9565), .ZN(n4557) );
  AOI21_X1 U5287 ( .B1(n8961), .B2(n8991), .A(n8960), .ZN(n4575) );
  NAND2_X1 U5288 ( .A1(n8968), .A2(n4573), .ZN(n4572) );
  AND2_X1 U5289 ( .A1(n8969), .A2(n4574), .ZN(n4573) );
  NAND2_X1 U5290 ( .A1(n7948), .A2(n8970), .ZN(n4574) );
  NOR2_X1 U5291 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6026) );
  NAND2_X1 U5292 ( .A1(n4968), .A2(n4969), .ZN(n4966) );
  OR2_X1 U5293 ( .A1(n9245), .A2(n9257), .ZN(n8991) );
  AOI21_X1 U5294 ( .B1(n4884), .B2(n4885), .A(n4883), .ZN(n4882) );
  INV_X1 U5295 ( .A(n8983), .ZN(n4883) );
  INV_X1 U5296 ( .A(n7913), .ZN(n4884) );
  NAND2_X1 U5297 ( .A1(n4505), .A2(n4885), .ZN(n4881) );
  NOR2_X1 U5298 ( .A1(n9524), .A2(n9360), .ZN(n4708) );
  OR2_X1 U5299 ( .A1(n9524), .A2(n8795), .ZN(n8995) );
  NOR2_X1 U5300 ( .A1(n9351), .A2(n4890), .ZN(n4889) );
  INV_X1 U5301 ( .A(n9096), .ZN(n4890) );
  OR2_X1 U5302 ( .A1(n9429), .A2(n9440), .ZN(n8919) );
  NOR2_X1 U5303 ( .A1(n9457), .A2(n4690), .ZN(n4689) );
  NAND2_X1 U5304 ( .A1(n7739), .A2(n8913), .ZN(n7740) );
  INV_X1 U5305 ( .A(n7666), .ZN(n4960) );
  INV_X1 U5306 ( .A(n4686), .ZN(n4685) );
  OAI21_X1 U5307 ( .B1(n7517), .B2(n4687), .A(n9551), .ZN(n4686) );
  INV_X1 U5308 ( .A(n9552), .ZN(n4687) );
  OR2_X1 U5309 ( .A1(n8711), .A2(n8828), .ZN(n9073) );
  NOR2_X1 U5310 ( .A1(n4952), .A2(n4949), .ZN(n4948) );
  NAND2_X1 U5311 ( .A1(n7627), .A2(n7518), .ZN(n8908) );
  NAND2_X1 U5312 ( .A1(n4456), .A2(n6991), .ZN(n4577) );
  INV_X1 U5313 ( .A(n7899), .ZN(n4777) );
  NOR2_X1 U5314 ( .A1(n6607), .A2(n6641), .ZN(n4531) );
  INV_X1 U5315 ( .A(n6581), .ZN(n4681) );
  OR2_X1 U5316 ( .A1(n9425), .A2(n7910), .ZN(n9406) );
  NOR2_X1 U5317 ( .A1(n5966), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4982) );
  NAND2_X1 U5318 ( .A1(n4715), .A2(n5147), .ZN(n5585) );
  NAND2_X1 U5319 ( .A1(n5576), .A2(n5575), .ZN(n4715) );
  NAND2_X1 U5320 ( .A1(n4735), .A2(n4733), .ZN(n5508) );
  AND2_X1 U5321 ( .A1(n4734), .A2(n5112), .ZN(n4733) );
  XNOR2_X1 U5322 ( .A(n5095), .B(SI_14_), .ZN(n5435) );
  NAND2_X1 U5323 ( .A1(n5093), .A2(n5092), .ZN(n5436) );
  INV_X1 U5324 ( .A(n5420), .ZN(n5090) );
  INV_X1 U5325 ( .A(n4722), .ZN(n4721) );
  OAI21_X1 U5326 ( .B1(n4725), .B2(n4449), .A(n5087), .ZN(n4722) );
  NOR2_X1 U5327 ( .A1(n5082), .A2(n4726), .ZN(n4725) );
  INV_X1 U5328 ( .A(n5391), .ZN(n5082) );
  NAND2_X1 U5329 ( .A1(n5371), .A2(n5076), .ZN(n5078) );
  NAND2_X1 U5330 ( .A1(n5080), .A2(SI_10_), .ZN(n5081) );
  NAND2_X1 U5331 ( .A1(n5087), .A2(n5086), .ZN(n5402) );
  INV_X1 U5332 ( .A(n7572), .ZN(n4985) );
  NAND2_X1 U5333 ( .A1(n8064), .A2(n8063), .ZN(n7838) );
  OR2_X1 U5334 ( .A1(n8622), .A2(n5636), .ZN(n5787) );
  OAI21_X1 U5335 ( .B1(n4658), .B2(n5625), .A(n5624), .ZN(n5945) );
  NAND2_X1 U5336 ( .A1(n7873), .A2(n7973), .ZN(n5624) );
  OAI211_X1 U5337 ( .C1(n4861), .C2(n7199), .A(n4858), .B(n4854), .ZN(n7290)
         );
  NOR2_X1 U5338 ( .A1(n4861), .A2(n7162), .ZN(n4855) );
  OR2_X1 U5339 ( .A1(n7357), .A2(n4813), .ZN(n4812) );
  AND2_X1 U5340 ( .A1(n7358), .A2(n7365), .ZN(n4813) );
  AND2_X1 U5341 ( .A1(n4812), .A2(n4811), .ZN(n9839) );
  INV_X1 U5342 ( .A(n9840), .ZN(n4811) );
  OAI21_X1 U5343 ( .B1(n7360), .B2(n7441), .A(n7454), .ZN(n7361) );
  NOR2_X1 U5344 ( .A1(n7371), .A2(n5365), .ZN(n7450) );
  NAND2_X1 U5345 ( .A1(n4841), .A2(n4839), .ZN(n7727) );
  AND2_X1 U5346 ( .A1(n4842), .A2(n4499), .ZN(n4839) );
  XNOR2_X1 U5347 ( .A(n7711), .B(n7729), .ZN(n7635) );
  OR2_X1 U5348 ( .A1(n7635), .A2(n5397), .ZN(n4851) );
  NOR2_X1 U5349 ( .A1(n7729), .A2(n7711), .ZN(n7713) );
  OR2_X1 U5350 ( .A1(n7788), .A2(n7794), .ZN(n4831) );
  OR2_X1 U5351 ( .A1(n8233), .A2(n8232), .ZN(n8234) );
  AND2_X1 U5352 ( .A1(n8260), .A2(n8267), .ZN(n4876) );
  NOR2_X1 U5353 ( .A1(n8257), .A2(n8536), .ZN(n4819) );
  NOR2_X1 U5354 ( .A1(n8277), .A2(n4532), .ZN(n8295) );
  NOR2_X1 U5355 ( .A1(n8266), .A2(n8518), .ZN(n4532) );
  NAND2_X1 U5356 ( .A1(n5784), .A2(n5783), .ZN(n5944) );
  NAND2_X1 U5357 ( .A1(n8369), .A2(n8500), .ZN(n5917) );
  AOI21_X1 U5358 ( .B1(n4795), .B2(n4797), .A(n4439), .ZN(n4793) );
  XNOR2_X1 U5359 ( .A(n7873), .B(n8369), .ZN(n7867) );
  AND3_X1 U5360 ( .A1(n5583), .A2(n5582), .A3(n5581), .ZN(n8402) );
  NOR2_X1 U5361 ( .A1(n5584), .A2(n4671), .ZN(n4670) );
  OAI21_X1 U5362 ( .B1(n5584), .B2(n4669), .A(n5772), .ZN(n4668) );
  NAND2_X1 U5363 ( .A1(n5766), .A2(n5825), .ZN(n4669) );
  NAND2_X1 U5364 ( .A1(n5217), .A2(n10012), .ZN(n5579) );
  INV_X1 U5365 ( .A(n5570), .ZN(n5217) );
  OR2_X1 U5366 ( .A1(n8646), .A2(n8189), .ZN(n5901) );
  AOI21_X1 U5367 ( .B1(n4656), .B2(n5896), .A(n4654), .ZN(n4653) );
  INV_X1 U5368 ( .A(n5803), .ZN(n4654) );
  INV_X1 U5369 ( .A(n4656), .ZN(n4655) );
  AND2_X1 U5370 ( .A1(n5804), .A2(n5803), .ZN(n8461) );
  AND4_X1 U5371 ( .A1(n5543), .A2(n5542), .A3(n5541), .A4(n5540), .ZN(n8464)
         );
  NAND2_X1 U5372 ( .A1(n8471), .A2(n5896), .ZN(n4800) );
  AND4_X1 U5373 ( .A1(n5490), .A2(n5489), .A3(n5488), .A4(n5487), .ZN(n8514)
         );
  OR2_X1 U5374 ( .A1(n9622), .A2(n8192), .ZN(n5887) );
  AND4_X1 U5375 ( .A1(n5461), .A2(n5460), .A3(n5459), .A4(n5458), .ZN(n8545)
         );
  AND2_X1 U5376 ( .A1(n5718), .A2(n5719), .ZN(n8551) );
  NAND2_X1 U5377 ( .A1(n4515), .A2(n4443), .ZN(n4805) );
  AND2_X1 U5378 ( .A1(n5419), .A2(n5704), .ZN(n4647) );
  INV_X1 U5379 ( .A(n7676), .ZN(n4646) );
  INV_X1 U5380 ( .A(n8193), .ZN(n8544) );
  NAND2_X1 U5381 ( .A1(n7677), .A2(n4421), .ZN(n7676) );
  INV_X1 U5382 ( .A(n8194), .ZN(n8137) );
  INV_X1 U5383 ( .A(n4790), .ZN(n4789) );
  OAI21_X1 U5384 ( .B1(n4791), .B2(n7586), .A(n5879), .ZN(n4790) );
  NAND2_X1 U5385 ( .A1(n5206), .A2(n5205), .ZN(n5379) );
  INV_X1 U5386 ( .A(n5363), .ZN(n5206) );
  AND4_X1 U5387 ( .A1(n5401), .A2(n5400), .A3(n5399), .A4(n5398), .ZN(n8038)
         );
  OR2_X1 U5388 ( .A1(n5350), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U5389 ( .A1(n5204), .A2(n5203), .ZN(n5350) );
  INV_X1 U5390 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5203) );
  INV_X1 U5391 ( .A(n5335), .ZN(n5204) );
  NAND2_X1 U5392 ( .A1(n5914), .A2(n6575), .ZN(n9863) );
  INV_X1 U5393 ( .A(n8500), .ZN(n9865) );
  INV_X1 U5394 ( .A(n8494), .ZN(n9869) );
  INV_X1 U5395 ( .A(n7012), .ZN(n5262) );
  INV_X1 U5396 ( .A(n7997), .ZN(n9910) );
  NAND2_X1 U5397 ( .A1(n5924), .A2(n5923), .ZN(n5925) );
  INV_X1 U5398 ( .A(n4673), .ZN(n5249) );
  INV_X1 U5399 ( .A(n7475), .ZN(n4929) );
  AND2_X1 U5400 ( .A1(n6139), .A2(n6138), .ZN(n7530) );
  NAND2_X1 U5401 ( .A1(n4927), .A2(n4926), .ZN(n8714) );
  AND2_X1 U5402 ( .A1(n5024), .A2(n6340), .ZN(n4926) );
  NAND2_X1 U5403 ( .A1(n6147), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6166) );
  NAND2_X1 U5404 ( .A1(n6277), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6313) );
  INV_X1 U5405 ( .A(n6293), .ZN(n6277) );
  OR2_X1 U5406 ( .A1(n6236), .A2(n6235), .ZN(n4918) );
  NAND2_X1 U5407 ( .A1(n4537), .A2(n6033), .ZN(n6034) );
  NAND2_X1 U5408 ( .A1(n4538), .A2(n6965), .ZN(n4537) );
  OR2_X1 U5409 ( .A1(n7310), .A2(n7309), .ZN(n4933) );
  NAND2_X1 U5410 ( .A1(n4436), .A2(n9109), .ZN(n4783) );
  NAND2_X1 U5411 ( .A1(n4547), .A2(n4546), .ZN(n9052) );
  AND2_X1 U5412 ( .A1(n4781), .A2(n9056), .ZN(n4780) );
  OR2_X1 U5413 ( .A1(n9055), .A2(n4539), .ZN(n4781) );
  OAI22_X1 U5414 ( .A1(n8871), .A2(n6640), .B1(n8873), .B2(n6030), .ZN(n4680)
         );
  AND2_X1 U5415 ( .A1(n7924), .A2(n6011), .ZN(n6041) );
  CLKBUF_X1 U5416 ( .A(n6026), .Z(n6027) );
  INV_X1 U5417 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4605) );
  OR2_X1 U5418 ( .A1(n6779), .A2(n6778), .ZN(n4600) );
  NOR2_X1 U5419 ( .A1(n9483), .A2(n7951), .ZN(n9231) );
  NAND2_X1 U5420 ( .A1(n4713), .A2(n7955), .ZN(n4712) );
  NAND2_X1 U5421 ( .A1(n9279), .A2(n9297), .ZN(n4973) );
  AND2_X1 U5422 ( .A1(n8990), .A2(n8965), .ZN(n9254) );
  NAND2_X1 U5423 ( .A1(n7890), .A2(n7889), .ZN(n9288) );
  OR2_X1 U5424 ( .A1(n4705), .A2(n8771), .ZN(n7889) );
  NAND2_X1 U5425 ( .A1(n9302), .A2(n7888), .ZN(n7890) );
  OR2_X1 U5426 ( .A1(n9514), .A2(n9322), .ZN(n7888) );
  NAND2_X1 U5427 ( .A1(n9318), .A2(n7913), .ZN(n9310) );
  NAND2_X1 U5428 ( .A1(n9320), .A2(n9319), .ZN(n9318) );
  AND2_X1 U5429 ( .A1(n9524), .A2(n9321), .ZN(n7886) );
  NAND2_X1 U5430 ( .A1(n8995), .A2(n8942), .ZN(n9339) );
  NAND2_X1 U5431 ( .A1(n9375), .A2(n4889), .ZN(n9353) );
  NAND2_X1 U5432 ( .A1(n9386), .A2(n7882), .ZN(n7883) );
  AND2_X1 U5433 ( .A1(n8936), .A2(n9096), .ZN(n9377) );
  NOR2_X1 U5434 ( .A1(n9467), .A2(n9452), .ZN(n9447) );
  OR2_X1 U5435 ( .A1(n9642), .A2(n8756), .ZN(n5028) );
  OR2_X1 U5436 ( .A1(n9452), .A2(n9459), .ZN(n7878) );
  NAND2_X1 U5437 ( .A1(n7909), .A2(n9082), .ZN(n9458) );
  OR2_X1 U5438 ( .A1(n6243), .A2(n8803), .ZN(n6260) );
  OR2_X1 U5439 ( .A1(n6166), .A2(n10217), .ZN(n6198) );
  AND2_X1 U5440 ( .A1(n9072), .A2(n4896), .ZN(n7516) );
  NAND2_X1 U5441 ( .A1(n7515), .A2(n7514), .ZN(n4896) );
  NAND2_X1 U5442 ( .A1(n7542), .A2(n7522), .ZN(n7523) );
  NAND2_X1 U5443 ( .A1(n7598), .A2(n8892), .ZN(n7597) );
  OAI21_X1 U5444 ( .B1(n7224), .B2(n7226), .A(n7223), .ZN(n7225) );
  NAND2_X1 U5445 ( .A1(n6981), .A2(n6980), .ZN(n6996) );
  OR2_X1 U5446 ( .A1(n9713), .A2(n6968), .ZN(n6969) );
  INV_X1 U5447 ( .A(n6964), .ZN(n4530) );
  NOR2_X1 U5448 ( .A1(n6974), .A2(n9739), .ZN(n9729) );
  NAND2_X1 U5449 ( .A1(n4420), .A2(n6000), .ZN(n7494) );
  NAND2_X1 U5450 ( .A1(n4776), .A2(n7898), .ZN(n9483) );
  INV_X1 U5451 ( .A(n8880), .ZN(n6342) );
  INV_X1 U5452 ( .A(n6607), .ZN(n6341) );
  AND2_X1 U5453 ( .A1(n6927), .A2(n9115), .ZN(n9629) );
  NAND2_X1 U5454 ( .A1(n5627), .A2(n5167), .ZN(n5198) );
  XNOR2_X1 U5455 ( .A(n5198), .B(n5197), .ZN(n8878) );
  NAND2_X1 U5456 ( .A1(n5626), .A2(SI_29_), .ZN(n5627) );
  NAND2_X1 U5457 ( .A1(n4772), .A2(n4773), .ZN(n4778) );
  INV_X1 U5458 ( .A(SI_29_), .ZN(n4773) );
  NAND2_X1 U5459 ( .A1(n5153), .A2(n5152), .ZN(n5597) );
  NAND2_X1 U5460 ( .A1(n5585), .A2(n5586), .ZN(n5153) );
  AND3_X1 U5461 ( .A1(n5972), .A2(n4983), .A3(n4982), .ZN(n5981) );
  XNOR2_X1 U5462 ( .A(n5576), .B(n5575), .ZN(n7765) );
  AND2_X1 U5463 ( .A1(n5136), .A2(n5135), .ZN(n5556) );
  OAI21_X1 U5464 ( .B1(n5535), .B2(n5126), .A(n5125), .ZN(n5545) );
  INV_X1 U5465 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4938) );
  NAND2_X1 U5466 ( .A1(n4732), .A2(n4737), .ZN(n5493) );
  OR2_X1 U5467 ( .A1(n5450), .A2(n4741), .ZN(n4732) );
  NAND2_X1 U5468 ( .A1(n4743), .A2(n4745), .ZN(n5477) );
  NAND2_X1 U5469 ( .A1(n5450), .A2(n4746), .ZN(n4743) );
  NAND2_X1 U5470 ( .A1(n5972), .A2(n4941), .ZN(n6271) );
  NAND2_X1 U5471 ( .A1(n4744), .A2(n5100), .ZN(n5465) );
  OR2_X1 U5472 ( .A1(n5450), .A2(n5101), .ZN(n4744) );
  OAI21_X1 U5473 ( .B1(n4629), .B2(n5370), .A(n4627), .ZN(n5392) );
  AOI21_X1 U5474 ( .B1(n5076), .B2(n4628), .A(n4726), .ZN(n4627) );
  INV_X1 U5475 ( .A(n5071), .ZN(n4628) );
  XNOR2_X1 U5476 ( .A(n5063), .B(SI_7_), .ZN(n5345) );
  XNOR2_X1 U5477 ( .A(n5041), .B(SI_1_), .ZN(n5247) );
  NAND2_X1 U5478 ( .A1(n7569), .A2(n4987), .ZN(n7571) );
  INV_X1 U5479 ( .A(n7865), .ZN(n4991) );
  AND4_X1 U5480 ( .A1(n5519), .A2(n5518), .A3(n5517), .A4(n5516), .ZN(n8463)
         );
  NAND2_X1 U5481 ( .A1(n7825), .A2(n4999), .ZN(n4998) );
  AND2_X1 U5482 ( .A1(n4997), .A2(n4995), .ZN(n4994) );
  INV_X1 U5483 ( .A(n7818), .ZN(n4999) );
  NAND2_X1 U5484 ( .A1(n5424), .A2(n5423), .ZN(n8117) );
  OR2_X1 U5485 ( .A1(n6812), .A2(n6886), .ZN(n8175) );
  NAND2_X1 U5486 ( .A1(n5455), .A2(n5454), .ZN(n8533) );
  NAND2_X1 U5487 ( .A1(n6819), .A2(n9860), .ZN(n8177) );
  AND2_X1 U5488 ( .A1(n5635), .A2(n5634), .ZN(n7871) );
  INV_X1 U5489 ( .A(n8463), .ZN(n8484) );
  NAND2_X1 U5490 ( .A1(n4823), .A2(n8246), .ZN(n4821) );
  INV_X1 U5491 ( .A(n8234), .ZN(n4823) );
  NAND2_X1 U5492 ( .A1(n8234), .A2(n8267), .ZN(n8254) );
  INV_X1 U5493 ( .A(n4873), .ZN(n8259) );
  AND3_X1 U5494 ( .A1(n4821), .A2(n8254), .A3(P2_REG2_REG_15__SCAN_IN), .ZN(
        n8255) );
  XNOR2_X1 U5495 ( .A(n8295), .B(n8307), .ZN(n8278) );
  NOR2_X1 U5496 ( .A1(n4835), .A2(n8325), .ZN(n4834) );
  INV_X1 U5497 ( .A(n4836), .ZN(n4835) );
  OR2_X1 U5498 ( .A1(n8278), .A2(n4837), .ZN(n4833) );
  NAND2_X1 U5499 ( .A1(n4838), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4837) );
  NOR2_X1 U5500 ( .A1(n8344), .A2(n8343), .ZN(n8346) );
  NAND2_X1 U5501 ( .A1(n4536), .A2(n4535), .ZN(n4534) );
  INV_X1 U5502 ( .A(n8347), .ZN(n4535) );
  NAND2_X1 U5503 ( .A1(n8348), .A2(n9821), .ZN(n4536) );
  NAND2_X1 U5504 ( .A1(n4514), .A2(n4513), .ZN(n4512) );
  NAND2_X1 U5505 ( .A1(n8389), .A2(n8500), .ZN(n4513) );
  INV_X1 U5506 ( .A(n9915), .ZN(n9927) );
  NAND2_X1 U5507 ( .A1(n5196), .A2(n5195), .ZN(n8555) );
  AND3_X1 U5508 ( .A1(n5377), .A2(n5376), .A3(n5375), .ZN(n7618) );
  INV_X1 U5509 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5039) );
  INV_X1 U5510 ( .A(n9580), .ZN(n9279) );
  NAND2_X1 U5511 ( .A1(n6422), .A2(n6421), .ZN(n9510) );
  AND2_X1 U5512 ( .A1(n6449), .A2(n6448), .ZN(n9256) );
  NAND2_X1 U5513 ( .A1(n6465), .A2(n6464), .ZN(n9275) );
  OR2_X1 U5514 ( .A1(n6683), .A2(n6682), .ZN(n4598) );
  AND2_X1 U5515 ( .A1(n4600), .A2(n4599), .ZN(n6683) );
  NAND2_X1 U5516 ( .A1(n6636), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4599) );
  NAND2_X1 U5517 ( .A1(n4893), .A2(n4892), .ZN(n4891) );
  NAND2_X1 U5518 ( .A1(n9132), .A2(n9225), .ZN(n4892) );
  OAI22_X1 U5519 ( .A1(n7950), .A2(n7897), .B1(n7955), .B2(n7914), .ZN(n7905)
         );
  AOI21_X1 U5520 ( .B1(n7958), .B2(n9715), .A(n4697), .ZN(n9492) );
  NAND2_X1 U5521 ( .A1(n4699), .A2(n4698), .ZN(n4697) );
  NAND2_X1 U5522 ( .A1(n9133), .A2(n9460), .ZN(n4698) );
  INV_X1 U5523 ( .A(n9740), .ZN(n9724) );
  AND2_X1 U5524 ( .A1(n6927), .A2(n6501), .ZN(n9736) );
  OR2_X1 U5525 ( .A1(n4419), .A2(n6935), .ZN(n9741) );
  OAI21_X1 U5526 ( .B1(n4618), .B2(n5720), .A(n4621), .ZN(n4616) );
  AND2_X1 U5527 ( .A1(n5735), .A2(n5721), .ZN(n4621) );
  OAI21_X1 U5528 ( .B1(n5717), .B2(n4622), .A(n4617), .ZN(n5734) );
  NAND2_X1 U5529 ( .A1(n4541), .A2(n4540), .ZN(n8907) );
  NAND2_X1 U5530 ( .A1(n8899), .A2(n8976), .ZN(n4540) );
  NAND2_X1 U5531 ( .A1(n4543), .A2(n4542), .ZN(n4541) );
  NAND2_X1 U5532 ( .A1(n8912), .A2(n9073), .ZN(n4568) );
  AOI21_X1 U5533 ( .B1(n5730), .B2(n5941), .A(n5744), .ZN(n4638) );
  NAND2_X1 U5534 ( .A1(n5729), .A2(n6575), .ZN(n4637) );
  AND2_X1 U5535 ( .A1(n5747), .A2(n5803), .ZN(n4635) );
  AND2_X1 U5536 ( .A1(n4565), .A2(n9084), .ZN(n4564) );
  NAND2_X1 U5537 ( .A1(n4585), .A2(n8953), .ZN(n8963) );
  NAND2_X1 U5538 ( .A1(n4588), .A2(n4586), .ZN(n4585) );
  NOR2_X1 U5539 ( .A1(n4587), .A2(n9287), .ZN(n4586) );
  INV_X1 U5540 ( .A(n7457), .ZN(n4843) );
  OR2_X1 U5541 ( .A1(n9510), .A2(n8952), .ZN(n8983) );
  NAND2_X1 U5542 ( .A1(n8908), .A2(n8883), .ZN(n8896) );
  OR2_X1 U5543 ( .A1(n9263), .A2(n9279), .ZN(n4714) );
  NOR2_X1 U5544 ( .A1(n8738), .A2(n4422), .ZN(n4704) );
  INV_X1 U5545 ( .A(n4753), .ZN(n4752) );
  OAI21_X1 U5546 ( .B1(n4754), .B2(n4756), .A(n5556), .ZN(n4753) );
  AND2_X1 U5547 ( .A1(n6761), .A2(n7334), .ZN(n5006) );
  OR4_X1 U5548 ( .A1(n5833), .A2(n5832), .A3(n5831), .A4(n5830), .ZN(n5837) );
  NOR2_X1 U5549 ( .A1(n4815), .A2(n9817), .ZN(n4814) );
  NAND2_X1 U5550 ( .A1(n4810), .A2(n4809), .ZN(n7360) );
  NAND2_X1 U5551 ( .A1(n9854), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4809) );
  INV_X1 U5552 ( .A(n9839), .ZN(n4810) );
  AOI21_X1 U5553 ( .B1(n8243), .B2(P2_REG1_REG_14__SCAN_IN), .A(n8242), .ZN(
        n8258) );
  INV_X1 U5554 ( .A(n4796), .ZN(n4795) );
  OAI21_X1 U5555 ( .B1(n4799), .B2(n4797), .A(n5907), .ZN(n4796) );
  NAND2_X1 U5556 ( .A1(n5906), .A2(n8378), .ZN(n5907) );
  INV_X1 U5557 ( .A(n4798), .ZN(n4797) );
  AND2_X1 U5558 ( .A1(n4437), .A2(n5905), .ZN(n4799) );
  NAND2_X1 U5559 ( .A1(n5860), .A2(n5251), .ZN(n5654) );
  NOR2_X1 U5560 ( .A1(n4912), .A2(n4909), .ZN(n4908) );
  INV_X1 U5561 ( .A(n6216), .ZN(n4909) );
  AND2_X1 U5562 ( .A1(n4480), .A2(n4907), .ZN(n4906) );
  OR2_X1 U5563 ( .A1(n4912), .A2(n4919), .ZN(n4907) );
  OR2_X1 U5564 ( .A1(n8873), .A2(n6040), .ZN(n6046) );
  NOR2_X1 U5565 ( .A1(n9245), .A2(n4714), .ZN(n4713) );
  AND2_X1 U5566 ( .A1(n9489), .A2(n7914), .ZN(n8959) );
  NOR2_X1 U5567 ( .A1(n9521), .A2(n4707), .ZN(n4706) );
  INV_X1 U5568 ( .A(n4708), .ZN(n4707) );
  AOI21_X1 U5569 ( .B1(n4961), .B2(n7517), .A(n4957), .ZN(n4956) );
  INV_X1 U5570 ( .A(n4959), .ZN(n4958) );
  INV_X1 U5571 ( .A(n8896), .ZN(n9025) );
  INV_X1 U5572 ( .A(n9730), .ZN(n9016) );
  NOR2_X1 U5573 ( .A1(n9289), .A2(n4714), .ZN(n9261) );
  NOR2_X1 U5574 ( .A1(n9289), .A2(n9279), .ZN(n9278) );
  NAND2_X1 U5575 ( .A1(n7669), .A2(n4704), .ZN(n7750) );
  AND2_X1 U5576 ( .A1(n7669), .A2(n9696), .ZN(n9548) );
  OR2_X1 U5577 ( .A1(n7545), .A2(n7627), .ZN(n7547) );
  AOI21_X1 U5578 ( .B1(n4769), .B2(n4771), .A(n4767), .ZN(n4766) );
  INV_X1 U5579 ( .A(n5163), .ZN(n4767) );
  XNOR2_X1 U5580 ( .A(n5166), .B(n5164), .ZN(n5626) );
  NAND2_X1 U5581 ( .A1(n4758), .A2(n5125), .ZN(n4757) );
  INV_X1 U5582 ( .A(n5544), .ZN(n4758) );
  AOI21_X1 U5583 ( .B1(n4740), .B2(n4739), .A(n4738), .ZN(n4737) );
  INV_X1 U5584 ( .A(n5108), .ZN(n4738) );
  INV_X1 U5585 ( .A(n4746), .ZN(n4739) );
  INV_X1 U5586 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4940) );
  AOI21_X1 U5587 ( .B1(n4746), .B2(n5101), .A(n4474), .ZN(n4745) );
  AND2_X1 U5588 ( .A1(n5972), .A2(n5973), .ZN(n6286) );
  XNOR2_X1 U5589 ( .A(n5091), .B(SI_13_), .ZN(n5420) );
  NAND2_X1 U5590 ( .A1(n4716), .A2(n4717), .ZN(n5421) );
  AOI21_X1 U5591 ( .B1(n4432), .B2(n4449), .A(n4475), .ZN(n4717) );
  OR2_X1 U5592 ( .A1(n6181), .A2(n6180), .ZN(n6193) );
  CLKBUF_X1 U5593 ( .A(n6115), .Z(n6116) );
  OAI21_X1 U5594 ( .B1(n5194), .B2(n4507), .A(n4506), .ZN(n5044) );
  NAND2_X1 U5595 ( .A1(n5194), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4506) );
  NAND2_X1 U5596 ( .A1(n5194), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5038) );
  NAND2_X1 U5597 ( .A1(n4988), .A2(n8200), .ZN(n4987) );
  OAI21_X1 U5598 ( .B1(n7819), .B2(n7818), .A(n4993), .ZN(n8034) );
  INV_X1 U5599 ( .A(n4996), .ZN(n4993) );
  AND2_X1 U5600 ( .A1(n7970), .A2(n7968), .ZN(n7865) );
  XNOR2_X1 U5601 ( .A(n9876), .B(n6880), .ZN(n6881) );
  NAND2_X1 U5602 ( .A1(n8095), .A2(n7846), .ZN(n8026) );
  INV_X1 U5603 ( .A(n8498), .ZN(n8078) );
  NOR2_X1 U5604 ( .A1(n8077), .A2(n5001), .ZN(n5000) );
  INV_X1 U5605 ( .A(n7837), .ZN(n5001) );
  NAND2_X1 U5606 ( .A1(n7286), .A2(n5201), .ZN(n5307) );
  INV_X1 U5607 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U5608 ( .A1(n8098), .A2(n4525), .ZN(n8095) );
  AND2_X1 U5609 ( .A1(n8096), .A2(n8097), .ZN(n4525) );
  AOI21_X1 U5610 ( .B1(n7825), .B2(n4996), .A(n4462), .ZN(n4995) );
  NAND2_X1 U5611 ( .A1(n7826), .A2(n7825), .ZN(n4997) );
  NAND2_X1 U5612 ( .A1(n5216), .A2(n5215), .ZN(n5548) );
  INV_X1 U5613 ( .A(n5538), .ZN(n5216) );
  OR2_X1 U5614 ( .A1(n5548), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5560) );
  AND2_X1 U5615 ( .A1(n6833), .A2(n6832), .ZN(n7065) );
  OR2_X1 U5616 ( .A1(n8555), .A2(n8353), .ZN(n5798) );
  NAND2_X1 U5617 ( .A1(n4425), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5242) );
  NAND2_X1 U5618 ( .A1(n7142), .A2(n7143), .ZN(n9816) );
  AND2_X1 U5619 ( .A1(n4816), .A2(n7143), .ZN(n7205) );
  NAND2_X1 U5620 ( .A1(n9828), .A2(n7161), .ZN(n7200) );
  INV_X1 U5621 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7286) );
  AND2_X1 U5622 ( .A1(n7144), .A2(n4861), .ZN(n7145) );
  NAND2_X1 U5623 ( .A1(n4857), .A2(n7287), .ZN(n7179) );
  NAND2_X1 U5624 ( .A1(n7199), .A2(n7162), .ZN(n4857) );
  NAND2_X1 U5625 ( .A1(n7149), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7246) );
  NAND3_X1 U5626 ( .A1(n4423), .A2(n4824), .A3(n4464), .ZN(n4825) );
  NAND2_X1 U5627 ( .A1(n7244), .A2(n4827), .ZN(n4826) );
  XNOR2_X1 U5628 ( .A(n7356), .B(n4533), .ZN(n7267) );
  INV_X1 U5629 ( .A(n7365), .ZN(n4533) );
  OR2_X1 U5630 ( .A1(n7271), .A2(n5337), .ZN(n4847) );
  NOR2_X1 U5631 ( .A1(n7450), .A2(n7449), .ZN(n7453) );
  NOR2_X1 U5632 ( .A1(n7453), .A2(n7452), .ZN(n7634) );
  NOR2_X1 U5633 ( .A1(n7361), .A2(n7362), .ZN(n7456) );
  NAND2_X1 U5634 ( .A1(n4841), .A2(n4842), .ZN(n7631) );
  INV_X1 U5635 ( .A(n7727), .ZN(n7728) );
  NOR2_X1 U5636 ( .A1(n8280), .A2(n8283), .ZN(n8301) );
  INV_X1 U5637 ( .A(n8298), .ZN(n4838) );
  NAND2_X1 U5638 ( .A1(n4864), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4863) );
  NAND2_X1 U5639 ( .A1(n8302), .A2(n4864), .ZN(n4862) );
  INV_X1 U5640 ( .A(n8304), .ZN(n4864) );
  NAND2_X1 U5641 ( .A1(n4660), .A2(n5775), .ZN(n4659) );
  INV_X1 U5642 ( .A(n4666), .ZN(n4664) );
  AOI21_X1 U5643 ( .B1(n4666), .B2(n4663), .A(n4472), .ZN(n4662) );
  INV_X1 U5644 ( .A(n4670), .ZN(n4663) );
  NAND2_X1 U5645 ( .A1(n8369), .A2(n8499), .ZN(n4514) );
  NAND2_X1 U5646 ( .A1(n5771), .A2(n5772), .ZN(n8394) );
  NAND2_X1 U5647 ( .A1(n5219), .A2(n5218), .ZN(n5589) );
  INV_X1 U5648 ( .A(n5579), .ZN(n5219) );
  INV_X1 U5649 ( .A(n8399), .ZN(n8411) );
  OR2_X1 U5650 ( .A1(n5560), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5570) );
  AOI21_X1 U5651 ( .B1(n4650), .B2(n4655), .A(n5752), .ZN(n4648) );
  NOR2_X1 U5652 ( .A1(n5756), .A2(n4651), .ZN(n4650) );
  NAND2_X1 U5653 ( .A1(n5214), .A2(n10033), .ZN(n5526) );
  INV_X1 U5654 ( .A(n5514), .ZN(n5214) );
  AND2_X1 U5655 ( .A1(n5738), .A2(n5725), .ZN(n8489) );
  NAND2_X1 U5656 ( .A1(n5213), .A2(n5212), .ZN(n5501) );
  INV_X1 U5657 ( .A(n5484), .ZN(n5213) );
  OR2_X1 U5658 ( .A1(n8533), .A2(n8545), .ZN(n5721) );
  OR2_X1 U5659 ( .A1(n5470), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U5660 ( .A1(n5211), .A2(n5210), .ZN(n5470) );
  INV_X1 U5661 ( .A(n5456), .ZN(n5211) );
  AND4_X1 U5662 ( .A1(n5475), .A2(n5474), .A3(n5473), .A4(n5472), .ZN(n8530)
         );
  NAND2_X1 U5663 ( .A1(n5209), .A2(n5208), .ZN(n5442) );
  INV_X1 U5664 ( .A(n5425), .ZN(n5209) );
  AOI21_X1 U5665 ( .B1(n7820), .B2(n4647), .A(n4643), .ZN(n4642) );
  INV_X1 U5666 ( .A(n4647), .ZN(n4644) );
  INV_X1 U5667 ( .A(n5710), .ZN(n4643) );
  NAND2_X1 U5668 ( .A1(n5207), .A2(n7721), .ZN(n5425) );
  INV_X1 U5669 ( .A(n5413), .ZN(n5207) );
  OR2_X1 U5670 ( .A1(n5395), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5413) );
  OR2_X1 U5671 ( .A1(n5379), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U5672 ( .A1(n4788), .A2(n5878), .ZN(n7652) );
  NAND2_X1 U5673 ( .A1(n7583), .A2(n7586), .ZN(n4788) );
  NAND2_X1 U5674 ( .A1(n5697), .A2(n5684), .ZN(n7586) );
  NAND2_X1 U5675 ( .A1(n5202), .A2(n10234), .ZN(n5321) );
  INV_X1 U5676 ( .A(n5307), .ZN(n5202) );
  OR2_X1 U5677 ( .A1(n5321), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U5678 ( .A1(n7052), .A2(n7054), .ZN(n7023) );
  AND2_X1 U5679 ( .A1(n7197), .A2(n8338), .ZN(n6875) );
  INV_X1 U5680 ( .A(n9863), .ZN(n8499) );
  AND2_X1 U5681 ( .A1(n6886), .A2(n5666), .ZN(n8500) );
  AND2_X1 U5682 ( .A1(n6822), .A2(n5940), .ZN(n6538) );
  AND2_X1 U5683 ( .A1(n5942), .A2(n5941), .ZN(n6533) );
  XNOR2_X1 U5684 ( .A(n5945), .B(n5944), .ZN(n6531) );
  NAND2_X1 U5685 ( .A1(n5588), .A2(n5587), .ZN(n7813) );
  NAND2_X1 U5686 ( .A1(n5578), .A2(n5577), .ZN(n8051) );
  NAND2_X1 U5687 ( .A1(n5537), .A2(n5536), .ZN(n8024) );
  NAND2_X1 U5688 ( .A1(n5525), .A2(n5524), .ZN(n8094) );
  NAND2_X1 U5689 ( .A1(n5440), .A2(n5439), .ZN(n9622) );
  AND2_X1 U5690 ( .A1(n9862), .A2(n9911), .ZN(n9922) );
  AND2_X1 U5691 ( .A1(n6831), .A2(n6721), .ZN(n6813) );
  NAND2_X1 U5692 ( .A1(n7334), .A2(n7484), .ZN(n9915) );
  AND3_X1 U5693 ( .A1(n5002), .A2(n4677), .A3(n5313), .ZN(n4676) );
  NOR2_X1 U5694 ( .A1(n4803), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4802) );
  NAND2_X1 U5695 ( .A1(n5188), .A2(n5192), .ZN(n4803) );
  NAND2_X1 U5696 ( .A1(n5640), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5645) );
  INV_X1 U5697 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5314) );
  INV_X1 U5698 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U5699 ( .A1(n6348), .A2(n6347), .ZN(n6361) );
  INV_X1 U5700 ( .A(n6349), .ZN(n6348) );
  NAND2_X1 U5701 ( .A1(n8837), .A2(n6339), .ZN(n4927) );
  AOI21_X1 U5702 ( .B1(n4922), .B2(n4921), .A(n4491), .ZN(n4920) );
  INV_X1 U5703 ( .A(n8742), .ZN(n4921) );
  INV_X1 U5704 ( .A(n6320), .ZN(n7926) );
  OR2_X1 U5705 ( .A1(n6361), .A2(n10016), .ZN(n6376) );
  INV_X1 U5706 ( .A(n9312), .ZN(n8952) );
  NAND2_X1 U5707 ( .A1(n6390), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6424) );
  INV_X1 U5708 ( .A(n6405), .ZN(n6390) );
  NOR2_X1 U5709 ( .A1(n4903), .A2(n4902), .ZN(n4901) );
  NOR2_X1 U5710 ( .A1(n8725), .A2(n4904), .ZN(n4902) );
  INV_X1 U5711 ( .A(n6416), .ZN(n4903) );
  NAND2_X1 U5712 ( .A1(n4901), .A2(n4904), .ZN(n4898) );
  INV_X1 U5714 ( .A(n6106), .ZN(n6104) );
  NAND2_X1 U5715 ( .A1(n8741), .A2(n8742), .ZN(n4925) );
  NAND2_X1 U5716 ( .A1(n4556), .A2(n4555), .ZN(n4554) );
  INV_X1 U5717 ( .A(n4557), .ZN(n4555) );
  INV_X1 U5718 ( .A(n4559), .ZN(n4556) );
  NAND2_X1 U5719 ( .A1(n4557), .A2(n4558), .ZN(n4552) );
  NAND2_X1 U5720 ( .A1(n4559), .A2(n8973), .ZN(n4553) );
  INV_X1 U5721 ( .A(n4561), .ZN(n4558) );
  NAND2_X1 U5722 ( .A1(n4729), .A2(n8971), .ZN(n8975) );
  OAI21_X1 U5723 ( .B1(n4575), .B2(n4572), .A(n4730), .ZN(n4729) );
  INV_X1 U5724 ( .A(n9046), .ZN(n4730) );
  AND3_X1 U5725 ( .A1(n6380), .A2(n6379), .A3(n6378), .ZN(n8795) );
  AND4_X1 U5726 ( .A1(n6204), .A2(n6203), .A3(n6202), .A4(n6201), .ZN(n8828)
         );
  AND4_X1 U5727 ( .A1(n6154), .A2(n6153), .A3(n6152), .A4(n6151), .ZN(n7548)
         );
  AND4_X1 U5728 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), .ZN(n7534)
         );
  NOR2_X1 U5729 ( .A1(n6709), .A2(n4601), .ZN(n6711) );
  AND2_X1 U5730 ( .A1(n6710), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4601) );
  NAND2_X1 U5731 ( .A1(n6711), .A2(n6712), .ZN(n6733) );
  NOR2_X1 U5732 ( .A1(n6852), .A2(n4602), .ZN(n6854) );
  AND2_X1 U5733 ( .A1(n6853), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4602) );
  NAND2_X1 U5734 ( .A1(n6854), .A2(n6855), .ZN(n6949) );
  NOR2_X1 U5735 ( .A1(n7379), .A2(n4596), .ZN(n7382) );
  AND2_X1 U5736 ( .A1(n7385), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4596) );
  NOR2_X1 U5737 ( .A1(n4595), .A2(n4594), .ZN(n9149) );
  INV_X1 U5738 ( .A(n7559), .ZN(n4594) );
  AOI21_X1 U5739 ( .B1(n7956), .B2(n8979), .A(n8959), .ZN(n4895) );
  NAND2_X1 U5740 ( .A1(n9240), .A2(n9461), .ZN(n4893) );
  INV_X1 U5741 ( .A(n9240), .ZN(n7914) );
  INV_X1 U5742 ( .A(n9489), .ZN(n7955) );
  NOR2_X1 U5743 ( .A1(n9289), .A2(n4711), .ZN(n9243) );
  INV_X1 U5744 ( .A(n4713), .ZN(n4711) );
  OR2_X1 U5745 ( .A1(n7948), .A2(n8959), .ZN(n9044) );
  NAND2_X1 U5746 ( .A1(n9134), .A2(n9461), .ZN(n4699) );
  NAND2_X1 U5747 ( .A1(n4970), .A2(n4434), .ZN(n4969) );
  INV_X1 U5748 ( .A(n4972), .ZN(n4970) );
  NAND2_X1 U5749 ( .A1(n4477), .A2(n4434), .ZN(n4968) );
  AND2_X1 U5750 ( .A1(n6514), .A2(n6460), .ZN(n9264) );
  AND2_X1 U5751 ( .A1(n6475), .A2(n6474), .ZN(n9257) );
  NAND2_X1 U5752 ( .A1(n4881), .A2(n4879), .ZN(n9273) );
  AND2_X1 U5753 ( .A1(n4880), .A2(n4882), .ZN(n4879) );
  NAND2_X1 U5754 ( .A1(n4881), .A2(n4882), .ZN(n9271) );
  NAND2_X1 U5755 ( .A1(n9368), .A2(n4706), .ZN(n9325) );
  OR2_X1 U5756 ( .A1(n6403), .A2(n6402), .ZN(n6405) );
  NAND2_X1 U5757 ( .A1(n6375), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6403) );
  INV_X1 U5758 ( .A(n6376), .ZN(n6375) );
  NAND2_X1 U5759 ( .A1(n4678), .A2(n4887), .ZN(n9320) );
  NAND2_X1 U5760 ( .A1(n4888), .A2(n8942), .ZN(n4887) );
  NAND2_X1 U5761 ( .A1(n9375), .A2(n4459), .ZN(n4678) );
  INV_X1 U5762 ( .A(n7912), .ZN(n4888) );
  NAND2_X1 U5763 ( .A1(n9368), .A2(n9588), .ZN(n9357) );
  NAND2_X1 U5764 ( .A1(n9375), .A2(n9096), .ZN(n9352) );
  OR2_X1 U5765 ( .A1(n6313), .A2(n10072), .ZN(n6349) );
  INV_X1 U5766 ( .A(n9422), .ZN(n9392) );
  NAND2_X1 U5767 ( .A1(n6312), .A2(n6311), .ZN(n7910) );
  AND2_X1 U5768 ( .A1(n8927), .A2(n8933), .ZN(n9402) );
  INV_X1 U5769 ( .A(n6291), .ZN(n6276) );
  NAND2_X1 U5770 ( .A1(n4688), .A2(n4440), .ZN(n9435) );
  AND2_X1 U5771 ( .A1(n4688), .A2(n8920), .ZN(n9436) );
  AND4_X1 U5772 ( .A1(n6282), .A2(n6281), .A3(n6280), .A4(n6279), .ZN(n9440)
         );
  NOR2_X1 U5773 ( .A1(n9473), .A2(n9437), .ZN(n4527) );
  INV_X1 U5774 ( .A(n9456), .ZN(n4528) );
  NAND2_X1 U5775 ( .A1(n7669), .A2(n4702), .ZN(n9467) );
  AND2_X1 U5776 ( .A1(n4435), .A2(n9790), .ZN(n4702) );
  NAND2_X1 U5777 ( .A1(n7669), .A2(n4435), .ZN(n9466) );
  INV_X1 U5778 ( .A(n9033), .ZN(n4877) );
  AND4_X1 U5779 ( .A1(n6231), .A2(n6230), .A3(n6229), .A4(n6228), .ZN(n8827)
         );
  INV_X1 U5780 ( .A(n6225), .ZN(n6223) );
  OR2_X1 U5781 ( .A1(n6200), .A2(n6801), .ZN(n6225) );
  AOI21_X1 U5782 ( .B1(n4685), .B2(n4687), .A(n4450), .ZN(n4684) );
  NAND2_X1 U5783 ( .A1(n7516), .A2(n4685), .ZN(n4683) );
  OAI21_X1 U5784 ( .B1(n7516), .B2(n4687), .A(n4685), .ZN(n9556) );
  NAND2_X1 U5785 ( .A1(n6185), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6200) );
  INV_X1 U5786 ( .A(n6198), .ZN(n6185) );
  AND4_X1 U5787 ( .A1(n6172), .A2(n6171), .A3(n6170), .A4(n6169), .ZN(n7518)
         );
  NAND2_X1 U5788 ( .A1(n7516), .A2(n7517), .ZN(n9554) );
  AOI21_X1 U5789 ( .B1(n7496), .B2(n4951), .A(n4471), .ZN(n4950) );
  INV_X1 U5790 ( .A(n7492), .ZN(n4951) );
  NAND2_X1 U5791 ( .A1(n9067), .A2(n8890), .ZN(n7600) );
  NAND2_X1 U5792 ( .A1(n4544), .A2(n4949), .ZN(n8886) );
  INV_X1 U5793 ( .A(n7600), .ZN(n4544) );
  AND2_X1 U5794 ( .A1(n7606), .A2(n7611), .ZN(n7604) );
  OAI21_X1 U5795 ( .B1(n4582), .B2(n4580), .A(n4579), .ZN(n7227) );
  INV_X1 U5796 ( .A(n9063), .ZN(n4580) );
  AND2_X1 U5797 ( .A1(n4576), .A2(n7226), .ZN(n4579) );
  OR2_X1 U5798 ( .A1(n7045), .A2(n7049), .ZN(n7232) );
  NAND2_X1 U5799 ( .A1(n6088), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6106) );
  INV_X1 U5800 ( .A(n6089), .ZN(n6088) );
  NAND2_X1 U5801 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6089) );
  NAND2_X1 U5802 ( .A1(n4578), .A2(n9063), .ZN(n8889) );
  NAND2_X1 U5803 ( .A1(n4582), .A2(n4581), .ZN(n4578) );
  INV_X1 U5804 ( .A(n4577), .ZN(n4581) );
  INV_X1 U5805 ( .A(n7039), .ZN(n4945) );
  NAND2_X1 U5806 ( .A1(n7000), .A2(n9762), .ZN(n7045) );
  INV_X1 U5807 ( .A(n8880), .ZN(n4682) );
  NAND2_X1 U5808 ( .A1(n7493), .A2(n7496), .ZN(n7521) );
  NAND2_X1 U5809 ( .A1(n7597), .A2(n7492), .ZN(n7493) );
  INV_X1 U5810 ( .A(n6973), .ZN(n9739) );
  AND2_X1 U5811 ( .A1(n4982), .A2(n4692), .ZN(n4691) );
  AND2_X1 U5812 ( .A1(n5967), .A2(n5970), .ZN(n4692) );
  NAND2_X1 U5813 ( .A1(n4693), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6006) );
  XNOR2_X1 U5814 ( .A(n5597), .B(n5596), .ZN(n7965) );
  INV_X1 U5815 ( .A(n5981), .ZN(n5982) );
  XNOR2_X1 U5816 ( .A(n5585), .B(n5586), .ZN(n7782) );
  INV_X1 U5817 ( .A(n4757), .ZN(n4756) );
  OAI21_X1 U5818 ( .B1(n4757), .B2(n4755), .A(n5131), .ZN(n4754) );
  INV_X1 U5819 ( .A(n5126), .ZN(n4755) );
  NAND2_X1 U5820 ( .A1(n4718), .A2(n4721), .ZN(n5408) );
  NAND2_X1 U5821 ( .A1(n4720), .A2(n4719), .ZN(n4718) );
  NAND2_X1 U5822 ( .A1(n4724), .A2(n5081), .ZN(n5403) );
  NAND2_X1 U5823 ( .A1(n5078), .A2(n4725), .ZN(n4724) );
  NAND2_X1 U5824 ( .A1(n5064), .A2(SI_7_), .ZN(n5065) );
  NAND2_X1 U5825 ( .A1(n5071), .A2(n5070), .ZN(n5357) );
  XNOR2_X1 U5826 ( .A(n5059), .B(SI_6_), .ZN(n5329) );
  XNOR2_X1 U5827 ( .A(n5055), .B(SI_5_), .ZN(n5316) );
  XNOR2_X1 U5828 ( .A(n5051), .B(SI_4_), .ZN(n5302) );
  AND2_X1 U5829 ( .A1(n6095), .A2(n6078), .ZN(n6636) );
  XNOR2_X1 U5830 ( .A(n5047), .B(SI_3_), .ZN(n5286) );
  OR2_X1 U5831 ( .A1(n6824), .A2(n6573), .ZN(n7124) );
  INV_X1 U5832 ( .A(n4984), .ZN(n7686) );
  AND2_X1 U5833 ( .A1(n5623), .A2(n5622), .ZN(n7973) );
  NAND2_X1 U5834 ( .A1(n8084), .A2(n5017), .ZN(n7987) );
  NAND2_X1 U5835 ( .A1(n5559), .A2(n5558), .ZN(n8420) );
  NOR2_X1 U5836 ( .A1(n8007), .A2(n8008), .ZN(n5013) );
  AND4_X1 U5837 ( .A1(n5531), .A2(n5530), .A3(n5529), .A4(n5528), .ZN(n8450)
         );
  AND3_X1 U5838 ( .A1(n5574), .A2(n5573), .A3(n5572), .ZN(n8417) );
  INV_X1 U5839 ( .A(n8175), .ZN(n8102) );
  AND2_X1 U5840 ( .A1(n6887), .A2(n6886), .ZN(n8172) );
  AND2_X1 U5841 ( .A1(n7401), .A2(n7398), .ZN(n7399) );
  INV_X1 U5842 ( .A(n8119), .ZN(n8170) );
  NAND2_X1 U5843 ( .A1(n7065), .A2(n7595), .ZN(n8179) );
  NAND2_X1 U5844 ( .A1(n5595), .A2(n5594), .ZN(n8389) );
  INV_X1 U5845 ( .A(n8417), .ZN(n8388) );
  INV_X1 U5846 ( .A(n8038), .ZN(n8195) );
  NAND4_X1 U5847 ( .A1(n5369), .A2(n5368), .A3(n5367), .A4(n5366), .ZN(n8197)
         );
  NAND4_X1 U5848 ( .A1(n5355), .A2(n5354), .A3(n5353), .A4(n5352), .ZN(n8198)
         );
  NAND4_X1 U5849 ( .A1(n5341), .A2(n5340), .A3(n5339), .A4(n5338), .ZN(n8199)
         );
  OR2_X1 U5850 ( .A1(n5291), .A2(n7141), .ZN(n5256) );
  AND2_X1 U5851 ( .A1(n5255), .A2(n5254), .ZN(n5258) );
  NAND2_X1 U5852 ( .A1(n4856), .A2(n4858), .ZN(n7288) );
  INV_X1 U5853 ( .A(n4853), .ZN(n4856) );
  INV_X1 U5854 ( .A(n4812), .ZN(n9841) );
  OR2_X1 U5855 ( .A1(P2_U3150), .A2(n7154), .ZN(n8341) );
  INV_X1 U5856 ( .A(n4851), .ZN(n7712) );
  XNOR2_X1 U5857 ( .A(n7727), .B(n7632), .ZN(n7633) );
  OAI21_X1 U5858 ( .B1(n7635), .B2(n4849), .A(n4848), .ZN(n7789) );
  NAND2_X1 U5859 ( .A1(n4852), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4849) );
  NAND2_X1 U5860 ( .A1(n7713), .A2(n4852), .ZN(n4848) );
  INV_X1 U5861 ( .A(n7715), .ZN(n4852) );
  INV_X1 U5862 ( .A(n7713), .ZN(n4850) );
  INV_X1 U5863 ( .A(n4868), .ZN(n8206) );
  INV_X1 U5864 ( .A(n4831), .ZN(n8212) );
  OR2_X1 U5865 ( .A1(n7790), .A2(n7793), .ZN(n4868) );
  INV_X1 U5866 ( .A(n8207), .ZN(n4867) );
  INV_X1 U5867 ( .A(n8211), .ZN(n4830) );
  OAI21_X1 U5868 ( .B1(n7790), .B2(n4866), .A(n4865), .ZN(n8242) );
  NAND2_X1 U5869 ( .A1(n4869), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4866) );
  NAND2_X1 U5870 ( .A1(n8207), .A2(n4869), .ZN(n4865) );
  INV_X1 U5871 ( .A(n8209), .ZN(n4869) );
  INV_X1 U5872 ( .A(n4876), .ZN(n4872) );
  NAND2_X1 U5873 ( .A1(n4820), .A2(n4818), .ZN(n8277) );
  INV_X1 U5874 ( .A(n8255), .ZN(n4817) );
  AOI21_X1 U5875 ( .B1(n4517), .B2(n4516), .A(n9844), .ZN(n8281) );
  NAND2_X1 U5876 ( .A1(n8280), .A2(n8283), .ZN(n4516) );
  INV_X1 U5877 ( .A(n8301), .ZN(n4517) );
  INV_X1 U5878 ( .A(n9855), .ZN(n9819) );
  NAND2_X1 U5879 ( .A1(n5917), .A2(n5916), .ZN(n5918) );
  NOR2_X1 U5880 ( .A1(n6560), .A2(n6559), .ZN(n6561) );
  NOR2_X1 U5881 ( .A1(n8378), .A2(n9865), .ZN(n6559) );
  INV_X1 U5882 ( .A(n4509), .ZN(n4508) );
  XNOR2_X1 U5883 ( .A(n8377), .B(n8379), .ZN(n4510) );
  OAI22_X1 U5884 ( .A1(n8378), .A2(n9863), .B1(n9865), .B2(n8402), .ZN(n4509)
         );
  NAND2_X1 U5885 ( .A1(n4667), .A2(n4665), .ZN(n8380) );
  INV_X1 U5886 ( .A(n4668), .ZN(n4665) );
  NAND2_X1 U5887 ( .A1(n8410), .A2(n4670), .ZN(n4667) );
  AND2_X1 U5888 ( .A1(n5569), .A2(n5568), .ZN(n8398) );
  NAND2_X1 U5889 ( .A1(n4652), .A2(n4653), .ZN(n8443) );
  OR2_X1 U5890 ( .A1(n8479), .A2(n4655), .ZN(n4652) );
  NAND2_X1 U5891 ( .A1(n8594), .A2(n5743), .ZN(n8457) );
  NAND2_X1 U5892 ( .A1(n4800), .A2(n5897), .ZN(n8460) );
  NAND2_X1 U5893 ( .A1(n8479), .A2(n8478), .ZN(n8594) );
  NAND2_X1 U5894 ( .A1(n5513), .A2(n5512), .ZN(n8477) );
  NAND2_X1 U5895 ( .A1(n5500), .A2(n5499), .ZN(n8599) );
  NAND2_X1 U5896 ( .A1(n5469), .A2(n5468), .ZN(n8609) );
  NAND2_X1 U5897 ( .A1(n4801), .A2(n5889), .ZN(n8512) );
  AND2_X1 U5898 ( .A1(n5434), .A2(n5433), .ZN(n8550) );
  INV_X1 U5899 ( .A(n8117), .ZN(n9623) );
  NAND2_X1 U5900 ( .A1(n4805), .A2(n5882), .ZN(n7807) );
  NOR2_X1 U5901 ( .A1(n4646), .A2(n4645), .ZN(n7757) );
  INV_X1 U5902 ( .A(n5704), .ZN(n4645) );
  NAND2_X1 U5903 ( .A1(n4626), .A2(n4625), .ZN(n7997) );
  AND2_X1 U5904 ( .A1(n5393), .A2(n4479), .ZN(n4625) );
  NAND2_X1 U5905 ( .A1(n6602), .A2(n5610), .ZN(n4626) );
  INV_X1 U5906 ( .A(n8524), .ZN(n8534) );
  INV_X1 U5907 ( .A(n5946), .ZN(n6841) );
  NAND2_X1 U5908 ( .A1(n5200), .A2(n5199), .ZN(n8622) );
  OR2_X1 U5909 ( .A1(n9611), .A2(n5288), .ZN(n5629) );
  NAND2_X1 U5910 ( .A1(n8564), .A2(n8563), .ZN(n8627) );
  INV_X1 U5911 ( .A(n8398), .ZN(n8638) );
  NAND2_X1 U5912 ( .A1(n5547), .A2(n5546), .ZN(n8646) );
  NAND2_X1 U5913 ( .A1(n5483), .A2(n5482), .ZN(n8660) );
  INV_X1 U5914 ( .A(n7343), .ZN(n7335) );
  AND2_X1 U5915 ( .A1(n5927), .A2(n5926), .ZN(n6616) );
  AND2_X1 U5916 ( .A1(n6824), .A2(n6834), .ZN(n6721) );
  AND2_X1 U5917 ( .A1(n6574), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6834) );
  INV_X1 U5918 ( .A(n5923), .ZN(n7784) );
  NOR2_X1 U5919 ( .A1(n4632), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6622) );
  INV_X1 U5920 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6603) );
  INV_X1 U5921 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6601) );
  AND2_X1 U5922 ( .A1(n5313), .A2(n5002), .ZN(n5372) );
  INV_X1 U5923 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10203) );
  INV_X1 U5924 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6593) );
  INV_X1 U5925 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6589) );
  INV_X1 U5926 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6588) );
  XNOR2_X1 U5927 ( .A(n5301), .B(n5300), .ZN(n7189) );
  OR2_X1 U5928 ( .A1(n6124), .A2(n6123), .ZN(n4931) );
  OR2_X1 U5929 ( .A1(n7475), .A2(n7309), .ZN(n4930) );
  NAND2_X1 U5930 ( .A1(n6103), .A2(n4465), .ZN(n4928) );
  NAND2_X1 U5931 ( .A1(n4927), .A2(n6340), .ZN(n8715) );
  NAND2_X1 U5932 ( .A1(n8790), .A2(n6372), .ZN(n8724) );
  NAND2_X1 U5933 ( .A1(n6374), .A2(n6373), .ZN(n9524) );
  NAND2_X1 U5934 ( .A1(n6274), .A2(n6273), .ZN(n9429) );
  NAND2_X1 U5935 ( .A1(n4489), .A2(n4918), .ZN(n8802) );
  NAND2_X1 U5936 ( .A1(n6328), .A2(n6327), .ZN(n9542) );
  NAND2_X1 U5937 ( .A1(n6103), .A2(n6102), .ZN(n4932) );
  NAND2_X1 U5938 ( .A1(n8845), .A2(n8844), .ZN(n4504) );
  NAND2_X1 U5939 ( .A1(n4925), .A2(n6455), .ZN(n8845) );
  NAND2_X1 U5940 ( .A1(n4925), .A2(n4922), .ZN(n8846) );
  INV_X1 U5941 ( .A(n8847), .ZN(n8858) );
  AOI21_X1 U5942 ( .B1(n8975), .B2(n4554), .A(n4551), .ZN(n9051) );
  NAND2_X1 U5943 ( .A1(n4779), .A2(n9119), .ZN(n9128) );
  NAND2_X1 U5944 ( .A1(n4782), .A2(n4780), .ZN(n4779) );
  INV_X1 U5945 ( .A(n9257), .ZN(n9134) );
  INV_X1 U5946 ( .A(n4680), .ZN(n4679) );
  NAND4_X2 U5947 ( .A1(n6017), .A2(n6016), .A3(n6015), .A4(n6014), .ZN(n6974)
         );
  OR2_X1 U5948 ( .A1(n8871), .A2(n6013), .ZN(n6014) );
  AND3_X1 U5949 ( .A1(n4606), .A2(n6028), .A3(n4604), .ZN(n9665) );
  NAND2_X1 U5950 ( .A1(n4476), .A2(P1_IR_REG_1__SCAN_IN), .ZN(n4606) );
  NAND2_X1 U5951 ( .A1(n4605), .A2(n5968), .ZN(n4604) );
  INV_X1 U5952 ( .A(n4600), .ZN(n6777) );
  AND2_X1 U5953 ( .A1(n4598), .A2(n4597), .ZN(n6695) );
  NAND2_X1 U5954 ( .A1(n6634), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4597) );
  NOR2_X1 U5955 ( .A1(n6668), .A2(n4488), .ZN(n6670) );
  NOR2_X1 U5956 ( .A1(n6670), .A2(n6669), .ZN(n6709) );
  NOR2_X1 U5957 ( .A1(n6791), .A2(n4603), .ZN(n6795) );
  AND2_X1 U5958 ( .A1(n6792), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4603) );
  NOR2_X1 U5959 ( .A1(n6795), .A2(n6794), .ZN(n6852) );
  XNOR2_X1 U5960 ( .A(n9149), .B(n9148), .ZN(n7560) );
  NAND2_X1 U5961 ( .A1(n4442), .A2(n9738), .ZN(n9477) );
  XNOR2_X1 U5962 ( .A(n4529), .B(n9254), .ZN(n9502) );
  NAND2_X1 U5963 ( .A1(n4971), .A2(n4973), .ZN(n4529) );
  NAND2_X1 U5964 ( .A1(n9310), .A2(n8981), .ZN(n9296) );
  NAND2_X1 U5965 ( .A1(n9353), .A2(n7912), .ZN(n9342) );
  AND2_X1 U5966 ( .A1(n4977), .A2(n4980), .ZN(n9350) );
  NAND2_X1 U5967 ( .A1(n7883), .A2(n5029), .ZN(n9367) );
  NAND2_X1 U5968 ( .A1(n6289), .A2(n6288), .ZN(n9452) );
  NAND2_X1 U5969 ( .A1(n6134), .A2(n6133), .ZN(n9705) );
  INV_X1 U5970 ( .A(n9736), .ZN(n9701) );
  NAND2_X1 U5971 ( .A1(n4582), .A2(n6991), .ZN(n7042) );
  NAND2_X1 U5972 ( .A1(n4944), .A2(n6998), .ZN(n7038) );
  NAND2_X1 U5973 ( .A1(n6969), .A2(n9061), .ZN(n6993) );
  AND2_X1 U5974 ( .A1(n9477), .A2(n9479), .ZN(n9562) );
  AND2_X1 U5975 ( .A1(n9492), .A2(n9491), .ZN(n9493) );
  AND2_X1 U5976 ( .A1(n6442), .A2(n6441), .ZN(n9580) );
  AOI211_X1 U5977 ( .C1(n9506), .C2(n9802), .A(n9505), .B(n9504), .ZN(n9577)
         );
  INV_X1 U5978 ( .A(n9705), .ZN(n7611) );
  INV_X1 U5979 ( .A(n7049), .ZN(n7322) );
  INV_X1 U5980 ( .A(n9788), .ZN(n9967) );
  OAI21_X1 U5981 ( .B1(n5198), .B2(n5197), .A(n5172), .ZN(n5175) );
  XNOR2_X1 U5982 ( .A(n5608), .B(n5609), .ZN(n8675) );
  NAND2_X1 U5983 ( .A1(n4768), .A2(n5158), .ZN(n5608) );
  XNOR2_X1 U5984 ( .A(n5557), .B(n5556), .ZN(n7594) );
  INV_X1 U5985 ( .A(n4751), .ZN(n5557) );
  AOI21_X1 U5986 ( .B1(n5535), .B2(n4756), .A(n4754), .ZN(n4751) );
  AND2_X1 U5987 ( .A1(P1_U3086), .A2(n4633), .ZN(n9608) );
  NAND2_X1 U5988 ( .A1(n5972), .A2(n5031), .ZN(n5978) );
  NAND2_X1 U5989 ( .A1(n5998), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4936) );
  INV_X1 U5990 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6605) );
  INV_X1 U5991 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6598) );
  INV_X1 U5992 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6594) );
  INV_X1 U5993 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9975) );
  INV_X1 U5994 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6591) );
  INV_X1 U5995 ( .A(n6636), .ZN(n6776) );
  INV_X1 U5996 ( .A(n9665), .ZN(n6641) );
  NAND2_X1 U5997 ( .A1(n4633), .A2(SI_0_), .ZN(n5957) );
  XNOR2_X1 U5998 ( .A(n4992), .B(n7868), .ZN(n7875) );
  NAND2_X1 U5999 ( .A1(n4520), .A2(n4518), .ZN(n5843) );
  NAND2_X1 U6000 ( .A1(n4821), .A2(n8254), .ZN(n8235) );
  AOI21_X1 U6001 ( .B1(n4438), .B2(n9830), .A(n4534), .ZN(n8349) );
  AND2_X1 U6002 ( .A1(n4833), .A2(n4834), .ZN(n8327) );
  OAI21_X1 U6003 ( .B1(n7962), .B2(n6581), .A(n4806), .ZN(P2_U3294) );
  INV_X1 U6004 ( .A(n4807), .ZN(n4806) );
  INV_X1 U6005 ( .A(n6529), .ZN(n4522) );
  INV_X1 U6006 ( .A(n4897), .ZN(n6766) );
  INV_X1 U6007 ( .A(n4598), .ZN(n6681) );
  OAI21_X1 U6008 ( .B1(n9492), .B2(n4419), .A(n4694), .ZN(P1_U3265) );
  INV_X1 U6009 ( .A(n4695), .ZN(n4694) );
  OAI21_X1 U6010 ( .B1(n9488), .B2(n9433), .A(n4696), .ZN(n4695) );
  AOI21_X1 U6011 ( .B1(n9490), .B2(n9348), .A(n7959), .ZN(n4696) );
  OAI21_X1 U6012 ( .B1(n9562), .B2(n9811), .A(n4700), .ZN(P1_U3553) );
  AOI21_X1 U6013 ( .B1(n9224), .B2(n9560), .A(n4701), .ZN(n4700) );
  NOR2_X1 U6014 ( .A1(n9814), .A2(n9478), .ZN(n4701) );
  AND2_X1 U6015 ( .A1(n4721), .A2(n5407), .ZN(n4432) );
  AND2_X1 U6016 ( .A1(n5890), .A2(n5889), .ZN(n4433) );
  OR2_X1 U6017 ( .A1(n9263), .A2(n9275), .ZN(n4434) );
  INV_X1 U6018 ( .A(n8892), .ZN(n4949) );
  AND2_X1 U6019 ( .A1(n4704), .A2(n4703), .ZN(n4435) );
  AND4_X1 U6020 ( .A1(n4728), .A2(n9048), .A3(n9108), .A4(n9047), .ZN(n4436)
         );
  OR2_X1 U6021 ( .A1(n7813), .A2(n8389), .ZN(n4437) );
  INV_X1 U6022 ( .A(n9318), .ZN(n4505) );
  XOR2_X1 U6023 ( .A(n8346), .B(n8345), .Z(n4438) );
  AND2_X1 U6024 ( .A1(n8561), .A2(n8186), .ZN(n4439) );
  AND2_X1 U6025 ( .A1(n9443), .A2(n8920), .ZN(n4440) );
  INV_X1 U6026 ( .A(n4449), .ZN(n4719) );
  NAND2_X1 U6027 ( .A1(n9223), .A2(n9132), .ZN(n4441) );
  XOR2_X1 U6028 ( .A(n9230), .B(n9224), .Z(n4442) );
  NAND2_X1 U6029 ( .A1(n9926), .A2(n8194), .ZN(n4443) );
  AND2_X1 U6030 ( .A1(n6031), .A2(n6032), .ZN(n4444) );
  OR2_X1 U6031 ( .A1(n9223), .A2(n9007), .ZN(n9108) );
  INV_X1 U6032 ( .A(n9108), .ZN(n4562) );
  AND2_X1 U6033 ( .A1(n8511), .A2(n5721), .ZN(n4445) );
  AND2_X1 U6034 ( .A1(n4802), .A2(n5226), .ZN(n4446) );
  AND2_X1 U6035 ( .A1(n9565), .A2(n9131), .ZN(n9012) );
  INV_X1 U6036 ( .A(n9012), .ZN(n4728) );
  NOR2_X1 U6037 ( .A1(n9370), .A2(n9135), .ZN(n7884) );
  AND2_X1 U6038 ( .A1(n4843), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4447) );
  INV_X1 U6039 ( .A(n5007), .ZN(n6872) );
  INV_X1 U6040 ( .A(n8511), .ZN(n5890) );
  INV_X1 U6041 ( .A(n8257), .ZN(n4822) );
  NAND2_X2 U6042 ( .A1(n5261), .A2(n5259), .ZN(n5288) );
  NAND2_X1 U6043 ( .A1(n6969), .A2(n4583), .ZN(n4582) );
  NAND2_X1 U6044 ( .A1(n5262), .A2(n6840), .ZN(n5656) );
  NAND2_X1 U6045 ( .A1(n5974), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6326) );
  NAND4_X1 U6046 ( .A1(n5384), .A2(n5383), .A3(n5382), .A4(n5381), .ZN(n8196)
         );
  INV_X1 U6047 ( .A(n8196), .ZN(n8036) );
  AND2_X1 U6048 ( .A1(n5314), .A2(n5005), .ZN(n4448) );
  NAND2_X1 U6049 ( .A1(n5313), .A2(n5004), .ZN(n5343) );
  INV_X1 U6050 ( .A(n8973), .ZN(n4731) );
  OR2_X1 U6051 ( .A1(n5402), .A2(n4723), .ZN(n4449) );
  AND2_X1 U6052 ( .A1(n5385), .A2(n5178), .ZN(n5388) );
  AOI21_X1 U6053 ( .B1(n8410), .B2(n4457), .A(n4659), .ZN(n4658) );
  OR2_X1 U6054 ( .A1(n7745), .A2(n7660), .ZN(n4450) );
  NAND2_X1 U6055 ( .A1(n5388), .A2(n5179), .ZN(n5409) );
  NAND2_X1 U6056 ( .A1(n5385), .A2(n5018), .ZN(n4451) );
  NAND2_X1 U6057 ( .A1(n6470), .A2(n6469), .ZN(n9245) );
  AND2_X1 U6058 ( .A1(n5923), .A2(n5009), .ZN(n4452) );
  AND4_X1 U6059 ( .A1(n5705), .A2(n5941), .A3(n5685), .A4(n5684), .ZN(n4453)
         );
  NAND2_X1 U6060 ( .A1(n6389), .A2(n6388), .ZN(n9514) );
  INV_X1 U6061 ( .A(n9514), .ZN(n4705) );
  OR2_X1 U6062 ( .A1(n5261), .A2(n4808), .ZN(n4454) );
  OR3_X1 U6063 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n4455) );
  OR2_X1 U6064 ( .A1(n9762), .A2(n9144), .ZN(n4456) );
  AND2_X1 U6065 ( .A1(n4662), .A2(n4661), .ZN(n4457) );
  INV_X1 U6066 ( .A(n7143), .ZN(n4815) );
  OR2_X1 U6067 ( .A1(n4846), .A2(n9843), .ZN(n4458) );
  AND2_X1 U6068 ( .A1(n8942), .A2(n4889), .ZN(n4459) );
  OR2_X1 U6069 ( .A1(n8638), .A2(n8417), .ZN(n5825) );
  INV_X1 U6070 ( .A(n5825), .ZN(n4671) );
  INV_X1 U6071 ( .A(n5896), .ZN(n8478) );
  NAND2_X1 U6072 ( .A1(n6401), .A2(n6400), .ZN(n9521) );
  OR2_X1 U6073 ( .A1(n8196), .A2(n7997), .ZN(n4460) );
  AND2_X1 U6074 ( .A1(n7813), .A2(n8389), .ZN(n4461) );
  NAND2_X1 U6075 ( .A1(n4946), .A2(n6027), .ZN(n6075) );
  NAND2_X1 U6076 ( .A1(n5313), .A2(n5314), .ZN(n5327) );
  AND2_X1 U6077 ( .A1(n7827), .A2(n8194), .ZN(n4462) );
  NOR2_X1 U6078 ( .A1(n8301), .A2(n8302), .ZN(n4463) );
  INV_X1 U6079 ( .A(n9223), .ZN(n8974) );
  NAND2_X1 U6080 ( .A1(n8882), .A2(n8881), .ZN(n9223) );
  XNOR2_X1 U6081 ( .A(n5088), .B(SI_12_), .ZN(n5407) );
  INV_X1 U6082 ( .A(n4741), .ZN(n4740) );
  NAND2_X1 U6083 ( .A1(n4745), .A2(n4742), .ZN(n4741) );
  INV_X1 U6084 ( .A(n9360), .ZN(n9588) );
  NAND2_X1 U6085 ( .A1(n6360), .A2(n6359), .ZN(n9360) );
  AND2_X1 U6086 ( .A1(n4827), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4464) );
  NAND2_X1 U6087 ( .A1(n9368), .A2(n4708), .ZN(n4709) );
  INV_X1 U6088 ( .A(n8738), .ZN(n9780) );
  NOR2_X1 U6089 ( .A1(n9287), .A2(n4886), .ZN(n4885) );
  AND2_X1 U6090 ( .A1(n9224), .A2(n9227), .ZN(n9053) );
  INV_X1 U6091 ( .A(n4962), .ZN(n4961) );
  NAND2_X1 U6092 ( .A1(n7666), .A2(n4422), .ZN(n4962) );
  AND2_X1 U6093 ( .A1(n4929), .A2(n6102), .ZN(n4465) );
  AND2_X1 U6094 ( .A1(n4873), .A2(n4872), .ZN(n4466) );
  AND2_X1 U6095 ( .A1(n4831), .A2(n4830), .ZN(n4467) );
  NOR2_X1 U6096 ( .A1(n9289), .A2(n4712), .ZN(n4710) );
  NAND2_X1 U6097 ( .A1(n5077), .A2(n5075), .ZN(n5370) );
  OR2_X1 U6098 ( .A1(n9790), .A2(n8861), .ZN(n4468) );
  OR2_X1 U6099 ( .A1(n9489), .A2(n7914), .ZN(n8979) );
  AND2_X1 U6100 ( .A1(n4817), .A2(n8254), .ZN(n4469) );
  OR2_X1 U6101 ( .A1(n8024), .A2(n8464), .ZN(n5802) );
  NAND3_X1 U6102 ( .A1(n5841), .A2(n5840), .A3(n5839), .ZN(n4470) );
  INV_X1 U6103 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5968) );
  NOR2_X1 U6104 ( .A1(n7779), .A2(n9140), .ZN(n4471) );
  NAND2_X1 U6105 ( .A1(n8869), .A2(n8868), .ZN(n9224) );
  NAND2_X1 U6106 ( .A1(n5073), .A2(n5072), .ZN(n5077) );
  INV_X1 U6107 ( .A(n5077), .ZN(n4726) );
  NOR2_X1 U6108 ( .A1(n7813), .A2(n7863), .ZN(n4472) );
  NAND2_X1 U6109 ( .A1(n5313), .A2(n4448), .ZN(n4473) );
  AND2_X1 U6110 ( .A1(n5102), .A2(SI_16_), .ZN(n4474) );
  INV_X1 U6111 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10001) );
  INV_X1 U6112 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5179) );
  INV_X1 U6113 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5178) );
  INV_X1 U6114 ( .A(n4923), .ZN(n4922) );
  OR2_X1 U6115 ( .A1(n8844), .A2(n4924), .ZN(n4923) );
  AND2_X1 U6116 ( .A1(n5089), .A2(SI_12_), .ZN(n4475) );
  OR2_X1 U6117 ( .A1(n9473), .A2(n8861), .ZN(n8920) );
  AND2_X1 U6118 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4476) );
  INV_X1 U6119 ( .A(n6476), .ZN(n4538) );
  INV_X1 U6120 ( .A(n9082), .ZN(n4690) );
  AND2_X1 U6121 ( .A1(n5735), .A2(n5733), .ZN(n8511) );
  NAND2_X1 U6122 ( .A1(n7893), .A2(n4973), .ZN(n4477) );
  NOR2_X1 U6123 ( .A1(n7891), .A2(n4974), .ZN(n4478) );
  OR2_X1 U6124 ( .A1(n4415), .A2(n7638), .ZN(n4479) );
  INV_X1 U6125 ( .A(n9270), .ZN(n4880) );
  INV_X2 U6126 ( .A(n6880), .ZN(n7069) );
  INV_X1 U6128 ( .A(n5695), .ZN(n4612) );
  AND2_X1 U6129 ( .A1(n4911), .A2(n8683), .ZN(n4480) );
  AND2_X1 U6130 ( .A1(n6420), .A2(n4898), .ZN(n4481) );
  INV_X1 U6131 ( .A(n9263), .ZN(n9576) );
  NAND2_X1 U6132 ( .A1(n6457), .A2(n6456), .ZN(n9263) );
  AND2_X1 U6133 ( .A1(n4706), .A2(n4705), .ZN(n4482) );
  AND2_X1 U6134 ( .A1(n8991), .A2(n8957), .ZN(n9238) );
  NAND2_X1 U6135 ( .A1(n6039), .A2(n6038), .ZN(n4483) );
  NAND2_X1 U6136 ( .A1(n5599), .A2(n5598), .ZN(n8561) );
  AND2_X1 U6137 ( .A1(n5898), .A2(n5897), .ZN(n4484) );
  AND2_X1 U6138 ( .A1(n4728), .A2(n4727), .ZN(n4485) );
  AND2_X1 U6139 ( .A1(n4985), .A2(n4987), .ZN(n4486) );
  NAND2_X1 U6140 ( .A1(n7268), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4487) );
  INV_X1 U6141 ( .A(n5016), .ZN(n5015) );
  NAND2_X1 U6142 ( .A1(n7068), .A2(n8203), .ZN(n5016) );
  INV_X1 U6143 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U6144 ( .A1(n5629), .A2(n5628), .ZN(n6554) );
  INV_X1 U6145 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4507) );
  AND2_X1 U6146 ( .A1(n6671), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4488) );
  INV_X1 U6147 ( .A(n4910), .ZN(n8681) );
  INV_X1 U6148 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5005) );
  NAND2_X1 U6149 ( .A1(n7676), .A2(n4647), .ZN(n7756) );
  OR2_X1 U6150 ( .A1(n8732), .A2(n8731), .ZN(n4489) );
  AND2_X1 U6151 ( .A1(n8920), .A2(n8915), .ZN(n4490) );
  INV_X1 U6152 ( .A(n8186), .ZN(n8378) );
  NAND2_X1 U6153 ( .A1(n5607), .A2(n5606), .ZN(n8186) );
  AND2_X1 U6154 ( .A1(n6468), .A2(n6467), .ZN(n4491) );
  NOR2_X1 U6155 ( .A1(n7456), .A2(n7455), .ZN(n4492) );
  INV_X1 U6156 ( .A(n9370), .ZN(n9592) );
  NAND2_X1 U6157 ( .A1(n6344), .A2(n6343), .ZN(n9370) );
  NAND2_X1 U6158 ( .A1(n6258), .A2(n6257), .ZN(n9473) );
  NOR2_X1 U6159 ( .A1(n9360), .A2(n9380), .ZN(n4493) );
  AND2_X1 U6160 ( .A1(n4868), .A2(n4867), .ZN(n4494) );
  AND2_X1 U6161 ( .A1(n4851), .A2(n4850), .ZN(n4495) );
  NOR2_X1 U6162 ( .A1(n7382), .A2(n7381), .ZN(n4595) );
  AND4_X1 U6163 ( .A1(n6191), .A2(n6190), .A3(n6189), .A4(n6188), .ZN(n7668)
         );
  INV_X1 U6164 ( .A(n7668), .ZN(n4957) );
  NAND2_X1 U6165 ( .A1(n5972), .A2(n4983), .ZN(n4496) );
  INV_X1 U6166 ( .A(n4975), .ZN(n4974) );
  NAND2_X1 U6167 ( .A1(n5972), .A2(n4939), .ZN(n4497) );
  AND2_X1 U6168 ( .A1(n7866), .A2(n8186), .ZN(n4498) );
  OR2_X1 U6169 ( .A1(n7461), .A2(n10185), .ZN(n4499) );
  NAND2_X1 U6170 ( .A1(n7838), .A2(n7837), .ZN(n8074) );
  AND2_X1 U6171 ( .A1(n5612), .A2(n5611), .ZN(n8362) );
  INV_X1 U6172 ( .A(n8362), .ZN(n7873) );
  INV_X1 U6173 ( .A(n7884), .ZN(n4980) );
  INV_X2 U6174 ( .A(n9929), .ZN(n9928) );
  INV_X1 U6175 ( .A(n7496), .ZN(n4952) );
  AND2_X2 U6176 ( .A1(n6538), .A2(n6537), .ZN(n9941) );
  INV_X2 U6177 ( .A(n7899), .ZN(n8877) );
  NAND2_X1 U6178 ( .A1(n6242), .A2(n6241), .ZN(n8807) );
  INV_X1 U6179 ( .A(n8807), .ZN(n4703) );
  NAND2_X1 U6180 ( .A1(n4954), .A2(n4953), .ZN(n7746) );
  NAND2_X1 U6181 ( .A1(n5008), .A2(n6761), .ZN(n5007) );
  INV_X1 U6182 ( .A(n5014), .ZN(n8006) );
  NAND2_X1 U6183 ( .A1(n5013), .A2(n5012), .ZN(n5014) );
  AND2_X1 U6184 ( .A1(n4933), .A2(n4932), .ZN(n4500) );
  AND2_X1 U6185 ( .A1(n4847), .A2(n4846), .ZN(n4501) );
  XNOR2_X1 U6186 ( .A(n6006), .B(n5969), .ZN(n6525) );
  OR2_X1 U6187 ( .A1(n6934), .A2(n9056), .ZN(n9549) );
  INV_X1 U6188 ( .A(n9549), .ZN(n9738) );
  AND2_X1 U6189 ( .A1(n4826), .A2(n4825), .ZN(n4502) );
  AND2_X1 U6190 ( .A1(n4632), .A2(P2_U3151), .ZN(n4503) );
  XNOR2_X1 U6191 ( .A(n5510), .B(n5509), .ZN(n8333) );
  INV_X1 U6192 ( .A(n8333), .ZN(n8338) );
  INV_X1 U6193 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5985) );
  INV_X1 U6194 ( .A(n7197), .ZN(n6873) );
  XNOR2_X1 U6195 ( .A(n5645), .B(n5644), .ZN(n7197) );
  INV_X1 U6196 ( .A(n7287), .ZN(n4861) );
  AND2_X1 U6197 ( .A1(n7035), .A2(n7279), .ZN(n6754) );
  XNOR2_X1 U6198 ( .A(n4936), .B(n5995), .ZN(n9062) );
  INV_X1 U6199 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4764) );
  XNOR2_X1 U6200 ( .A(n8210), .B(n8216), .ZN(n7788) );
  INV_X1 U6201 ( .A(n8853), .ZN(n8864) );
  NAND2_X1 U6202 ( .A1(n4899), .A2(n4481), .ZN(n8769) );
  AOI21_X2 U6203 ( .B1(n8749), .B2(n6309), .A(n6308), .ZN(n8763) );
  NOR2_X2 U6204 ( .A1(n7771), .A2(n6159), .ZN(n8780) );
  NAND2_X1 U6205 ( .A1(n6157), .A2(n6156), .ZN(n6158) );
  XNOR2_X1 U6206 ( .A(n6050), .B(n4429), .ZN(n6052) );
  NAND2_X4 U6207 ( .A1(n6525), .A2(n9651), .ZN(n6607) );
  NAND3_X1 U6208 ( .A1(n4504), .A2(n8846), .A3(n8817), .ZN(n8852) );
  NAND2_X1 U6209 ( .A1(n8724), .A2(n8725), .ZN(n4900) );
  NAND2_X1 U6210 ( .A1(n4524), .A2(n8817), .ZN(n4523) );
  NAND2_X1 U6211 ( .A1(n9273), .A2(n9000), .ZN(n9253) );
  NAND2_X1 U6212 ( .A1(n9236), .A2(n8957), .ZN(n7956) );
  INV_X1 U6213 ( .A(n5078), .ZN(n4720) );
  NAND2_X1 U6214 ( .A1(n4684), .A2(n4683), .ZN(n7739) );
  INV_X1 U6215 ( .A(n7740), .ZN(n4878) );
  XNOR2_X1 U6216 ( .A(n4895), .B(n9046), .ZN(n4894) );
  NAND2_X1 U6217 ( .A1(n5270), .A2(n5269), .ZN(n5046) );
  INV_X1 U6218 ( .A(n7758), .ZN(n4515) );
  AOI21_X2 U6219 ( .B1(n8415), .B2(n5903), .A(n5902), .ZN(n8400) );
  NOR2_X1 U6220 ( .A1(n7204), .A2(n7205), .ZN(n7203) );
  NAND2_X1 U6221 ( .A1(n8256), .A2(n4822), .ZN(n4820) );
  AOI21_X1 U6222 ( .B1(n7284), .B2(n7184), .A(n7185), .ZN(n7183) );
  INV_X1 U6223 ( .A(n7148), .ZN(n4824) );
  NOR2_X1 U6224 ( .A1(n7146), .A2(n7145), .ZN(n7285) );
  NAND2_X1 U6225 ( .A1(n8211), .A2(n4832), .ZN(n4828) );
  AOI21_X1 U6226 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7795), .A(n7787), .ZN(
        n8210) );
  NOR2_X1 U6227 ( .A1(n7731), .A2(n7730), .ZN(n7734) );
  INV_X1 U6228 ( .A(n5229), .ZN(n5230) );
  NAND2_X1 U6229 ( .A1(n5872), .A2(n5871), .ZN(n7414) );
  NAND2_X1 U6230 ( .A1(n4794), .A2(n4798), .ZN(n8368) );
  AOI21_X1 U6231 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n7795), .A(n7789), .ZN(
        n8205) );
  OAI211_X2 U6232 ( .C1(n7310), .C2(n4930), .A(n4928), .B(n4931), .ZN(n7533)
         );
  NOR2_X1 U6233 ( .A1(n7772), .A2(n7773), .ZN(n7771) );
  AOI21_X1 U6234 ( .B1(n6894), .B2(n6893), .A(n5026), .ZN(n6941) );
  AOI21_X1 U6235 ( .B1(n8732), .B2(n4914), .A(n4912), .ZN(n4910) );
  NAND2_X1 U6236 ( .A1(n7946), .A2(n6499), .ZN(n4524) );
  NAND3_X1 U6237 ( .A1(n4946), .A2(n6026), .A3(n5958), .ZN(n6112) );
  NAND2_X1 U6238 ( .A1(n8791), .A2(n8792), .ZN(n8790) );
  NAND2_X1 U6239 ( .A1(n4523), .A2(n4522), .ZN(P1_U3214) );
  MUX2_X1 U6240 ( .A(n5761), .B(n5760), .S(n5666), .Z(n5765) );
  NAND2_X1 U6241 ( .A1(n8526), .A2(n4619), .ZN(n4618) );
  INV_X1 U6242 ( .A(n4616), .ZN(n4615) );
  NAND2_X1 U6243 ( .A1(n4636), .A2(n4635), .ZN(n4634) );
  NAND2_X1 U6244 ( .A1(n5303), .A2(n5302), .ZN(n5054) );
  INV_X1 U6245 ( .A(n5742), .ZN(n4639) );
  INV_X2 U6246 ( .A(n5194), .ZN(n5259) );
  INV_X1 U6247 ( .A(n6500), .ZN(n6000) );
  NAND2_X1 U6248 ( .A1(n6326), .A2(n5994), .ZN(n5996) );
  NAND2_X1 U6249 ( .A1(n4943), .A2(n5028), .ZN(n9414) );
  OAI21_X2 U6250 ( .B1(n4528), .B2(n4527), .A(n4468), .ZN(n9444) );
  NAND2_X1 U6251 ( .A1(n4963), .A2(n4968), .ZN(n9235) );
  AOI211_X1 U6252 ( .C1(n9497), .C2(n9802), .A(n9496), .B(n9495), .ZN(n9571)
         );
  NAND2_X1 U6253 ( .A1(n9444), .A2(n7878), .ZN(n4943) );
  XNOR2_X2 U6254 ( .A(n6965), .B(n4530), .ZN(n9730) );
  AOI21_X2 U6255 ( .B1(n4777), .B2(n4681), .A(n4531), .ZN(n4593) );
  NAND2_X1 U6256 ( .A1(n7285), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7284) );
  AOI21_X1 U6257 ( .B1(n6143), .B2(n6142), .A(n5027), .ZN(n6157) );
  NAND2_X1 U6258 ( .A1(n6996), .A2(n9015), .ZN(n4944) );
  AOI211_X1 U6259 ( .C1(n9502), .C2(n9802), .A(n9501), .B(n9500), .ZN(n9574)
         );
  INV_X2 U6260 ( .A(n6965), .ZN(n9749) );
  NAND2_X2 U6261 ( .A1(n4593), .A2(n4592), .ZN(n6965) );
  OAI21_X2 U6262 ( .B1(n8741), .B2(n4923), .A(n4920), .ZN(n6481) );
  NAND2_X1 U6263 ( .A1(n5981), .A2(n5967), .ZN(n4545) );
  NAND2_X1 U6264 ( .A1(n6973), .A2(n4538), .ZN(n6019) );
  NAND2_X1 U6265 ( .A1(n8724), .A2(n4901), .ZN(n4899) );
  NAND2_X1 U6266 ( .A1(n8975), .A2(n4548), .ZN(n4547) );
  NAND2_X1 U6267 ( .A1(n4563), .A2(n4564), .ZN(n8903) );
  NAND3_X1 U6268 ( .A1(n8902), .A2(n4490), .A3(n4567), .ZN(n4563) );
  NAND2_X1 U6269 ( .A1(n8910), .A2(n9081), .ZN(n4571) );
  MUX2_X1 U6270 ( .A(n6030), .B(P1_REG2_REG_1__SCAN_IN), .S(n9665), .Z(n9662)
         );
  NAND2_X1 U6271 ( .A1(n4607), .A2(n5712), .ZN(n5714) );
  NAND2_X1 U6272 ( .A1(n4608), .A2(n5419), .ZN(n4607) );
  NAND3_X1 U6273 ( .A1(n4613), .A2(n5709), .A3(n4609), .ZN(n4608) );
  NAND2_X1 U6274 ( .A1(n4453), .A2(n4610), .ZN(n4609) );
  NAND2_X1 U6275 ( .A1(n4612), .A2(n4611), .ZN(n4610) );
  NAND2_X1 U6276 ( .A1(n5699), .A2(n5700), .ZN(n4613) );
  NAND2_X1 U6277 ( .A1(n5717), .A2(n4617), .ZN(n4614) );
  NAND2_X1 U6278 ( .A1(n4614), .A2(n4615), .ZN(n5722) );
  INV_X1 U6279 ( .A(n5720), .ZN(n4622) );
  AOI21_X2 U6280 ( .B1(n5799), .B2(n5798), .A(n5832), .ZN(n4624) );
  NAND2_X1 U6281 ( .A1(n4629), .A2(n5071), .ZN(n5371) );
  NAND2_X1 U6282 ( .A1(n5066), .A2(n5065), .ZN(n5359) );
  MUX2_X1 U6283 ( .A(n6591), .B(n6589), .S(n5259), .Z(n5055) );
  MUX2_X1 U6284 ( .A(n9975), .B(n6593), .S(n5259), .Z(n5059) );
  MUX2_X1 U6285 ( .A(n6594), .B(n10203), .S(n5259), .Z(n5063) );
  MUX2_X1 U6286 ( .A(n6598), .B(n6596), .S(n5259), .Z(n5068) );
  MUX2_X1 U6287 ( .A(n6605), .B(n6603), .S(n5259), .Z(n5079) );
  MUX2_X1 U6288 ( .A(n6612), .B(n10163), .S(n5259), .Z(n5084) );
  MUX2_X1 U6289 ( .A(n6599), .B(n6601), .S(n5259), .Z(n5073) );
  MUX2_X1 U6290 ( .A(n10178), .B(n6619), .S(n4632), .Z(n5088) );
  MUX2_X1 U6291 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n4632), .Z(n5448) );
  MUX2_X1 U6292 ( .A(n10042), .B(n6765), .S(n4632), .Z(n5463) );
  MUX2_X1 U6293 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n4632), .Z(n5091) );
  MUX2_X1 U6294 ( .A(n10187), .B(n6838), .S(n4632), .Z(n5105) );
  MUX2_X1 U6295 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n4632), .Z(n5095) );
  MUX2_X1 U6296 ( .A(n5109), .B(n6901), .S(n4632), .Z(n5110) );
  MUX2_X1 U6297 ( .A(n7487), .B(n7485), .S(n4632), .Z(n5128) );
  MUX2_X1 U6298 ( .A(n10232), .B(n9971), .S(n4632), .Z(n5533) );
  MUX2_X1 U6299 ( .A(n7037), .B(n7034), .S(n4632), .Z(n5114) );
  MUX2_X1 U6300 ( .A(n7593), .B(n9986), .S(n4632), .Z(n5133) );
  MUX2_X1 U6301 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n4632), .Z(n5521) );
  MUX2_X1 U6302 ( .A(n7683), .B(n7769), .S(n4632), .Z(n5138) );
  MUX2_X1 U6303 ( .A(n10015), .B(n7766), .S(n4632), .Z(n5144) );
  MUX2_X1 U6304 ( .A(n9615), .B(n7966), .S(n4632), .Z(n5155) );
  MUX2_X1 U6305 ( .A(n10008), .B(n7783), .S(n4632), .Z(n5149) );
  MUX2_X1 U6306 ( .A(n7894), .B(n8678), .S(n4632), .Z(n5160) );
  MUX2_X1 U6307 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n4632), .Z(n5164) );
  MUX2_X1 U6308 ( .A(n8879), .B(n7960), .S(n4632), .Z(n5169) );
  MUX2_X1 U6309 ( .A(n9604), .B(n8671), .S(n4632), .Z(n5173) );
  NAND2_X2 U6310 ( .A1(n6607), .A2(n4633), .ZN(n7899) );
  NAND3_X1 U6311 ( .A1(n4639), .A2(n4638), .A3(n4637), .ZN(n4636) );
  NAND2_X2 U6312 ( .A1(n5654), .A2(n5657), .ZN(n5859) );
  INV_X1 U6313 ( .A(n4641), .ZN(n5251) );
  OR2_X1 U6314 ( .A1(n5288), .A2(n6581), .ZN(n5861) );
  OR2_X1 U6315 ( .A1(n4430), .A2(n5039), .ZN(n5862) );
  NAND3_X1 U6316 ( .A1(n5434), .A2(n5433), .A3(n8551), .ZN(n8549) );
  NAND2_X1 U6317 ( .A1(n5462), .A2(n4445), .ZN(n8519) );
  NAND2_X1 U6318 ( .A1(n8519), .A2(n5733), .ZN(n8508) );
  NAND2_X1 U6319 ( .A1(n5462), .A2(n5721), .ZN(n8521) );
  OAI21_X2 U6320 ( .B1(n7677), .B2(n4644), .A(n4642), .ZN(n7805) );
  NAND2_X1 U6321 ( .A1(n8479), .A2(n4650), .ZN(n4649) );
  INV_X1 U6322 ( .A(n4658), .ZN(n6557) );
  NAND3_X1 U6323 ( .A1(n4662), .A2(n4664), .A3(n4661), .ZN(n4660) );
  NAND2_X1 U6324 ( .A1(n4673), .A2(n5271), .ZN(n5283) );
  NAND2_X1 U6325 ( .A1(n5249), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6326 ( .A1(n4673), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7161) );
  NAND2_X1 U6327 ( .A1(n4673), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7143) );
  NAND2_X1 U6328 ( .A1(n4675), .A2(n5018), .ZN(n5191) );
  INV_X1 U6329 ( .A(n5189), .ZN(n5851) );
  NAND2_X2 U6330 ( .A1(n9376), .A2(n9377), .ZN(n9375) );
  NAND2_X1 U6331 ( .A1(n7909), .A2(n4689), .ZN(n4688) );
  NAND3_X1 U6332 ( .A1(n4983), .A2(n4691), .A3(n5972), .ZN(n4693) );
  INV_X1 U6333 ( .A(n4693), .ZN(n6003) );
  NOR2_X2 U6334 ( .A1(n9721), .A2(n6987), .ZN(n7000) );
  NAND2_X1 U6335 ( .A1(n9368), .A2(n4482), .ZN(n9303) );
  INV_X1 U6336 ( .A(n4709), .ZN(n9334) );
  INV_X1 U6337 ( .A(n4710), .ZN(n7951) );
  NAND2_X1 U6338 ( .A1(n5142), .A2(n5141), .ZN(n5576) );
  NAND2_X1 U6339 ( .A1(n5078), .A2(n4432), .ZN(n4716) );
  NAND2_X1 U6340 ( .A1(n5450), .A2(n4736), .ZN(n4735) );
  NAND3_X1 U6341 ( .A1(n4737), .A2(n4741), .A3(n5492), .ZN(n4734) );
  INV_X1 U6342 ( .A(n4748), .ZN(n5567) );
  MUX2_X1 U6343 ( .A(n6586), .B(n6588), .S(n5259), .Z(n5051) );
  NAND2_X1 U6344 ( .A1(n5597), .A2(n4769), .ZN(n4765) );
  NAND2_X1 U6345 ( .A1(n4765), .A2(n4766), .ZN(n5166) );
  NAND2_X1 U6346 ( .A1(n5597), .A2(n5596), .ZN(n4768) );
  INV_X1 U6347 ( .A(n5626), .ZN(n4772) );
  NAND2_X1 U6348 ( .A1(n4778), .A2(n5627), .ZN(n9611) );
  NAND2_X1 U6349 ( .A1(n4776), .A2(n4774), .ZN(n8980) );
  NOR2_X1 U6350 ( .A1(n7957), .A2(n4775), .ZN(n4774) );
  INV_X1 U6351 ( .A(n7898), .ZN(n4775) );
  NAND3_X1 U6352 ( .A1(n9052), .A2(n4539), .A3(n4783), .ZN(n4782) );
  OAI21_X1 U6353 ( .B1(n7583), .B2(n4791), .A(n4789), .ZN(n7674) );
  NAND2_X1 U6354 ( .A1(n4787), .A2(n4786), .ZN(n5881) );
  NAND2_X1 U6355 ( .A1(n7583), .A2(n4789), .ZN(n4787) );
  NAND2_X1 U6356 ( .A1(n8386), .A2(n4795), .ZN(n4792) );
  NAND2_X1 U6357 ( .A1(n4792), .A2(n4793), .ZN(n6558) );
  NAND2_X1 U6358 ( .A1(n8386), .A2(n4799), .ZN(n4794) );
  NAND2_X1 U6359 ( .A1(n8386), .A2(n5905), .ZN(n8377) );
  NAND2_X1 U6360 ( .A1(n4800), .A2(n4484), .ZN(n8444) );
  NAND2_X1 U6361 ( .A1(n4801), .A2(n4433), .ZN(n8513) );
  OAI22_X2 U6362 ( .A1(n7414), .A2(n5873), .B1(n8200), .B2(n7404), .ZN(n7433)
         );
  AND2_X1 U6363 ( .A1(n5189), .A2(n4802), .ZN(n5225) );
  NAND2_X1 U6364 ( .A1(n5189), .A2(n4446), .ZN(n8669) );
  AND2_X1 U6365 ( .A1(n5884), .A2(n5882), .ZN(n4804) );
  AND3_X2 U6366 ( .A1(n5313), .A2(n5002), .A3(n5373), .ZN(n5385) );
  NAND2_X1 U6367 ( .A1(n5859), .A2(n7010), .ZN(n5864) );
  NOR2_X4 U6368 ( .A1(n5299), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U6369 ( .A1(n5250), .A2(n5249), .ZN(n4808) );
  INV_X1 U6370 ( .A(n4808), .ZN(n9818) );
  OAI21_X1 U6371 ( .B1(n4808), .B2(n7160), .A(n7161), .ZN(n9829) );
  OAI22_X1 U6372 ( .A1(n8679), .A2(n5039), .B1(P2_U3151), .B2(n4808), .ZN(
        n4807) );
  XNOR2_X1 U6373 ( .A(n7126), .B(n4808), .ZN(n9823) );
  NAND2_X1 U6374 ( .A1(n7142), .A2(n4814), .ZN(n4816) );
  INV_X1 U6375 ( .A(n4816), .ZN(n9815) );
  NAND3_X1 U6376 ( .A1(n4821), .A2(n8254), .A3(n4819), .ZN(n4818) );
  NOR2_X1 U6377 ( .A1(n7244), .A2(n7148), .ZN(n7149) );
  OAI21_X1 U6378 ( .B1(n4829), .B2(n7788), .A(n4828), .ZN(n8233) );
  NAND2_X1 U6379 ( .A1(n8297), .A2(n4838), .ZN(n4836) );
  NOR2_X1 U6380 ( .A1(n8278), .A2(n8505), .ZN(n8296) );
  NAND2_X1 U6381 ( .A1(n4833), .A2(n4836), .ZN(n8326) );
  NOR2_X1 U6382 ( .A1(n8296), .A2(n8297), .ZN(n8299) );
  NAND2_X1 U6383 ( .A1(n7455), .A2(n4843), .ZN(n4842) );
  INV_X1 U6384 ( .A(n4847), .ZN(n7363) );
  NAND2_X1 U6385 ( .A1(n7364), .A2(n7365), .ZN(n4846) );
  XNOR2_X1 U6386 ( .A(n7364), .B(n7365), .ZN(n7271) );
  INV_X1 U6387 ( .A(n7162), .ZN(n4860) );
  AOI21_X1 U6388 ( .B1(n7199), .B2(n7162), .A(n4861), .ZN(n4853) );
  NOR2_X1 U6389 ( .A1(n4855), .A2(n5277), .ZN(n4854) );
  OAI21_X1 U6390 ( .B1(n8280), .B2(n4863), .A(n4862), .ZN(n8344) );
  XNOR2_X1 U6391 ( .A(n8205), .B(n8216), .ZN(n7790) );
  OAI22_X2 U6392 ( .A1(n6862), .A2(n6863), .B1(n6052), .B2(n6051), .ZN(n6894)
         );
  AND2_X2 U6393 ( .A1(n4897), .A2(n4483), .ZN(n6862) );
  OR2_X1 U6394 ( .A1(n6768), .A2(n6767), .ZN(n4897) );
  NAND2_X1 U6395 ( .A1(n4905), .A2(n4906), .ZN(n6267) );
  NAND2_X1 U6396 ( .A1(n8821), .A2(n4908), .ZN(n4905) );
  NAND2_X1 U6397 ( .A1(n6254), .A2(n6253), .ZN(n4917) );
  INV_X1 U6398 ( .A(n6215), .ZN(n4919) );
  INV_X1 U6399 ( .A(n4933), .ZN(n7308) );
  NAND2_X1 U6400 ( .A1(n5972), .A2(n4937), .ZN(n5974) );
  AOI21_X2 U6401 ( .B1(n9414), .B2(n9416), .A(n4942), .ZN(n9401) );
  NAND3_X1 U6402 ( .A1(n4945), .A2(n6998), .A3(n4944), .ZN(n7041) );
  NAND2_X1 U6403 ( .A1(n4947), .A2(n4950), .ZN(n7544) );
  NAND2_X1 U6404 ( .A1(n7598), .A2(n4948), .ZN(n4947) );
  NAND2_X1 U6405 ( .A1(n7523), .A2(n4955), .ZN(n4954) );
  AOI22_X1 U6406 ( .A1(n4956), .A2(n4962), .B1(n4958), .B2(n4960), .ZN(n4953)
         );
  OR2_X1 U6407 ( .A1(n4958), .A2(n4956), .ZN(n4955) );
  NAND2_X1 U6408 ( .A1(n7523), .A2(n9028), .ZN(n7667) );
  OAI21_X1 U6409 ( .B1(n9028), .B2(n4960), .A(n9696), .ZN(n4959) );
  NAND2_X1 U6410 ( .A1(n7667), .A2(n7666), .ZN(n9547) );
  OR2_X1 U6411 ( .A1(n7891), .A2(n4969), .ZN(n4963) );
  NAND3_X1 U6412 ( .A1(n7891), .A2(n4968), .A3(n9043), .ZN(n4967) );
  NAND2_X1 U6413 ( .A1(n9294), .A2(n8952), .ZN(n4975) );
  NAND2_X1 U6414 ( .A1(n4977), .A2(n4976), .ZN(n7885) );
  NAND2_X1 U6415 ( .A1(n7883), .A2(n4978), .ZN(n4977) );
  NAND3_X1 U6416 ( .A1(n5972), .A2(n4983), .A3(n10001), .ZN(n5984) );
  NAND2_X1 U6417 ( .A1(n7569), .A2(n4486), .ZN(n4984) );
  NAND2_X1 U6418 ( .A1(n7400), .A2(n7399), .ZN(n7569) );
  AND2_X2 U6419 ( .A1(n4984), .A2(n4986), .ZN(n7703) );
  INV_X1 U6420 ( .A(n7570), .ZN(n4988) );
  NAND2_X1 U6421 ( .A1(n8157), .A2(n8158), .ZN(n8156) );
  AOI21_X1 U6422 ( .B1(n7865), .B2(n4990), .A(n4498), .ZN(n4989) );
  INV_X1 U6423 ( .A(n8158), .ZN(n4990) );
  NAND2_X1 U6424 ( .A1(n8156), .A2(n7865), .ZN(n7969) );
  INV_X1 U6425 ( .A(n8111), .ZN(n7830) );
  NAND2_X2 U6426 ( .A1(n8075), .A2(n7840), .ZN(n8147) );
  NAND2_X1 U6427 ( .A1(n7838), .A2(n5000), .ZN(n8075) );
  AND2_X2 U6428 ( .A1(n5004), .A2(n5003), .ZN(n5002) );
  NAND2_X1 U6429 ( .A1(n5008), .A2(n5006), .ZN(n6874) );
  INV_X1 U6430 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5009) );
  AND2_X1 U6431 ( .A1(n7072), .A2(n5016), .ZN(n5011) );
  INV_X1 U6432 ( .A(n8009), .ZN(n5012) );
  NAND2_X1 U6433 ( .A1(n5014), .A2(n5011), .ZN(n7338) );
  NOR2_X1 U6434 ( .A1(n8006), .A2(n5015), .ZN(n7073) );
  NAND2_X1 U6435 ( .A1(n7338), .A2(n7337), .ZN(n7339) );
  NAND3_X1 U6436 ( .A1(n8084), .A2(n5017), .A3(n8401), .ZN(n7986) );
  NAND2_X1 U6437 ( .A1(n7853), .A2(n7852), .ZN(n5017) );
  OR2_X2 U6438 ( .A1(n7853), .A2(n7852), .ZN(n8084) );
  AND2_X2 U6439 ( .A1(n5385), .A2(n5019), .ZN(n5648) );
  OR2_X1 U6440 ( .A1(n9488), .A2(n9544), .ZN(n9494) );
  NAND2_X1 U6441 ( .A1(n7885), .A2(n5022), .ZN(n9333) );
  OR2_X1 U6442 ( .A1(n6275), .A2(n6042), .ZN(n6043) );
  INV_X1 U6443 ( .A(n6008), .ZN(n6010) );
  XNOR2_X1 U6444 ( .A(n7905), .B(n9046), .ZN(n9487) );
  XNOR2_X1 U6445 ( .A(n6558), .B(n5625), .ZN(n6562) );
  OR2_X1 U6446 ( .A1(n5848), .A2(n5847), .ZN(n5850) );
  OAI21_X2 U6447 ( .B1(n5844), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U6448 ( .A1(n5652), .A2(n5651), .ZN(n5844) );
  OAI222_X1 U6449 ( .A1(P2_U3151), .A2(n7963), .B1(n7962), .B2(n7961), .C1(
        n7960), .C2(n8679), .ZN(P2_U3265) );
  NAND2_X1 U6450 ( .A1(n7963), .A2(n5230), .ZN(n5278) );
  OR2_X1 U6451 ( .A1(n9588), .A2(n8930), .ZN(n5022) );
  OR2_X1 U6452 ( .A1(n6572), .A2(n9666), .ZN(n5023) );
  OR2_X1 U6453 ( .A1(n6358), .A2(n6357), .ZN(n5024) );
  OR2_X1 U6454 ( .A1(n5646), .A2(n7334), .ZN(n5025) );
  AND2_X1 U6455 ( .A1(n6067), .A2(n6066), .ZN(n5026) );
  AND2_X1 U6456 ( .A1(n6141), .A2(n6140), .ZN(n5027) );
  OR2_X1 U6457 ( .A1(n7881), .A2(n7880), .ZN(n5029) );
  OR2_X1 U6458 ( .A1(n6325), .A2(n6324), .ZN(n5030) );
  INV_X1 U6459 ( .A(n7867), .ZN(n5625) );
  NAND2_X1 U6460 ( .A1(n9857), .A2(n5655), .ZN(n9856) );
  INV_X1 U6461 ( .A(P2_U3893), .ZN(n8187) );
  INV_X1 U6462 ( .A(n9379), .ZN(n7880) );
  AND2_X1 U6463 ( .A1(n9024), .A2(n9023), .ZN(n5032) );
  NAND2_X1 U6464 ( .A1(n7054), .A2(n5870), .ZN(n5033) );
  OR2_X1 U6465 ( .A1(n8201), .A2(n7343), .ZN(n5034) );
  AND2_X1 U6466 ( .A1(n6020), .A2(n5023), .ZN(n5035) );
  AND2_X1 U6467 ( .A1(n6554), .A2(n8524), .ZN(n5036) );
  INV_X1 U6468 ( .A(n7759), .ZN(n5419) );
  AND3_X1 U6469 ( .A1(n5842), .A2(n5949), .A3(n5834), .ZN(n5037) );
  NAND2_X1 U6470 ( .A1(n8549), .A2(n5718), .ZN(n8531) );
  INV_X1 U6471 ( .A(n7813), .ZN(n8631) );
  INV_X1 U6472 ( .A(n9542), .ZN(n7881) );
  NAND2_X1 U6473 ( .A1(n5034), .A2(n5033), .ZN(n5871) );
  AND4_X1 U6474 ( .A1(n5186), .A2(n5185), .A3(n5184), .A4(n5642), .ZN(n5187)
         );
  MUX2_X1 U6475 ( .A(n9008), .B(n8980), .S(n8970), .Z(n8971) );
  INV_X1 U6476 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10217) );
  INV_X1 U6477 ( .A(n8110), .ZN(n7829) );
  OR2_X1 U6478 ( .A1(n8051), .A2(n8188), .ZN(n5905) );
  NAND2_X1 U6479 ( .A1(n5664), .A2(n5665), .ZN(n5865) );
  OR2_X1 U6480 ( .A1(n8834), .A2(n8835), .ZN(n6339) );
  NAND2_X1 U6481 ( .A1(n6754), .A2(n9050), .ZN(n6001) );
  OR2_X1 U6482 ( .A1(n9053), .A2(n8972), .ZN(n8973) );
  INV_X1 U6483 ( .A(n6424), .ZN(n6423) );
  NAND2_X1 U6484 ( .A1(n9253), .A2(n9254), .ZN(n9252) );
  NAND2_X1 U6485 ( .A1(n7881), .A2(n7880), .ZN(n7882) );
  INV_X1 U6486 ( .A(n6149), .ZN(n6147) );
  NAND2_X1 U6487 ( .A1(n9054), .A2(n7279), .ZN(n6500) );
  INV_X1 U6488 ( .A(n5463), .ZN(n5102) );
  INV_X1 U6489 ( .A(n5370), .ZN(n5076) );
  INV_X1 U6490 ( .A(n8389), .ZN(n7863) );
  OR2_X1 U6491 ( .A1(n5613), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U6492 ( .A1(n7202), .A2(n5264), .ZN(n7158) );
  AND2_X1 U6493 ( .A1(n7147), .A2(n7241), .ZN(n7148) );
  NAND2_X1 U6494 ( .A1(n8185), .A2(n8351), .ZN(n5916) );
  NOR2_X1 U6495 ( .A1(n8561), .A2(n8378), .ZN(n5778) );
  INV_X1 U6496 ( .A(n6616), .ZN(n6543) );
  NAND2_X1 U6497 ( .A1(n5333), .A2(n5691), .ZN(n7432) );
  INV_X1 U6498 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6499 ( .A1(n6084), .A2(n6086), .ZN(n6087) );
  OR2_X1 U6500 ( .A1(n6459), .A2(n6458), .ZN(n6514) );
  NAND2_X1 U6501 ( .A1(n6423), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6443) );
  OR2_X1 U6502 ( .A1(n6260), .A2(n8685), .ZN(n6291) );
  NAND2_X1 U6503 ( .A1(n8987), .A2(n9000), .ZN(n9270) );
  NAND2_X1 U6504 ( .A1(n6276), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U6505 ( .A1(n6223), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U6506 ( .A1(n6104), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U6507 ( .A1(n9800), .A2(n9145), .ZN(n9064) );
  OR2_X1 U6508 ( .A1(n5166), .A2(n5165), .ZN(n5167) );
  NOR2_X1 U6509 ( .A1(n5099), .A2(n5098), .ZN(n5101) );
  AND2_X1 U6510 ( .A1(n7862), .A2(n7860), .ZN(n8054) );
  AND2_X1 U6511 ( .A1(n8053), .A2(n7856), .ZN(n8085) );
  INV_X1 U6512 ( .A(n8431), .ZN(n8401) );
  INV_X1 U6513 ( .A(n5615), .ZN(n5951) );
  OAI21_X1 U6514 ( .B1(n4417), .B2(n5264), .A(n7158), .ZN(n7201) );
  INV_X1 U6515 ( .A(n7729), .ZN(n7632) );
  INV_X1 U6516 ( .A(n8371), .ZN(n8367) );
  INV_X1 U6517 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6539) );
  INV_X1 U6518 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6551) );
  AOI21_X1 U6519 ( .B1(n8508), .B2(n5737), .A(n5491), .ZN(n8490) );
  INV_X1 U6520 ( .A(n8192), .ZN(n8529) );
  INV_X1 U6521 ( .A(n6879), .ZN(n9876) );
  NAND2_X1 U6522 ( .A1(n5849), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5846) );
  INV_X1 U6523 ( .A(n9275), .ZN(n8744) );
  INV_X1 U6524 ( .A(n9322), .ZN(n8771) );
  INV_X1 U6525 ( .A(n9437), .ZN(n8861) );
  INV_X1 U6526 ( .A(n6069), .ZN(n6070) );
  INV_X1 U6527 ( .A(n8871), .ZN(n6517) );
  INV_X1 U6528 ( .A(n9510), .ZN(n9294) );
  INV_X1 U6529 ( .A(n9521), .ZN(n9330) );
  AND2_X1 U6530 ( .A1(n8888), .A2(n8887), .ZN(n7226) );
  OR2_X1 U6531 ( .A1(n9013), .A2(n6785), .ZN(n9439) );
  AND2_X1 U6532 ( .A1(n8918), .A2(n9415), .ZN(n9443) );
  INV_X1 U6533 ( .A(n7779), .ZN(n9768) );
  AND2_X1 U6534 ( .A1(n5147), .A2(n5146), .ZN(n5575) );
  AND2_X1 U6535 ( .A1(n5635), .A2(n5240), .ZN(n8353) );
  AND4_X1 U6536 ( .A1(n5555), .A2(n5554), .A3(n5553), .A4(n5552), .ZN(n8451)
         );
  NAND2_X1 U6537 ( .A1(n4426), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5267) );
  OR2_X1 U6538 ( .A1(n5291), .A2(n5263), .ZN(n5268) );
  AND2_X1 U6539 ( .A1(P2_U3893), .A2(n5855), .ZN(n9821) );
  INV_X1 U6540 ( .A(n8552), .ZN(n8539) );
  NAND2_X1 U6541 ( .A1(n6721), .A2(n6532), .ZN(n9860) );
  INV_X1 U6542 ( .A(n7618), .ZN(n7706) );
  AND2_X1 U6543 ( .A1(n9941), .A2(n9927), .ZN(n8607) );
  INV_X1 U6544 ( .A(n9922), .ZN(n9920) );
  INV_X1 U6545 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6546 ( .A1(n6021), .A2(n5035), .ZN(n6723) );
  AND2_X1 U6547 ( .A1(n6509), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8847) );
  AND2_X1 U6548 ( .A1(n9118), .A2(n9117), .ZN(n9119) );
  OR2_X1 U6549 ( .A1(n7937), .A2(n6516), .ZN(n6523) );
  AND4_X1 U6550 ( .A1(n6248), .A2(n6247), .A3(n6246), .A4(n6245), .ZN(n8686)
         );
  INV_X1 U6551 ( .A(n9213), .ZN(n9684) );
  OR2_X1 U6552 ( .A1(n9659), .A2(n6629), .ZN(n9660) );
  INV_X1 U6553 ( .A(n9044), .ZN(n7949) );
  AOI22_X1 U6554 ( .A1(n9401), .A2(n7879), .B1(n9631), .B2(n9392), .ZN(n9386)
         );
  AND2_X1 U6555 ( .A1(n6526), .A2(n6785), .ZN(n9461) );
  INV_X1 U6556 ( .A(n9439), .ZN(n9460) );
  AND2_X1 U6557 ( .A1(n6486), .A2(n9602), .ZN(n6807) );
  AND2_X1 U6558 ( .A1(n7599), .A2(n9546), .ZN(n9544) );
  INV_X1 U6559 ( .A(n9544), .ZN(n9802) );
  AND2_X1 U6560 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n9945), .ZN(n9942) );
  INV_X1 U6561 ( .A(n5261), .ZN(n6577) );
  AND2_X1 U6562 ( .A1(n6817), .A2(n6816), .ZN(n8119) );
  INV_X1 U6563 ( .A(n8179), .ZN(n8150) );
  INV_X1 U6564 ( .A(n8402), .ZN(n8188) );
  AND2_X1 U6565 ( .A1(n7156), .A2(n7155), .ZN(n9855) );
  NAND2_X1 U6566 ( .A1(n9872), .A2(n5950), .ZN(n8552) );
  INV_X2 U6567 ( .A(n9872), .ZN(n9874) );
  NAND2_X2 U6568 ( .A1(n5953), .A2(n9860), .ZN(n9872) );
  INV_X1 U6569 ( .A(n8607), .ZN(n8617) );
  INV_X1 U6570 ( .A(n9941), .ZN(n9939) );
  NAND2_X1 U6571 ( .A1(n6554), .A2(n8661), .ZN(n6555) );
  OR2_X1 U6572 ( .A1(n9929), .A2(n9915), .ZN(n8667) );
  AND2_X1 U6573 ( .A1(n6550), .A2(n6549), .ZN(n9929) );
  INV_X1 U6574 ( .A(n6760), .ZN(n6731) );
  AND2_X1 U6575 ( .A1(n6721), .A2(n5925), .ZN(n6760) );
  INV_X1 U6576 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10163) );
  INV_X1 U6577 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6596) );
  INV_X1 U6578 ( .A(n7910), .ZN(n9631) );
  NAND2_X1 U6579 ( .A1(n6503), .A2(n6498), .ZN(n8866) );
  NAND2_X1 U6580 ( .A1(n6523), .A2(n6522), .ZN(n9240) );
  INV_X1 U6581 ( .A(n8795), .ZN(n9321) );
  INV_X1 U6582 ( .A(n6979), .ZN(n9146) );
  OR2_X1 U6583 ( .A1(n9659), .A2(n6785), .ZN(n9212) );
  OR2_X1 U6584 ( .A1(n4419), .A2(n4539), .ZN(n9740) );
  OR2_X1 U6585 ( .A1(n4419), .A2(n6972), .ZN(n9433) );
  INV_X1 U6586 ( .A(n9814), .ZN(n9811) );
  INV_X1 U6587 ( .A(n9245), .ZN(n9573) );
  INV_X1 U6588 ( .A(n9747), .ZN(n9746) );
  INV_X1 U6589 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10178) );
  INV_X1 U6590 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6599) );
  INV_X1 U6591 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6586) );
  INV_X1 U6592 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10013) );
  OAI21_X1 U6593 ( .B1(n6530), .B2(n9874), .A(n5956), .ZN(P2_U3204) );
  MUX2_X1 U6594 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(P2_DATAO_REG_0__SCAN_IN), 
        .S(n5194), .Z(n5040) );
  NAND2_X1 U6595 ( .A1(n5040), .A2(SI_0_), .ZN(n5246) );
  NAND2_X1 U6596 ( .A1(n5041), .A2(SI_1_), .ZN(n5042) );
  INV_X1 U6597 ( .A(SI_2_), .ZN(n5043) );
  XNOR2_X1 U6598 ( .A(n5044), .B(n5043), .ZN(n5269) );
  NAND2_X1 U6599 ( .A1(n5044), .A2(SI_2_), .ZN(n5045) );
  NAND2_X1 U6600 ( .A1(n5046), .A2(n5045), .ZN(n5287) );
  INV_X1 U6601 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6578) );
  INV_X1 U6602 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6580) );
  MUX2_X1 U6603 ( .A(n6578), .B(n6580), .S(n5194), .Z(n5047) );
  NAND2_X1 U6604 ( .A1(n5287), .A2(n5286), .ZN(n5050) );
  INV_X1 U6605 ( .A(n5047), .ZN(n5048) );
  NAND2_X1 U6606 ( .A1(n5048), .A2(SI_3_), .ZN(n5049) );
  NAND2_X1 U6607 ( .A1(n5050), .A2(n5049), .ZN(n5303) );
  INV_X1 U6608 ( .A(n5051), .ZN(n5052) );
  NAND2_X1 U6609 ( .A1(n5052), .A2(SI_4_), .ZN(n5053) );
  NAND2_X1 U6610 ( .A1(n5054), .A2(n5053), .ZN(n5317) );
  NAND2_X1 U6611 ( .A1(n5317), .A2(n5316), .ZN(n5058) );
  INV_X1 U6612 ( .A(n5055), .ZN(n5056) );
  NAND2_X1 U6613 ( .A1(n5056), .A2(SI_5_), .ZN(n5057) );
  NAND2_X1 U6614 ( .A1(n5058), .A2(n5057), .ZN(n5330) );
  NAND2_X1 U6615 ( .A1(n5330), .A2(n5329), .ZN(n5062) );
  INV_X1 U6616 ( .A(n5059), .ZN(n5060) );
  NAND2_X1 U6617 ( .A1(n5060), .A2(SI_6_), .ZN(n5061) );
  NAND2_X1 U6618 ( .A1(n5062), .A2(n5061), .ZN(n5346) );
  NAND2_X1 U6619 ( .A1(n5346), .A2(n5345), .ZN(n5066) );
  INV_X1 U6620 ( .A(n5063), .ZN(n5064) );
  INV_X1 U6621 ( .A(SI_8_), .ZN(n5067) );
  INV_X1 U6622 ( .A(n5068), .ZN(n5069) );
  NAND2_X1 U6623 ( .A1(n5069), .A2(SI_8_), .ZN(n5070) );
  INV_X1 U6624 ( .A(SI_9_), .ZN(n5072) );
  INV_X1 U6625 ( .A(n5073), .ZN(n5074) );
  NAND2_X1 U6626 ( .A1(n5074), .A2(SI_9_), .ZN(n5075) );
  INV_X1 U6627 ( .A(n5079), .ZN(n5080) );
  INV_X1 U6628 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6612) );
  INV_X1 U6629 ( .A(SI_11_), .ZN(n5083) );
  INV_X1 U6630 ( .A(n5084), .ZN(n5085) );
  NAND2_X1 U6631 ( .A1(n5085), .A2(SI_11_), .ZN(n5086) );
  INV_X1 U6632 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6619) );
  INV_X1 U6633 ( .A(n5088), .ZN(n5089) );
  NAND2_X1 U6634 ( .A1(n5421), .A2(n5090), .ZN(n5093) );
  NAND2_X1 U6635 ( .A1(n5091), .A2(SI_13_), .ZN(n5092) );
  NAND2_X1 U6636 ( .A1(n5436), .A2(n5094), .ZN(n5097) );
  NAND2_X1 U6637 ( .A1(n5095), .A2(SI_14_), .ZN(n5096) );
  INV_X1 U6638 ( .A(SI_15_), .ZN(n5098) );
  NAND2_X1 U6639 ( .A1(n5099), .A2(n5098), .ZN(n5100) );
  INV_X1 U6640 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6765) );
  INV_X1 U6641 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10042) );
  INV_X1 U6642 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6838) );
  INV_X1 U6643 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10187) );
  INV_X1 U6644 ( .A(SI_17_), .ZN(n5104) );
  NAND2_X1 U6645 ( .A1(n5105), .A2(n5104), .ZN(n5108) );
  INV_X1 U6646 ( .A(n5105), .ZN(n5106) );
  NAND2_X1 U6647 ( .A1(n5106), .A2(SI_17_), .ZN(n5107) );
  NAND2_X1 U6648 ( .A1(n5108), .A2(n5107), .ZN(n5476) );
  INV_X1 U6649 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6901) );
  INV_X1 U6650 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5109) );
  XNOR2_X1 U6651 ( .A(n5110), .B(SI_18_), .ZN(n5492) );
  INV_X1 U6652 ( .A(n5110), .ZN(n5111) );
  NAND2_X1 U6653 ( .A1(n5111), .A2(SI_18_), .ZN(n5112) );
  INV_X1 U6654 ( .A(n5508), .ZN(n5118) );
  INV_X1 U6655 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7034) );
  INV_X1 U6656 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7037) );
  INV_X1 U6657 ( .A(SI_19_), .ZN(n5113) );
  NAND2_X1 U6658 ( .A1(n5114), .A2(n5113), .ZN(n5119) );
  INV_X1 U6659 ( .A(n5114), .ZN(n5115) );
  NAND2_X1 U6660 ( .A1(n5115), .A2(SI_19_), .ZN(n5116) );
  NAND2_X1 U6661 ( .A1(n5119), .A2(n5116), .ZN(n5507) );
  INV_X1 U6662 ( .A(n5507), .ZN(n5117) );
  NAND2_X1 U6663 ( .A1(n5118), .A2(n5117), .ZN(n5120) );
  INV_X1 U6664 ( .A(SI_20_), .ZN(n5520) );
  INV_X1 U6665 ( .A(n5521), .ZN(n5121) );
  OAI21_X1 U6666 ( .B1(n5523), .B2(n5520), .A(n5121), .ZN(n5123) );
  NAND2_X1 U6667 ( .A1(n5123), .A2(n5122), .ZN(n5535) );
  INV_X1 U6668 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n9971) );
  INV_X1 U6669 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10232) );
  INV_X1 U6670 ( .A(n5533), .ZN(n5124) );
  NOR2_X1 U6671 ( .A1(n5124), .A2(SI_21_), .ZN(n5126) );
  NAND2_X1 U6672 ( .A1(n5124), .A2(SI_21_), .ZN(n5125) );
  INV_X1 U6673 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7485) );
  INV_X1 U6674 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7487) );
  INV_X1 U6675 ( .A(SI_22_), .ZN(n5127) );
  NAND2_X1 U6676 ( .A1(n5128), .A2(n5127), .ZN(n5131) );
  INV_X1 U6677 ( .A(n5128), .ZN(n5129) );
  NAND2_X1 U6678 ( .A1(n5129), .A2(SI_22_), .ZN(n5130) );
  NAND2_X1 U6679 ( .A1(n5131), .A2(n5130), .ZN(n5544) );
  INV_X1 U6680 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9986) );
  INV_X1 U6681 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7593) );
  INV_X1 U6682 ( .A(SI_23_), .ZN(n5132) );
  NAND2_X1 U6683 ( .A1(n5133), .A2(n5132), .ZN(n5136) );
  INV_X1 U6684 ( .A(n5133), .ZN(n5134) );
  NAND2_X1 U6685 ( .A1(n5134), .A2(SI_23_), .ZN(n5135) );
  INV_X1 U6686 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7769) );
  INV_X1 U6687 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7683) );
  INV_X1 U6688 ( .A(SI_24_), .ZN(n5137) );
  NAND2_X1 U6689 ( .A1(n5138), .A2(n5137), .ZN(n5141) );
  INV_X1 U6690 ( .A(n5138), .ZN(n5139) );
  NAND2_X1 U6691 ( .A1(n5139), .A2(SI_24_), .ZN(n5140) );
  NAND2_X1 U6692 ( .A1(n5567), .A2(n5566), .ZN(n5142) );
  INV_X1 U6693 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7766) );
  INV_X1 U6694 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10015) );
  INV_X1 U6695 ( .A(SI_25_), .ZN(n5143) );
  NAND2_X1 U6696 ( .A1(n5144), .A2(n5143), .ZN(n5147) );
  INV_X1 U6697 ( .A(n5144), .ZN(n5145) );
  NAND2_X1 U6698 ( .A1(n5145), .A2(SI_25_), .ZN(n5146) );
  INV_X1 U6699 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7783) );
  INV_X1 U6700 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10008) );
  INV_X1 U6701 ( .A(SI_26_), .ZN(n5148) );
  NAND2_X1 U6702 ( .A1(n5149), .A2(n5148), .ZN(n5152) );
  INV_X1 U6703 ( .A(n5149), .ZN(n5150) );
  NAND2_X1 U6704 ( .A1(n5150), .A2(SI_26_), .ZN(n5151) );
  AND2_X1 U6705 ( .A1(n5152), .A2(n5151), .ZN(n5586) );
  INV_X1 U6706 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7966) );
  INV_X1 U6707 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9615) );
  INV_X1 U6708 ( .A(SI_27_), .ZN(n5154) );
  NAND2_X1 U6709 ( .A1(n5155), .A2(n5154), .ZN(n5158) );
  INV_X1 U6710 ( .A(n5155), .ZN(n5156) );
  NAND2_X1 U6711 ( .A1(n5156), .A2(SI_27_), .ZN(n5157) );
  AND2_X1 U6712 ( .A1(n5158), .A2(n5157), .ZN(n5596) );
  INV_X1 U6713 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8678) );
  INV_X1 U6714 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7894) );
  INV_X1 U6715 ( .A(SI_28_), .ZN(n5159) );
  NAND2_X1 U6716 ( .A1(n5160), .A2(n5159), .ZN(n5163) );
  INV_X1 U6717 ( .A(n5160), .ZN(n5161) );
  NAND2_X1 U6718 ( .A1(n5161), .A2(SI_28_), .ZN(n5162) );
  AND2_X1 U6719 ( .A1(n5163), .A2(n5162), .ZN(n5609) );
  INV_X1 U6720 ( .A(n5164), .ZN(n5165) );
  INV_X1 U6721 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7960) );
  INV_X1 U6722 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8879) );
  INV_X1 U6723 ( .A(SI_30_), .ZN(n5168) );
  NAND2_X1 U6724 ( .A1(n5169), .A2(n5168), .ZN(n5172) );
  INV_X1 U6725 ( .A(n5169), .ZN(n5170) );
  NAND2_X1 U6726 ( .A1(n5170), .A2(SI_30_), .ZN(n5171) );
  NAND2_X1 U6727 ( .A1(n5172), .A2(n5171), .ZN(n5197) );
  INV_X1 U6728 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8671) );
  INV_X1 U6729 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9604) );
  XNOR2_X1 U6730 ( .A(n5173), .B(SI_31_), .ZN(n5174) );
  NOR2_X1 U6731 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5494) );
  NOR2_X1 U6732 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5182) );
  NOR2_X1 U6733 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5181) );
  INV_X1 U6734 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5180) );
  NAND4_X1 U6735 ( .A1(n5494), .A2(n5182), .A3(n5181), .A4(n5180), .ZN(n5183)
         );
  NOR2_X1 U6736 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5186) );
  NOR2_X1 U6737 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n5185) );
  NOR2_X1 U6738 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5184) );
  INV_X1 U6739 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5642) );
  INV_X1 U6740 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5188) );
  INV_X1 U6741 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5190) );
  INV_X1 U6742 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U6743 ( .A1(n9609), .A2(n5610), .ZN(n5196) );
  OR2_X1 U6744 ( .A1(n4431), .A2(n8671), .ZN(n5195) );
  NAND2_X1 U6745 ( .A1(n8878), .A2(n5610), .ZN(n5200) );
  OR2_X1 U6746 ( .A1(n5285), .A2(n7960), .ZN(n5199) );
  INV_X1 U6747 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5205) );
  INV_X1 U6748 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7721) );
  INV_X1 U6749 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5208) );
  INV_X1 U6750 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5210) );
  INV_X1 U6751 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5212) );
  INV_X1 U6752 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10033) );
  INV_X1 U6753 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5215) );
  INV_X1 U6754 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10012) );
  INV_X1 U6755 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5218) );
  INV_X1 U6756 ( .A(n5600), .ZN(n5221) );
  INV_X1 U6757 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U6758 ( .A1(n5221), .A2(n5220), .ZN(n5613) );
  INV_X1 U6759 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5226) );
  INV_X1 U6760 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8670) );
  OR2_X2 U6761 ( .A1(n5225), .A2(n5190), .ZN(n5227) );
  XNOR2_X2 U6762 ( .A(n5227), .B(n5226), .ZN(n5229) );
  NAND2_X1 U6763 ( .A1(n5951), .A2(n4511), .ZN(n5635) );
  INV_X1 U6764 ( .A(n7963), .ZN(n5228) );
  INV_X1 U6765 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n10060) );
  INV_X1 U6766 ( .A(n5620), .ZN(n5630) );
  NAND2_X1 U6767 ( .A1(n5630), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5232) );
  NAND2_X1 U6768 ( .A1(n5617), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5231) );
  OAI211_X1 U6769 ( .C1(n5291), .C2(n10060), .A(n5232), .B(n5231), .ZN(n5233)
         );
  INV_X1 U6770 ( .A(n5233), .ZN(n5234) );
  NAND2_X1 U6771 ( .A1(n5635), .A2(n5234), .ZN(n8185) );
  INV_X1 U6772 ( .A(n8185), .ZN(n5636) );
  INV_X1 U6773 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6774 ( .A1(n5617), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5237) );
  INV_X1 U6775 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n5235) );
  OR2_X1 U6776 ( .A1(n5291), .A2(n5235), .ZN(n5236) );
  OAI211_X1 U6777 ( .C1(n5238), .C2(n5620), .A(n5237), .B(n5236), .ZN(n5239)
         );
  INV_X1 U6778 ( .A(n5239), .ZN(n5240) );
  INV_X1 U6779 ( .A(n8353), .ZN(n8184) );
  NAND2_X1 U6780 ( .A1(n5787), .A2(n8184), .ZN(n5639) );
  INV_X1 U6781 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7015) );
  NAND2_X1 U6782 ( .A1(n5253), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5241) );
  INV_X1 U6783 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7125) );
  OR2_X1 U6784 ( .A1(n5278), .A2(n7125), .ZN(n5244) );
  XNOR2_X1 U6785 ( .A(n5247), .B(n5246), .ZN(n6581) );
  NAND2_X1 U6786 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5248) );
  MUX2_X1 U6787 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5248), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5250) );
  INV_X1 U6788 ( .A(n5859), .ZN(n5806) );
  INV_X1 U6789 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7330) );
  OR2_X1 U6790 ( .A1(n5252), .A2(n7330), .ZN(n5255) );
  NAND2_X1 U6791 ( .A1(n4426), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5254) );
  INV_X1 U6792 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7159) );
  OR2_X1 U6793 ( .A1(n5278), .A2(n7159), .ZN(n5257) );
  INV_X1 U6794 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7141) );
  NAND2_X1 U6795 ( .A1(n5259), .A2(SI_0_), .ZN(n5260) );
  XNOR2_X1 U6796 ( .A(n5260), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8680) );
  MUX2_X1 U6797 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8680), .S(n4415), .Z(n6840) );
  INV_X1 U6798 ( .A(n5656), .ZN(n6878) );
  NAND2_X1 U6799 ( .A1(n5806), .A2(n6878), .ZN(n7009) );
  NAND2_X1 U6800 ( .A1(n7009), .A2(n5657), .ZN(n9857) );
  INV_X1 U6801 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5263) );
  INV_X1 U6802 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9859) );
  OR2_X1 U6803 ( .A1(n5486), .A2(n9859), .ZN(n5266) );
  INV_X1 U6804 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5264) );
  OR2_X1 U6805 ( .A1(n5278), .A2(n5264), .ZN(n5265) );
  OR2_X1 U6806 ( .A1(n4431), .A2(n4507), .ZN(n5275) );
  XNOR2_X1 U6807 ( .A(n5270), .B(n5269), .ZN(n6584) );
  OR2_X1 U6808 ( .A1(n5288), .A2(n6584), .ZN(n5274) );
  OR2_X1 U6809 ( .A1(n5261), .A2(n4417), .ZN(n5273) );
  NAND2_X1 U6810 ( .A1(n8204), .A2(n9882), .ZN(n5665) );
  INV_X1 U6811 ( .A(n5865), .ZN(n5655) );
  NAND2_X1 U6812 ( .A1(n9856), .A2(n5664), .ZN(n7298) );
  NAND2_X1 U6813 ( .A1(n4426), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5282) );
  INV_X1 U6814 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5276) );
  OR2_X1 U6815 ( .A1(n5291), .A2(n5276), .ZN(n5281) );
  OR2_X1 U6816 ( .A1(n5486), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5280) );
  INV_X1 U6817 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5277) );
  OR2_X1 U6818 ( .A1(n5278), .A2(n5277), .ZN(n5279) );
  NAND4_X1 U6819 ( .A1(n5282), .A2(n5281), .A3(n5280), .A4(n5279), .ZN(n8203)
         );
  NAND2_X1 U6820 ( .A1(n5283), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5284) );
  XNOR2_X1 U6821 ( .A(n5284), .B(n5176), .ZN(n7287) );
  XNOR2_X1 U6822 ( .A(n5287), .B(n5286), .ZN(n6579) );
  OR2_X1 U6823 ( .A1(n5288), .A2(n6579), .ZN(n5289) );
  OAI211_X1 U6824 ( .C1(n5261), .C2(n7287), .A(n5290), .B(n5289), .ZN(n8011)
         );
  OR2_X1 U6825 ( .A1(n8203), .A2(n9888), .ZN(n7024) );
  NAND2_X1 U6826 ( .A1(n8203), .A2(n9888), .ZN(n5674) );
  AND2_X1 U6827 ( .A1(n7024), .A2(n5674), .ZN(n7299) );
  NAND2_X1 U6828 ( .A1(n7298), .A2(n7299), .ZN(n7022) );
  NAND2_X1 U6829 ( .A1(n7022), .A2(n7024), .ZN(n5306) );
  NAND2_X1 U6830 ( .A1(n5616), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5298) );
  INV_X1 U6831 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5292) );
  OR2_X1 U6832 ( .A1(n5602), .A2(n5292), .ZN(n5297) );
  NAND2_X1 U6833 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5293) );
  AND2_X1 U6834 ( .A1(n5307), .A2(n5293), .ZN(n7079) );
  OR2_X1 U6835 ( .A1(n5486), .A2(n7079), .ZN(n5296) );
  INV_X1 U6836 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5294) );
  OR2_X1 U6837 ( .A1(n5620), .A2(n5294), .ZN(n5295) );
  NAND2_X1 U6838 ( .A1(n5299), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5301) );
  INV_X1 U6839 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5300) );
  OR2_X1 U6840 ( .A1(n4431), .A2(n6588), .ZN(n5305) );
  XNOR2_X1 U6841 ( .A(n5303), .B(n5302), .ZN(n6587) );
  OR2_X1 U6842 ( .A1(n5288), .A2(n6587), .ZN(n5304) );
  OAI211_X1 U6843 ( .C1(n5261), .C2(n7189), .A(n5305), .B(n5304), .ZN(n7070)
         );
  OR2_X1 U6844 ( .A1(n8202), .A2(n7070), .ZN(n7052) );
  NAND2_X1 U6845 ( .A1(n8202), .A2(n7070), .ZN(n7054) );
  NAND2_X1 U6846 ( .A1(n5306), .A2(n7023), .ZN(n7027) );
  INV_X1 U6847 ( .A(n7070), .ZN(n9892) );
  OR2_X1 U6848 ( .A1(n8202), .A2(n9892), .ZN(n5675) );
  NAND2_X1 U6849 ( .A1(n7027), .A2(n5675), .ZN(n7060) );
  NAND2_X1 U6850 ( .A1(n4426), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5312) );
  INV_X1 U6851 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7137) );
  OR2_X1 U6852 ( .A1(n5291), .A2(n7137), .ZN(n5311) );
  NAND2_X1 U6853 ( .A1(n5307), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5308) );
  AND2_X1 U6854 ( .A1(n5321), .A2(n5308), .ZN(n7349) );
  OR2_X1 U6855 ( .A1(n5486), .A2(n7349), .ZN(n5310) );
  INV_X1 U6856 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7136) );
  OR2_X1 U6857 ( .A1(n5620), .A2(n7136), .ZN(n5309) );
  OR2_X1 U6858 ( .A1(n5313), .A2(n5190), .ZN(n5315) );
  XNOR2_X1 U6859 ( .A(n5315), .B(n5314), .ZN(n7165) );
  XNOR2_X1 U6860 ( .A(n5317), .B(n5316), .ZN(n6590) );
  OR2_X1 U6861 ( .A1(n5288), .A2(n6590), .ZN(n5319) );
  OR2_X1 U6862 ( .A1(n4431), .A2(n6589), .ZN(n5318) );
  OAI211_X1 U6863 ( .C1(n5261), .C2(n7165), .A(n5319), .B(n5318), .ZN(n7343)
         );
  NAND2_X1 U6864 ( .A1(n8201), .A2(n7335), .ZN(n5805) );
  NAND2_X1 U6865 ( .A1(n7060), .A2(n5805), .ZN(n7410) );
  OR2_X1 U6866 ( .A1(n8201), .A2(n7335), .ZN(n7411) );
  NAND2_X1 U6867 ( .A1(n5616), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5326) );
  INV_X1 U6868 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5320) );
  OR2_X1 U6869 ( .A1(n5602), .A2(n5320), .ZN(n5325) );
  NAND2_X1 U6870 ( .A1(n5321), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5322) );
  AND2_X1 U6871 ( .A1(n5335), .A2(n5322), .ZN(n7413) );
  OR2_X1 U6872 ( .A1(n5486), .A2(n7413), .ZN(n5324) );
  INV_X1 U6873 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7248) );
  OR2_X1 U6874 ( .A1(n5620), .A2(n7248), .ZN(n5323) );
  NAND4_X1 U6875 ( .A1(n5326), .A2(n5325), .A3(n5324), .A4(n5323), .ZN(n8200)
         );
  NAND2_X1 U6876 ( .A1(n5327), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5328) );
  XNOR2_X1 U6877 ( .A(n5328), .B(n5005), .ZN(n7268) );
  XNOR2_X1 U6878 ( .A(n5330), .B(n5329), .ZN(n6592) );
  OR2_X1 U6879 ( .A1(n5288), .A2(n6592), .ZN(n5332) );
  OR2_X1 U6880 ( .A1(n4431), .A2(n6593), .ZN(n5331) );
  OAI211_X1 U6881 ( .C1(n4415), .C2(n7268), .A(n5332), .B(n5331), .ZN(n7404)
         );
  INV_X1 U6882 ( .A(n7404), .ZN(n9896) );
  OR2_X1 U6883 ( .A1(n8200), .A2(n9896), .ZN(n5678) );
  AND2_X1 U6884 ( .A1(n7411), .A2(n5678), .ZN(n5689) );
  NAND2_X1 U6885 ( .A1(n7410), .A2(n5689), .ZN(n5333) );
  NAND2_X1 U6886 ( .A1(n8200), .A2(n9896), .ZN(n5691) );
  NAND2_X1 U6887 ( .A1(n5617), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5341) );
  INV_X1 U6888 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5334) );
  OR2_X1 U6889 ( .A1(n5291), .A2(n5334), .ZN(n5340) );
  NAND2_X1 U6890 ( .A1(n5335), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5336) );
  AND2_X1 U6891 ( .A1(n5350), .A2(n5336), .ZN(n7573) );
  OR2_X1 U6892 ( .A1(n5486), .A2(n7573), .ZN(n5339) );
  INV_X1 U6893 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5337) );
  OR2_X1 U6894 ( .A1(n5620), .A2(n5337), .ZN(n5338) );
  NAND2_X1 U6895 ( .A1(n4473), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5342) );
  MUX2_X1 U6896 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5342), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5344) );
  NAND2_X1 U6897 ( .A1(n5344), .A2(n5343), .ZN(n7365) );
  XNOR2_X1 U6898 ( .A(n5346), .B(n5345), .ZN(n6595) );
  OR2_X1 U6899 ( .A1(n5288), .A2(n6595), .ZN(n5348) );
  OR2_X1 U6900 ( .A1(n4431), .A2(n10203), .ZN(n5347) );
  OAI211_X1 U6901 ( .C1(n4415), .C2(n7365), .A(n5348), .B(n5347), .ZN(n7576)
         );
  INV_X1 U6902 ( .A(n7576), .ZN(n9900) );
  OR2_X1 U6903 ( .A1(n8199), .A2(n9900), .ZN(n5693) );
  NAND2_X1 U6904 ( .A1(n8199), .A2(n9900), .ZN(n7464) );
  NAND2_X1 U6905 ( .A1(n7432), .A2(n7434), .ZN(n7431) );
  NAND2_X1 U6906 ( .A1(n5616), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5355) );
  INV_X1 U6907 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5349) );
  OR2_X1 U6908 ( .A1(n5602), .A2(n5349), .ZN(n5354) );
  NAND2_X1 U6909 ( .A1(n5350), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5351) );
  AND2_X1 U6910 ( .A1(n5363), .A2(n5351), .ZN(n7698) );
  OR2_X1 U6911 ( .A1(n5486), .A2(n7698), .ZN(n5353) );
  INV_X1 U6912 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7368) );
  OR2_X1 U6913 ( .A1(n5620), .A2(n7368), .ZN(n5352) );
  NAND2_X1 U6914 ( .A1(n5343), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5356) );
  XNOR2_X1 U6915 ( .A(n5356), .B(n5003), .ZN(n9854) );
  INV_X1 U6916 ( .A(n5357), .ZN(n5358) );
  XNOR2_X1 U6917 ( .A(n5359), .B(n5358), .ZN(n6597) );
  OR2_X1 U6918 ( .A1(n5288), .A2(n6597), .ZN(n5361) );
  OR2_X1 U6919 ( .A1(n4431), .A2(n6596), .ZN(n5360) );
  OAI211_X1 U6920 ( .C1(n5261), .C2(n9854), .A(n5361), .B(n5360), .ZN(n7692)
         );
  NAND2_X1 U6921 ( .A1(n8198), .A2(n9905), .ZN(n5810) );
  AND2_X1 U6922 ( .A1(n5810), .A2(n7464), .ZN(n5682) );
  NAND2_X1 U6923 ( .A1(n7431), .A2(n5682), .ZN(n5362) );
  NAND2_X1 U6924 ( .A1(n5362), .A2(n5811), .ZN(n7585) );
  NAND2_X1 U6925 ( .A1(n5617), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5369) );
  OR2_X1 U6926 ( .A1(n5291), .A2(n7362), .ZN(n5368) );
  NAND2_X1 U6927 ( .A1(n5363), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5364) );
  AND2_X1 U6928 ( .A1(n5379), .A2(n5364), .ZN(n7587) );
  OR2_X1 U6929 ( .A1(n5252), .A2(n7587), .ZN(n5367) );
  INV_X1 U6930 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5365) );
  OR2_X1 U6931 ( .A1(n5620), .A2(n5365), .ZN(n5366) );
  XNOR2_X1 U6932 ( .A(n5371), .B(n5370), .ZN(n6600) );
  OR2_X1 U6933 ( .A1(n5288), .A2(n6600), .ZN(n5377) );
  OR2_X1 U6934 ( .A1(n4431), .A2(n6601), .ZN(n5376) );
  OR2_X1 U6935 ( .A1(n5372), .A2(n5190), .ZN(n5374) );
  XNOR2_X1 U6936 ( .A(n5374), .B(n5373), .ZN(n7441) );
  OR2_X1 U6937 ( .A1(n4415), .A2(n7441), .ZN(n5375) );
  NAND2_X1 U6938 ( .A1(n8197), .A2(n7618), .ZN(n5684) );
  NAND2_X1 U6939 ( .A1(n5616), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5384) );
  INV_X1 U6940 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5378) );
  OR2_X1 U6941 ( .A1(n5602), .A2(n5378), .ZN(n5383) );
  NAND2_X1 U6942 ( .A1(n5379), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5380) );
  AND2_X1 U6943 ( .A1(n5395), .A2(n5380), .ZN(n7998) );
  OR2_X1 U6944 ( .A1(n5252), .A2(n7998), .ZN(n5382) );
  INV_X1 U6945 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7451) );
  OR2_X1 U6946 ( .A1(n5620), .A2(n7451), .ZN(n5381) );
  NOR2_X1 U6947 ( .A1(n5385), .A2(n5190), .ZN(n5386) );
  MUX2_X1 U6948 ( .A(n5190), .B(n5386), .S(P2_IR_REG_10__SCAN_IN), .Z(n5387)
         );
  INV_X1 U6949 ( .A(n5387), .ZN(n5390) );
  INV_X1 U6950 ( .A(n5388), .ZN(n5389) );
  NAND2_X1 U6951 ( .A1(n5390), .A2(n5389), .ZN(n7638) );
  XNOR2_X1 U6952 ( .A(n5392), .B(n5391), .ZN(n6602) );
  OR2_X1 U6953 ( .A1(n4431), .A2(n6603), .ZN(n5393) );
  NAND2_X1 U6954 ( .A1(n8196), .A2(n9910), .ZN(n5685) );
  NAND2_X1 U6955 ( .A1(n5698), .A2(n5685), .ZN(n7651) );
  NAND2_X1 U6956 ( .A1(n5617), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5401) );
  INV_X1 U6957 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5394) );
  OR2_X1 U6958 ( .A1(n5291), .A2(n5394), .ZN(n5400) );
  NAND2_X1 U6959 ( .A1(n5395), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5396) );
  AND2_X1 U6960 ( .A1(n5413), .A2(n5396), .ZN(n8140) );
  OR2_X1 U6961 ( .A1(n5486), .A2(n8140), .ZN(n5399) );
  INV_X1 U6962 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5397) );
  OR2_X1 U6963 ( .A1(n5620), .A2(n5397), .ZN(n5398) );
  NAND2_X1 U6964 ( .A1(n6611), .A2(n5610), .ZN(n5406) );
  OR2_X1 U6965 ( .A1(n5388), .A2(n5190), .ZN(n5404) );
  XNOR2_X1 U6966 ( .A(n5404), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7729) );
  AOI22_X1 U6967 ( .A1(n5511), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6577), .B2(
        n7729), .ZN(n5405) );
  NAND2_X1 U6968 ( .A1(n5406), .A2(n5405), .ZN(n8139) );
  NAND2_X1 U6969 ( .A1(n8038), .A2(n8139), .ZN(n5704) );
  INV_X1 U6970 ( .A(n8139), .ZN(n9916) );
  NAND2_X1 U6971 ( .A1(n9916), .A2(n8195), .ZN(n5705) );
  NAND2_X1 U6972 ( .A1(n6618), .A2(n5610), .ZN(n5412) );
  NAND2_X1 U6973 ( .A1(n5409), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5410) );
  XNOR2_X1 U6974 ( .A(n5410), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7732) );
  AOI22_X1 U6975 ( .A1(n5511), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6577), .B2(
        n7732), .ZN(n5411) );
  NAND2_X1 U6976 ( .A1(n5617), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5418) );
  INV_X1 U6977 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7761) );
  OR2_X1 U6978 ( .A1(n5291), .A2(n7761), .ZN(n5417) );
  NAND2_X1 U6979 ( .A1(n5413), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5414) );
  AND2_X1 U6980 ( .A1(n5425), .A2(n5414), .ZN(n8042) );
  OR2_X1 U6981 ( .A1(n5252), .A2(n8042), .ZN(n5416) );
  INV_X1 U6982 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7714) );
  OR2_X1 U6983 ( .A1(n5620), .A2(n7714), .ZN(n5415) );
  NAND4_X1 U6984 ( .A1(n5418), .A2(n5417), .A3(n5416), .A4(n5415), .ZN(n8194)
         );
  NAND2_X1 U6985 ( .A1(n9926), .A2(n8137), .ZN(n5711) );
  NAND2_X1 U6986 ( .A1(n5710), .A2(n5711), .ZN(n7759) );
  XNOR2_X1 U6987 ( .A(n5421), .B(n5420), .ZN(n6621) );
  NAND2_X1 U6988 ( .A1(n6621), .A2(n5610), .ZN(n5424) );
  OR2_X1 U6989 ( .A1(n5409), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U6990 ( .A1(n5437), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5422) );
  XNOR2_X1 U6991 ( .A(n5422), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8216) );
  AOI22_X1 U6992 ( .A1(n5511), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6577), .B2(
        n8216), .ZN(n5423) );
  NAND2_X1 U6993 ( .A1(n7805), .A2(n9623), .ZN(n5431) );
  NAND2_X1 U6994 ( .A1(n5617), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5430) );
  INV_X1 U6995 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7794) );
  OR2_X1 U6996 ( .A1(n5291), .A2(n7794), .ZN(n5429) );
  NAND2_X1 U6997 ( .A1(n5425), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5426) );
  AND2_X1 U6998 ( .A1(n5442), .A2(n5426), .ZN(n8115) );
  OR2_X1 U6999 ( .A1(n5252), .A2(n8115), .ZN(n5428) );
  INV_X1 U7000 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7793) );
  OR2_X1 U7001 ( .A1(n5620), .A2(n7793), .ZN(n5427) );
  NAND4_X1 U7002 ( .A1(n5430), .A2(n5429), .A3(n5428), .A4(n5427), .ZN(n8193)
         );
  NAND2_X1 U7003 ( .A1(n5431), .A2(n8544), .ZN(n5434) );
  INV_X1 U7004 ( .A(n7805), .ZN(n5432) );
  NAND2_X1 U7005 ( .A1(n5432), .A2(n8117), .ZN(n5433) );
  XNOR2_X1 U7006 ( .A(n5436), .B(n5435), .ZN(n6727) );
  NAND2_X1 U7007 ( .A1(n6727), .A2(n5610), .ZN(n5440) );
  NOR2_X1 U7008 ( .A1(n5437), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5452) );
  OR2_X1 U7009 ( .A1(n5452), .A2(n5190), .ZN(n5438) );
  XNOR2_X1 U7010 ( .A(n5438), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8231) );
  AOI22_X1 U7011 ( .A1(n5511), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6577), .B2(
        n8231), .ZN(n5439) );
  NAND2_X1 U7012 ( .A1(n5616), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5447) );
  INV_X1 U7013 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n5441) );
  OR2_X1 U7014 ( .A1(n5602), .A2(n5441), .ZN(n5446) );
  NAND2_X1 U7015 ( .A1(n5442), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5443) );
  AND2_X1 U7016 ( .A1(n5456), .A2(n5443), .ZN(n8546) );
  OR2_X1 U7017 ( .A1(n5252), .A2(n8546), .ZN(n5445) );
  INV_X1 U7018 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8208) );
  OR2_X1 U7019 ( .A1(n5620), .A2(n8208), .ZN(n5444) );
  NAND4_X1 U7020 ( .A1(n5447), .A2(n5446), .A3(n5445), .A4(n5444), .ZN(n8192)
         );
  NAND2_X1 U7021 ( .A1(n9622), .A2(n8529), .ZN(n5719) );
  XNOR2_X1 U7022 ( .A(n5448), .B(SI_15_), .ZN(n5449) );
  XNOR2_X1 U7023 ( .A(n5450), .B(n5449), .ZN(n6747) );
  NAND2_X1 U7024 ( .A1(n6747), .A2(n5610), .ZN(n5455) );
  INV_X1 U7025 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5451) );
  AND2_X1 U7026 ( .A1(n5452), .A2(n5451), .ZN(n5467) );
  OR2_X1 U7027 ( .A1(n5467), .A2(n5190), .ZN(n5453) );
  XNOR2_X1 U7028 ( .A(n5453), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8246) );
  AOI22_X1 U7029 ( .A1(n5511), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6577), .B2(
        n8246), .ZN(n5454) );
  NAND2_X1 U7030 ( .A1(n5617), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5461) );
  INV_X1 U7031 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8536) );
  OR2_X1 U7032 ( .A1(n5291), .A2(n8536), .ZN(n5460) );
  NAND2_X1 U7033 ( .A1(n5456), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5457) );
  AND2_X1 U7034 ( .A1(n5470), .A2(n5457), .ZN(n8535) );
  OR2_X1 U7035 ( .A1(n5252), .A2(n8535), .ZN(n5459) );
  INV_X1 U7036 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8615) );
  OR2_X1 U7037 ( .A1(n5620), .A2(n8615), .ZN(n5458) );
  NAND2_X1 U7038 ( .A1(n8533), .A2(n8545), .ZN(n5732) );
  NAND2_X1 U7039 ( .A1(n8531), .A2(n5732), .ZN(n5462) );
  XNOR2_X1 U7040 ( .A(n5463), .B(SI_16_), .ZN(n5464) );
  XNOR2_X1 U7041 ( .A(n5465), .B(n5464), .ZN(n6763) );
  NAND2_X1 U7042 ( .A1(n6763), .A2(n5610), .ZN(n5469) );
  INV_X1 U7043 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U7044 ( .A1(n5467), .A2(n5466), .ZN(n5496) );
  NAND2_X1 U7045 ( .A1(n5496), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5479) );
  XNOR2_X1 U7046 ( .A(n5479), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8266) );
  AOI22_X1 U7047 ( .A1(n5511), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6577), .B2(
        n8266), .ZN(n5468) );
  INV_X1 U7048 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8518) );
  OR2_X1 U7049 ( .A1(n5291), .A2(n8518), .ZN(n5475) );
  INV_X1 U7050 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n10025) );
  OR2_X1 U7051 ( .A1(n5602), .A2(n10025), .ZN(n5474) );
  NAND2_X1 U7052 ( .A1(n5470), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5471) );
  AND2_X1 U7053 ( .A1(n5484), .A2(n5471), .ZN(n8517) );
  OR2_X1 U7054 ( .A1(n5252), .A2(n8517), .ZN(n5473) );
  INV_X1 U7055 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8261) );
  OR2_X1 U7056 ( .A1(n5620), .A2(n8261), .ZN(n5472) );
  NAND2_X1 U7057 ( .A1(n8609), .A2(n8530), .ZN(n5733) );
  XNOR2_X1 U7058 ( .A(n5477), .B(n5476), .ZN(n6837) );
  NAND2_X1 U7059 ( .A1(n6837), .A2(n5610), .ZN(n5483) );
  INV_X1 U7060 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U7061 ( .A1(n5479), .A2(n5478), .ZN(n5480) );
  NAND2_X1 U7062 ( .A1(n5480), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5481) );
  XNOR2_X1 U7063 ( .A(n5481), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8307) );
  AOI22_X1 U7064 ( .A1(n5511), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8307), .B2(
        n6577), .ZN(n5482) );
  NAND2_X1 U7065 ( .A1(n5617), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5490) );
  INV_X1 U7066 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8505) );
  OR2_X1 U7067 ( .A1(n5291), .A2(n8505), .ZN(n5489) );
  NAND2_X1 U7068 ( .A1(n5484), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5485) );
  AND2_X1 U7069 ( .A1(n5501), .A2(n5485), .ZN(n8504) );
  OR2_X1 U7070 ( .A1(n5252), .A2(n8504), .ZN(n5488) );
  INV_X1 U7071 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8283) );
  OR2_X1 U7072 ( .A1(n5620), .A2(n8283), .ZN(n5487) );
  NAND2_X1 U7073 ( .A1(n8660), .A2(n8514), .ZN(n5724) );
  INV_X1 U7074 ( .A(n5724), .ZN(n5491) );
  XNOR2_X1 U7075 ( .A(n5493), .B(n5492), .ZN(n6869) );
  NAND2_X1 U7076 ( .A1(n6869), .A2(n5610), .ZN(n5500) );
  INV_X1 U7077 ( .A(n5494), .ZN(n5495) );
  OAI21_X1 U7078 ( .B1(n5496), .B2(n5495), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5497) );
  MUX2_X1 U7079 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5497), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n5498) );
  AND2_X1 U7080 ( .A1(n5498), .A2(n4451), .ZN(n8328) );
  AOI22_X1 U7081 ( .A1(n5511), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6577), .B2(
        n8328), .ZN(n5499) );
  NAND2_X1 U7082 ( .A1(n5616), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5506) );
  INV_X1 U7083 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n10171) );
  OR2_X1 U7084 ( .A1(n5602), .A2(n10171), .ZN(n5505) );
  NAND2_X1 U7085 ( .A1(n5501), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5502) );
  AND2_X1 U7086 ( .A1(n5514), .A2(n5502), .ZN(n8486) );
  OR2_X1 U7087 ( .A1(n5252), .A2(n8486), .ZN(n5504) );
  INV_X1 U7088 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n10233) );
  OR2_X1 U7089 ( .A1(n5620), .A2(n10233), .ZN(n5503) );
  NAND4_X1 U7090 ( .A1(n5506), .A2(n5505), .A3(n5504), .A4(n5503), .ZN(n8498)
         );
  NAND2_X1 U7091 ( .A1(n8599), .A2(n8078), .ZN(n5725) );
  NAND2_X1 U7092 ( .A1(n8490), .A2(n8489), .ZN(n8488) );
  NAND2_X1 U7093 ( .A1(n8488), .A2(n5738), .ZN(n8479) );
  XNOR2_X1 U7094 ( .A(n5508), .B(n5507), .ZN(n7033) );
  NAND2_X1 U7095 ( .A1(n7033), .A2(n5610), .ZN(n5513) );
  NAND2_X1 U7096 ( .A1(n4451), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5510) );
  INV_X1 U7097 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5509) );
  AOI22_X1 U7098 ( .A1(n5511), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8338), .B2(
        n6577), .ZN(n5512) );
  NAND2_X1 U7099 ( .A1(n5617), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5519) );
  INV_X1 U7100 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8332) );
  OR2_X1 U7101 ( .A1(n5620), .A2(n8332), .ZN(n5518) );
  NAND2_X1 U7102 ( .A1(n5514), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5515) );
  AND2_X1 U7103 ( .A1(n5526), .A2(n5515), .ZN(n8474) );
  OR2_X1 U7104 ( .A1(n5252), .A2(n8474), .ZN(n5517) );
  INV_X1 U7105 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8475) );
  OR2_X1 U7106 ( .A1(n4416), .A2(n8475), .ZN(n5516) );
  NAND2_X1 U7107 ( .A1(n8477), .A2(n8463), .ZN(n5731) );
  NAND2_X1 U7108 ( .A1(n5743), .A2(n5731), .ZN(n5896) );
  XNOR2_X1 U7109 ( .A(n5521), .B(n5520), .ZN(n5522) );
  XNOR2_X1 U7110 ( .A(n5523), .B(n5522), .ZN(n7196) );
  NAND2_X1 U7111 ( .A1(n7196), .A2(n5610), .ZN(n5525) );
  INV_X1 U7112 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7198) );
  OR2_X1 U7113 ( .A1(n4431), .A2(n7198), .ZN(n5524) );
  NAND2_X1 U7114 ( .A1(n5616), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5531) );
  INV_X1 U7115 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8653) );
  OR2_X1 U7116 ( .A1(n5602), .A2(n8653), .ZN(n5530) );
  NAND2_X1 U7117 ( .A1(n5526), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5527) );
  AND2_X1 U7118 ( .A1(n5538), .A2(n5527), .ZN(n8101) );
  OR2_X1 U7119 ( .A1(n5252), .A2(n8101), .ZN(n5529) );
  INV_X1 U7120 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8592) );
  OR2_X1 U7121 ( .A1(n5620), .A2(n8592), .ZN(n5528) );
  INV_X1 U7122 ( .A(n5804), .ZN(n5532) );
  NAND2_X1 U7123 ( .A1(n8094), .A2(n8450), .ZN(n5803) );
  XNOR2_X1 U7124 ( .A(n5533), .B(SI_21_), .ZN(n5534) );
  XNOR2_X1 U7125 ( .A(n5535), .B(n5534), .ZN(n7333) );
  NAND2_X1 U7126 ( .A1(n7333), .A2(n5610), .ZN(n5537) );
  OR2_X1 U7127 ( .A1(n4431), .A2(n9971), .ZN(n5536) );
  NAND2_X1 U7128 ( .A1(n5616), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5543) );
  INV_X1 U7129 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8649) );
  OR2_X1 U7130 ( .A1(n5602), .A2(n8649), .ZN(n5542) );
  NAND2_X1 U7131 ( .A1(n5538), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5539) );
  AND2_X1 U7132 ( .A1(n5548), .A2(n5539), .ZN(n8029) );
  OR2_X1 U7133 ( .A1(n5252), .A2(n8029), .ZN(n5541) );
  INV_X1 U7134 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8588) );
  OR2_X1 U7135 ( .A1(n5620), .A2(n8588), .ZN(n5540) );
  NAND2_X1 U7136 ( .A1(n8024), .A2(n8464), .ZN(n5801) );
  INV_X1 U7137 ( .A(n5801), .ZN(n5756) );
  XNOR2_X1 U7138 ( .A(n5545), .B(n5544), .ZN(n7483) );
  NAND2_X1 U7139 ( .A1(n7483), .A2(n5610), .ZN(n5547) );
  OR2_X1 U7140 ( .A1(n4431), .A2(n7485), .ZN(n5546) );
  NAND2_X1 U7141 ( .A1(n5548), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U7142 ( .A1(n5560), .A2(n5549), .ZN(n8435) );
  NAND2_X1 U7143 ( .A1(n4511), .A2(n8435), .ZN(n5555) );
  INV_X1 U7144 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8437) );
  OR2_X1 U7145 ( .A1(n5291), .A2(n8437), .ZN(n5554) );
  INV_X1 U7146 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n5550) );
  OR2_X1 U7147 ( .A1(n5602), .A2(n5550), .ZN(n5553) );
  INV_X1 U7148 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n5551) );
  OR2_X1 U7149 ( .A1(n5620), .A2(n5551), .ZN(n5552) );
  NAND2_X1 U7150 ( .A1(n8646), .A2(n8451), .ZN(n5753) );
  INV_X1 U7151 ( .A(n5751), .ZN(n5757) );
  AOI21_X1 U7152 ( .B1(n8440), .B2(n5753), .A(n5757), .ZN(n8419) );
  NAND2_X1 U7153 ( .A1(n7594), .A2(n5610), .ZN(n5559) );
  OR2_X1 U7154 ( .A1(n4431), .A2(n9986), .ZN(n5558) );
  NAND2_X1 U7155 ( .A1(n5560), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7156 ( .A1(n5570), .A2(n5561), .ZN(n8421) );
  NAND2_X1 U7157 ( .A1(n8421), .A2(n4511), .ZN(n5565) );
  NAND2_X1 U7158 ( .A1(n5617), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7159 ( .A1(n5630), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U7160 ( .A1(n5616), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5562) );
  NAND4_X1 U7161 ( .A1(n5565), .A2(n5564), .A3(n5563), .A4(n5562), .ZN(n8431)
         );
  XNOR2_X1 U7162 ( .A(n5567), .B(n5566), .ZN(n7682) );
  NAND2_X1 U7163 ( .A1(n7682), .A2(n5610), .ZN(n5569) );
  OR2_X1 U7164 ( .A1(n4431), .A2(n7769), .ZN(n5568) );
  NAND2_X1 U7165 ( .A1(n5570), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U7166 ( .A1(n5579), .A2(n5571), .ZN(n8407) );
  NAND2_X1 U7167 ( .A1(n8407), .A2(n4511), .ZN(n5574) );
  AOI22_X1 U7168 ( .A1(n5630), .A2(P2_REG1_REG_24__SCAN_IN), .B1(n5617), .B2(
        P2_REG0_REG_24__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7169 ( .A1(n5616), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7170 ( .A1(n8638), .A2(n8417), .ZN(n5824) );
  NAND2_X1 U7171 ( .A1(n8420), .A2(n8401), .ZN(n8408) );
  NAND2_X1 U7172 ( .A1(n5824), .A2(n8408), .ZN(n5766) );
  NAND2_X1 U7173 ( .A1(n7765), .A2(n5610), .ZN(n5578) );
  OR2_X1 U7174 ( .A1(n4431), .A2(n7766), .ZN(n5577) );
  NAND2_X1 U7175 ( .A1(n5579), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7176 ( .A1(n5589), .A2(n5580), .ZN(n8393) );
  NAND2_X1 U7177 ( .A1(n8393), .A2(n4511), .ZN(n5583) );
  AOI22_X1 U7178 ( .A1(n5630), .A2(P2_REG1_REG_25__SCAN_IN), .B1(n5617), .B2(
        P2_REG0_REG_25__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7179 ( .A1(n5616), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5581) );
  INV_X1 U7180 ( .A(n5771), .ZN(n5584) );
  NAND2_X1 U7181 ( .A1(n7782), .A2(n5610), .ZN(n5588) );
  OR2_X1 U7182 ( .A1(n4431), .A2(n7783), .ZN(n5587) );
  NAND2_X1 U7183 ( .A1(n5589), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U7184 ( .A1(n5600), .A2(n5590), .ZN(n8381) );
  NAND2_X1 U7185 ( .A1(n8381), .A2(n4511), .ZN(n5595) );
  INV_X1 U7186 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n10188) );
  NAND2_X1 U7187 ( .A1(n5616), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7188 ( .A1(n5617), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5591) );
  OAI211_X1 U7189 ( .C1(n10188), .C2(n5620), .A(n5592), .B(n5591), .ZN(n5593)
         );
  INV_X1 U7190 ( .A(n5593), .ZN(n5594) );
  NAND2_X1 U7191 ( .A1(n7965), .A2(n5610), .ZN(n5599) );
  OR2_X1 U7192 ( .A1(n4431), .A2(n7966), .ZN(n5598) );
  NAND2_X1 U7193 ( .A1(n5600), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U7194 ( .A1(n5613), .A2(n5601), .ZN(n8373) );
  NAND2_X1 U7195 ( .A1(n8373), .A2(n4511), .ZN(n5607) );
  INV_X1 U7196 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10041) );
  NAND2_X1 U7197 ( .A1(n5616), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5604) );
  INV_X1 U7198 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n10068) );
  OR2_X1 U7199 ( .A1(n5602), .A2(n10068), .ZN(n5603) );
  OAI211_X1 U7200 ( .C1(n5620), .C2(n10041), .A(n5604), .B(n5603), .ZN(n5605)
         );
  INV_X1 U7201 ( .A(n5605), .ZN(n5606) );
  NAND2_X1 U7202 ( .A1(n8561), .A2(n8378), .ZN(n5775) );
  NAND2_X1 U7203 ( .A1(n8675), .A2(n5610), .ZN(n5612) );
  OR2_X1 U7204 ( .A1(n4431), .A2(n8678), .ZN(n5611) );
  NAND2_X1 U7205 ( .A1(n5613), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U7206 ( .A1(n5615), .A2(n5614), .ZN(n8360) );
  NAND2_X1 U7207 ( .A1(n8360), .A2(n4511), .ZN(n5623) );
  INV_X1 U7208 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U7209 ( .A1(n5616), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U7210 ( .A1(n5617), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5618) );
  OAI211_X1 U7211 ( .C1(n6563), .C2(n5620), .A(n5619), .B(n5618), .ZN(n5621)
         );
  INV_X1 U7212 ( .A(n5621), .ZN(n5622) );
  INV_X1 U7213 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7967) );
  OR2_X1 U7214 ( .A1(n4431), .A2(n7967), .ZN(n5628) );
  INV_X1 U7215 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n10201) );
  NAND2_X1 U7216 ( .A1(n5617), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U7217 ( .A1(n5630), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5631) );
  OAI211_X1 U7218 ( .C1(n10201), .C2(n4416), .A(n5632), .B(n5631), .ZN(n5633)
         );
  INV_X1 U7219 ( .A(n5633), .ZN(n5634) );
  INV_X1 U7220 ( .A(n8622), .ZN(n8358) );
  NOR2_X1 U7221 ( .A1(n8555), .A2(n8358), .ZN(n5637) );
  NAND2_X1 U7222 ( .A1(n8622), .A2(n5636), .ZN(n5789) );
  NAND2_X1 U7223 ( .A1(n6554), .A2(n7871), .ZN(n5783) );
  AND2_X1 U7224 ( .A1(n5789), .A2(n5783), .ZN(n5793) );
  NAND2_X1 U7225 ( .A1(n5798), .A2(n5793), .ZN(n5833) );
  AOI211_X1 U7226 ( .C1(n5945), .C2(n5784), .A(n5637), .B(n5833), .ZN(n5638)
         );
  AOI21_X1 U7227 ( .B1(n8555), .B2(n5639), .A(n5638), .ZN(n5842) );
  INV_X1 U7228 ( .A(n5648), .ZN(n5640) );
  INV_X1 U7229 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7230 ( .A1(n5645), .A2(n5644), .ZN(n5641) );
  NAND2_X1 U7231 ( .A1(n5641), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5643) );
  INV_X1 U7232 ( .A(n7334), .ZN(n5949) );
  NOR2_X1 U7233 ( .A1(n7197), .A2(n8333), .ZN(n5834) );
  NOR2_X1 U7234 ( .A1(n7197), .A2(n8338), .ZN(n5836) );
  INV_X1 U7235 ( .A(n5836), .ZN(n5646) );
  INV_X1 U7236 ( .A(n5725), .ZN(n5730) );
  NOR2_X1 U7237 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5647) );
  AND2_X2 U7238 ( .A1(n5648), .A2(n5647), .ZN(n5652) );
  INV_X1 U7239 ( .A(n5652), .ZN(n5649) );
  NAND2_X1 U7240 ( .A1(n5649), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5650) );
  MUX2_X1 U7241 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5650), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n5653) );
  INV_X1 U7242 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U7243 ( .A1(n5653), .A2(n5844), .ZN(n7484) );
  MUX2_X1 U7244 ( .A(n5657), .B(n5654), .S(n5941), .Z(n5663) );
  INV_X1 U7245 ( .A(n6840), .ZN(n6917) );
  NAND2_X1 U7246 ( .A1(n7012), .A2(n6917), .ZN(n5807) );
  INV_X1 U7247 ( .A(n7484), .ZN(n5910) );
  NAND2_X1 U7248 ( .A1(n5807), .A2(n5910), .ZN(n5660) );
  NAND2_X1 U7249 ( .A1(n5807), .A2(n5949), .ZN(n5658) );
  NAND3_X1 U7250 ( .A1(n5658), .A2(n5941), .A3(n5657), .ZN(n5659) );
  OAI21_X1 U7251 ( .B1(n5859), .B2(n5660), .A(n5659), .ZN(n5661) );
  OAI21_X1 U7252 ( .B1(n5949), .B2(n5656), .A(n5661), .ZN(n5662) );
  NAND3_X1 U7253 ( .A1(n5663), .A2(n5655), .A3(n5662), .ZN(n5671) );
  NAND2_X1 U7254 ( .A1(n7024), .A2(n5664), .ZN(n5668) );
  NAND2_X1 U7255 ( .A1(n5674), .A2(n5665), .ZN(n5667) );
  MUX2_X1 U7256 ( .A(n5668), .B(n5667), .S(n5666), .Z(n5669) );
  INV_X1 U7257 ( .A(n5669), .ZN(n5670) );
  NAND2_X1 U7258 ( .A1(n5671), .A2(n5670), .ZN(n5673) );
  NAND2_X1 U7259 ( .A1(n8202), .A2(n9892), .ZN(n5686) );
  MUX2_X1 U7260 ( .A(n5686), .B(n5675), .S(n6575), .Z(n5672) );
  NAND2_X1 U7261 ( .A1(n5673), .A2(n5672), .ZN(n5688) );
  INV_X1 U7262 ( .A(n5674), .ZN(n5676) );
  OAI211_X1 U7263 ( .C1(n5688), .C2(n5676), .A(n7411), .B(n5675), .ZN(n5677)
         );
  NAND3_X1 U7264 ( .A1(n5677), .A2(n5691), .A3(n5805), .ZN(n5679) );
  NAND3_X1 U7265 ( .A1(n5679), .A2(n7434), .A3(n5678), .ZN(n5683) );
  NAND2_X1 U7266 ( .A1(n5811), .A2(n5697), .ZN(n5681) );
  NAND2_X1 U7267 ( .A1(n5684), .A2(n5810), .ZN(n5680) );
  MUX2_X1 U7268 ( .A(n5681), .B(n5680), .S(n6575), .Z(n5695) );
  INV_X1 U7269 ( .A(n7024), .ZN(n5687) );
  OAI211_X1 U7270 ( .C1(n5688), .C2(n5687), .A(n5805), .B(n5686), .ZN(n5690)
         );
  NAND2_X1 U7271 ( .A1(n5690), .A2(n5689), .ZN(n5692) );
  NAND3_X1 U7272 ( .A1(n5692), .A2(n7434), .A3(n5691), .ZN(n5694) );
  NAND3_X1 U7273 ( .A1(n5694), .A2(n5811), .A3(n5693), .ZN(n5696) );
  NAND2_X1 U7274 ( .A1(n5696), .A2(n4612), .ZN(n5700) );
  AND4_X1 U7275 ( .A1(n5704), .A2(n5698), .A3(n5697), .A4(n6575), .ZN(n5699)
         );
  OAI21_X1 U7276 ( .B1(n8038), .B2(n5941), .A(n9916), .ZN(n5703) );
  NAND2_X1 U7277 ( .A1(n8038), .A2(n5941), .ZN(n5701) );
  NAND2_X1 U7278 ( .A1(n5701), .A2(n8139), .ZN(n5702) );
  NAND2_X1 U7279 ( .A1(n5703), .A2(n5702), .ZN(n5708) );
  NAND4_X1 U7280 ( .A1(n5704), .A2(n6575), .A3(n9910), .A4(n8196), .ZN(n5707)
         );
  NAND4_X1 U7281 ( .A1(n5705), .A2(n8036), .A3(n5941), .A4(n7997), .ZN(n5706)
         );
  AND3_X1 U7282 ( .A1(n5708), .A2(n5707), .A3(n5706), .ZN(n5709) );
  MUX2_X1 U7283 ( .A(n5711), .B(n5710), .S(n6575), .Z(n5712) );
  INV_X1 U7284 ( .A(n5714), .ZN(n5716) );
  NAND2_X1 U7285 ( .A1(n8117), .A2(n8193), .ZN(n5885) );
  NOR2_X1 U7286 ( .A1(n8117), .A2(n8193), .ZN(n5883) );
  MUX2_X1 U7287 ( .A(n8544), .B(n9623), .S(n6575), .Z(n5713) );
  OAI21_X1 U7288 ( .B1(n5714), .B2(n5884), .A(n5713), .ZN(n5715) );
  OAI21_X1 U7289 ( .B1(n5716), .B2(n5885), .A(n5715), .ZN(n5717) );
  MUX2_X1 U7290 ( .A(n5719), .B(n5718), .S(n6575), .Z(n5720) );
  NAND2_X1 U7291 ( .A1(n5721), .A2(n5732), .ZN(n8532) );
  INV_X1 U7292 ( .A(n8532), .ZN(n8526) );
  NAND3_X1 U7293 ( .A1(n5722), .A2(n5666), .A3(n5733), .ZN(n5723) );
  NAND2_X1 U7294 ( .A1(n5737), .A2(n5724), .ZN(n8497) );
  INV_X1 U7295 ( .A(n8497), .ZN(n8507) );
  NAND2_X1 U7296 ( .A1(n5723), .A2(n8507), .ZN(n5728) );
  AND2_X1 U7297 ( .A1(n5725), .A2(n5724), .ZN(n5818) );
  INV_X1 U7298 ( .A(n5818), .ZN(n5726) );
  INV_X2 U7299 ( .A(n5941), .ZN(n6575) );
  NAND2_X1 U7300 ( .A1(n5726), .A2(n6575), .ZN(n5727) );
  NAND2_X1 U7301 ( .A1(n5728), .A2(n5727), .ZN(n5741) );
  NAND3_X1 U7302 ( .A1(n5741), .A2(n5743), .A3(n5738), .ZN(n5729) );
  INV_X1 U7303 ( .A(n5731), .ZN(n5744) );
  NAND3_X1 U7304 ( .A1(n5734), .A2(n5733), .A3(n5732), .ZN(n5736) );
  NAND3_X1 U7305 ( .A1(n5736), .A2(n5941), .A3(n5735), .ZN(n5740) );
  AND2_X1 U7306 ( .A1(n5738), .A2(n5737), .ZN(n5819) );
  INV_X1 U7307 ( .A(n5819), .ZN(n5739) );
  AOI21_X1 U7308 ( .B1(n5741), .B2(n5740), .A(n5739), .ZN(n5742) );
  NAND2_X1 U7309 ( .A1(n5804), .A2(n5743), .ZN(n5745) );
  MUX2_X1 U7310 ( .A(n5745), .B(n5744), .S(n6575), .Z(n5746) );
  INV_X1 U7311 ( .A(n5746), .ZN(n5747) );
  AND2_X1 U7312 ( .A1(n5801), .A2(n5803), .ZN(n5749) );
  AND2_X1 U7313 ( .A1(n5802), .A2(n5804), .ZN(n5748) );
  MUX2_X1 U7314 ( .A(n5749), .B(n5748), .S(n6575), .Z(n5750) );
  NAND2_X1 U7315 ( .A1(n5751), .A2(n5753), .ZN(n8439) );
  INV_X1 U7316 ( .A(n5802), .ZN(n5752) );
  NOR2_X1 U7317 ( .A1(n8439), .A2(n5752), .ZN(n5755) );
  NAND2_X1 U7318 ( .A1(n8408), .A2(n5753), .ZN(n5754) );
  AOI21_X1 U7319 ( .B1(n5759), .B2(n5755), .A(n5754), .ZN(n5761) );
  NOR2_X1 U7320 ( .A1(n8439), .A2(n5756), .ZN(n5758) );
  AOI21_X1 U7321 ( .B1(n5759), .B2(n5758), .A(n5757), .ZN(n5760) );
  INV_X1 U7322 ( .A(n5765), .ZN(n5764) );
  AND2_X1 U7323 ( .A1(n5825), .A2(n5800), .ZN(n5763) );
  INV_X1 U7324 ( .A(n5824), .ZN(n5762) );
  AOI21_X1 U7325 ( .B1(n5764), .B2(n5763), .A(n5762), .ZN(n5770) );
  NAND2_X1 U7326 ( .A1(n5765), .A2(n5800), .ZN(n5768) );
  INV_X1 U7327 ( .A(n5766), .ZN(n5767) );
  AOI21_X1 U7328 ( .B1(n5768), .B2(n5767), .A(n4671), .ZN(n5769) );
  MUX2_X1 U7329 ( .A(n5770), .B(n5769), .S(n5666), .Z(n5774) );
  MUX2_X1 U7330 ( .A(n5772), .B(n5771), .S(n6575), .Z(n5773) );
  OAI211_X1 U7331 ( .C1(n5774), .C2(n8394), .A(n8379), .B(n5773), .ZN(n5782)
         );
  INV_X1 U7332 ( .A(n5775), .ZN(n5779) );
  MUX2_X1 U7333 ( .A(n5776), .B(n4472), .S(n5941), .Z(n5777) );
  NOR2_X1 U7334 ( .A1(n8371), .A2(n5777), .ZN(n5781) );
  MUX2_X1 U7335 ( .A(n5779), .B(n5778), .S(n6575), .Z(n5780) );
  MUX2_X1 U7336 ( .A(n7973), .B(n8362), .S(n5941), .Z(n5785) );
  AOI21_X1 U7337 ( .B1(n5786), .B2(n5785), .A(n5944), .ZN(n5790) );
  NAND2_X1 U7338 ( .A1(n5787), .A2(n5784), .ZN(n5831) );
  AOI211_X1 U7339 ( .C1(n5790), .C2(n8362), .A(n5831), .B(n5791), .ZN(n5797)
         );
  INV_X1 U7340 ( .A(n5787), .ZN(n5788) );
  AOI21_X1 U7341 ( .B1(n6575), .B2(n5789), .A(n5788), .ZN(n5796) );
  NAND2_X1 U7342 ( .A1(n5790), .A2(n7973), .ZN(n5794) );
  INV_X1 U7343 ( .A(n5791), .ZN(n5792) );
  NAND4_X1 U7344 ( .A1(n5794), .A2(n5793), .A3(n5941), .A4(n5792), .ZN(n5795)
         );
  OAI21_X1 U7345 ( .B1(n5797), .B2(n5796), .A(n5795), .ZN(n5799) );
  AND2_X1 U7346 ( .A1(n8555), .A2(n8353), .ZN(n5832) );
  AND2_X1 U7347 ( .A1(n5800), .A2(n8408), .ZN(n8418) );
  INV_X1 U7348 ( .A(n8439), .ZN(n8429) );
  NAND2_X1 U7349 ( .A1(n5802), .A2(n5801), .ZN(n8445) );
  AND2_X1 U7350 ( .A1(n7411), .A2(n5805), .ZN(n7059) );
  NAND4_X1 U7351 ( .A1(n5806), .A2(n5655), .A3(n7059), .A4(n7023), .ZN(n5809)
         );
  AND2_X1 U7352 ( .A1(n5656), .A2(n5807), .ZN(n6842) );
  NAND2_X1 U7353 ( .A1(n7299), .A2(n6842), .ZN(n5808) );
  NOR2_X1 U7354 ( .A1(n5809), .A2(n5808), .ZN(n5812) );
  AND2_X1 U7355 ( .A1(n5811), .A2(n5810), .ZN(n7466) );
  XNOR2_X1 U7356 ( .A(n8200), .B(n7404), .ZN(n7415) );
  NAND4_X1 U7357 ( .A1(n5812), .A2(n7466), .A3(n7434), .A4(n7415), .ZN(n5813)
         );
  NOR4_X1 U7358 ( .A1(n5813), .A2(n7820), .A3(n7651), .A4(n7586), .ZN(n5815)
         );
  INV_X1 U7359 ( .A(n5885), .ZN(n5814) );
  OR2_X1 U7360 ( .A1(n5883), .A2(n5814), .ZN(n7806) );
  NAND4_X1 U7361 ( .A1(n5815), .A2(n5419), .A3(n8551), .A4(n7806), .ZN(n5816)
         );
  NOR2_X1 U7362 ( .A1(n5816), .A2(n8532), .ZN(n5817) );
  NAND4_X1 U7363 ( .A1(n5819), .A2(n5818), .A3(n8511), .A4(n5817), .ZN(n5820)
         );
  NOR2_X1 U7364 ( .A1(n5896), .A2(n5820), .ZN(n5821) );
  NAND2_X1 U7365 ( .A1(n8461), .A2(n5821), .ZN(n5822) );
  NOR2_X1 U7366 ( .A1(n8445), .A2(n5822), .ZN(n5823) );
  NAND3_X1 U7367 ( .A1(n8418), .A2(n8429), .A3(n5823), .ZN(n5826) );
  NAND2_X1 U7368 ( .A1(n5825), .A2(n5824), .ZN(n8399) );
  OR3_X1 U7369 ( .A1(n8394), .A2(n5826), .A3(n8399), .ZN(n5827) );
  NOR2_X1 U7370 ( .A1(n5828), .A2(n5827), .ZN(n5829) );
  NAND3_X1 U7371 ( .A1(n8367), .A2(n7867), .A3(n5829), .ZN(n5830) );
  INV_X1 U7372 ( .A(n5837), .ZN(n5835) );
  NAND3_X1 U7373 ( .A1(n5835), .A2(n5834), .A3(n7334), .ZN(n5841) );
  NAND3_X1 U7374 ( .A1(n5837), .A2(n5836), .A3(n7334), .ZN(n5840) );
  NAND2_X1 U7375 ( .A1(n5844), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5838) );
  INV_X1 U7376 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n10028) );
  XNOR2_X1 U7377 ( .A(n5838), .B(n10028), .ZN(n6574) );
  OR2_X1 U7378 ( .A1(n6574), .A2(P2_U3151), .ZN(n7595) );
  INV_X1 U7379 ( .A(n7595), .ZN(n5839) );
  INV_X1 U7380 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U7381 ( .A1(n5848), .A2(n5847), .ZN(n5849) );
  INV_X1 U7382 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5845) );
  INV_X1 U7383 ( .A(n5921), .ZN(n5854) );
  NAND2_X1 U7384 ( .A1(n5850), .A2(n5849), .ZN(n5920) );
  NAND2_X1 U7385 ( .A1(n5851), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5852) );
  XNOR2_X1 U7386 ( .A(n5852), .B(P2_IR_REG_26__SCAN_IN), .ZN(n5923) );
  NOR2_X1 U7387 ( .A1(n5920), .A2(n7784), .ZN(n5853) );
  NAND2_X1 U7388 ( .A1(n5854), .A2(n5853), .ZN(n6824) );
  NAND2_X1 U7389 ( .A1(n7197), .A2(n8333), .ZN(n5939) );
  INV_X1 U7390 ( .A(n5939), .ZN(n5948) );
  NAND2_X1 U7391 ( .A1(n6575), .A2(n5948), .ZN(n5946) );
  NAND2_X1 U7392 ( .A1(n6721), .A2(n6841), .ZN(n6829) );
  NOR3_X1 U7393 ( .A1(n6829), .A2(n7135), .A3(n5855), .ZN(n5857) );
  OAI21_X1 U7394 ( .B1(n7595), .B2(n5910), .A(P2_B_REG_SCAN_IN), .ZN(n5856) );
  OR2_X1 U7395 ( .A1(n5857), .A2(n5856), .ZN(n5858) );
  OAI21_X1 U7396 ( .B1(n5037), .B2(n5843), .A(n5858), .ZN(P2_U3296) );
  NAND2_X1 U7397 ( .A1(n7012), .A2(n6840), .ZN(n7010) );
  NAND3_X1 U7398 ( .A1(n5862), .A2(n5861), .A3(n4454), .ZN(n6879) );
  OR2_X1 U7399 ( .A1(n5860), .A2(n6879), .ZN(n5863) );
  NAND2_X1 U7400 ( .A1(n5864), .A2(n5863), .ZN(n9861) );
  NAND2_X1 U7401 ( .A1(n9861), .A2(n5865), .ZN(n5867) );
  INV_X1 U7402 ( .A(n9882), .ZN(n6908) );
  OR2_X1 U7403 ( .A1(n8204), .A2(n6908), .ZN(n5866) );
  NOR2_X1 U7404 ( .A1(n8203), .A2(n8011), .ZN(n5868) );
  INV_X1 U7405 ( .A(n8203), .ZN(n9864) );
  AND2_X1 U7406 ( .A1(n7052), .A2(n5034), .ZN(n5869) );
  NAND2_X1 U7407 ( .A1(n7053), .A2(n5869), .ZN(n5872) );
  NAND2_X1 U7408 ( .A1(n8201), .A2(n7343), .ZN(n5870) );
  AND2_X1 U7409 ( .A1(n8200), .A2(n7404), .ZN(n5873) );
  NOR2_X1 U7410 ( .A1(n8199), .A2(n7576), .ZN(n5874) );
  NAND2_X1 U7411 ( .A1(n8199), .A2(n7576), .ZN(n5875) );
  AND2_X1 U7412 ( .A1(n8198), .A2(n7692), .ZN(n5877) );
  OR2_X1 U7413 ( .A1(n8198), .A2(n7692), .ZN(n5876) );
  OR2_X1 U7414 ( .A1(n8197), .A2(n7706), .ZN(n5878) );
  NAND2_X1 U7415 ( .A1(n8196), .A2(n7997), .ZN(n5879) );
  NAND2_X1 U7416 ( .A1(n8139), .A2(n8195), .ZN(n5880) );
  NAND2_X1 U7417 ( .A1(n5881), .A2(n5880), .ZN(n7758) );
  OR2_X1 U7418 ( .A1(n9926), .A2(n8194), .ZN(n5882) );
  INV_X1 U7419 ( .A(n5883), .ZN(n5884) );
  AND2_X1 U7420 ( .A1(n9622), .A2(n8192), .ZN(n5888) );
  OAI21_X2 U7421 ( .B1(n8542), .B2(n5888), .A(n5887), .ZN(n8527) );
  INV_X1 U7422 ( .A(n8545), .ZN(n8191) );
  OR2_X1 U7423 ( .A1(n8533), .A2(n8191), .ZN(n5889) );
  INV_X1 U7424 ( .A(n8530), .ZN(n8501) );
  NAND2_X1 U7425 ( .A1(n8609), .A2(n8501), .ZN(n5891) );
  NAND2_X1 U7426 ( .A1(n8513), .A2(n5891), .ZN(n8496) );
  NAND2_X1 U7427 ( .A1(n8496), .A2(n8497), .ZN(n8495) );
  INV_X1 U7428 ( .A(n8514), .ZN(n8483) );
  NAND2_X1 U7429 ( .A1(n8660), .A2(n8483), .ZN(n5892) );
  NAND2_X1 U7430 ( .A1(n8495), .A2(n5892), .ZN(n8482) );
  OR2_X1 U7431 ( .A1(n8599), .A2(n8498), .ZN(n5893) );
  NAND2_X1 U7432 ( .A1(n8482), .A2(n5893), .ZN(n5895) );
  NAND2_X1 U7433 ( .A1(n8599), .A2(n8498), .ZN(n5894) );
  NAND2_X1 U7434 ( .A1(n5895), .A2(n5894), .ZN(n8471) );
  NAND2_X1 U7435 ( .A1(n8477), .A2(n8484), .ZN(n5897) );
  INV_X1 U7436 ( .A(n8450), .ZN(n8472) );
  OR2_X1 U7437 ( .A1(n8094), .A2(n8472), .ZN(n8446) );
  NAND2_X1 U7438 ( .A1(n8444), .A2(n8446), .ZN(n5899) );
  NAND2_X1 U7439 ( .A1(n5899), .A2(n8445), .ZN(n8427) );
  INV_X1 U7440 ( .A(n8464), .ZN(n8190) );
  NAND2_X1 U7441 ( .A1(n8427), .A2(n8428), .ZN(n5900) );
  INV_X1 U7442 ( .A(n8451), .ZN(n8189) );
  NAND2_X1 U7443 ( .A1(n8420), .A2(n8431), .ZN(n5903) );
  NOR2_X1 U7444 ( .A1(n8420), .A2(n8431), .ZN(n5902) );
  NAND2_X1 U7445 ( .A1(n8398), .A2(n8417), .ZN(n5904) );
  INV_X1 U7446 ( .A(n8561), .ZN(n5906) );
  NOR2_X1 U7447 ( .A1(n8362), .A2(n7973), .ZN(n5908) );
  XNOR2_X1 U7448 ( .A(n5909), .B(n5944), .ZN(n5919) );
  NAND2_X1 U7449 ( .A1(n5910), .A2(n8338), .ZN(n6546) );
  NAND2_X1 U7450 ( .A1(n5949), .A2(n6873), .ZN(n5911) );
  INV_X1 U7451 ( .A(n5855), .ZN(n5912) );
  INV_X1 U7452 ( .A(n7140), .ZN(n7135) );
  NAND2_X1 U7453 ( .A1(n5912), .A2(n7135), .ZN(n5913) );
  NAND2_X1 U7454 ( .A1(n5261), .A2(n5913), .ZN(n5914) );
  INV_X1 U7455 ( .A(n5914), .ZN(n6886) );
  AND2_X1 U7456 ( .A1(n5261), .A2(P2_B_REG_SCAN_IN), .ZN(n5915) );
  NOR2_X1 U7457 ( .A1(n9863), .A2(n5915), .ZN(n8351) );
  XNOR2_X1 U7458 ( .A(n5920), .B(P2_B_REG_SCAN_IN), .ZN(n5922) );
  NAND2_X1 U7459 ( .A1(n5920), .A2(n7784), .ZN(n6761) );
  OR2_X1 U7460 ( .A1(n5925), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U7461 ( .A1(n5921), .A2(n7784), .ZN(n5926) );
  NAND2_X1 U7462 ( .A1(n6872), .A2(n6616), .ZN(n6822) );
  NOR2_X1 U7463 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .ZN(
        n5931) );
  NOR4_X1 U7464 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5930) );
  NOR4_X1 U7465 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5929) );
  NOR4_X1 U7466 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5928) );
  NAND4_X1 U7467 ( .A1(n5931), .A2(n5930), .A3(n5929), .A4(n5928), .ZN(n5937)
         );
  NOR4_X1 U7468 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n5935) );
  NOR4_X1 U7469 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5934) );
  NOR4_X1 U7470 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5933) );
  NOR4_X1 U7471 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n5932) );
  NAND4_X1 U7472 ( .A1(n5935), .A2(n5934), .A3(n5933), .A4(n5932), .ZN(n5936)
         );
  NOR2_X1 U7473 ( .A1(n5937), .A2(n5936), .ZN(n5938) );
  OR2_X1 U7474 ( .A1(n5925), .A2(n5938), .ZN(n6547) );
  NAND2_X1 U7475 ( .A1(n6575), .A2(n5939), .ZN(n6823) );
  AND3_X1 U7476 ( .A1(n6547), .A2(n6721), .A3(n6823), .ZN(n5940) );
  NOR2_X1 U7477 ( .A1(n7484), .A2(n8338), .ZN(n5947) );
  NAND2_X1 U7478 ( .A1(n5947), .A2(n6873), .ZN(n5942) );
  MUX2_X1 U7479 ( .A(n6872), .B(n6616), .S(n6533), .Z(n5943) );
  NAND2_X1 U7480 ( .A1(n6538), .A2(n5943), .ZN(n5953) );
  NAND2_X1 U7481 ( .A1(n6875), .A2(n7484), .ZN(n9911) );
  NOR2_X1 U7482 ( .A1(n9911), .A2(n5949), .ZN(n6532) );
  OAI211_X1 U7483 ( .C1(n5948), .C2(n5947), .A(n5946), .B(n9915), .ZN(n9862)
         );
  NAND2_X1 U7484 ( .A1(n5949), .A2(n6875), .ZN(n7648) );
  NAND2_X1 U7485 ( .A1(n9862), .A2(n7648), .ZN(n5950) );
  NOR2_X1 U7486 ( .A1(n6531), .A2(n8552), .ZN(n5955) );
  INV_X1 U7487 ( .A(n9860), .ZN(n8466) );
  NAND2_X1 U7488 ( .A1(n5951), .A2(n8466), .ZN(n8354) );
  OAI21_X1 U7489 ( .B1(n9872), .B2(n10201), .A(n8354), .ZN(n5954) );
  INV_X1 U7490 ( .A(n6875), .ZN(n5952) );
  NAND2_X1 U7491 ( .A1(n9927), .A2(n5952), .ZN(n9858) );
  XNOR2_X1 U7492 ( .A(n5957), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9617) );
  NOR2_X2 U7493 ( .A1(n6112), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6115) );
  NOR2_X1 U7494 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5961) );
  NOR2_X1 U7495 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5960) );
  NOR2_X1 U7496 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5959) );
  NOR2_X1 U7497 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5965) );
  NOR2_X1 U7498 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5964) );
  NOR2_X1 U7499 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5963) );
  INV_X1 U7500 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7501 ( .A1(n5985), .A2(n5987), .ZN(n5966) );
  INV_X1 U7502 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5967) );
  INV_X1 U7503 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5969) );
  INV_X1 U7504 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5970) );
  XNOR2_X2 U7505 ( .A(n5971), .B(n5970), .ZN(n9651) );
  MUX2_X1 U7506 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9617), .S(n6607), .Z(n6973) );
  INV_X1 U7507 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5973) );
  INV_X1 U7508 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n10189) );
  INV_X1 U7509 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7510 ( .A1(n6326), .A2(n5975), .ZN(n5976) );
  NAND2_X1 U7511 ( .A1(n5978), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5980) );
  INV_X1 U7512 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5979) );
  XNOR2_X1 U7513 ( .A(n5980), .B(n5979), .ZN(n9050) );
  NAND2_X1 U7514 ( .A1(n5982), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5983) );
  XNOR2_X1 U7515 ( .A(n5983), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6484) );
  NAND2_X1 U7516 ( .A1(n5984), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7517 ( .A1(n5988), .A2(n5987), .ZN(n5990) );
  OR2_X1 U7518 ( .A1(n5988), .A2(n5987), .ZN(n5989) );
  NAND2_X1 U7519 ( .A1(n5990), .A2(n5989), .ZN(n7684) );
  NAND2_X2 U7520 ( .A1(n5991), .A2(n6484), .ZN(n6572) );
  INV_X1 U7521 ( .A(n5992), .ZN(n5993) );
  NAND2_X1 U7522 ( .A1(n5993), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5994) );
  INV_X1 U7523 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7524 ( .A1(n5996), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n5997) );
  NAND2_X2 U7525 ( .A1(n4420), .A2(n7279), .ZN(n9125) );
  NOR2_X1 U7526 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n6002) );
  NAND2_X1 U7527 ( .A1(n6003), .A2(n6002), .ZN(n9606) );
  INV_X1 U7528 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9603) );
  NAND2_X1 U7529 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n6005) );
  NAND2_X1 U7530 ( .A1(n6006), .A2(n6005), .ZN(n6007) );
  XNOR2_X2 U7531 ( .A(n6007), .B(P1_IR_REG_29__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7532 ( .A1(n6041), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7533 ( .A1(n6010), .A2(n6012), .ZN(n6069) );
  INV_X1 U7534 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6009) );
  OR2_X1 U7535 ( .A1(n6069), .A2(n6009), .ZN(n6016) );
  NAND2_X2 U7536 ( .A1(n6011), .A2(n6010), .ZN(n8873) );
  INV_X1 U7537 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6938) );
  OR2_X1 U7538 ( .A1(n8873), .A2(n6938), .ZN(n6015) );
  NAND2_X4 U7539 ( .A1(n6012), .A2(n7924), .ZN(n8871) );
  INV_X1 U7540 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6013) );
  INV_X2 U7541 ( .A(n6062), .ZN(n6333) );
  NAND2_X1 U7542 ( .A1(n6974), .A2(n6333), .ZN(n6018) );
  AND2_X1 U7543 ( .A1(n6019), .A2(n6018), .ZN(n6024) );
  INV_X1 U7544 ( .A(n6024), .ZN(n6025) );
  NAND2_X1 U7545 ( .A1(n6974), .A2(n7927), .ZN(n6021) );
  NAND2_X1 U7546 ( .A1(n6973), .A2(n6333), .ZN(n6020) );
  INV_X1 U7547 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9666) );
  NAND2_X1 U7548 ( .A1(n6022), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7549 ( .A1(n6024), .A2(n6023), .ZN(n6724) );
  OAI21_X1 U7550 ( .B1(n6025), .B2(n4429), .A(n6722), .ZN(n6767) );
  INV_X1 U7551 ( .A(n6027), .ZN(n6028) );
  NAND2_X4 U7552 ( .A1(n6607), .A2(n5259), .ZN(n8880) );
  INV_X1 U7553 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6582) );
  NAND2_X1 U7554 ( .A1(n6041), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6032) );
  INV_X1 U7555 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6029) );
  OR2_X1 U7556 ( .A1(n6069), .A2(n6029), .ZN(n6031) );
  INV_X1 U7557 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6030) );
  INV_X1 U7558 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U7559 ( .A1(n6964), .A2(n6333), .ZN(n6033) );
  INV_X1 U7560 ( .A(n6964), .ZN(n6975) );
  OAI22_X1 U7561 ( .A1(n6975), .A2(n4418), .B1(n9749), .B2(n6320), .ZN(n6037)
         );
  XNOR2_X1 U7562 ( .A(n6036), .B(n6037), .ZN(n6768) );
  INV_X1 U7563 ( .A(n6036), .ZN(n6039) );
  INV_X1 U7564 ( .A(n6037), .ZN(n6038) );
  INV_X1 U7565 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6040) );
  INV_X1 U7566 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6867) );
  OR2_X1 U7567 ( .A1(n6069), .A2(n6867), .ZN(n6045) );
  INV_X1 U7568 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6639) );
  OR2_X1 U7569 ( .A1(n8871), .A2(n6639), .ZN(n6044) );
  INV_X1 U7570 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6042) );
  OR2_X1 U7571 ( .A1(n6027), .A2(n5968), .ZN(n6047) );
  XNOR2_X1 U7572 ( .A(n6047), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9676) );
  INV_X1 U7573 ( .A(n9676), .ZN(n6583) );
  OR2_X1 U7574 ( .A1(n7899), .A2(n6584), .ZN(n6049) );
  INV_X1 U7575 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6585) );
  OR2_X1 U7576 ( .A1(n8880), .A2(n6585), .ZN(n6048) );
  OAI211_X1 U7577 ( .C1(n6607), .C2(n6583), .A(n6049), .B(n6048), .ZN(n6982)
         );
  OAI22_X1 U7578 ( .A1(n6979), .A2(n4418), .B1(n9756), .B2(n6320), .ZN(n6051)
         );
  XNOR2_X1 U7579 ( .A(n6052), .B(n6051), .ZN(n6863) );
  NAND2_X1 U7580 ( .A1(n8870), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6056) );
  OR2_X1 U7581 ( .A1(n6069), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6055) );
  INV_X1 U7582 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6985) );
  OR2_X1 U7583 ( .A1(n8873), .A2(n6985), .ZN(n6054) );
  INV_X1 U7584 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6638) );
  OR2_X1 U7585 ( .A1(n8871), .A2(n6638), .ZN(n6053) );
  OR2_X1 U7586 ( .A1(n6997), .A2(n4418), .ZN(n6061) );
  NAND2_X1 U7587 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4455), .ZN(n6057) );
  XNOR2_X1 U7588 ( .A(n6057), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6637) );
  INV_X1 U7589 ( .A(n6637), .ZN(n6665) );
  OR2_X1 U7590 ( .A1(n7899), .A2(n6579), .ZN(n6059) );
  OR2_X1 U7591 ( .A1(n8880), .A2(n6580), .ZN(n6058) );
  OAI211_X1 U7592 ( .C1(n6607), .C2(n6665), .A(n6059), .B(n6058), .ZN(n6987)
         );
  NAND2_X1 U7593 ( .A1(n6987), .A2(n6333), .ZN(n6060) );
  NAND2_X1 U7594 ( .A1(n6061), .A2(n6060), .ZN(n6065) );
  OAI22_X1 U7595 ( .A1(n6997), .A2(n6320), .B1(n9800), .B2(n6476), .ZN(n6063)
         );
  XNOR2_X1 U7596 ( .A(n6063), .B(n4429), .ZN(n6064) );
  XOR2_X1 U7597 ( .A(n6065), .B(n6064), .Z(n6893) );
  INV_X1 U7598 ( .A(n6064), .ZN(n6067) );
  INV_X1 U7599 ( .A(n6065), .ZN(n6066) );
  NAND2_X1 U7600 ( .A1(n8870), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6074) );
  INV_X1 U7601 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6068) );
  OR2_X1 U7602 ( .A1(n8871), .A2(n6068), .ZN(n6073) );
  OAI21_X1 U7603 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n6089), .ZN(n7001) );
  OR2_X1 U7604 ( .A1(n6516), .A2(n7001), .ZN(n6072) );
  INV_X1 U7605 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7002) );
  OR2_X1 U7606 ( .A1(n8873), .A2(n7002), .ZN(n6071) );
  NAND4_X1 U7607 ( .A1(n6074), .A2(n6073), .A3(n6072), .A4(n6071), .ZN(n9144)
         );
  NAND2_X1 U7608 ( .A1(n9144), .A2(n6333), .ZN(n6082) );
  NAND2_X1 U7609 ( .A1(n6075), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6077) );
  INV_X1 U7610 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7611 ( .A1(n6077), .A2(n6076), .ZN(n6095) );
  OR2_X1 U7612 ( .A1(n6077), .A2(n6076), .ZN(n6078) );
  OR2_X1 U7613 ( .A1(n7899), .A2(n6587), .ZN(n6080) );
  OR2_X1 U7614 ( .A1(n8880), .A2(n6586), .ZN(n6079) );
  OAI211_X1 U7615 ( .C1(n6607), .C2(n6776), .A(n6080), .B(n6079), .ZN(n7004)
         );
  NAND2_X1 U7616 ( .A1(n7004), .A2(n7931), .ZN(n6081) );
  NAND2_X1 U7617 ( .A1(n6082), .A2(n6081), .ZN(n6083) );
  XNOR2_X1 U7618 ( .A(n6083), .B(n4429), .ZN(n6084) );
  AOI22_X1 U7619 ( .A1(n9144), .A2(n7927), .B1(n7004), .B2(n6333), .ZN(n6085)
         );
  XNOR2_X1 U7620 ( .A(n6084), .B(n6085), .ZN(n6940) );
  NAND2_X1 U7621 ( .A1(n6941), .A2(n6940), .ZN(n6939) );
  INV_X1 U7622 ( .A(n6085), .ZN(n6086) );
  INV_X1 U7623 ( .A(n6101), .ZN(n6103) );
  NAND2_X1 U7624 ( .A1(n8870), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6094) );
  INV_X1 U7625 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6635) );
  OR2_X1 U7626 ( .A1(n8871), .A2(n6635), .ZN(n6093) );
  INV_X1 U7627 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10045) );
  NAND2_X1 U7628 ( .A1(n6089), .A2(n10045), .ZN(n6090) );
  NAND2_X1 U7629 ( .A1(n6106), .A2(n6090), .ZN(n7311) );
  OR2_X1 U7630 ( .A1(n6516), .A2(n7311), .ZN(n6092) );
  INV_X1 U7631 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7044) );
  OR2_X1 U7632 ( .A1(n8873), .A2(n7044), .ZN(n6091) );
  NAND2_X1 U7633 ( .A1(n6095), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6096) );
  XNOR2_X1 U7634 ( .A(n6096), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6634) );
  INV_X1 U7635 ( .A(n6634), .ZN(n6690) );
  OR2_X1 U7636 ( .A1(n7899), .A2(n6590), .ZN(n6098) );
  OR2_X1 U7637 ( .A1(n8880), .A2(n6591), .ZN(n6097) );
  OAI211_X1 U7638 ( .C1(n6607), .C2(n6690), .A(n6098), .B(n6097), .ZN(n7049)
         );
  OAI22_X1 U7639 ( .A1(n7229), .A2(n6320), .B1(n7322), .B2(n4521), .ZN(n6099)
         );
  XNOR2_X1 U7640 ( .A(n6099), .B(n4429), .ZN(n6100) );
  INV_X1 U7641 ( .A(n6100), .ZN(n6102) );
  OAI22_X1 U7642 ( .A1(n7229), .A2(n4418), .B1(n7322), .B2(n6320), .ZN(n7309)
         );
  NAND2_X1 U7643 ( .A1(n8870), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6111) );
  INV_X1 U7644 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6633) );
  OR2_X1 U7645 ( .A1(n8871), .A2(n6633), .ZN(n6110) );
  INV_X1 U7646 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7647 ( .A1(n6106), .A2(n6105), .ZN(n6107) );
  NAND2_X1 U7648 ( .A1(n6126), .A2(n6107), .ZN(n7478) );
  OR2_X1 U7649 ( .A1(n6516), .A2(n7478), .ZN(n6109) );
  INV_X1 U7650 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7233) );
  OR2_X1 U7651 ( .A1(n8873), .A2(n7233), .ZN(n6108) );
  NAND2_X1 U7652 ( .A1(n6112), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6113) );
  MUX2_X1 U7653 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6113), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n6114) );
  INV_X1 U7654 ( .A(n6114), .ZN(n6117) );
  NOR2_X1 U7655 ( .A1(n6117), .A2(n6116), .ZN(n6632) );
  INV_X1 U7656 ( .A(n6632), .ZN(n6702) );
  OR2_X1 U7657 ( .A1(n7899), .A2(n6592), .ZN(n6119) );
  OR2_X1 U7658 ( .A1(n8880), .A2(n9975), .ZN(n6118) );
  OAI211_X1 U7659 ( .C1(n6607), .C2(n6702), .A(n6119), .B(n6118), .ZN(n7480)
         );
  INV_X1 U7660 ( .A(n7480), .ZN(n7488) );
  OAI22_X1 U7661 ( .A1(n7534), .A2(n6320), .B1(n7488), .B2(n4521), .ZN(n6120)
         );
  XNOR2_X1 U7662 ( .A(n6120), .B(n4429), .ZN(n6124) );
  OR2_X1 U7663 ( .A1(n7534), .A2(n4418), .ZN(n6122) );
  NAND2_X1 U7664 ( .A1(n7480), .A2(n6333), .ZN(n6121) );
  NAND2_X1 U7665 ( .A1(n6122), .A2(n6121), .ZN(n6123) );
  XNOR2_X1 U7666 ( .A(n6124), .B(n6123), .ZN(n7475) );
  INV_X1 U7667 ( .A(n7533), .ZN(n6143) );
  NAND2_X1 U7668 ( .A1(n8870), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6131) );
  INV_X1 U7669 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9703) );
  OR2_X1 U7670 ( .A1(n8873), .A2(n9703), .ZN(n6130) );
  INV_X1 U7671 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6648) );
  NAND2_X1 U7672 ( .A1(n6126), .A2(n6648), .ZN(n6127) );
  NAND2_X1 U7673 ( .A1(n6149), .A2(n6127), .ZN(n9702) );
  OR2_X1 U7674 ( .A1(n6516), .A2(n9702), .ZN(n6129) );
  INV_X1 U7675 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6645) );
  OR2_X1 U7676 ( .A1(n8871), .A2(n6645), .ZN(n6128) );
  OR2_X1 U7677 ( .A1(n6116), .A2(n5968), .ZN(n6132) );
  XNOR2_X1 U7678 ( .A(n6132), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6671) );
  AOI22_X1 U7679 ( .A1(n6342), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6341), .B2(
        n6671), .ZN(n6134) );
  OR2_X1 U7680 ( .A1(n6595), .A2(n7899), .ZN(n6133) );
  NAND2_X1 U7681 ( .A1(n9705), .A2(n7931), .ZN(n6135) );
  OAI21_X1 U7682 ( .B1(n7491), .B2(n6320), .A(n6135), .ZN(n6137) );
  XNOR2_X1 U7683 ( .A(n6137), .B(n6136), .ZN(n7531) );
  OR2_X1 U7684 ( .A1(n7491), .A2(n4418), .ZN(n6139) );
  NAND2_X1 U7685 ( .A1(n9705), .A2(n6333), .ZN(n6138) );
  NAND2_X1 U7686 ( .A1(n7531), .A2(n7530), .ZN(n6142) );
  INV_X1 U7687 ( .A(n7531), .ZN(n6141) );
  INV_X1 U7688 ( .A(n7530), .ZN(n6140) );
  OR2_X1 U7689 ( .A1(n6597), .A2(n7899), .ZN(n6146) );
  INV_X1 U7690 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7691 ( .A1(n6116), .A2(n6144), .ZN(n6181) );
  NAND2_X1 U7692 ( .A1(n6181), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6160) );
  XNOR2_X1 U7693 ( .A(n6160), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6710) );
  AOI22_X1 U7694 ( .A1(n6342), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6341), .B2(
        n6710), .ZN(n6145) );
  NAND2_X1 U7695 ( .A1(n6146), .A2(n6145), .ZN(n7779) );
  NAND2_X1 U7696 ( .A1(n8870), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6154) );
  INV_X1 U7697 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6674) );
  OR2_X1 U7698 ( .A1(n8871), .A2(n6674), .ZN(n6153) );
  INV_X1 U7699 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7700 ( .A1(n6149), .A2(n6148), .ZN(n6150) );
  NAND2_X1 U7701 ( .A1(n6166), .A2(n6150), .ZN(n7777) );
  OR2_X1 U7702 ( .A1(n6516), .A2(n7777), .ZN(n6152) );
  INV_X1 U7703 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7502) );
  OR2_X1 U7704 ( .A1(n8873), .A2(n7502), .ZN(n6151) );
  OAI22_X1 U7705 ( .A1(n9768), .A2(n4521), .B1(n7548), .B2(n6320), .ZN(n6155)
         );
  XOR2_X1 U7706 ( .A(n4429), .B(n6155), .Z(n6156) );
  OAI21_X1 U7707 ( .B1(n6157), .B2(n6156), .A(n6158), .ZN(n7772) );
  OAI22_X1 U7708 ( .A1(n9768), .A2(n6320), .B1(n7548), .B2(n4418), .ZN(n7773)
         );
  INV_X1 U7709 ( .A(n6158), .ZN(n6159) );
  OR2_X1 U7710 ( .A1(n6600), .A2(n7899), .ZN(n6164) );
  INV_X1 U7711 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7712 ( .A1(n6160), .A2(n6178), .ZN(n6161) );
  NAND2_X1 U7713 ( .A1(n6161), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6162) );
  XNOR2_X1 U7714 ( .A(n6162), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6736) );
  AOI22_X1 U7715 ( .A1(n6342), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6341), .B2(
        n6736), .ZN(n6163) );
  NAND2_X1 U7716 ( .A1(n8870), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6172) );
  INV_X1 U7717 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6165) );
  OR2_X1 U7718 ( .A1(n8871), .A2(n6165), .ZN(n6171) );
  NAND2_X1 U7719 ( .A1(n6166), .A2(n10217), .ZN(n6167) );
  NAND2_X1 U7720 ( .A1(n6198), .A2(n6167), .ZN(n7553) );
  OR2_X1 U7721 ( .A1(n6516), .A2(n7553), .ZN(n6170) );
  INV_X1 U7722 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6168) );
  OR2_X1 U7723 ( .A1(n8873), .A2(n6168), .ZN(n6169) );
  NOR2_X1 U7724 ( .A1(n7518), .A2(n6320), .ZN(n6173) );
  AOI21_X1 U7725 ( .B1(n7627), .B2(n7931), .A(n6173), .ZN(n6174) );
  XNOR2_X1 U7726 ( .A(n6174), .B(n4429), .ZN(n6177) );
  NOR2_X1 U7727 ( .A1(n7518), .A2(n4418), .ZN(n6175) );
  AOI21_X1 U7728 ( .B1(n7627), .B2(n7926), .A(n6175), .ZN(n6176) );
  NOR2_X1 U7729 ( .A1(n6177), .A2(n6176), .ZN(n8776) );
  NAND2_X1 U7730 ( .A1(n6177), .A2(n6176), .ZN(n8777) );
  NAND2_X1 U7731 ( .A1(n6611), .A2(n8877), .ZN(n6184) );
  NAND2_X1 U7732 ( .A1(n6179), .A2(n6178), .ZN(n6180) );
  NOR2_X1 U7733 ( .A1(n6193), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6218) );
  OR2_X1 U7734 ( .A1(n6218), .A2(n5968), .ZN(n6182) );
  XNOR2_X1 U7735 ( .A(n6182), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6853) );
  AOI22_X1 U7736 ( .A1(n6342), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6341), .B2(
        n6853), .ZN(n6183) );
  AND2_X2 U7737 ( .A1(n6184), .A2(n6183), .ZN(n9696) );
  NAND2_X1 U7738 ( .A1(n8870), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6191) );
  INV_X1 U7739 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6798) );
  OR2_X1 U7740 ( .A1(n8871), .A2(n6798), .ZN(n6190) );
  INV_X1 U7741 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6801) );
  NAND2_X1 U7742 ( .A1(n6200), .A2(n6801), .ZN(n6186) );
  NAND2_X1 U7743 ( .A1(n6225), .A2(n6186), .ZN(n9692) );
  OR2_X1 U7744 ( .A1(n6516), .A2(n9692), .ZN(n6189) );
  INV_X1 U7745 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6187) );
  OR2_X1 U7746 ( .A1(n8873), .A2(n6187), .ZN(n6188) );
  OAI22_X1 U7747 ( .A1(n9696), .A2(n4521), .B1(n7668), .B2(n6320), .ZN(n6192)
         );
  XNOR2_X1 U7748 ( .A(n6192), .B(n4429), .ZN(n8824) );
  AOI22_X1 U7749 ( .A1(n4422), .A2(n7926), .B1(n7927), .B2(n4957), .ZN(n8823)
         );
  INV_X1 U7750 ( .A(n8823), .ZN(n6210) );
  NAND2_X1 U7751 ( .A1(n6602), .A2(n8877), .ZN(n6196) );
  NAND2_X1 U7752 ( .A1(n6193), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6194) );
  XNOR2_X1 U7753 ( .A(n6194), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6792) );
  AOI22_X1 U7754 ( .A1(n6342), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6341), .B2(
        n6792), .ZN(n6195) );
  NAND2_X1 U7755 ( .A1(n8711), .A2(n7931), .ZN(n6206) );
  NAND2_X1 U7756 ( .A1(n8870), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6204) );
  INV_X1 U7757 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6739) );
  OR2_X1 U7758 ( .A1(n8871), .A2(n6739), .ZN(n6203) );
  INV_X1 U7759 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7760 ( .A1(n6198), .A2(n6197), .ZN(n6199) );
  NAND2_X1 U7761 ( .A1(n6200), .A2(n6199), .ZN(n8709) );
  OR2_X1 U7762 ( .A1(n6516), .A2(n8709), .ZN(n6202) );
  INV_X1 U7763 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7524) );
  OR2_X1 U7764 ( .A1(n8873), .A2(n7524), .ZN(n6201) );
  OR2_X1 U7765 ( .A1(n8828), .A2(n6320), .ZN(n6205) );
  NAND2_X1 U7766 ( .A1(n6206), .A2(n6205), .ZN(n6208) );
  XNOR2_X1 U7767 ( .A(n6208), .B(n6136), .ZN(n8822) );
  INV_X1 U7768 ( .A(n8822), .ZN(n6213) );
  NOR2_X1 U7769 ( .A1(n8828), .A2(n4418), .ZN(n6209) );
  AOI21_X1 U7770 ( .B1(n8711), .B2(n7926), .A(n6209), .ZN(n6211) );
  INV_X1 U7771 ( .A(n6211), .ZN(n8705) );
  AOI22_X1 U7772 ( .A1(n8824), .A2(n6210), .B1(n6213), .B2(n8705), .ZN(n6216)
         );
  AOI21_X1 U7773 ( .B1(n8822), .B2(n6211), .A(n8823), .ZN(n6214) );
  NAND2_X1 U7774 ( .A1(n8823), .A2(n6211), .ZN(n6212) );
  OAI22_X1 U7775 ( .A1(n6214), .A2(n8824), .B1(n6213), .B2(n6212), .ZN(n6215)
         );
  NAND2_X1 U7776 ( .A1(n6618), .A2(n8877), .ZN(n6221) );
  INV_X1 U7777 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7778 ( .A1(n6218), .A2(n6217), .ZN(n6219) );
  NAND2_X1 U7779 ( .A1(n6219), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6238) );
  XNOR2_X1 U7780 ( .A(n6238), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6952) );
  AOI22_X1 U7781 ( .A1(n6342), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6341), .B2(
        n6952), .ZN(n6220) );
  NAND2_X1 U7782 ( .A1(n8738), .A2(n7931), .ZN(n6233) );
  NAND2_X1 U7783 ( .A1(n8870), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6231) );
  INV_X1 U7784 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6222) );
  OR2_X1 U7785 ( .A1(n8871), .A2(n6222), .ZN(n6230) );
  INV_X1 U7786 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7787 ( .A1(n6225), .A2(n6224), .ZN(n6226) );
  NAND2_X1 U7788 ( .A1(n6243), .A2(n6226), .ZN(n8736) );
  OR2_X1 U7789 ( .A1(n6516), .A2(n8736), .ZN(n6229) );
  INV_X1 U7790 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6227) );
  OR2_X1 U7791 ( .A1(n8873), .A2(n6227), .ZN(n6228) );
  OR2_X1 U7792 ( .A1(n8827), .A2(n6320), .ZN(n6232) );
  NAND2_X1 U7793 ( .A1(n6233), .A2(n6232), .ZN(n6234) );
  XNOR2_X1 U7794 ( .A(n6234), .B(n4429), .ZN(n6236) );
  OAI22_X1 U7795 ( .A1(n9780), .A2(n6320), .B1(n8827), .B2(n4418), .ZN(n6235)
         );
  XNOR2_X1 U7796 ( .A(n6236), .B(n6235), .ZN(n8731) );
  NAND2_X1 U7797 ( .A1(n6621), .A2(n8877), .ZN(n6242) );
  INV_X1 U7798 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7799 ( .A1(n6238), .A2(n6237), .ZN(n6239) );
  NAND2_X1 U7800 ( .A1(n6239), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6240) );
  XNOR2_X1 U7801 ( .A(n6240), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7385) );
  AOI22_X1 U7802 ( .A1(n6342), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6341), .B2(
        n7385), .ZN(n6241) );
  NAND2_X1 U7803 ( .A1(n8807), .A2(n7931), .ZN(n6250) );
  NAND2_X1 U7804 ( .A1(n8870), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6248) );
  INV_X1 U7805 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7749) );
  OR2_X1 U7806 ( .A1(n8873), .A2(n7749), .ZN(n6247) );
  INV_X1 U7807 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8803) );
  NAND2_X1 U7808 ( .A1(n6243), .A2(n8803), .ZN(n6244) );
  NAND2_X1 U7809 ( .A1(n6260), .A2(n6244), .ZN(n8804) );
  OR2_X1 U7810 ( .A1(n6516), .A2(n8804), .ZN(n6246) );
  INV_X1 U7811 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6955) );
  OR2_X1 U7812 ( .A1(n8871), .A2(n6955), .ZN(n6245) );
  OR2_X1 U7813 ( .A1(n8686), .A2(n6320), .ZN(n6249) );
  NAND2_X1 U7814 ( .A1(n6250), .A2(n6249), .ZN(n6251) );
  XNOR2_X1 U7815 ( .A(n6251), .B(n4429), .ZN(n6252) );
  INV_X1 U7816 ( .A(n8686), .ZN(n9462) );
  AOI22_X1 U7817 ( .A1(n8807), .A2(n7926), .B1(n7927), .B2(n9462), .ZN(n6253)
         );
  XNOR2_X1 U7818 ( .A(n6252), .B(n6253), .ZN(n8801) );
  INV_X1 U7819 ( .A(n6252), .ZN(n6254) );
  NAND2_X1 U7820 ( .A1(n6727), .A2(n8877), .ZN(n6258) );
  NOR2_X1 U7821 ( .A1(n5972), .A2(n5968), .ZN(n6255) );
  MUX2_X1 U7822 ( .A(n5968), .B(n6255), .S(P1_IR_REG_14__SCAN_IN), .Z(n6256)
         );
  NOR2_X1 U7823 ( .A1(n6256), .A2(n6286), .ZN(n7391) );
  AOI22_X1 U7824 ( .A1(n6342), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6341), .B2(
        n7391), .ZN(n6257) );
  INV_X1 U7825 ( .A(n9473), .ZN(n9790) );
  NAND2_X1 U7826 ( .A1(n6517), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6265) );
  INV_X1 U7827 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n6259) );
  OR2_X1 U7828 ( .A1(n6275), .A2(n6259), .ZN(n6264) );
  INV_X1 U7829 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8685) );
  NAND2_X1 U7830 ( .A1(n6260), .A2(n8685), .ZN(n6261) );
  NAND2_X1 U7831 ( .A1(n6291), .A2(n6261), .ZN(n9469) );
  OR2_X1 U7832 ( .A1(n6516), .A2(n9469), .ZN(n6263) );
  INV_X1 U7833 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9470) );
  OR2_X1 U7834 ( .A1(n8873), .A2(n9470), .ZN(n6262) );
  NAND4_X1 U7835 ( .A1(n6265), .A2(n6264), .A3(n6263), .A4(n6262), .ZN(n9437)
         );
  OAI22_X1 U7836 ( .A1(n9790), .A2(n4521), .B1(n8861), .B2(n6320), .ZN(n6266)
         );
  XNOR2_X1 U7837 ( .A(n6266), .B(n4429), .ZN(n8683) );
  AOI22_X1 U7838 ( .A1(n9473), .A2(n7926), .B1(n7927), .B2(n9437), .ZN(n8682)
         );
  NAND2_X1 U7839 ( .A1(n6267), .A2(n8682), .ZN(n6270) );
  INV_X1 U7840 ( .A(n8683), .ZN(n6268) );
  NAND2_X1 U7841 ( .A1(n4910), .A2(n6268), .ZN(n6269) );
  NAND2_X1 U7842 ( .A1(n6270), .A2(n6269), .ZN(n8749) );
  NAND2_X1 U7843 ( .A1(n6763), .A2(n8877), .ZN(n6274) );
  NAND2_X1 U7844 ( .A1(n6271), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6272) );
  XNOR2_X1 U7845 ( .A(n6272), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9170) );
  AOI22_X1 U7846 ( .A1(n6342), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6341), .B2(
        n9170), .ZN(n6273) );
  NAND2_X1 U7847 ( .A1(n9429), .A2(n7931), .ZN(n6284) );
  NAND2_X1 U7848 ( .A1(n8870), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6282) );
  INV_X1 U7849 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9159) );
  OR2_X1 U7850 ( .A1(n8871), .A2(n9159), .ZN(n6281) );
  INV_X1 U7851 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U7852 ( .A1(n6293), .A2(n8755), .ZN(n6278) );
  NAND2_X1 U7853 ( .A1(n6313), .A2(n6278), .ZN(n9426) );
  OR2_X1 U7854 ( .A1(n6516), .A2(n9426), .ZN(n6280) );
  INV_X1 U7855 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9427) );
  OR2_X1 U7856 ( .A1(n8873), .A2(n9427), .ZN(n6279) );
  OR2_X1 U7857 ( .A1(n9440), .A2(n6320), .ZN(n6283) );
  NAND2_X1 U7858 ( .A1(n6284), .A2(n6283), .ZN(n6285) );
  XNOR2_X1 U7859 ( .A(n6285), .B(n4428), .ZN(n8752) );
  INV_X1 U7860 ( .A(n9440), .ZN(n9136) );
  AOI22_X1 U7861 ( .A1(n9429), .A2(n7926), .B1(n7927), .B2(n9136), .ZN(n8751)
         );
  INV_X1 U7862 ( .A(n8751), .ZN(n6303) );
  NAND2_X1 U7863 ( .A1(n6747), .A2(n8877), .ZN(n6289) );
  OR2_X1 U7864 ( .A1(n6286), .A2(n5968), .ZN(n6287) );
  XNOR2_X1 U7865 ( .A(n6287), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9156) );
  AOI22_X1 U7866 ( .A1(n6342), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6341), .B2(
        n9156), .ZN(n6288) );
  NAND2_X1 U7867 ( .A1(n9452), .A2(n7931), .ZN(n6299) );
  NAND2_X1 U7868 ( .A1(n8870), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6297) );
  INV_X1 U7869 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6290) );
  OR2_X1 U7870 ( .A1(n8871), .A2(n6290), .ZN(n6296) );
  INV_X1 U7871 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8857) );
  NAND2_X1 U7872 ( .A1(n6291), .A2(n8857), .ZN(n6292) );
  NAND2_X1 U7873 ( .A1(n6293), .A2(n6292), .ZN(n9445) );
  OR2_X1 U7874 ( .A1(n6516), .A2(n9445), .ZN(n6295) );
  INV_X1 U7875 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9446) );
  OR2_X1 U7876 ( .A1(n8873), .A2(n9446), .ZN(n6294) );
  NAND4_X1 U7877 ( .A1(n6297), .A2(n6296), .A3(n6295), .A4(n6294), .ZN(n9459)
         );
  NAND2_X1 U7878 ( .A1(n9459), .A2(n7926), .ZN(n6298) );
  NAND2_X1 U7879 ( .A1(n6299), .A2(n6298), .ZN(n6300) );
  XNOR2_X1 U7880 ( .A(n6300), .B(n6136), .ZN(n8750) );
  INV_X1 U7881 ( .A(n8750), .ZN(n6306) );
  NAND2_X1 U7882 ( .A1(n9452), .A2(n7926), .ZN(n6302) );
  NAND2_X1 U7883 ( .A1(n9459), .A2(n7927), .ZN(n6301) );
  AND2_X1 U7884 ( .A1(n6302), .A2(n6301), .ZN(n6304) );
  INV_X1 U7885 ( .A(n6304), .ZN(n8855) );
  AOI22_X1 U7886 ( .A1(n8752), .A2(n6303), .B1(n6306), .B2(n8855), .ZN(n6309)
         );
  AOI21_X1 U7887 ( .B1(n8750), .B2(n6304), .A(n8751), .ZN(n6307) );
  NAND2_X1 U7888 ( .A1(n8751), .A2(n6304), .ZN(n6305) );
  OAI22_X1 U7889 ( .A1(n6307), .A2(n8752), .B1(n6306), .B2(n6305), .ZN(n6308)
         );
  NAND2_X1 U7890 ( .A1(n6837), .A2(n8877), .ZN(n6312) );
  NAND2_X1 U7891 ( .A1(n4497), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6310) );
  XNOR2_X1 U7892 ( .A(n6310), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9188) );
  AOI22_X1 U7893 ( .A1(n6342), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6341), .B2(
        n9188), .ZN(n6311) );
  INV_X1 U7894 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n10072) );
  NAND2_X1 U7895 ( .A1(n6313), .A2(n10072), .ZN(n6314) );
  AND2_X1 U7896 ( .A1(n6349), .A2(n6314), .ZN(n9408) );
  NAND2_X1 U7897 ( .A1(n6070), .A2(n9408), .ZN(n6319) );
  INV_X1 U7898 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n6315) );
  OR2_X1 U7899 ( .A1(n6275), .A2(n6315), .ZN(n6318) );
  INV_X1 U7900 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9192) );
  OR2_X1 U7901 ( .A1(n8873), .A2(n9192), .ZN(n6317) );
  INV_X1 U7902 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9175) );
  OR2_X1 U7903 ( .A1(n8871), .A2(n9175), .ZN(n6316) );
  NAND4_X1 U7904 ( .A1(n6319), .A2(n6318), .A3(n6317), .A4(n6316), .ZN(n9422)
         );
  OAI22_X1 U7905 ( .A1(n9631), .A2(n6320), .B1(n9392), .B2(n4418), .ZN(n6323)
         );
  OAI22_X1 U7906 ( .A1(n9631), .A2(n4521), .B1(n9392), .B2(n6320), .ZN(n6321)
         );
  XNOR2_X1 U7907 ( .A(n6321), .B(n4429), .ZN(n6322) );
  XOR2_X1 U7908 ( .A(n6323), .B(n6322), .Z(n8762) );
  NAND2_X1 U7909 ( .A1(n8763), .A2(n8762), .ZN(n8761) );
  INV_X1 U7910 ( .A(n6322), .ZN(n6325) );
  INV_X1 U7911 ( .A(n6323), .ZN(n6324) );
  NAND2_X1 U7912 ( .A1(n8761), .A2(n5030), .ZN(n8837) );
  NAND2_X1 U7913 ( .A1(n6869), .A2(n8877), .ZN(n6328) );
  XNOR2_X1 U7914 ( .A(n6326), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9210) );
  AOI22_X1 U7915 ( .A1(n6342), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6341), .B2(
        n9210), .ZN(n6327) );
  NAND2_X1 U7916 ( .A1(n9542), .A2(n7931), .ZN(n6335) );
  XNOR2_X1 U7917 ( .A(n6349), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n9396) );
  NAND2_X1 U7918 ( .A1(n9396), .A2(n6070), .ZN(n6332) );
  INV_X1 U7919 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9988) );
  OR2_X1 U7920 ( .A1(n8871), .A2(n9988), .ZN(n6331) );
  NAND2_X1 U7921 ( .A1(n8870), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U7922 ( .A1(n7915), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6329) );
  NAND4_X1 U7923 ( .A1(n6332), .A2(n6331), .A3(n6330), .A4(n6329), .ZN(n9379)
         );
  NAND2_X1 U7924 ( .A1(n9379), .A2(n6333), .ZN(n6334) );
  NAND2_X1 U7925 ( .A1(n6335), .A2(n6334), .ZN(n6336) );
  XNOR2_X1 U7926 ( .A(n6336), .B(n4429), .ZN(n8834) );
  NAND2_X1 U7927 ( .A1(n9542), .A2(n7926), .ZN(n6338) );
  NAND2_X1 U7928 ( .A1(n9379), .A2(n7927), .ZN(n6337) );
  NAND2_X1 U7929 ( .A1(n6338), .A2(n6337), .ZN(n8835) );
  NAND2_X1 U7930 ( .A1(n8834), .A2(n8835), .ZN(n6340) );
  NAND2_X1 U7931 ( .A1(n7033), .A2(n8877), .ZN(n6344) );
  AOI22_X1 U7932 ( .A1(n6342), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6341), .B2(
        n4539), .ZN(n6343) );
  NAND2_X1 U7933 ( .A1(n9370), .A2(n7931), .ZN(n6354) );
  INV_X1 U7934 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9372) );
  INV_X1 U7935 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9537) );
  OR2_X1 U7936 ( .A1(n8871), .A2(n9537), .ZN(n6346) );
  INV_X1 U7937 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9590) );
  OR2_X1 U7938 ( .A1(n6275), .A2(n9590), .ZN(n6345) );
  AND2_X1 U7939 ( .A1(n6346), .A2(n6345), .ZN(n6352) );
  AND2_X1 U7940 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n6347) );
  INV_X1 U7941 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8838) );
  INV_X1 U7942 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8719) );
  OAI21_X1 U7943 ( .B1(n6349), .B2(n8838), .A(n8719), .ZN(n6350) );
  NAND2_X1 U7944 ( .A1(n6361), .A2(n6350), .ZN(n9371) );
  OR2_X1 U7945 ( .A1(n9371), .A2(n6516), .ZN(n6351) );
  OAI211_X1 U7946 ( .C1(n8873), .C2(n9372), .A(n6352), .B(n6351), .ZN(n9135)
         );
  NAND2_X1 U7947 ( .A1(n9135), .A2(n7926), .ZN(n6353) );
  NAND2_X1 U7948 ( .A1(n6354), .A2(n6353), .ZN(n6355) );
  XNOR2_X1 U7949 ( .A(n6355), .B(n6136), .ZN(n6358) );
  AND2_X1 U7950 ( .A1(n9135), .A2(n7927), .ZN(n6356) );
  AOI21_X1 U7951 ( .B1(n9370), .B2(n7926), .A(n6356), .ZN(n6357) );
  NAND2_X1 U7952 ( .A1(n6358), .A2(n6357), .ZN(n8717) );
  NAND2_X1 U7953 ( .A1(n8714), .A2(n8717), .ZN(n8791) );
  NAND2_X1 U7954 ( .A1(n7196), .A2(n8877), .ZN(n6360) );
  INV_X1 U7955 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7280) );
  OR2_X1 U7956 ( .A1(n8880), .A2(n7280), .ZN(n6359) );
  INV_X1 U7957 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n10016) );
  NAND2_X1 U7958 ( .A1(n6361), .A2(n10016), .ZN(n6362) );
  NAND2_X1 U7959 ( .A1(n6376), .A2(n6362), .ZN(n8794) );
  AOI22_X1 U7960 ( .A1(n7915), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n8870), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n6364) );
  NAND2_X1 U7961 ( .A1(n6517), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6363) );
  OAI211_X1 U7962 ( .C1(n8794), .C2(n6516), .A(n6364), .B(n6363), .ZN(n9380)
         );
  INV_X1 U7963 ( .A(n9380), .ZN(n8930) );
  OAI22_X1 U7964 ( .A1(n9588), .A2(n6062), .B1(n8930), .B2(n4418), .ZN(n6369)
         );
  NAND2_X1 U7965 ( .A1(n9360), .A2(n7931), .ZN(n6366) );
  NAND2_X1 U7966 ( .A1(n9380), .A2(n7926), .ZN(n6365) );
  NAND2_X1 U7967 ( .A1(n6366), .A2(n6365), .ZN(n6367) );
  XNOR2_X1 U7968 ( .A(n6367), .B(n4429), .ZN(n6368) );
  XOR2_X1 U7969 ( .A(n6369), .B(n6368), .Z(n8792) );
  INV_X1 U7970 ( .A(n6368), .ZN(n6371) );
  INV_X1 U7971 ( .A(n6369), .ZN(n6370) );
  NAND2_X1 U7972 ( .A1(n6371), .A2(n6370), .ZN(n6372) );
  NAND2_X1 U7973 ( .A1(n7333), .A2(n8877), .ZN(n6374) );
  OR2_X1 U7974 ( .A1(n8880), .A2(n10232), .ZN(n6373) );
  NAND2_X1 U7975 ( .A1(n9524), .A2(n7931), .ZN(n6382) );
  INV_X1 U7976 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8726) );
  NAND2_X1 U7977 ( .A1(n6376), .A2(n8726), .ZN(n6377) );
  NAND2_X1 U7978 ( .A1(n6403), .A2(n6377), .ZN(n9335) );
  OR2_X1 U7979 ( .A1(n9335), .A2(n6516), .ZN(n6380) );
  AOI22_X1 U7980 ( .A1(n7915), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n8870), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U7981 ( .A1(n6517), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U7982 ( .A1(n9321), .A2(n7926), .ZN(n6381) );
  NAND2_X1 U7983 ( .A1(n6382), .A2(n6381), .ZN(n6383) );
  XNOR2_X1 U7984 ( .A(n6383), .B(n4428), .ZN(n6384) );
  AOI22_X1 U7985 ( .A1(n9524), .A2(n7926), .B1(n7927), .B2(n9321), .ZN(n6385)
         );
  XNOR2_X1 U7986 ( .A(n6384), .B(n6385), .ZN(n8725) );
  INV_X1 U7987 ( .A(n6384), .ZN(n6386) );
  NAND2_X1 U7988 ( .A1(n6386), .A2(n6385), .ZN(n6387) );
  NAND2_X1 U7989 ( .A1(n7594), .A2(n8877), .ZN(n6389) );
  OR2_X1 U7990 ( .A1(n8880), .A2(n7593), .ZN(n6388) );
  NAND2_X1 U7991 ( .A1(n9514), .A2(n7931), .ZN(n6398) );
  INV_X1 U7992 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6402) );
  INV_X1 U7993 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8699) );
  NAND2_X1 U7994 ( .A1(n6405), .A2(n8699), .ZN(n6391) );
  NAND2_X1 U7995 ( .A1(n6424), .A2(n6391), .ZN(n9305) );
  OR2_X1 U7996 ( .A1(n9305), .A2(n6516), .ZN(n6396) );
  INV_X1 U7997 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10221) );
  NAND2_X1 U7998 ( .A1(n7915), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U7999 ( .A1(n8870), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6392) );
  OAI211_X1 U8000 ( .C1(n8871), .C2(n10221), .A(n6393), .B(n6392), .ZN(n6394)
         );
  INV_X1 U8001 ( .A(n6394), .ZN(n6395) );
  NAND2_X1 U8002 ( .A1(n6396), .A2(n6395), .ZN(n9322) );
  NAND2_X1 U8003 ( .A1(n9322), .A2(n7926), .ZN(n6397) );
  NAND2_X1 U8004 ( .A1(n6398), .A2(n6397), .ZN(n6399) );
  XNOR2_X1 U8005 ( .A(n6399), .B(n4429), .ZN(n8696) );
  OAI22_X1 U8006 ( .A1(n4705), .A2(n6062), .B1(n8771), .B2(n4418), .ZN(n8695)
         );
  NAND2_X1 U8007 ( .A1(n7483), .A2(n8877), .ZN(n6401) );
  OR2_X1 U8008 ( .A1(n8880), .A2(n7487), .ZN(n6400) );
  NAND2_X1 U8009 ( .A1(n9521), .A2(n7926), .ZN(n6412) );
  NAND2_X1 U8010 ( .A1(n6403), .A2(n6402), .ZN(n6404) );
  AND2_X1 U8011 ( .A1(n6405), .A2(n6404), .ZN(n9327) );
  NAND2_X1 U8012 ( .A1(n9327), .A2(n6070), .ZN(n6410) );
  INV_X1 U8013 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9996) );
  NAND2_X1 U8014 ( .A1(n8870), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U8015 ( .A1(n7915), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6406) );
  OAI211_X1 U8016 ( .C1(n8871), .C2(n9996), .A(n6407), .B(n6406), .ZN(n6408)
         );
  INV_X1 U8017 ( .A(n6408), .ZN(n6409) );
  NAND2_X1 U8018 ( .A1(n6410), .A2(n6409), .ZN(n9344) );
  NAND2_X1 U8019 ( .A1(n9344), .A2(n7927), .ZN(n6411) );
  NAND2_X1 U8020 ( .A1(n6412), .A2(n6411), .ZN(n8692) );
  NAND2_X1 U8021 ( .A1(n9521), .A2(n7931), .ZN(n6414) );
  NAND2_X1 U8022 ( .A1(n9344), .A2(n7926), .ZN(n6413) );
  NAND2_X1 U8023 ( .A1(n6414), .A2(n6413), .ZN(n6415) );
  XNOR2_X1 U8024 ( .A(n6415), .B(n4429), .ZN(n8693) );
  AOI22_X1 U8025 ( .A1(n8696), .A2(n8695), .B1(n8692), .B2(n8693), .ZN(n6416)
         );
  INV_X1 U8026 ( .A(n8696), .ZN(n6419) );
  OAI21_X1 U8027 ( .B1(n8693), .B2(n8692), .A(n8695), .ZN(n6418) );
  NOR3_X1 U8028 ( .A1(n8695), .A2(n8692), .A3(n8693), .ZN(n6417) );
  AOI21_X1 U8029 ( .B1(n6419), .B2(n6418), .A(n6417), .ZN(n6420) );
  NAND2_X1 U8030 ( .A1(n7682), .A2(n8877), .ZN(n6422) );
  OR2_X1 U8031 ( .A1(n8880), .A2(n7683), .ZN(n6421) );
  INV_X1 U8032 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n10044) );
  NAND2_X1 U8033 ( .A1(n6424), .A2(n10044), .ZN(n6425) );
  NAND2_X1 U8034 ( .A1(n6443), .A2(n6425), .ZN(n9291) );
  OR2_X1 U8035 ( .A1(n9291), .A2(n6516), .ZN(n6431) );
  INV_X1 U8036 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U8037 ( .A1(n7915), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6427) );
  NAND2_X1 U8038 ( .A1(n8870), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6426) );
  OAI211_X1 U8039 ( .C1(n8871), .C2(n6428), .A(n6427), .B(n6426), .ZN(n6429)
         );
  INV_X1 U8040 ( .A(n6429), .ZN(n6430) );
  NAND2_X1 U8041 ( .A1(n6431), .A2(n6430), .ZN(n9312) );
  OAI22_X1 U8042 ( .A1(n9294), .A2(n6062), .B1(n8952), .B2(n4418), .ZN(n6436)
         );
  NAND2_X1 U8043 ( .A1(n9510), .A2(n7931), .ZN(n6433) );
  NAND2_X1 U8044 ( .A1(n9312), .A2(n7926), .ZN(n6432) );
  NAND2_X1 U8045 ( .A1(n6433), .A2(n6432), .ZN(n6434) );
  XNOR2_X1 U8046 ( .A(n6434), .B(n4429), .ZN(n6435) );
  XOR2_X1 U8047 ( .A(n6436), .B(n6435), .Z(n8770) );
  NAND2_X1 U8048 ( .A1(n8769), .A2(n8770), .ZN(n6440) );
  INV_X1 U8049 ( .A(n6435), .ZN(n6438) );
  INV_X1 U8050 ( .A(n6436), .ZN(n6437) );
  NAND2_X1 U8051 ( .A1(n6438), .A2(n6437), .ZN(n6439) );
  NAND2_X1 U8052 ( .A1(n7765), .A2(n8877), .ZN(n6442) );
  OR2_X1 U8053 ( .A1(n8880), .A2(n10015), .ZN(n6441) );
  INV_X1 U8054 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U8055 ( .A1(n6443), .A2(n8743), .ZN(n6444) );
  NAND2_X1 U8056 ( .A1(n6459), .A2(n6444), .ZN(n9280) );
  OR2_X1 U8057 ( .A1(n9280), .A2(n6516), .ZN(n6449) );
  INV_X1 U8058 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9507) );
  NAND2_X1 U8059 ( .A1(n7915), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6446) );
  NAND2_X1 U8060 ( .A1(n8870), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6445) );
  OAI211_X1 U8061 ( .C1(n8871), .C2(n9507), .A(n6446), .B(n6445), .ZN(n6447)
         );
  INV_X1 U8062 ( .A(n6447), .ZN(n6448) );
  OAI22_X1 U8063 ( .A1(n9580), .A2(n6062), .B1(n9256), .B2(n4418), .ZN(n6452)
         );
  OAI22_X1 U8064 ( .A1(n9580), .A2(n4521), .B1(n9256), .B2(n6320), .ZN(n6450)
         );
  XNOR2_X1 U8065 ( .A(n6450), .B(n4428), .ZN(n6451) );
  XOR2_X1 U8066 ( .A(n6452), .B(n6451), .Z(n8742) );
  INV_X1 U8067 ( .A(n6451), .ZN(n6454) );
  INV_X1 U8068 ( .A(n6452), .ZN(n6453) );
  NAND2_X1 U8069 ( .A1(n6454), .A2(n6453), .ZN(n6455) );
  NAND2_X1 U8070 ( .A1(n7782), .A2(n8877), .ZN(n6457) );
  OR2_X1 U8071 ( .A1(n8880), .A2(n10008), .ZN(n6456) );
  INV_X1 U8072 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U8073 ( .A1(n6459), .A2(n6458), .ZN(n6460) );
  NAND2_X1 U8074 ( .A1(n9264), .A2(n6070), .ZN(n6465) );
  INV_X1 U8075 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10059) );
  NAND2_X1 U8076 ( .A1(n7915), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6462) );
  INV_X1 U8077 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9997) );
  OR2_X1 U8078 ( .A1(n6275), .A2(n9997), .ZN(n6461) );
  OAI211_X1 U8079 ( .C1(n8871), .C2(n10059), .A(n6462), .B(n6461), .ZN(n6463)
         );
  INV_X1 U8080 ( .A(n6463), .ZN(n6464) );
  OAI22_X1 U8081 ( .A1(n9576), .A2(n4521), .B1(n8744), .B2(n6062), .ZN(n6466)
         );
  XNOR2_X1 U8082 ( .A(n6466), .B(n4429), .ZN(n6468) );
  OAI22_X1 U8083 ( .A1(n9576), .A2(n6062), .B1(n8744), .B2(n4418), .ZN(n6467)
         );
  XNOR2_X1 U8084 ( .A(n6468), .B(n6467), .ZN(n8844) );
  INV_X1 U8085 ( .A(n6481), .ZN(n6479) );
  NAND2_X1 U8086 ( .A1(n7965), .A2(n8877), .ZN(n6470) );
  OR2_X1 U8087 ( .A1(n8880), .A2(n9615), .ZN(n6469) );
  XNOR2_X1 U8088 ( .A(n6514), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9246) );
  NAND2_X1 U8089 ( .A1(n9246), .A2(n6070), .ZN(n6475) );
  INV_X1 U8090 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10035) );
  NAND2_X1 U8091 ( .A1(n6517), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6472) );
  NAND2_X1 U8092 ( .A1(n7915), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6471) );
  OAI211_X1 U8093 ( .C1(n6275), .C2(n10035), .A(n6472), .B(n6471), .ZN(n6473)
         );
  INV_X1 U8094 ( .A(n6473), .ZN(n6474) );
  OAI22_X1 U8095 ( .A1(n9573), .A2(n4521), .B1(n9257), .B2(n6320), .ZN(n6477)
         );
  XNOR2_X1 U8096 ( .A(n6477), .B(n4429), .ZN(n7936) );
  OAI22_X1 U8097 ( .A1(n9573), .A2(n6062), .B1(n9257), .B2(n4418), .ZN(n7935)
         );
  XNOR2_X1 U8098 ( .A(n7936), .B(n7935), .ZN(n6480) );
  INV_X1 U8099 ( .A(n6480), .ZN(n6478) );
  NAND2_X1 U8100 ( .A1(n6481), .A2(n6480), .ZN(n6499) );
  NAND2_X1 U8101 ( .A1(n7768), .A2(P1_B_REG_SCAN_IN), .ZN(n6482) );
  MUX2_X1 U8102 ( .A(P1_B_REG_SCAN_IN), .B(n6482), .S(n7684), .Z(n6483) );
  NAND2_X1 U8103 ( .A1(n6483), .A2(n6484), .ZN(n9600) );
  OR2_X1 U8104 ( .A1(n9600), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6485) );
  INV_X1 U8105 ( .A(n6484), .ZN(n7786) );
  NAND2_X1 U8106 ( .A1(n7768), .A2(n7786), .ZN(n9601) );
  NAND2_X1 U8107 ( .A1(n6485), .A2(n9601), .ZN(n6752) );
  INV_X1 U8108 ( .A(n6752), .ZN(n6924) );
  OR2_X1 U8109 ( .A1(n9600), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U8110 ( .A1(n7786), .A2(n7684), .ZN(n9602) );
  NOR4_X1 U8111 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6495) );
  NOR4_X1 U8112 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6494) );
  INV_X1 U8113 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10078) );
  INV_X1 U8114 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10056) );
  INV_X1 U8115 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10160) );
  INV_X1 U8116 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10173) );
  NAND4_X1 U8117 ( .A1(n10078), .A2(n10056), .A3(n10160), .A4(n10173), .ZN(
        n6492) );
  NOR4_X1 U8118 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6490) );
  NOR4_X1 U8119 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6489) );
  NOR4_X1 U8120 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6488) );
  NOR4_X1 U8121 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6487) );
  NAND4_X1 U8122 ( .A1(n6490), .A2(n6489), .A3(n6488), .A4(n6487), .ZN(n6491)
         );
  NOR4_X1 U8123 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6492), .A4(n6491), .ZN(n6493) );
  AND3_X1 U8124 ( .A1(n6495), .A2(n6494), .A3(n6493), .ZN(n6496) );
  OR2_X1 U8125 ( .A1(n9600), .A2(n6496), .ZN(n6922) );
  NAND3_X1 U8126 ( .A1(n6924), .A2(n6807), .A3(n6922), .ZN(n6504) );
  NAND2_X1 U8127 ( .A1(n4496), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6497) );
  XNOR2_X1 U8128 ( .A(n6497), .B(n10001), .ZN(n6609) );
  AND2_X1 U8129 ( .A1(n6609), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6570) );
  NAND2_X1 U8130 ( .A1(n6572), .A2(n6570), .ZN(n9120) );
  OR2_X1 U8131 ( .A1(n6504), .A2(n9120), .ZN(n6524) );
  INV_X1 U8132 ( .A(n6524), .ZN(n6503) );
  NAND2_X1 U8133 ( .A1(n9062), .A2(n9050), .ZN(n6934) );
  INV_X1 U8134 ( .A(n6934), .ZN(n6927) );
  INV_X1 U8135 ( .A(n6754), .ZN(n9115) );
  NAND2_X1 U8136 ( .A1(n4420), .A2(n4550), .ZN(n9013) );
  INV_X1 U8137 ( .A(n9013), .ZN(n6526) );
  NOR2_X1 U8138 ( .A1(n9629), .A2(n6526), .ZN(n6498) );
  OR2_X1 U8139 ( .A1(n6934), .A2(n7279), .ZN(n6935) );
  INV_X1 U8140 ( .A(n6935), .ZN(n6502) );
  NOR2_X1 U8141 ( .A1(n9120), .A2(n6500), .ZN(n6501) );
  AOI21_X1 U8142 ( .B1(n6503), .B2(n6502), .A(n9736), .ZN(n8853) );
  OR2_X1 U8143 ( .A1(n6934), .A2(n6500), .ZN(n6751) );
  NAND2_X1 U8144 ( .A1(n6504), .A2(n6751), .ZN(n6508) );
  OR2_X1 U8145 ( .A1(n9013), .A2(n6754), .ZN(n6506) );
  AND2_X1 U8146 ( .A1(n6572), .A2(n6609), .ZN(n6505) );
  NAND2_X1 U8147 ( .A1(n6506), .A2(n6505), .ZN(n6753) );
  INV_X1 U8148 ( .A(n6753), .ZN(n6507) );
  NAND2_X1 U8149 ( .A1(n6508), .A2(n6507), .ZN(n6509) );
  AOI22_X1 U8150 ( .A1(n9246), .A2(n8847), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6528) );
  INV_X1 U8151 ( .A(n6514), .ZN(n6511) );
  AND2_X1 U8152 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6510) );
  NAND2_X1 U8153 ( .A1(n6511), .A2(n6510), .ZN(n7900) );
  INV_X1 U8154 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6513) );
  INV_X1 U8155 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6512) );
  OAI21_X1 U8156 ( .B1(n6514), .B2(n6513), .A(n6512), .ZN(n6515) );
  NAND2_X1 U8157 ( .A1(n7900), .A2(n6515), .ZN(n7937) );
  INV_X1 U8158 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U8159 ( .A1(n6517), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6519) );
  NAND2_X1 U8160 ( .A1(n8870), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6518) );
  OAI211_X1 U8161 ( .C1(n6520), .C2(n8873), .A(n6519), .B(n6518), .ZN(n6521)
         );
  INV_X1 U8162 ( .A(n6521), .ZN(n6522) );
  NOR2_X1 U8163 ( .A1(n6524), .A2(n9115), .ZN(n8829) );
  INV_X1 U8164 ( .A(n6525), .ZN(n6785) );
  AND2_X1 U8165 ( .A1(n8829), .A2(n9460), .ZN(n8850) );
  AND2_X1 U8166 ( .A1(n8829), .A2(n9461), .ZN(n8813) );
  AOI22_X1 U8167 ( .A1(n9240), .A2(n8850), .B1(n8813), .B2(n9275), .ZN(n6527)
         );
  OAI211_X1 U8168 ( .C1(n9573), .C2(n8853), .A(n6528), .B(n6527), .ZN(n6529)
         );
  OAI21_X1 U8169 ( .B1(n5007), .B2(n6532), .A(n6533), .ZN(n6536) );
  INV_X1 U8170 ( .A(n6533), .ZN(n6534) );
  NAND2_X1 U8171 ( .A1(n6543), .A2(n6534), .ZN(n6535) );
  AND2_X1 U8172 ( .A1(n6536), .A2(n6535), .ZN(n6537) );
  NAND2_X1 U8173 ( .A1(n9939), .A2(n6539), .ZN(n6540) );
  OAI21_X1 U8174 ( .B1(n6553), .B2(n9939), .A(n6540), .ZN(n6542) );
  NAND2_X1 U8175 ( .A1(n6554), .A2(n8607), .ZN(n6541) );
  NAND2_X1 U8176 ( .A1(n6542), .A2(n6541), .ZN(P2_U3488) );
  INV_X1 U8177 ( .A(n6547), .ZN(n6821) );
  NOR2_X1 U8178 ( .A1(n6872), .A2(n6821), .ZN(n6544) );
  AND2_X1 U8179 ( .A1(n6544), .A2(n6543), .ZN(n6831) );
  OAI211_X1 U8180 ( .C1(n7197), .C2(n6546), .A(n5941), .B(n9915), .ZN(n6814)
         );
  NAND2_X1 U8181 ( .A1(n6814), .A2(n9858), .ZN(n6820) );
  NAND2_X1 U8182 ( .A1(n6813), .A2(n6820), .ZN(n6550) );
  NAND2_X1 U8183 ( .A1(n7334), .A2(n6873), .ZN(n6545) );
  NOR2_X1 U8184 ( .A1(n6546), .A2(n6545), .ZN(n6827) );
  NAND2_X1 U8185 ( .A1(n6547), .A2(n6721), .ZN(n6548) );
  NOR2_X1 U8186 ( .A1(n6822), .A2(n6548), .ZN(n6818) );
  OAI21_X1 U8187 ( .B1(n6841), .B2(n6827), .A(n6818), .ZN(n6549) );
  NAND2_X1 U8188 ( .A1(n9929), .A2(n6551), .ZN(n6552) );
  OAI21_X1 U8189 ( .B1(n6553), .B2(n9929), .A(n6552), .ZN(n6556) );
  NAND2_X1 U8190 ( .A1(n6556), .A2(n6555), .ZN(P2_U3456) );
  XNOR2_X1 U8191 ( .A(n6557), .B(n7867), .ZN(n8364) );
  NOR2_X1 U8192 ( .A1(n7871), .A2(n9863), .ZN(n6560) );
  OAI21_X2 U8193 ( .B1(n6562), .B2(n9869), .A(n6561), .ZN(n8359) );
  AOI21_X1 U8194 ( .B1(n9920), .B2(n8364), .A(n8359), .ZN(n6566) );
  NAND2_X1 U8195 ( .A1(n7873), .A2(n8607), .ZN(n6564) );
  NAND2_X1 U8196 ( .A1(n6565), .A2(n6564), .ZN(P2_U3487) );
  INV_X1 U8197 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6567) );
  MUX2_X1 U8198 ( .A(n6567), .B(n6566), .S(n9928), .Z(n6569) );
  NAND2_X1 U8199 ( .A1(n7873), .A2(n8661), .ZN(n6568) );
  NAND2_X1 U8200 ( .A1(n6569), .A2(n6568), .ZN(P2_U3455) );
  INV_X1 U8201 ( .A(n6570), .ZN(n6571) );
  NOR2_X1 U8202 ( .A1(n6572), .A2(n6571), .ZN(n9147) );
  INV_X1 U8203 ( .A(n6574), .ZN(n6573) );
  NOR2_X4 U8204 ( .A1(n7124), .A2(P2_U3151), .ZN(P2_U3893) );
  NAND2_X1 U8205 ( .A1(n6575), .A2(n6574), .ZN(n6576) );
  NAND2_X1 U8206 ( .A1(n7124), .A2(n6576), .ZN(n7152) );
  OAI21_X1 U8207 ( .B1(n7152), .B2(n6577), .A(P2_STATE_REG_SCAN_IN), .ZN(
        P2_U3150) );
  INV_X2 U8208 ( .A(n6622), .ZN(n8679) );
  OAI222_X1 U8209 ( .A1(n8679), .A2(n4507), .B1(n7962), .B2(n6584), .C1(
        P2_U3151), .C2(n4417), .ZN(P2_U3293) );
  OAI222_X1 U8210 ( .A1(n8679), .A2(n6578), .B1(n7962), .B2(n6579), .C1(
        P2_U3151), .C2(n7287), .ZN(P2_U3292) );
  AND2_X1 U8211 ( .A1(n5259), .A2(P1_U3086), .ZN(n6870) );
  INV_X2 U8212 ( .A(n6870), .ZN(n9616) );
  OAI222_X1 U8213 ( .A1(n9616), .A2(n6580), .B1(n7925), .B2(n6579), .C1(
        P1_U3086), .C2(n6665), .ZN(P1_U3352) );
  OAI222_X1 U8214 ( .A1(n9616), .A2(n6582), .B1(n7925), .B2(n6581), .C1(n6641), 
        .C2(P1_U3086), .ZN(P1_U3354) );
  OAI222_X1 U8215 ( .A1(n9616), .A2(n6585), .B1(n7925), .B2(n6584), .C1(
        P1_U3086), .C2(n6583), .ZN(P1_U3353) );
  OAI222_X1 U8216 ( .A1(n9616), .A2(n6586), .B1(n7925), .B2(n6587), .C1(
        P1_U3086), .C2(n6776), .ZN(P1_U3351) );
  OAI222_X1 U8217 ( .A1(n8679), .A2(n6588), .B1(n7962), .B2(n6587), .C1(
        P2_U3151), .C2(n7189), .ZN(P2_U3291) );
  OAI222_X1 U8218 ( .A1(n8679), .A2(n6589), .B1(n7962), .B2(n6590), .C1(
        P2_U3151), .C2(n7165), .ZN(P2_U3290) );
  OAI222_X1 U8219 ( .A1(n9616), .A2(n6591), .B1(n7925), .B2(n6590), .C1(
        P1_U3086), .C2(n6690), .ZN(P1_U3350) );
  OAI222_X1 U8220 ( .A1(n9616), .A2(n9975), .B1(n7925), .B2(n6592), .C1(
        P1_U3086), .C2(n6702), .ZN(P1_U3349) );
  OAI222_X1 U8221 ( .A1(n8679), .A2(n6593), .B1(n7962), .B2(n6592), .C1(
        P2_U3151), .C2(n7268), .ZN(P2_U3289) );
  INV_X1 U8222 ( .A(n6671), .ZN(n6652) );
  OAI222_X1 U8223 ( .A1(n9616), .A2(n6594), .B1(n7925), .B2(n6595), .C1(
        P1_U3086), .C2(n6652), .ZN(P1_U3348) );
  OAI222_X1 U8224 ( .A1(n8679), .A2(n10203), .B1(n7962), .B2(n6595), .C1(
        P2_U3151), .C2(n7365), .ZN(P2_U3288) );
  OAI222_X1 U8225 ( .A1(n8679), .A2(n6596), .B1(n7962), .B2(n6597), .C1(
        P2_U3151), .C2(n9854), .ZN(P2_U3287) );
  INV_X1 U8226 ( .A(n6710), .ZN(n6706) );
  OAI222_X1 U8227 ( .A1(n9616), .A2(n6598), .B1(n7925), .B2(n6597), .C1(
        P1_U3086), .C2(n6706), .ZN(P1_U3347) );
  INV_X1 U8228 ( .A(n6736), .ZN(n6714) );
  OAI222_X1 U8229 ( .A1(n9616), .A2(n6599), .B1(n7925), .B2(n6600), .C1(n6714), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  OAI222_X1 U8230 ( .A1(n8679), .A2(n6601), .B1(n7962), .B2(n6600), .C1(n7441), 
        .C2(P2_U3151), .ZN(P2_U3286) );
  INV_X1 U8231 ( .A(n6602), .ZN(n6604) );
  OAI222_X1 U8232 ( .A1(n8679), .A2(n6603), .B1(n7962), .B2(n6604), .C1(n7638), 
        .C2(P2_U3151), .ZN(P2_U3285) );
  INV_X1 U8233 ( .A(n6792), .ZN(n6797) );
  OAI222_X1 U8234 ( .A1(n9616), .A2(n6605), .B1(n7925), .B2(n6604), .C1(n6797), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U8235 ( .A(n6609), .ZN(n6606) );
  OR2_X1 U8236 ( .A1(n9013), .A2(n6606), .ZN(n6608) );
  AND2_X1 U8237 ( .A1(n6608), .A2(n6607), .ZN(n6628) );
  OR2_X1 U8238 ( .A1(n6609), .A2(P1_U3086), .ZN(n9113) );
  NAND2_X1 U8239 ( .A1(n9120), .A2(n9113), .ZN(n6627) );
  INV_X1 U8240 ( .A(n6627), .ZN(n6610) );
  NOR2_X2 U8241 ( .A1(n6628), .A2(n6610), .ZN(n9673) );
  NOR2_X1 U8242 ( .A1(n9673), .A2(n9147), .ZN(P1_U3085) );
  INV_X1 U8243 ( .A(n6611), .ZN(n6613) );
  INV_X1 U8244 ( .A(n6853), .ZN(n6848) );
  OAI222_X1 U8245 ( .A1(n9616), .A2(n6612), .B1(n7925), .B2(n6613), .C1(
        P1_U3086), .C2(n6848), .ZN(P1_U3344) );
  OAI222_X1 U8246 ( .A1(n8679), .A2(n10163), .B1(n7962), .B2(n6613), .C1(
        P2_U3151), .C2(n7632), .ZN(P2_U3284) );
  INV_X1 U8247 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6615) );
  NAND2_X1 U8248 ( .A1(n6974), .A2(n9147), .ZN(n6614) );
  OAI21_X1 U8249 ( .B1(n9147), .B2(n6615), .A(n6614), .ZN(P1_U3554) );
  INV_X1 U8250 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10219) );
  NAND2_X1 U8251 ( .A1(n6616), .A2(n6721), .ZN(n6617) );
  OAI21_X1 U8252 ( .B1(n6721), .B2(n10219), .A(n6617), .ZN(P2_U3377) );
  INV_X1 U8253 ( .A(n6618), .ZN(n6620) );
  INV_X1 U8254 ( .A(n7732), .ZN(n7795) );
  OAI222_X1 U8255 ( .A1(n8679), .A2(n6619), .B1(n7962), .B2(n6620), .C1(n7795), 
        .C2(P2_U3151), .ZN(P2_U3283) );
  INV_X1 U8256 ( .A(n6952), .ZN(n6851) );
  OAI222_X1 U8257 ( .A1(n9616), .A2(n10178), .B1(n7925), .B2(n6620), .C1(n6851), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8258 ( .A(n6621), .ZN(n6719) );
  AOI22_X1 U8259 ( .A1(n8216), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n6622), .ZN(n6623) );
  OAI21_X1 U8260 ( .B1(n6719), .B2(n7962), .A(n6623), .ZN(P2_U3282) );
  NAND2_X1 U8261 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9663) );
  NOR2_X1 U8262 ( .A1(n9662), .A2(n9663), .ZN(n9661) );
  AOI21_X1 U8263 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n9665), .A(n9661), .ZN(
        n9679) );
  NAND2_X1 U8264 ( .A1(n9676), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6624) );
  OAI21_X1 U8265 ( .B1(n9676), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6624), .ZN(
        n9680) );
  NOR2_X1 U8266 ( .A1(n9679), .A2(n9680), .ZN(n9678) );
  AOI21_X1 U8267 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n9676), .A(n9678), .ZN(
        n6657) );
  NAND2_X1 U8268 ( .A1(n6637), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6625) );
  OAI21_X1 U8269 ( .B1(n6637), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6625), .ZN(
        n6656) );
  NOR2_X1 U8270 ( .A1(n6657), .A2(n6656), .ZN(n6655) );
  AOI21_X1 U8271 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n6637), .A(n6655), .ZN(
        n6779) );
  AOI22_X1 U8272 ( .A1(n6636), .A2(n7002), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n6776), .ZN(n6778) );
  AOI22_X1 U8273 ( .A1(n6634), .A2(n7044), .B1(P1_REG2_REG_5__SCAN_IN), .B2(
        n6690), .ZN(n6682) );
  AOI22_X1 U8274 ( .A1(n6632), .A2(n7233), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n6702), .ZN(n6694) );
  NOR2_X1 U8275 ( .A1(n6695), .A2(n6694), .ZN(n6693) );
  AOI21_X1 U8276 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6632), .A(n6693), .ZN(
        n6631) );
  NAND2_X1 U8277 ( .A1(n6671), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6626) );
  OAI21_X1 U8278 ( .B1(n6671), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6626), .ZN(
        n6630) );
  NOR2_X1 U8279 ( .A1(n6631), .A2(n6630), .ZN(n6668) );
  NAND2_X1 U8280 ( .A1(n6628), .A2(n6627), .ZN(n9659) );
  NOR2_X1 U8281 ( .A1(n6525), .A2(n9651), .ZN(n9122) );
  INV_X1 U8282 ( .A(n9122), .ZN(n6629) );
  AOI211_X1 U8283 ( .C1(n6631), .C2(n6630), .A(n6668), .B(n9660), .ZN(n6654)
         );
  MUX2_X1 U8284 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6633), .S(n6632), .Z(n6697)
         );
  MUX2_X1 U8285 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6635), .S(n6634), .Z(n6685)
         );
  AOI22_X1 U8286 ( .A1(n6636), .A2(P1_REG1_REG_4__SCAN_IN), .B1(n6068), .B2(
        n6776), .ZN(n6774) );
  NAND2_X1 U8287 ( .A1(n6637), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6643) );
  MUX2_X1 U8288 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6638), .S(n6637), .Z(n6659)
         );
  NAND2_X1 U8289 ( .A1(n9676), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6642) );
  MUX2_X1 U8290 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6639), .S(n9676), .Z(n9685)
         );
  MUX2_X1 U8291 ( .A(n6640), .B(P1_REG1_REG_1__SCAN_IN), .S(n6641), .Z(n9668)
         );
  NAND3_X1 U8292 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .A3(n9668), .ZN(n9667) );
  OAI21_X1 U8293 ( .B1(n6641), .B2(n6640), .A(n9667), .ZN(n9686) );
  NAND2_X1 U8294 ( .A1(n9685), .A2(n9686), .ZN(n9683) );
  NAND2_X1 U8295 ( .A1(n6642), .A2(n9683), .ZN(n6660) );
  NAND2_X1 U8296 ( .A1(n6659), .A2(n6660), .ZN(n6658) );
  NAND2_X1 U8297 ( .A1(n6643), .A2(n6658), .ZN(n6773) );
  NAND2_X1 U8298 ( .A1(n6774), .A2(n6773), .ZN(n6644) );
  OAI21_X1 U8299 ( .B1(n6068), .B2(n6776), .A(n6644), .ZN(n6686) );
  NAND2_X1 U8300 ( .A1(n6685), .A2(n6686), .ZN(n6684) );
  OAI21_X1 U8301 ( .B1(n6690), .B2(n6635), .A(n6684), .ZN(n6698) );
  NAND2_X1 U8302 ( .A1(n6697), .A2(n6698), .ZN(n6696) );
  OAI21_X1 U8303 ( .B1(n6702), .B2(n6633), .A(n6696), .ZN(n6647) );
  MUX2_X1 U8304 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6645), .S(n6671), .Z(n6646)
         );
  INV_X1 U8305 ( .A(n9651), .ZN(n7919) );
  OR2_X1 U8306 ( .A1(n9659), .A2(n7919), .ZN(n9213) );
  NAND2_X1 U8307 ( .A1(n6646), .A2(n6647), .ZN(n6672) );
  OAI211_X1 U8308 ( .C1(n6647), .C2(n6646), .A(n9684), .B(n6672), .ZN(n6651)
         );
  NOR2_X1 U8309 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6648), .ZN(n6649) );
  AOI21_X1 U8310 ( .B1(n9673), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n6649), .ZN(
        n6650) );
  OAI211_X1 U8311 ( .C1(n9212), .C2(n6652), .A(n6651), .B(n6650), .ZN(n6653)
         );
  OR2_X1 U8312 ( .A1(n6654), .A2(n6653), .ZN(P1_U3250) );
  AOI211_X1 U8313 ( .C1(n6657), .C2(n6656), .A(n6655), .B(n9660), .ZN(n6667)
         );
  OAI211_X1 U8314 ( .C1(n6660), .C2(n6659), .A(n9684), .B(n6658), .ZN(n6664)
         );
  INV_X1 U8315 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6661) );
  NOR2_X1 U8316 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6661), .ZN(n6662) );
  AOI21_X1 U8317 ( .B1(n9673), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6662), .ZN(
        n6663) );
  OAI211_X1 U8318 ( .C1(n9212), .C2(n6665), .A(n6664), .B(n6663), .ZN(n6666)
         );
  OR2_X1 U8319 ( .A1(n6667), .A2(n6666), .ZN(P1_U3246) );
  AOI22_X1 U8320 ( .A1(n6710), .A2(n7502), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n6706), .ZN(n6669) );
  AOI211_X1 U8321 ( .C1(n6670), .C2(n6669), .A(n6709), .B(n9660), .ZN(n6680)
         );
  NAND2_X1 U8322 ( .A1(n6671), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U8323 ( .A1(n6673), .A2(n6672), .ZN(n6676) );
  MUX2_X1 U8324 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6674), .S(n6710), .Z(n6675)
         );
  NAND2_X1 U8325 ( .A1(n6675), .A2(n6676), .ZN(n6705) );
  OAI211_X1 U8326 ( .C1(n6676), .C2(n6675), .A(n9684), .B(n6705), .ZN(n6678)
         );
  AND2_X1 U8327 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7774) );
  AOI21_X1 U8328 ( .B1(n9673), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n7774), .ZN(
        n6677) );
  OAI211_X1 U8329 ( .C1(n9212), .C2(n6706), .A(n6678), .B(n6677), .ZN(n6679)
         );
  OR2_X1 U8330 ( .A1(n6680), .A2(n6679), .ZN(P1_U3251) );
  AOI211_X1 U8331 ( .C1(n6683), .C2(n6682), .A(n6681), .B(n9660), .ZN(n6692)
         );
  OAI211_X1 U8332 ( .C1(n6686), .C2(n6685), .A(n9684), .B(n6684), .ZN(n6689)
         );
  NOR2_X1 U8333 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10045), .ZN(n6687) );
  AOI21_X1 U8334 ( .B1(n9673), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n6687), .ZN(
        n6688) );
  OAI211_X1 U8335 ( .C1(n9212), .C2(n6690), .A(n6689), .B(n6688), .ZN(n6691)
         );
  OR2_X1 U8336 ( .A1(n6692), .A2(n6691), .ZN(P1_U3248) );
  AOI211_X1 U8337 ( .C1(n6695), .C2(n6694), .A(n6693), .B(n9660), .ZN(n6704)
         );
  OAI211_X1 U8338 ( .C1(n6698), .C2(n6697), .A(n9684), .B(n6696), .ZN(n6701)
         );
  AND2_X1 U8339 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6699) );
  AOI21_X1 U8340 ( .B1(n9673), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n6699), .ZN(
        n6700) );
  OAI211_X1 U8341 ( .C1(n9212), .C2(n6702), .A(n6701), .B(n6700), .ZN(n6703)
         );
  OR2_X1 U8342 ( .A1(n6704), .A2(n6703), .ZN(P1_U3249) );
  AOI22_X1 U8343 ( .A1(n6736), .A2(n6165), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6714), .ZN(n6708) );
  OAI21_X1 U8344 ( .B1(n6674), .B2(n6706), .A(n6705), .ZN(n6707) );
  NOR2_X1 U8345 ( .A1(n6708), .A2(n6707), .ZN(n6738) );
  AOI21_X1 U8346 ( .B1(n6708), .B2(n6707), .A(n6738), .ZN(n6718) );
  AOI22_X1 U8347 ( .A1(n6736), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n6168), .B2(
        n6714), .ZN(n6712) );
  OAI21_X1 U8348 ( .B1(n6712), .B2(n6711), .A(n6733), .ZN(n6713) );
  INV_X1 U8349 ( .A(n9660), .ZN(n9682) );
  NAND2_X1 U8350 ( .A1(n6713), .A2(n9682), .ZN(n6717) );
  AND2_X1 U8351 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8781) );
  NOR2_X1 U8352 ( .A1(n9212), .A2(n6714), .ZN(n6715) );
  AOI211_X1 U8353 ( .C1(n9673), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n8781), .B(
        n6715), .ZN(n6716) );
  OAI211_X1 U8354 ( .C1(n6718), .C2(n9213), .A(n6717), .B(n6716), .ZN(P1_U3252) );
  INV_X1 U8355 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6720) );
  INV_X1 U8356 ( .A(n7385), .ZN(n6961) );
  OAI222_X1 U8357 ( .A1(n9616), .A2(n6720), .B1(n7925), .B2(n6719), .C1(
        P1_U3086), .C2(n6961), .ZN(P1_U3342) );
  INV_X1 U8358 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10069) );
  NOR2_X1 U8359 ( .A1(n6760), .A2(n10069), .ZN(P2_U3242) );
  INV_X1 U8360 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10263) );
  NOR2_X1 U8361 ( .A1(n6760), .A2(n10263), .ZN(P2_U3243) );
  INV_X1 U8362 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n10243) );
  NOR2_X1 U8363 ( .A1(n6760), .A2(n10243), .ZN(P2_U3246) );
  INV_X1 U8364 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10159) );
  NOR2_X1 U8365 ( .A1(n6760), .A2(n10159), .ZN(P2_U3254) );
  INV_X1 U8366 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n9973) );
  NOR2_X1 U8367 ( .A1(n6760), .A2(n9973), .ZN(P2_U3261) );
  OAI21_X1 U8368 ( .B1(n6724), .B2(n6723), .A(n6722), .ZN(n6784) );
  NOR2_X1 U8369 ( .A1(n8847), .A2(P1_U3086), .ZN(n6868) );
  INV_X1 U8370 ( .A(n6868), .ZN(n6770) );
  AOI22_X1 U8371 ( .A1(n6770), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n8850), .B2(
        n6964), .ZN(n6726) );
  NAND2_X1 U8372 ( .A1(n8864), .A2(n6973), .ZN(n6725) );
  OAI211_X1 U8373 ( .C1(n6784), .C2(n8866), .A(n6726), .B(n6725), .ZN(P1_U3232) );
  INV_X1 U8374 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6728) );
  INV_X1 U8375 ( .A(n6727), .ZN(n6729) );
  INV_X1 U8376 ( .A(n8231), .ZN(n8243) );
  OAI222_X1 U8377 ( .A1(n8679), .A2(n6728), .B1(n7962), .B2(n6729), .C1(
        P2_U3151), .C2(n8243), .ZN(P2_U3281) );
  INV_X1 U8378 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6730) );
  INV_X1 U8379 ( .A(n7391), .ZN(n7562) );
  OAI222_X1 U8380 ( .A1(n9616), .A2(n6730), .B1(n7925), .B2(n6729), .C1(
        P1_U3086), .C2(n7562), .ZN(P1_U3341) );
  AND2_X1 U8381 ( .A1(n6731), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8382 ( .A1(n6731), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8383 ( .A1(n6731), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8384 ( .A1(n6731), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8385 ( .A1(n6731), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8386 ( .A1(n6731), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8387 ( .A1(n6731), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8388 ( .A1(n6731), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  NAND2_X1 U8389 ( .A1(n6792), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6732) );
  OAI21_X1 U8390 ( .B1(n6792), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6732), .ZN(
        n6735) );
  OAI21_X1 U8391 ( .B1(n6736), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6733), .ZN(
        n6734) );
  NOR2_X1 U8392 ( .A1(n6735), .A2(n6734), .ZN(n6791) );
  AOI211_X1 U8393 ( .C1(n6735), .C2(n6734), .A(n6791), .B(n9660), .ZN(n6746)
         );
  NOR2_X1 U8394 ( .A1(n6736), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6737) );
  NOR2_X1 U8395 ( .A1(n6738), .A2(n6737), .ZN(n6741) );
  MUX2_X1 U8396 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6739), .S(n6792), .Z(n6740)
         );
  NAND2_X1 U8397 ( .A1(n6740), .A2(n6741), .ZN(n6796) );
  OAI211_X1 U8398 ( .C1(n6741), .C2(n6740), .A(n6796), .B(n9684), .ZN(n6744)
         );
  AND2_X1 U8399 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6742) );
  AOI21_X1 U8400 ( .B1(n9673), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n6742), .ZN(
        n6743) );
  OAI211_X1 U8401 ( .C1(n9212), .C2(n6797), .A(n6744), .B(n6743), .ZN(n6745)
         );
  OR2_X1 U8402 ( .A1(n6746), .A2(n6745), .ZN(P1_U3253) );
  INV_X1 U8403 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6748) );
  INV_X1 U8404 ( .A(n6747), .ZN(n6749) );
  INV_X1 U8405 ( .A(n8246), .ZN(n8267) );
  OAI222_X1 U8406 ( .A1(n8679), .A2(n6748), .B1(n7962), .B2(n6749), .C1(
        P2_U3151), .C2(n8267), .ZN(P2_U3280) );
  INV_X1 U8407 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6750) );
  INV_X1 U8408 ( .A(n9156), .ZN(n9148) );
  OAI222_X1 U8409 ( .A1(n9616), .A2(n6750), .B1(n7925), .B2(n6749), .C1(
        P1_U3086), .C2(n9148), .ZN(P1_U3340) );
  AND3_X1 U8410 ( .A1(n6752), .A2(n6922), .A3(n6751), .ZN(n6808) );
  NOR2_X1 U8411 ( .A1(n6753), .A2(P1_U3086), .ZN(n6925) );
  AND3_X2 U8412 ( .A1(n6808), .A2(n6807), .A3(n6925), .ZN(n9814) );
  MUX2_X1 U8413 ( .A(n6754), .B(n9125), .S(n9121), .Z(n6755) );
  NAND2_X1 U8414 ( .A1(n6755), .A2(n6934), .ZN(n7599) );
  OR2_X1 U8415 ( .A1(n6500), .A2(n4550), .ZN(n9546) );
  INV_X1 U8416 ( .A(n7279), .ZN(n9056) );
  NAND2_X1 U8417 ( .A1(n4420), .A2(n9056), .ZN(n8977) );
  NAND2_X1 U8418 ( .A1(n4539), .A2(n4550), .ZN(n6756) );
  NAND2_X1 U8419 ( .A1(n8977), .A2(n6756), .ZN(n9715) );
  AND2_X1 U8420 ( .A1(n9739), .A2(n6974), .ZN(n9059) );
  NOR2_X1 U8421 ( .A1(n9729), .A2(n9059), .ZN(n9018) );
  INV_X1 U8422 ( .A(n9018), .ZN(n6757) );
  OAI21_X1 U8423 ( .B1(n9802), .B2(n9715), .A(n6757), .ZN(n6758) );
  NAND2_X1 U8424 ( .A1(n6964), .A2(n9460), .ZN(n6928) );
  OAI211_X1 U8425 ( .C1(n6934), .C2(n9739), .A(n6758), .B(n6928), .ZN(n6809)
         );
  NAND2_X1 U8426 ( .A1(n6809), .A2(n9814), .ZN(n6759) );
  OAI21_X1 U8427 ( .B1(n9814), .B2(n6013), .A(n6759), .ZN(P1_U3522) );
  AND2_X1 U8428 ( .A1(n6731), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8429 ( .A1(n6731), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8430 ( .A1(n6731), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8431 ( .A1(n6731), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8432 ( .A1(n6731), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8433 ( .A1(n6731), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8434 ( .A1(n6731), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8435 ( .A1(n6731), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8436 ( .A1(n6731), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8437 ( .A1(n6731), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8438 ( .A1(n6731), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8439 ( .A1(n6731), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8440 ( .A1(n6731), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8441 ( .A1(n6731), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8442 ( .A1(n6731), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8443 ( .A1(n6731), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8444 ( .A1(n6731), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  INV_X1 U8445 ( .A(n6761), .ZN(n6762) );
  AOI22_X1 U8446 ( .A1(n6731), .A2(n5009), .B1(n6762), .B2(n6834), .ZN(
        P2_U3376) );
  INV_X1 U8447 ( .A(n6763), .ZN(n6764) );
  INV_X1 U8448 ( .A(n9170), .ZN(n9177) );
  OAI222_X1 U8449 ( .A1(n9616), .A2(n10042), .B1(n7925), .B2(n6764), .C1(n9177), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U8450 ( .A(n8266), .ZN(n8285) );
  OAI222_X1 U8451 ( .A1(n8679), .A2(n6765), .B1(n7962), .B2(n6764), .C1(n8285), 
        .C2(P2_U3151), .ZN(P2_U3279) );
  AOI21_X1 U8452 ( .B1(n6768), .B2(n6767), .A(n6766), .ZN(n6772) );
  AOI22_X1 U8453 ( .A1(n9146), .A2(n9460), .B1(n9461), .B2(n6974), .ZN(n9731)
         );
  INV_X1 U8454 ( .A(n8829), .ZN(n8797) );
  OAI22_X1 U8455 ( .A1(n9731), .A2(n8797), .B1(n8853), .B2(n9749), .ZN(n6769)
         );
  AOI21_X1 U8456 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6770), .A(n6769), .ZN(
        n6771) );
  OAI21_X1 U8457 ( .B1(n6772), .B2(n8866), .A(n6771), .ZN(P1_U3222) );
  XOR2_X1 U8458 ( .A(n6774), .B(n6773), .Z(n6782) );
  NAND2_X1 U8459 ( .A1(n9673), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n6775) );
  NAND2_X1 U8460 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n6942) );
  OAI211_X1 U8461 ( .C1(n9212), .C2(n6776), .A(n6775), .B(n6942), .ZN(n6781)
         );
  AOI211_X1 U8462 ( .C1(n6779), .C2(n6778), .A(n6777), .B(n9660), .ZN(n6780)
         );
  AOI211_X1 U8463 ( .C1(n9684), .C2(n6782), .A(n6781), .B(n6780), .ZN(n6790)
         );
  INV_X1 U8464 ( .A(n9663), .ZN(n6783) );
  MUX2_X1 U8465 ( .A(n6784), .B(n6783), .S(n7919), .Z(n6786) );
  NAND2_X1 U8466 ( .A1(n6786), .A2(n6785), .ZN(n6789) );
  NOR2_X1 U8467 ( .A1(n9651), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6787) );
  OR2_X1 U8468 ( .A1(n6525), .A2(n6787), .ZN(n9650) );
  NAND2_X1 U8469 ( .A1(n9650), .A2(n9666), .ZN(n9655) );
  AND2_X1 U8470 ( .A1(n9655), .A2(P1_U3973), .ZN(n6788) );
  NAND2_X1 U8471 ( .A1(n6789), .A2(n6788), .ZN(n9674) );
  NAND2_X1 U8472 ( .A1(n6790), .A2(n9674), .ZN(P1_U3247) );
  NAND2_X1 U8473 ( .A1(n6853), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6793) );
  OAI21_X1 U8474 ( .B1(n6853), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6793), .ZN(
        n6794) );
  AOI211_X1 U8475 ( .C1(n6795), .C2(n6794), .A(n6852), .B(n9660), .ZN(n6806)
         );
  OAI21_X1 U8476 ( .B1(n6797), .B2(n6739), .A(n6796), .ZN(n6800) );
  MUX2_X1 U8477 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6798), .S(n6853), .Z(n6799)
         );
  NAND2_X1 U8478 ( .A1(n6799), .A2(n6800), .ZN(n6847) );
  OAI211_X1 U8479 ( .C1(n6800), .C2(n6799), .A(n9684), .B(n6847), .ZN(n6804)
         );
  NOR2_X1 U8480 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6801), .ZN(n6802) );
  AOI21_X1 U8481 ( .B1(n9673), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n6802), .ZN(
        n6803) );
  OAI211_X1 U8482 ( .C1(n9212), .C2(n6848), .A(n6804), .B(n6803), .ZN(n6805)
         );
  OR2_X1 U8483 ( .A1(n6806), .A2(n6805), .ZN(P1_U3254) );
  INV_X1 U8484 ( .A(n6807), .ZN(n6923) );
  INV_X1 U8485 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6811) );
  NAND2_X1 U8486 ( .A1(n6809), .A2(n9788), .ZN(n6810) );
  OAI21_X1 U8487 ( .B1(n9788), .B2(n6811), .A(n6810), .ZN(P1_U3453) );
  AND2_X1 U8488 ( .A1(n6813), .A2(n6841), .ZN(n6887) );
  INV_X1 U8489 ( .A(n6887), .ZN(n6812) );
  NAND2_X1 U8490 ( .A1(n6813), .A2(n6827), .ZN(n6817) );
  INV_X1 U8491 ( .A(n6814), .ZN(n6815) );
  NAND2_X1 U8492 ( .A1(n6818), .A2(n6815), .ZN(n6816) );
  INV_X1 U8493 ( .A(n6842), .ZN(n6914) );
  NAND2_X1 U8494 ( .A1(n6818), .A2(n9927), .ZN(n6819) );
  AOI22_X1 U8495 ( .A1(n8170), .A2(n6914), .B1(n6840), .B2(n8177), .ZN(n6836)
         );
  OAI21_X1 U8496 ( .B1(n6822), .B2(n6821), .A(n6820), .ZN(n6825) );
  NAND3_X1 U8497 ( .A1(n6825), .A2(n6824), .A3(n6823), .ZN(n6826) );
  NAND2_X1 U8498 ( .A1(n6826), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6833) );
  NAND2_X1 U8499 ( .A1(n6827), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6828) );
  AND2_X1 U8500 ( .A1(n6829), .A2(n6828), .ZN(n6830) );
  OR2_X1 U8501 ( .A1(n6831), .A2(n6830), .ZN(n6832) );
  NAND2_X1 U8502 ( .A1(n7065), .A2(n6834), .ZN(n6911) );
  NAND2_X1 U8503 ( .A1(n6911), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6835) );
  OAI211_X1 U8504 ( .C1(n4640), .C2(n8175), .A(n6836), .B(n6835), .ZN(P2_U3172) );
  INV_X1 U8505 ( .A(n6837), .ZN(n6839) );
  INV_X1 U8506 ( .A(n8307), .ZN(n8284) );
  OAI222_X1 U8507 ( .A1(n8679), .A2(n6838), .B1(n7962), .B2(n6839), .C1(
        P2_U3151), .C2(n8284), .ZN(P2_U3278) );
  INV_X1 U8508 ( .A(n9188), .ZN(n9193) );
  OAI222_X1 U8509 ( .A1(n9616), .A2(n10187), .B1(n7925), .B2(n6839), .C1(
        P1_U3086), .C2(n9193), .ZN(P1_U3338) );
  AOI22_X1 U8510 ( .A1(n8524), .A2(n6840), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8466), .ZN(n6846) );
  NOR3_X1 U8511 ( .A1(n6842), .A2(n6841), .A3(n9927), .ZN(n6844) );
  NAND2_X1 U8512 ( .A1(n5860), .A2(n8499), .ZN(n6915) );
  INV_X1 U8513 ( .A(n6915), .ZN(n6843) );
  OAI21_X1 U8514 ( .B1(n6844), .B2(n6843), .A(n9872), .ZN(n6845) );
  OAI211_X1 U8515 ( .C1(n7141), .C2(n9872), .A(n6846), .B(n6845), .ZN(P2_U3233) );
  OAI21_X1 U8516 ( .B1(n6798), .B2(n6848), .A(n6847), .ZN(n6850) );
  AOI22_X1 U8517 ( .A1(n6952), .A2(n6222), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n6851), .ZN(n6849) );
  NOR2_X1 U8518 ( .A1(n6850), .A2(n6849), .ZN(n6954) );
  AOI21_X1 U8519 ( .B1(n6850), .B2(n6849), .A(n6954), .ZN(n6861) );
  AOI22_X1 U8520 ( .A1(n6952), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n6227), .B2(
        n6851), .ZN(n6855) );
  OAI21_X1 U8521 ( .B1(n6855), .B2(n6854), .A(n6949), .ZN(n6856) );
  NAND2_X1 U8522 ( .A1(n6856), .A2(n9682), .ZN(n6860) );
  INV_X1 U8523 ( .A(n9212), .ZN(n9677) );
  INV_X1 U8524 ( .A(n9673), .ZN(n9222) );
  INV_X1 U8525 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6857) );
  NAND2_X1 U8526 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8735) );
  OAI21_X1 U8527 ( .B1(n9222), .B2(n6857), .A(n8735), .ZN(n6858) );
  AOI21_X1 U8528 ( .B1(n6952), .B2(n9677), .A(n6858), .ZN(n6859) );
  OAI211_X1 U8529 ( .C1(n6861), .C2(n9213), .A(n6860), .B(n6859), .ZN(P1_U3255) );
  XNOR2_X1 U8530 ( .A(n6862), .B(n6863), .ZN(n6864) );
  INV_X1 U8531 ( .A(n8866), .ZN(n8817) );
  NAND2_X1 U8532 ( .A1(n6864), .A2(n8817), .ZN(n6866) );
  INV_X1 U8533 ( .A(n9461), .ZN(n9393) );
  OAI22_X1 U8534 ( .A1(n6975), .A2(n9393), .B1(n6997), .B2(n9439), .ZN(n9714)
         );
  AOI22_X1 U8535 ( .A1(n8864), .A2(n6982), .B1(n8829), .B2(n9714), .ZN(n6865)
         );
  OAI211_X1 U8536 ( .C1(n6868), .C2(n6867), .A(n6866), .B(n6865), .ZN(P1_U3237) );
  INV_X1 U8537 ( .A(n6869), .ZN(n6902) );
  AOI22_X1 U8538 ( .A1(n9210), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n6870), .ZN(n6871) );
  OAI21_X1 U8539 ( .B1(n6902), .B2(n7925), .A(n6871), .ZN(P1_U3337) );
  NAND2_X1 U8540 ( .A1(n6874), .A2(n6873), .ZN(n6877) );
  NAND2_X1 U8541 ( .A1(n6875), .A2(n7334), .ZN(n6876) );
  NAND2_X2 U8542 ( .A1(n6877), .A2(n6876), .ZN(n6880) );
  NAND2_X1 U8543 ( .A1(n6881), .A2(n4640), .ZN(n6903) );
  INV_X1 U8544 ( .A(n6881), .ZN(n6882) );
  NAND2_X1 U8545 ( .A1(n6882), .A2(n5860), .ZN(n6883) );
  NAND2_X1 U8546 ( .A1(n6903), .A2(n6883), .ZN(n6884) );
  NOR2_X2 U8547 ( .A1(n6884), .A2(n6885), .ZN(n6905) );
  AOI21_X1 U8548 ( .B1(n6885), .B2(n6884), .A(n6905), .ZN(n6892) );
  INV_X1 U8549 ( .A(n8204), .ZN(n6889) );
  AOI22_X1 U8550 ( .A1(n8172), .A2(n7012), .B1(n6879), .B2(n8177), .ZN(n6888)
         );
  OAI21_X1 U8551 ( .B1(n6889), .B2(n8175), .A(n6888), .ZN(n6890) );
  AOI21_X1 U8552 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n6911), .A(n6890), .ZN(
        n6891) );
  OAI21_X1 U8553 ( .B1(n8119), .B2(n6892), .A(n6891), .ZN(P2_U3162) );
  XOR2_X1 U8554 ( .A(n6894), .B(n6893), .Z(n6900) );
  OR2_X1 U8555 ( .A1(n6979), .A2(n9393), .ZN(n6896) );
  NAND2_X1 U8556 ( .A1(n9144), .A2(n9460), .ZN(n6895) );
  NAND2_X1 U8557 ( .A1(n6896), .A2(n6895), .ZN(n6970) );
  MUX2_X1 U8558 ( .A(n8847), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n6898) );
  NOR2_X1 U8559 ( .A1(n8853), .A2(n9800), .ZN(n6897) );
  AOI211_X1 U8560 ( .C1(n8829), .C2(n6970), .A(n6898), .B(n6897), .ZN(n6899)
         );
  OAI21_X1 U8561 ( .B1(n6900), .B2(n8866), .A(n6899), .ZN(P1_U3218) );
  INV_X1 U8562 ( .A(n8328), .ZN(n8303) );
  OAI222_X1 U8563 ( .A1(P2_U3151), .A2(n8303), .B1(n7962), .B2(n6902), .C1(
        n6901), .C2(n8679), .ZN(P2_U3277) );
  INV_X1 U8564 ( .A(n6903), .ZN(n6904) );
  XNOR2_X1 U8565 ( .A(n6880), .B(n6908), .ZN(n7066) );
  XNOR2_X1 U8566 ( .A(n7066), .B(n8204), .ZN(n6906) );
  AOI21_X1 U8567 ( .B1(n6907), .B2(n6906), .A(n8009), .ZN(n6913) );
  AOI22_X1 U8568 ( .A1(n8172), .A2(n5860), .B1(n6908), .B2(n8177), .ZN(n6909)
         );
  OAI21_X1 U8569 ( .B1(n9864), .B2(n8175), .A(n6909), .ZN(n6910) );
  AOI21_X1 U8570 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n6911), .A(n6910), .ZN(
        n6912) );
  OAI21_X1 U8571 ( .B1(n6913), .B2(n8119), .A(n6912), .ZN(P2_U3177) );
  INV_X1 U8572 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6919) );
  OAI21_X1 U8573 ( .B1(n8494), .B2(n9920), .A(n6914), .ZN(n6916) );
  OAI211_X1 U8574 ( .C1(n6917), .C2(n9915), .A(n6916), .B(n6915), .ZN(n8618)
         );
  NAND2_X1 U8575 ( .A1(n9928), .A2(n8618), .ZN(n6918) );
  OAI21_X1 U8576 ( .B1(n9928), .B2(n6919), .A(n6918), .ZN(P2_U3390) );
  INV_X1 U8577 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6921) );
  NAND2_X1 U8578 ( .A1(P2_U3893), .A2(n7012), .ZN(n6920) );
  OAI21_X1 U8579 ( .B1(P2_U3893), .B2(n6921), .A(n6920), .ZN(P2_U3491) );
  NAND4_X1 U8580 ( .A1(n6925), .A2(n6924), .A3(n6923), .A4(n6922), .ZN(n6926)
         );
  NOR2_X1 U8581 ( .A1(n9018), .A2(n6927), .ZN(n6930) );
  INV_X1 U8582 ( .A(n6930), .ZN(n6932) );
  OAI21_X1 U8583 ( .B1(n6009), .B2(n9701), .A(n6928), .ZN(n6929) );
  AOI21_X1 U8584 ( .B1(n6930), .B2(n9125), .A(n6929), .ZN(n6931) );
  OAI21_X1 U8585 ( .B1(n9121), .B2(n6932), .A(n6931), .ZN(n6933) );
  NAND2_X1 U8586 ( .A1(n6933), .A2(n9471), .ZN(n6937) );
  NOR2_X1 U8587 ( .A1(n9740), .A2(n9549), .ZN(n9348) );
  INV_X1 U8588 ( .A(n9741), .ZN(n9706) );
  OAI21_X1 U8589 ( .B1(n9348), .B2(n9706), .A(n6973), .ZN(n6936) );
  OAI211_X1 U8590 ( .C1(n9471), .C2(n6938), .A(n6937), .B(n6936), .ZN(P1_U3293) );
  OAI211_X1 U8591 ( .C1(n6941), .C2(n6940), .A(n6939), .B(n8817), .ZN(n6946)
         );
  INV_X1 U8592 ( .A(n6997), .ZN(n9145) );
  OAI21_X1 U8593 ( .B1(n8858), .B2(n7001), .A(n6942), .ZN(n6944) );
  INV_X1 U8594 ( .A(n8850), .ZN(n8859) );
  INV_X1 U8595 ( .A(n7004), .ZN(n9762) );
  OAI22_X1 U8596 ( .A1(n8859), .A2(n7229), .B1(n9762), .B2(n8853), .ZN(n6943)
         );
  AOI211_X1 U8597 ( .C1(n8813), .C2(n9145), .A(n6944), .B(n6943), .ZN(n6945)
         );
  NAND2_X1 U8598 ( .A1(n6946), .A2(n6945), .ZN(P1_U3230) );
  NAND2_X1 U8599 ( .A1(n8187), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6947) );
  OAI21_X1 U8600 ( .B1(n7871), .B2(n8187), .A(n6947), .ZN(P2_U3520) );
  NAND2_X1 U8601 ( .A1(n7385), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6948) );
  OAI21_X1 U8602 ( .B1(n7385), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6948), .ZN(
        n6951) );
  OAI21_X1 U8603 ( .B1(n6952), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6949), .ZN(
        n6950) );
  NOR2_X1 U8604 ( .A1(n6951), .A2(n6950), .ZN(n7379) );
  AOI211_X1 U8605 ( .C1(n6951), .C2(n6950), .A(n7379), .B(n9660), .ZN(n6963)
         );
  NOR2_X1 U8606 ( .A1(n6952), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6953) );
  NOR2_X1 U8607 ( .A1(n6954), .A2(n6953), .ZN(n6957) );
  MUX2_X1 U8608 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6955), .S(n7385), .Z(n6956)
         );
  NAND2_X1 U8609 ( .A1(n6956), .A2(n6957), .ZN(n7387) );
  OAI211_X1 U8610 ( .C1(n6957), .C2(n6956), .A(n7387), .B(n9684), .ZN(n6960)
         );
  NOR2_X1 U8611 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8803), .ZN(n6958) );
  AOI21_X1 U8612 ( .B1(n9673), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n6958), .ZN(
        n6959) );
  OAI211_X1 U8613 ( .C1(n9212), .C2(n6961), .A(n6960), .B(n6959), .ZN(n6962)
         );
  OR2_X1 U8614 ( .A1(n6963), .A2(n6962), .ZN(P1_U3256) );
  NAND2_X1 U8615 ( .A1(n9016), .A2(n9729), .ZN(n6967) );
  NAND2_X1 U8616 ( .A1(n6975), .A2(n6965), .ZN(n6966) );
  NAND2_X1 U8617 ( .A1(n6967), .A2(n6966), .ZN(n9713) );
  NAND2_X1 U8618 ( .A1(n6979), .A2(n6982), .ZN(n6978) );
  INV_X1 U8619 ( .A(n6978), .ZN(n6968) );
  NAND2_X1 U8620 ( .A1(n6997), .A2(n6987), .ZN(n6991) );
  NAND2_X1 U8621 ( .A1(n6991), .A2(n9064), .ZN(n9015) );
  XNOR2_X1 U8622 ( .A(n6993), .B(n9015), .ZN(n6971) );
  AOI21_X1 U8623 ( .B1(n6971), .B2(n9715), .A(n6970), .ZN(n9804) );
  AND2_X1 U8624 ( .A1(n7599), .A2(n7494), .ZN(n6972) );
  INV_X1 U8625 ( .A(n9433), .ZN(n9725) );
  NAND2_X1 U8626 ( .A1(n6974), .A2(n6973), .ZN(n9728) );
  NAND2_X1 U8627 ( .A1(n6975), .A2(n9749), .ZN(n6976) );
  NAND2_X1 U8628 ( .A1(n6977), .A2(n6976), .ZN(n9719) );
  NAND2_X1 U8629 ( .A1(n9719), .A2(n9720), .ZN(n6981) );
  NAND2_X1 U8630 ( .A1(n6979), .A2(n9756), .ZN(n6980) );
  XNOR2_X1 U8631 ( .A(n6996), .B(n9015), .ZN(n9803) );
  NAND2_X1 U8632 ( .A1(n9749), .A2(n9739), .ZN(n9737) );
  OR2_X1 U8633 ( .A1(n9737), .A2(n6982), .ZN(n9721) );
  NAND2_X1 U8634 ( .A1(n9721), .A2(n6987), .ZN(n6983) );
  NAND2_X1 U8635 ( .A1(n6983), .A2(n9738), .ZN(n6984) );
  OR2_X1 U8636 ( .A1(n6984), .A2(n7000), .ZN(n9798) );
  OAI22_X1 U8637 ( .A1(n9471), .A2(n6985), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9701), .ZN(n6986) );
  AOI21_X1 U8638 ( .B1(n9706), .B2(n6987), .A(n6986), .ZN(n6988) );
  OAI21_X1 U8639 ( .B1(n9740), .B2(n9798), .A(n6988), .ZN(n6989) );
  AOI21_X1 U8640 ( .B1(n9725), .B2(n9803), .A(n6989), .ZN(n6990) );
  OAI21_X1 U8641 ( .B1(n9804), .B2(n4419), .A(n6990), .ZN(P1_U3290) );
  INV_X1 U8642 ( .A(n9064), .ZN(n6992) );
  NAND2_X1 U8643 ( .A1(n9144), .A2(n7004), .ZN(n7040) );
  INV_X1 U8644 ( .A(n7040), .ZN(n6994) );
  NOR2_X1 U8645 ( .A1(n9144), .A2(n7004), .ZN(n7039) );
  OR2_X1 U8646 ( .A1(n6994), .A2(n7039), .ZN(n6999) );
  XNOR2_X1 U8647 ( .A(n7042), .B(n6999), .ZN(n6995) );
  INV_X1 U8648 ( .A(n7229), .ZN(n9143) );
  AOI222_X1 U8649 ( .A1(n9715), .A2(n6995), .B1(n9143), .B2(n9460), .C1(n9145), 
        .C2(n9461), .ZN(n9763) );
  NAND2_X1 U8650 ( .A1(n6997), .A2(n9800), .ZN(n6998) );
  INV_X1 U8651 ( .A(n6999), .ZN(n9020) );
  XNOR2_X1 U8652 ( .A(n7038), .B(n9020), .ZN(n9766) );
  OAI211_X1 U8653 ( .C1(n7000), .C2(n9762), .A(n7045), .B(n9738), .ZN(n9761)
         );
  OAI22_X1 U8654 ( .A1(n9471), .A2(n7002), .B1(n7001), .B2(n9701), .ZN(n7003)
         );
  AOI21_X1 U8655 ( .B1(n9706), .B2(n7004), .A(n7003), .ZN(n7005) );
  OAI21_X1 U8656 ( .B1(n9761), .B2(n9740), .A(n7005), .ZN(n7006) );
  AOI21_X1 U8657 ( .B1(n9766), .B2(n9725), .A(n7006), .ZN(n7007) );
  OAI21_X1 U8658 ( .B1(n9763), .B2(n4419), .A(n7007), .ZN(P1_U3289) );
  NAND2_X1 U8659 ( .A1(n5859), .A2(n5656), .ZN(n7008) );
  NAND2_X1 U8660 ( .A1(n7009), .A2(n7008), .ZN(n9879) );
  XNOR2_X1 U8661 ( .A(n5859), .B(n7010), .ZN(n7011) );
  NAND2_X1 U8662 ( .A1(n7011), .A2(n8494), .ZN(n7014) );
  AOI22_X1 U8663 ( .A1(n8500), .A2(n7012), .B1(n8204), .B2(n8499), .ZN(n7013)
         );
  NAND2_X1 U8664 ( .A1(n7014), .A2(n7013), .ZN(n9878) );
  MUX2_X1 U8665 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n9878), .S(n9872), .Z(n7017)
         );
  OAI22_X1 U8666 ( .A1(n8534), .A2(n9876), .B1(n7015), .B2(n9860), .ZN(n7016)
         );
  AOI211_X1 U8667 ( .C1(n8539), .C2(n9879), .A(n7017), .B(n7016), .ZN(n7018)
         );
  INV_X1 U8668 ( .A(n7018), .ZN(P2_U3232) );
  XNOR2_X1 U8669 ( .A(n7053), .B(n7023), .ZN(n7019) );
  NAND2_X1 U8670 ( .A1(n7019), .A2(n8494), .ZN(n7021) );
  AOI22_X1 U8671 ( .A1(n8500), .A2(n8203), .B1(n8201), .B2(n8499), .ZN(n7020)
         );
  NAND2_X1 U8672 ( .A1(n7021), .A2(n7020), .ZN(n9893) );
  INV_X1 U8673 ( .A(n9893), .ZN(n7032) );
  INV_X1 U8674 ( .A(n7023), .ZN(n7025) );
  NAND3_X1 U8675 ( .A1(n7022), .A2(n7025), .A3(n7024), .ZN(n7026) );
  NAND2_X1 U8676 ( .A1(n7027), .A2(n7026), .ZN(n9895) );
  INV_X1 U8677 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7028) );
  NOR2_X1 U8678 ( .A1(n9872), .A2(n7028), .ZN(n7030) );
  OAI22_X1 U8679 ( .A1(n8534), .A2(n9892), .B1(n7079), .B2(n9860), .ZN(n7029)
         );
  AOI211_X1 U8680 ( .C1(n8539), .C2(n9895), .A(n7030), .B(n7029), .ZN(n7031)
         );
  OAI21_X1 U8681 ( .B1(n9874), .B2(n7032), .A(n7031), .ZN(P2_U3229) );
  INV_X1 U8682 ( .A(n7033), .ZN(n7036) );
  OAI222_X1 U8683 ( .A1(n8679), .A2(n7034), .B1(n7962), .B2(n7036), .C1(
        P2_U3151), .C2(n8333), .ZN(P2_U3276) );
  OAI222_X1 U8684 ( .A1(n9616), .A2(n7037), .B1(n7925), .B2(n7036), .C1(
        P1_U3086), .C2(n7035), .ZN(P1_U3336) );
  NAND2_X1 U8685 ( .A1(n7041), .A2(n7040), .ZN(n7224) );
  NAND2_X1 U8686 ( .A1(n7229), .A2(n7049), .ZN(n8888) );
  NAND2_X1 U8687 ( .A1(n7322), .A2(n9143), .ZN(n8887) );
  INV_X1 U8688 ( .A(n7226), .ZN(n9021) );
  XNOR2_X1 U8689 ( .A(n7224), .B(n9021), .ZN(n7318) );
  NAND2_X1 U8690 ( .A1(n9762), .A2(n9144), .ZN(n9063) );
  XNOR2_X1 U8691 ( .A(n8889), .B(n9021), .ZN(n7043) );
  INV_X1 U8692 ( .A(n7534), .ZN(n9142) );
  AOI222_X1 U8693 ( .A1(n9715), .A2(n7043), .B1(n9142), .B2(n9460), .C1(n9144), 
        .C2(n9461), .ZN(n7317) );
  OR2_X1 U8694 ( .A1(n7317), .A2(n4419), .ZN(n7051) );
  OAI22_X1 U8695 ( .A1(n9471), .A2(n7044), .B1(n7311), .B2(n9701), .ZN(n7048)
         );
  INV_X1 U8696 ( .A(n7045), .ZN(n7046) );
  OAI211_X1 U8697 ( .C1(n7046), .C2(n7322), .A(n9738), .B(n7232), .ZN(n7316)
         );
  NOR2_X1 U8698 ( .A1(n7316), .A2(n9740), .ZN(n7047) );
  AOI211_X1 U8699 ( .C1(n9706), .C2(n7049), .A(n7048), .B(n7047), .ZN(n7050)
         );
  OAI211_X1 U8700 ( .C1(n7318), .C2(n9433), .A(n7051), .B(n7050), .ZN(P1_U3288) );
  INV_X1 U8701 ( .A(n8200), .ZN(n7578) );
  INV_X1 U8702 ( .A(n8202), .ZN(n7058) );
  NAND2_X1 U8703 ( .A1(n7053), .A2(n7052), .ZN(n7055) );
  NAND2_X1 U8704 ( .A1(n7055), .A2(n7054), .ZN(n7056) );
  XOR2_X1 U8705 ( .A(n7059), .B(n7056), .Z(n7057) );
  OAI222_X1 U8706 ( .A1(n9863), .A2(n7578), .B1(n9865), .B2(n7058), .C1(n7057), 
        .C2(n9869), .ZN(n7216) );
  INV_X1 U8707 ( .A(n7216), .ZN(n7064) );
  XNOR2_X1 U8708 ( .A(n7060), .B(n7059), .ZN(n7217) );
  NOR2_X1 U8709 ( .A1(n9872), .A2(n7137), .ZN(n7062) );
  OAI22_X1 U8710 ( .A1(n8534), .A2(n7335), .B1(n7349), .B2(n9860), .ZN(n7061)
         );
  AOI211_X1 U8711 ( .C1(n7217), .C2(n8539), .A(n7062), .B(n7061), .ZN(n7063)
         );
  OAI21_X1 U8712 ( .B1(n7064), .B2(n9874), .A(n7063), .ZN(P2_U3228) );
  INV_X2 U8713 ( .A(n7069), .ZN(n7847) );
  XNOR2_X1 U8714 ( .A(n7847), .B(n9888), .ZN(n7067) );
  INV_X1 U8715 ( .A(n7067), .ZN(n7068) );
  NOR2_X1 U8716 ( .A1(n7066), .A2(n8204), .ZN(n8008) );
  XNOR2_X1 U8717 ( .A(n7067), .B(n9864), .ZN(n8007) );
  XNOR2_X1 U8718 ( .A(n7847), .B(n7070), .ZN(n7071) );
  NOR2_X1 U8719 ( .A1(n7071), .A2(n8202), .ZN(n7336) );
  AOI21_X1 U8720 ( .B1(n8202), .B2(n7071), .A(n7336), .ZN(n7072) );
  OAI21_X1 U8721 ( .B1(n7073), .B2(n7072), .A(n7338), .ZN(n7074) );
  NAND2_X1 U8722 ( .A1(n7074), .A2(n8170), .ZN(n7078) );
  INV_X1 U8723 ( .A(n8177), .ZN(n8164) );
  NAND2_X1 U8724 ( .A1(n8172), .A2(n8203), .ZN(n7075) );
  NAND2_X1 U8725 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7188) );
  OAI211_X1 U8726 ( .C1(n9892), .C2(n8164), .A(n7075), .B(n7188), .ZN(n7076)
         );
  AOI21_X1 U8727 ( .B1(n8102), .B2(n8201), .A(n7076), .ZN(n7077) );
  OAI211_X1 U8728 ( .C1(n7079), .C2(n8150), .A(n7078), .B(n7077), .ZN(P2_U3170) );
  INV_X1 U8729 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8319) );
  NOR2_X1 U8730 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7120) );
  NOR2_X1 U8731 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7117) );
  NOR2_X1 U8732 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7113) );
  NOR2_X1 U8733 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7111) );
  NOR2_X1 U8734 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7109) );
  NOR2_X1 U8735 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7106) );
  NOR2_X1 U8736 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7104) );
  NOR2_X1 U8737 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7100) );
  NOR2_X1 U8738 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7097) );
  NOR2_X1 U8739 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7094) );
  NOR2_X1 U8740 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7092) );
  NOR2_X1 U8741 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7090) );
  NOR2_X1 U8742 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7088) );
  NOR2_X1 U8743 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7086) );
  NAND2_X1 U8744 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7084) );
  XOR2_X1 U8745 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10295) );
  NAND2_X1 U8746 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7082) );
  AOI21_X1 U8747 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9943) );
  INV_X1 U8748 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9946) );
  NOR2_X1 U8749 ( .A1(n9946), .A2(n10013), .ZN(n9945) );
  NOR2_X1 U8750 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n9942), .ZN(n7080) );
  NOR2_X1 U8751 ( .A1(n9943), .A2(n7080), .ZN(n10293) );
  XOR2_X1 U8752 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10292) );
  NAND2_X1 U8753 ( .A1(n10293), .A2(n10292), .ZN(n7081) );
  NAND2_X1 U8754 ( .A1(n7082), .A2(n7081), .ZN(n10294) );
  NAND2_X1 U8755 ( .A1(n10295), .A2(n10294), .ZN(n7083) );
  NAND2_X1 U8756 ( .A1(n7084), .A2(n7083), .ZN(n10297) );
  XNOR2_X1 U8757 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10296) );
  NOR2_X1 U8758 ( .A1(n10297), .A2(n10296), .ZN(n7085) );
  NOR2_X1 U8759 ( .A1(n7086), .A2(n7085), .ZN(n10283) );
  XNOR2_X1 U8760 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10282) );
  NOR2_X1 U8761 ( .A1(n10283), .A2(n10282), .ZN(n7087) );
  NOR2_X1 U8762 ( .A1(n7088), .A2(n7087), .ZN(n10291) );
  XNOR2_X1 U8763 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10290) );
  NOR2_X1 U8764 ( .A1(n10291), .A2(n10290), .ZN(n7089) );
  NOR2_X1 U8765 ( .A1(n7090), .A2(n7089), .ZN(n10287) );
  XNOR2_X1 U8766 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10286) );
  NOR2_X1 U8767 ( .A1(n10287), .A2(n10286), .ZN(n7091) );
  NOR2_X1 U8768 ( .A1(n7092), .A2(n7091), .ZN(n10289) );
  XNOR2_X1 U8769 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10288) );
  NOR2_X1 U8770 ( .A1(n10289), .A2(n10288), .ZN(n7093) );
  NOR2_X1 U8771 ( .A1(n7094), .A2(n7093), .ZN(n10285) );
  INV_X1 U8772 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7095) );
  INV_X1 U8773 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7378) );
  AOI22_X1 U8774 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7095), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n7378), .ZN(n10284) );
  NOR2_X1 U8775 ( .A1(n10285), .A2(n10284), .ZN(n7096) );
  NOR2_X1 U8776 ( .A1(n7097), .A2(n7096), .ZN(n9965) );
  INV_X1 U8777 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7098) );
  INV_X1 U8778 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10000) );
  AOI22_X1 U8779 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n7098), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n10000), .ZN(n9964) );
  NOR2_X1 U8780 ( .A1(n9965), .A2(n9964), .ZN(n7099) );
  NOR2_X1 U8781 ( .A1(n7100), .A2(n7099), .ZN(n9963) );
  INV_X1 U8782 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7102) );
  INV_X1 U8783 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7101) );
  AOI22_X1 U8784 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n7102), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n7101), .ZN(n9962) );
  NOR2_X1 U8785 ( .A1(n9963), .A2(n9962), .ZN(n7103) );
  NOR2_X1 U8786 ( .A1(n7104), .A2(n7103), .ZN(n9961) );
  INV_X1 U8787 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7723) );
  AOI22_X1 U8788 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n6857), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n7723), .ZN(n9960) );
  NOR2_X1 U8789 ( .A1(n9961), .A2(n9960), .ZN(n7105) );
  NOR2_X1 U8790 ( .A1(n7106), .A2(n7105), .ZN(n9959) );
  INV_X1 U8791 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10246) );
  INV_X1 U8792 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7107) );
  AOI22_X1 U8793 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n10246), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n7107), .ZN(n9958) );
  NOR2_X1 U8794 ( .A1(n9959), .A2(n9958), .ZN(n7108) );
  NOR2_X1 U8795 ( .A1(n7109), .A2(n7108), .ZN(n9957) );
  XNOR2_X1 U8796 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9956) );
  NOR2_X1 U8797 ( .A1(n9957), .A2(n9956), .ZN(n7110) );
  NOR2_X1 U8798 ( .A1(n7111), .A2(n7110), .ZN(n9955) );
  INV_X1 U8799 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10245) );
  INV_X1 U8800 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8241) );
  AOI22_X1 U8801 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n10245), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8241), .ZN(n9954) );
  NOR2_X1 U8802 ( .A1(n9955), .A2(n9954), .ZN(n7112) );
  NOR2_X1 U8803 ( .A1(n7113), .A2(n7112), .ZN(n9953) );
  INV_X1 U8804 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7115) );
  INV_X1 U8805 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7114) );
  AOI22_X1 U8806 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n7115), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n7114), .ZN(n9952) );
  NOR2_X1 U8807 ( .A1(n9953), .A2(n9952), .ZN(n7116) );
  NOR2_X1 U8808 ( .A1(n7117), .A2(n7116), .ZN(n9951) );
  INV_X1 U8809 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7118) );
  INV_X1 U8810 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10027) );
  AOI22_X1 U8811 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n7118), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n10027), .ZN(n9950) );
  NOR2_X1 U8812 ( .A1(n9951), .A2(n9950), .ZN(n7119) );
  NOR2_X1 U8813 ( .A1(n7120), .A2(n7119), .ZN(n9948) );
  NOR2_X1 U8814 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9948), .ZN(n7121) );
  NAND2_X1 U8815 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9948), .ZN(n9947) );
  OAI21_X1 U8816 ( .B1(n8319), .B2(n7121), .A(n9947), .ZN(n7123) );
  XNOR2_X1 U8817 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7122) );
  XNOR2_X1 U8818 ( .A(n7123), .B(n7122), .ZN(ADD_1068_U4) );
  INV_X1 U8819 ( .A(n7124), .ZN(n7154) );
  INV_X1 U8820 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7174) );
  INV_X1 U8821 ( .A(n7189), .ZN(n7134) );
  MUX2_X1 U8822 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8334), .Z(n7132) );
  INV_X1 U8823 ( .A(n7132), .ZN(n7133) );
  MUX2_X1 U8824 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8334), .Z(n7130) );
  INV_X1 U8825 ( .A(n7130), .ZN(n7131) );
  INV_X1 U8826 ( .A(n4417), .ZN(n7129) );
  MUX2_X1 U8827 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8334), .Z(n7127) );
  INV_X1 U8828 ( .A(n7127), .ZN(n7128) );
  MUX2_X1 U8829 ( .A(n9817), .B(n7125), .S(n7140), .Z(n7126) );
  MUX2_X1 U8830 ( .A(n7141), .B(n7159), .S(n7140), .Z(n7326) );
  NAND2_X1 U8831 ( .A1(n7326), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9822) );
  NAND2_X1 U8832 ( .A1(n9823), .A2(n9822), .ZN(n9820) );
  OAI21_X1 U8833 ( .B1(n9818), .B2(n7126), .A(n9820), .ZN(n7211) );
  XOR2_X1 U8834 ( .A(n4417), .B(n7127), .Z(n7212) );
  NAND2_X1 U8835 ( .A1(n7211), .A2(n7212), .ZN(n7210) );
  OAI21_X1 U8836 ( .B1(n7129), .B2(n7128), .A(n7210), .ZN(n7282) );
  XNOR2_X1 U8837 ( .A(n7130), .B(n7287), .ZN(n7283) );
  NOR2_X1 U8838 ( .A1(n7282), .A2(n7283), .ZN(n7281) );
  AOI21_X1 U8839 ( .B1(n4861), .B2(n7131), .A(n7281), .ZN(n7177) );
  XOR2_X1 U8840 ( .A(n7189), .B(n7132), .Z(n7176) );
  NAND2_X1 U8841 ( .A1(n7177), .A2(n7176), .ZN(n7175) );
  OAI21_X1 U8842 ( .B1(n7134), .B2(n7133), .A(n7175), .ZN(n7139) );
  MUX2_X1 U8843 ( .A(n7137), .B(n7136), .S(n8334), .Z(n7240) );
  XNOR2_X1 U8844 ( .A(n7240), .B(n7165), .ZN(n7138) );
  NAND2_X1 U8845 ( .A1(n7139), .A2(n7138), .ZN(n7239) );
  OAI211_X1 U8846 ( .C1(n7139), .C2(n7138), .A(n7239), .B(n9821), .ZN(n7173)
         );
  NOR2_X1 U8847 ( .A1(n5855), .A2(P2_U3151), .ZN(n7153) );
  INV_X1 U8848 ( .A(n7153), .ZN(n8676) );
  NOR2_X1 U8849 ( .A1(n7152), .A2(n8676), .ZN(n7328) );
  NAND2_X1 U8850 ( .A1(n7328), .A2(n7135), .ZN(n9846) );
  INV_X1 U8851 ( .A(n9846), .ZN(n7294) );
  OAI21_X1 U8852 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7141), .A(n9818), .ZN(n7142) );
  INV_X1 U8853 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9817) );
  MUX2_X1 U8854 ( .A(n5263), .B(P2_REG2_REG_2__SCAN_IN), .S(n7202), .Z(n7204)
         );
  AOI21_X1 U8855 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n4417), .A(n7203), .ZN(
        n7144) );
  INV_X1 U8856 ( .A(n7146), .ZN(n7184) );
  MUX2_X1 U8857 ( .A(n7028), .B(P2_REG2_REG_4__SCAN_IN), .S(n7189), .Z(n7185)
         );
  AOI21_X1 U8858 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n7189), .A(n7183), .ZN(
        n7147) );
  INV_X1 U8859 ( .A(n7165), .ZN(n7241) );
  OAI21_X1 U8860 ( .B1(n7149), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7246), .ZN(
        n7171) );
  NOR2_X1 U8861 ( .A1(n8334), .A2(P2_U3151), .ZN(n7150) );
  NAND2_X1 U8862 ( .A1(n7150), .A2(n5855), .ZN(n7151) );
  OR2_X1 U8863 ( .A1(n7152), .A2(n7151), .ZN(n7156) );
  NAND2_X1 U8864 ( .A1(n7154), .A2(n7153), .ZN(n7155) );
  INV_X1 U8865 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10234) );
  NOR2_X1 U8866 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10234), .ZN(n7342) );
  INV_X1 U8867 ( .A(n7342), .ZN(n7157) );
  OAI21_X1 U8868 ( .B1(n9855), .B2(n7165), .A(n7157), .ZN(n7170) );
  NOR2_X1 U8869 ( .A1(n7159), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7160) );
  OR2_X1 U8870 ( .A1(n9829), .A2(n7125), .ZN(n9828) );
  NAND2_X1 U8871 ( .A1(n4417), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7162) );
  NAND2_X1 U8872 ( .A1(n7290), .A2(n7179), .ZN(n7163) );
  MUX2_X1 U8873 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n5294), .S(n7189), .Z(n7178)
         );
  NAND2_X1 U8874 ( .A1(n7163), .A2(n7178), .ZN(n7182) );
  NAND2_X1 U8875 ( .A1(n7189), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7164) );
  NAND2_X1 U8876 ( .A1(n7182), .A2(n7164), .ZN(n7166) );
  OAI21_X1 U8877 ( .B1(n7166), .B2(n7165), .A(n7251), .ZN(n7167) );
  NAND2_X1 U8878 ( .A1(n7167), .A2(n7136), .ZN(n7168) );
  NAND2_X1 U8879 ( .A1(n7328), .A2(n8334), .ZN(n9844) );
  AOI21_X1 U8880 ( .B1(n7253), .B2(n7168), .A(n9844), .ZN(n7169) );
  AOI211_X1 U8881 ( .C1(n7294), .C2(n7171), .A(n7170), .B(n7169), .ZN(n7172)
         );
  OAI211_X1 U8882 ( .C1(n8341), .C2(n7174), .A(n7173), .B(n7172), .ZN(P2_U3187) );
  INV_X1 U8883 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7195) );
  OAI211_X1 U8884 ( .C1(n7177), .C2(n7176), .A(n7175), .B(n9821), .ZN(n7194)
         );
  INV_X1 U8885 ( .A(n7178), .ZN(n7180) );
  NAND3_X1 U8886 ( .A1(n7290), .A2(n7180), .A3(n7179), .ZN(n7181) );
  AOI21_X1 U8887 ( .B1(n7182), .B2(n7181), .A(n9844), .ZN(n7192) );
  INV_X1 U8888 ( .A(n7183), .ZN(n7187) );
  NAND3_X1 U8889 ( .A1(n7284), .A2(n7185), .A3(n7184), .ZN(n7186) );
  AOI21_X1 U8890 ( .B1(n7187), .B2(n7186), .A(n9846), .ZN(n7191) );
  OAI21_X1 U8891 ( .B1(n9855), .B2(n7189), .A(n7188), .ZN(n7190) );
  NOR3_X1 U8892 ( .A1(n7192), .A2(n7191), .A3(n7190), .ZN(n7193) );
  OAI211_X1 U8893 ( .C1(n8341), .C2(n7195), .A(n7194), .B(n7193), .ZN(P2_U3186) );
  INV_X1 U8894 ( .A(n7196), .ZN(n7278) );
  OAI222_X1 U8895 ( .A1(n8679), .A2(n7198), .B1(n7962), .B2(n7278), .C1(n7197), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  INV_X1 U8896 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7215) );
  INV_X1 U8897 ( .A(n9844), .ZN(n9830) );
  OAI21_X1 U8898 ( .B1(n7201), .B2(n7200), .A(n7199), .ZN(n7209) );
  OAI22_X1 U8899 ( .A1(n9855), .A2(n4417), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9859), .ZN(n7208) );
  AOI21_X1 U8900 ( .B1(n7205), .B2(n7204), .A(n7203), .ZN(n7206) );
  NOR2_X1 U8901 ( .A1(n9846), .A2(n7206), .ZN(n7207) );
  AOI211_X1 U8902 ( .C1(n9830), .C2(n7209), .A(n7208), .B(n7207), .ZN(n7214)
         );
  OAI211_X1 U8903 ( .C1(n7212), .C2(n7211), .A(n9821), .B(n7210), .ZN(n7213)
         );
  OAI211_X1 U8904 ( .C1(n8341), .C2(n7215), .A(n7214), .B(n7213), .ZN(P2_U3184) );
  AOI21_X1 U8905 ( .B1(n7217), .B2(n9920), .A(n7216), .ZN(n7222) );
  INV_X1 U8906 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7218) );
  OAI22_X1 U8907 ( .A1(n7335), .A2(n8667), .B1(n9928), .B2(n7218), .ZN(n7219)
         );
  INV_X1 U8908 ( .A(n7219), .ZN(n7220) );
  OAI21_X1 U8909 ( .B1(n7222), .B2(n9929), .A(n7220), .ZN(P2_U3405) );
  AOI22_X1 U8910 ( .A1(n8607), .A2(n7343), .B1(n9939), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n7221) );
  OAI21_X1 U8911 ( .B1(n7222), .B2(n9939), .A(n7221), .ZN(P2_U3464) );
  NAND2_X1 U8912 ( .A1(n7229), .A2(n7322), .ZN(n7223) );
  NAND2_X1 U8913 ( .A1(n7534), .A2(n7480), .ZN(n9024) );
  NAND2_X1 U8914 ( .A1(n7488), .A2(n9142), .ZN(n8890) );
  NAND2_X1 U8915 ( .A1(n9024), .A2(n8890), .ZN(n7228) );
  NAND2_X1 U8916 ( .A1(n7225), .A2(n7228), .ZN(n7490) );
  OAI21_X1 U8917 ( .B1(n7225), .B2(n7228), .A(n7490), .ZN(n7424) );
  INV_X1 U8918 ( .A(n7424), .ZN(n7238) );
  NAND2_X1 U8919 ( .A1(n7227), .A2(n8887), .ZN(n7515) );
  XOR2_X1 U8920 ( .A(n7228), .B(n7515), .Z(n7231) );
  INV_X1 U8921 ( .A(n9715), .ZN(n9732) );
  OAI22_X1 U8922 ( .A1(n7229), .A2(n9393), .B1(n7491), .B2(n9439), .ZN(n7476)
         );
  INV_X1 U8923 ( .A(n7476), .ZN(n7230) );
  OAI21_X1 U8924 ( .B1(n7231), .B2(n9732), .A(n7230), .ZN(n7422) );
  NAND2_X1 U8925 ( .A1(n7422), .A2(n9471), .ZN(n7237) );
  AOI211_X1 U8926 ( .C1(n7480), .C2(n7232), .A(n9549), .B(n7606), .ZN(n7423)
         );
  NOR2_X1 U8927 ( .A1(n9741), .A2(n7488), .ZN(n7235) );
  OAI22_X1 U8928 ( .A1(n9471), .A2(n7233), .B1(n7478), .B2(n9701), .ZN(n7234)
         );
  AOI211_X1 U8929 ( .C1(n7423), .C2(n9724), .A(n7235), .B(n7234), .ZN(n7236)
         );
  OAI211_X1 U8930 ( .C1(n7238), .C2(n9433), .A(n7237), .B(n7236), .ZN(P1_U3287) );
  MUX2_X1 U8931 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8334), .Z(n7263) );
  XNOR2_X1 U8932 ( .A(n7263), .B(n7268), .ZN(n7243) );
  OAI21_X1 U8933 ( .B1(n7241), .B2(n7240), .A(n7239), .ZN(n7242) );
  NOR2_X1 U8934 ( .A1(n7242), .A2(n7243), .ZN(n7264) );
  AOI21_X1 U8935 ( .B1(n7243), .B2(n7242), .A(n7264), .ZN(n7262) );
  INV_X1 U8936 ( .A(n9821), .ZN(n9837) );
  INV_X1 U8937 ( .A(n8341), .ZN(n9850) );
  XNOR2_X1 U8938 ( .A(n7268), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7245) );
  NAND3_X1 U8939 ( .A1(n7246), .A2(n7245), .A3(n4423), .ZN(n7247) );
  AOI21_X1 U8940 ( .B1(n4502), .B2(n7247), .A(n9846), .ZN(n7256) );
  NAND2_X1 U8941 ( .A1(n7253), .A2(n7251), .ZN(n7249) );
  XNOR2_X1 U8942 ( .A(n7268), .B(n7248), .ZN(n7250) );
  NAND2_X1 U8943 ( .A1(n7249), .A2(n7250), .ZN(n7270) );
  INV_X1 U8944 ( .A(n7250), .ZN(n7252) );
  NAND3_X1 U8945 ( .A1(n7253), .A2(n7252), .A3(n7251), .ZN(n7254) );
  AOI21_X1 U8946 ( .B1(n7270), .B2(n7254), .A(n9844), .ZN(n7255) );
  NOR2_X1 U8947 ( .A1(n7256), .A2(n7255), .ZN(n7259) );
  INV_X1 U8948 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7257) );
  NOR2_X1 U8949 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7257), .ZN(n7403) );
  INV_X1 U8950 ( .A(n7403), .ZN(n7258) );
  OAI211_X1 U8951 ( .C1(n9855), .C2(n7268), .A(n7259), .B(n7258), .ZN(n7260)
         );
  AOI21_X1 U8952 ( .B1(n9850), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7260), .ZN(
        n7261) );
  OAI21_X1 U8953 ( .B1(n7262), .B2(n9837), .A(n7261), .ZN(P2_U3188) );
  MUX2_X1 U8954 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8334), .Z(n7350) );
  XNOR2_X1 U8955 ( .A(n7350), .B(n7365), .ZN(n7351) );
  INV_X1 U8956 ( .A(n7268), .ZN(n7266) );
  INV_X1 U8957 ( .A(n7263), .ZN(n7265) );
  AOI21_X1 U8958 ( .B1(n7266), .B2(n7265), .A(n7264), .ZN(n7352) );
  XOR2_X1 U8959 ( .A(n7351), .B(n7352), .Z(n7277) );
  NAND2_X1 U8960 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7574) );
  OAI21_X1 U8961 ( .B1(n9855), .B2(n7365), .A(n7574), .ZN(n7275) );
  NOR2_X1 U8962 ( .A1(n7267), .A2(n5334), .ZN(n7357) );
  AOI21_X1 U8963 ( .B1(n5334), .B2(n7267), .A(n7357), .ZN(n7273) );
  NAND2_X1 U8964 ( .A1(n7268), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7269) );
  NAND2_X1 U8965 ( .A1(n7270), .A2(n7269), .ZN(n7364) );
  AOI21_X1 U8966 ( .B1(n5337), .B2(n7271), .A(n7363), .ZN(n7272) );
  OAI22_X1 U8967 ( .A1(n7273), .A2(n9846), .B1(n7272), .B2(n9844), .ZN(n7274)
         );
  AOI211_X1 U8968 ( .C1(n9850), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7275), .B(
        n7274), .ZN(n7276) );
  OAI21_X1 U8969 ( .B1(n7277), .B2(n9837), .A(n7276), .ZN(P2_U3189) );
  OAI222_X1 U8970 ( .A1(n9616), .A2(n7280), .B1(P1_U3086), .B2(n7279), .C1(
        n7925), .C2(n7278), .ZN(P1_U3335) );
  AOI21_X1 U8971 ( .B1(n7283), .B2(n7282), .A(n7281), .ZN(n7297) );
  OAI21_X1 U8972 ( .B1(n7285), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7284), .ZN(
        n7293) );
  OAI22_X1 U8973 ( .A1(n9855), .A2(n7287), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7286), .ZN(n7292) );
  NAND2_X1 U8974 ( .A1(n7288), .A2(n5277), .ZN(n7289) );
  AOI21_X1 U8975 ( .B1(n7290), .B2(n7289), .A(n9844), .ZN(n7291) );
  AOI211_X1 U8976 ( .C1(n7294), .C2(n7293), .A(n7292), .B(n7291), .ZN(n7296)
         );
  NAND2_X1 U8977 ( .A1(n9850), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n7295) );
  OAI211_X1 U8978 ( .C1(n7297), .C2(n9837), .A(n7296), .B(n7295), .ZN(P2_U3185) );
  OAI21_X1 U8979 ( .B1(n7298), .B2(n7299), .A(n7022), .ZN(n9891) );
  OAI22_X1 U8980 ( .A1(n8534), .A2(n9888), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9860), .ZN(n7306) );
  INV_X1 U8981 ( .A(n7299), .ZN(n7300) );
  XNOR2_X1 U8982 ( .A(n7301), .B(n7300), .ZN(n7302) );
  NAND2_X1 U8983 ( .A1(n7302), .A2(n8494), .ZN(n7304) );
  AOI22_X1 U8984 ( .A1(n8500), .A2(n8204), .B1(n8202), .B2(n8499), .ZN(n7303)
         );
  NAND2_X1 U8985 ( .A1(n7304), .A2(n7303), .ZN(n9889) );
  MUX2_X1 U8986 ( .A(n9889), .B(P2_REG2_REG_3__SCAN_IN), .S(n9874), .Z(n7305)
         );
  AOI211_X1 U8987 ( .C1(n8539), .C2(n9891), .A(n7306), .B(n7305), .ZN(n7307)
         );
  INV_X1 U8988 ( .A(n7307), .ZN(P2_U3230) );
  AOI21_X1 U8989 ( .B1(n7310), .B2(n7309), .A(n7308), .ZN(n7315) );
  OAI22_X1 U8990 ( .A1(n8858), .A2(n7311), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10045), .ZN(n7313) );
  OAI22_X1 U8991 ( .A1(n8859), .A2(n7534), .B1(n7322), .B2(n8853), .ZN(n7312)
         );
  AOI211_X1 U8992 ( .C1(n8813), .C2(n9144), .A(n7313), .B(n7312), .ZN(n7314)
         );
  OAI21_X1 U8993 ( .B1(n7315), .B2(n8866), .A(n7314), .ZN(P1_U3227) );
  OAI211_X1 U8994 ( .C1(n9544), .C2(n7318), .A(n7317), .B(n7316), .ZN(n7324)
         );
  NAND2_X1 U8995 ( .A1(n9814), .A2(n9629), .ZN(n9539) );
  OAI22_X1 U8996 ( .A1(n9539), .A2(n7322), .B1(n9814), .B2(n6635), .ZN(n7319)
         );
  AOI21_X1 U8997 ( .B1(n7324), .B2(n9814), .A(n7319), .ZN(n7320) );
  INV_X1 U8998 ( .A(n7320), .ZN(P1_U3527) );
  NAND2_X1 U8999 ( .A1(n9788), .A2(n9629), .ZN(n9595) );
  INV_X1 U9000 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7321) );
  OAI22_X1 U9001 ( .A1(n9595), .A2(n7322), .B1(n9788), .B2(n7321), .ZN(n7323)
         );
  AOI21_X1 U9002 ( .B1(n7324), .B2(n9788), .A(n7323), .ZN(n7325) );
  INV_X1 U9003 ( .A(n7325), .ZN(P1_U3468) );
  OAI21_X1 U9004 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7326), .A(n9822), .ZN(n7327) );
  OAI21_X1 U9005 ( .B1(n9821), .B2(n7328), .A(n7327), .ZN(n7329) );
  OAI21_X1 U9006 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7330), .A(n7329), .ZN(n7331) );
  AOI21_X1 U9007 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9819), .A(n7331), .ZN(n7332) );
  OAI21_X1 U9008 ( .B1(n8341), .B2(n10013), .A(n7332), .ZN(P2_U3182) );
  INV_X1 U9009 ( .A(n7333), .ZN(n7430) );
  OAI222_X1 U9010 ( .A1(n8679), .A2(n9971), .B1(n7962), .B2(n7430), .C1(n7334), 
        .C2(P2_U3151), .ZN(P2_U3274) );
  XNOR2_X1 U9011 ( .A(n4526), .B(n7335), .ZN(n7397) );
  XNOR2_X1 U9012 ( .A(n7397), .B(n8201), .ZN(n7340) );
  INV_X1 U9013 ( .A(n7336), .ZN(n7337) );
  NAND2_X1 U9014 ( .A1(n7339), .A2(n7340), .ZN(n7400) );
  OAI21_X1 U9015 ( .B1(n7340), .B2(n7339), .A(n7400), .ZN(n7341) );
  NAND2_X1 U9016 ( .A1(n7341), .A2(n8170), .ZN(n7348) );
  NAND2_X1 U9017 ( .A1(n8172), .A2(n8202), .ZN(n7345) );
  AOI21_X1 U9018 ( .B1(n8177), .B2(n7343), .A(n7342), .ZN(n7344) );
  OAI211_X1 U9019 ( .C1(n7578), .C2(n8175), .A(n7345), .B(n7344), .ZN(n7346)
         );
  INV_X1 U9020 ( .A(n7346), .ZN(n7347) );
  OAI211_X1 U9021 ( .C1(n7349), .C2(n8150), .A(n7348), .B(n7347), .ZN(P2_U3167) );
  OAI22_X1 U9022 ( .A1(n7352), .A2(n7351), .B1(n7350), .B2(n7365), .ZN(n9835)
         );
  MUX2_X1 U9023 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8334), .Z(n7353) );
  XOR2_X1 U9024 ( .A(n9854), .B(n7353), .Z(n9836) );
  INV_X1 U9025 ( .A(n9854), .ZN(n7369) );
  INV_X1 U9026 ( .A(n7353), .ZN(n7354) );
  AOI22_X1 U9027 ( .A1(n9835), .A2(n9836), .B1(n7369), .B2(n7354), .ZN(n7444)
         );
  MUX2_X1 U9028 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8334), .Z(n7442) );
  XNOR2_X1 U9029 ( .A(n7442), .B(n7441), .ZN(n7443) );
  XNOR2_X1 U9030 ( .A(n7444), .B(n7443), .ZN(n7355) );
  NAND2_X1 U9031 ( .A1(n7355), .A2(n9821), .ZN(n7377) );
  INV_X1 U9032 ( .A(n7441), .ZN(n7375) );
  AND2_X1 U9033 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7705) );
  INV_X1 U9034 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7362) );
  INV_X1 U9035 ( .A(n7356), .ZN(n7358) );
  NAND2_X1 U9036 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n9854), .ZN(n7359) );
  OAI21_X1 U9037 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n9854), .A(n7359), .ZN(
        n9840) );
  NAND2_X1 U9038 ( .A1(n7360), .A2(n7441), .ZN(n7454) );
  AOI21_X1 U9039 ( .B1(n7362), .B2(n7361), .A(n7456), .ZN(n7373) );
  NAND2_X1 U9040 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n9854), .ZN(n7366) );
  OAI21_X1 U9041 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n9854), .A(n7366), .ZN(
        n9843) );
  INV_X1 U9042 ( .A(n9842), .ZN(n7367) );
  OAI21_X1 U9043 ( .B1(n7369), .B2(n7368), .A(n7367), .ZN(n7370) );
  NAND2_X1 U9044 ( .A1(n7370), .A2(n7441), .ZN(n7448) );
  OAI21_X1 U9045 ( .B1(n7370), .B2(n7441), .A(n7448), .ZN(n7371) );
  AOI21_X1 U9046 ( .B1(n5365), .B2(n7371), .A(n7450), .ZN(n7372) );
  OAI22_X1 U9047 ( .A1(n7373), .A2(n9846), .B1(n9844), .B2(n7372), .ZN(n7374)
         );
  AOI211_X1 U9048 ( .C1(n7375), .C2(n9819), .A(n7705), .B(n7374), .ZN(n7376)
         );
  OAI211_X1 U9049 ( .C1(n7378), .C2(n8341), .A(n7377), .B(n7376), .ZN(P2_U3191) );
  NOR2_X1 U9050 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8685), .ZN(n7384) );
  NAND2_X1 U9051 ( .A1(n7391), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7559) );
  OR2_X1 U9052 ( .A1(n7391), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7380) );
  NAND2_X1 U9053 ( .A1(n7559), .A2(n7380), .ZN(n7381) );
  AOI211_X1 U9054 ( .C1(n7382), .C2(n7381), .A(n4595), .B(n9660), .ZN(n7383)
         );
  AOI211_X1 U9055 ( .C1(n9673), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n7384), .B(
        n7383), .ZN(n7395) );
  NAND2_X1 U9056 ( .A1(n7385), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7388) );
  INV_X1 U9057 ( .A(n7388), .ZN(n7393) );
  INV_X1 U9058 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9812) );
  OR2_X1 U9059 ( .A1(n7391), .A2(n9812), .ZN(n7386) );
  OAI211_X1 U9060 ( .C1(n7562), .C2(P1_REG1_REG_14__SCAN_IN), .A(n7387), .B(
        n7386), .ZN(n7392) );
  NAND2_X1 U9061 ( .A1(n7388), .A2(n7387), .ZN(n7390) );
  NAND2_X1 U9062 ( .A1(n7391), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7389) );
  OAI211_X1 U9063 ( .C1(n7391), .C2(P1_REG1_REG_14__SCAN_IN), .A(n7390), .B(
        n7389), .ZN(n7561) );
  OAI211_X1 U9064 ( .C1(n7393), .C2(n7392), .A(n9684), .B(n7561), .ZN(n7394)
         );
  OAI211_X1 U9065 ( .C1(n9212), .C2(n7562), .A(n7395), .B(n7394), .ZN(P1_U3257) );
  INV_X1 U9066 ( .A(n8201), .ZN(n7396) );
  NAND2_X1 U9067 ( .A1(n7397), .A2(n7396), .ZN(n7398) );
  AND2_X1 U9068 ( .A1(n7400), .A2(n7398), .ZN(n7402) );
  XNOR2_X1 U9069 ( .A(n4526), .B(n9896), .ZN(n7570) );
  XNOR2_X1 U9070 ( .A(n7570), .B(n8200), .ZN(n7401) );
  OAI211_X1 U9071 ( .C1(n7402), .C2(n7401), .A(n8170), .B(n7569), .ZN(n7409)
         );
  INV_X1 U9072 ( .A(n8199), .ZN(n7687) );
  NAND2_X1 U9073 ( .A1(n8172), .A2(n8201), .ZN(n7406) );
  AOI21_X1 U9074 ( .B1(n8177), .B2(n7404), .A(n7403), .ZN(n7405) );
  OAI211_X1 U9075 ( .C1(n7687), .C2(n8175), .A(n7406), .B(n7405), .ZN(n7407)
         );
  INV_X1 U9076 ( .A(n7407), .ZN(n7408) );
  OAI211_X1 U9077 ( .C1(n7413), .C2(n8150), .A(n7409), .B(n7408), .ZN(P2_U3179) );
  NAND2_X1 U9078 ( .A1(n7410), .A2(n7411), .ZN(n7412) );
  XNOR2_X1 U9079 ( .A(n7412), .B(n7415), .ZN(n9899) );
  OAI22_X1 U9080 ( .A1(n8534), .A2(n9896), .B1(n7413), .B2(n9860), .ZN(n7420)
         );
  XNOR2_X1 U9081 ( .A(n7414), .B(n7415), .ZN(n7416) );
  NAND2_X1 U9082 ( .A1(n7416), .A2(n8494), .ZN(n7418) );
  AOI22_X1 U9083 ( .A1(n8500), .A2(n8201), .B1(n8199), .B2(n8499), .ZN(n7417)
         );
  NAND2_X1 U9084 ( .A1(n7418), .A2(n7417), .ZN(n9897) );
  MUX2_X1 U9085 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n9897), .S(n9872), .Z(n7419)
         );
  AOI211_X1 U9086 ( .C1(n8539), .C2(n9899), .A(n7420), .B(n7419), .ZN(n7421)
         );
  INV_X1 U9087 ( .A(n7421), .ZN(P2_U3227) );
  AOI211_X1 U9088 ( .C1(n9802), .C2(n7424), .A(n7423), .B(n7422), .ZN(n7429)
         );
  INV_X1 U9089 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10262) );
  OAI22_X1 U9090 ( .A1(n9595), .A2(n7488), .B1(n9788), .B2(n10262), .ZN(n7425)
         );
  INV_X1 U9091 ( .A(n7425), .ZN(n7426) );
  OAI21_X1 U9092 ( .B1(n7429), .B2(n9967), .A(n7426), .ZN(P1_U3471) );
  OAI22_X1 U9093 ( .A1(n9539), .A2(n7488), .B1(n9814), .B2(n6633), .ZN(n7427)
         );
  INV_X1 U9094 ( .A(n7427), .ZN(n7428) );
  OAI21_X1 U9095 ( .B1(n7429), .B2(n9811), .A(n7428), .ZN(P1_U3528) );
  OAI222_X1 U9096 ( .A1(P1_U3086), .A2(n9062), .B1(n7925), .B2(n7430), .C1(
        n10232), .C2(n9616), .ZN(P1_U3334) );
  OAI21_X1 U9097 ( .B1(n7432), .B2(n7434), .A(n7431), .ZN(n9901) );
  XOR2_X1 U9098 ( .A(n7434), .B(n7433), .Z(n7435) );
  NAND2_X1 U9099 ( .A1(n7435), .A2(n8494), .ZN(n7437) );
  AOI22_X1 U9100 ( .A1(n8500), .A2(n8200), .B1(n8198), .B2(n8499), .ZN(n7436)
         );
  OAI211_X1 U9101 ( .C1(n9862), .C2(n9901), .A(n7437), .B(n7436), .ZN(n9903)
         );
  OAI22_X1 U9102 ( .A1(n9901), .A2(n7648), .B1(n7573), .B2(n9860), .ZN(n7438)
         );
  OAI21_X1 U9103 ( .B1(n9903), .B2(n7438), .A(n9872), .ZN(n7440) );
  NAND2_X1 U9104 ( .A1(n8524), .A2(n7576), .ZN(n7439) );
  OAI211_X1 U9105 ( .C1(n5334), .C2(n9872), .A(n7440), .B(n7439), .ZN(P2_U3226) );
  OAI22_X1 U9106 ( .A1(n7444), .A2(n7443), .B1(n7442), .B2(n7441), .ZN(n7446)
         );
  MUX2_X1 U9107 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8334), .Z(n7639) );
  XOR2_X1 U9108 ( .A(n7638), .B(n7639), .Z(n7445) );
  NAND2_X1 U9109 ( .A1(n7445), .A2(n7446), .ZN(n7640) );
  OAI21_X1 U9110 ( .B1(n7446), .B2(n7445), .A(n7640), .ZN(n7447) );
  NAND2_X1 U9111 ( .A1(n7447), .A2(n9821), .ZN(n7463) );
  INV_X1 U9112 ( .A(n7638), .ZN(n7461) );
  INV_X1 U9113 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9999) );
  NOR2_X1 U9114 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9999), .ZN(n7996) );
  INV_X1 U9115 ( .A(n7448), .ZN(n7449) );
  MUX2_X1 U9116 ( .A(n7451), .B(P2_REG1_REG_10__SCAN_IN), .S(n7638), .Z(n7452)
         );
  AOI21_X1 U9117 ( .B1(n7453), .B2(n7452), .A(n7634), .ZN(n7459) );
  INV_X1 U9118 ( .A(n7454), .ZN(n7455) );
  MUX2_X1 U9119 ( .A(n10185), .B(P2_REG2_REG_10__SCAN_IN), .S(n7638), .Z(n7457) );
  AOI21_X1 U9120 ( .B1(n4492), .B2(n7457), .A(n7631), .ZN(n7458) );
  OAI22_X1 U9121 ( .A1(n7459), .A2(n9844), .B1(n9846), .B2(n7458), .ZN(n7460)
         );
  AOI211_X1 U9122 ( .C1(n7461), .C2(n9819), .A(n7996), .B(n7460), .ZN(n7462)
         );
  OAI211_X1 U9123 ( .C1(n10000), .C2(n8341), .A(n7463), .B(n7462), .ZN(
        P2_U3192) );
  NAND2_X1 U9124 ( .A1(n7431), .A2(n7464), .ZN(n7465) );
  XNOR2_X1 U9125 ( .A(n7465), .B(n7466), .ZN(n9906) );
  INV_X1 U9126 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7471) );
  XNOR2_X1 U9127 ( .A(n7467), .B(n7466), .ZN(n7468) );
  NAND2_X1 U9128 ( .A1(n7468), .A2(n8494), .ZN(n7470) );
  AOI22_X1 U9129 ( .A1(n8500), .A2(n8199), .B1(n8197), .B2(n8499), .ZN(n7469)
         );
  AND2_X1 U9130 ( .A1(n7470), .A2(n7469), .ZN(n9908) );
  MUX2_X1 U9131 ( .A(n7471), .B(n9908), .S(n9872), .Z(n7474) );
  INV_X1 U9132 ( .A(n7698), .ZN(n7472) );
  AOI22_X1 U9133 ( .A1(n8524), .A2(n7692), .B1(n8466), .B2(n7472), .ZN(n7473)
         );
  OAI211_X1 U9134 ( .C1(n9906), .C2(n8552), .A(n7474), .B(n7473), .ZN(P2_U3225) );
  XOR2_X1 U9135 ( .A(n7475), .B(n4500), .Z(n7482) );
  AOI22_X1 U9136 ( .A1(n7476), .A2(n8829), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7477) );
  OAI21_X1 U9137 ( .B1(n7478), .B2(n8858), .A(n7477), .ZN(n7479) );
  AOI21_X1 U9138 ( .B1(n7480), .B2(n8864), .A(n7479), .ZN(n7481) );
  OAI21_X1 U9139 ( .B1(n7482), .B2(n8866), .A(n7481), .ZN(P1_U3239) );
  INV_X1 U9140 ( .A(n7483), .ZN(n7486) );
  OAI222_X1 U9141 ( .A1(n8679), .A2(n7485), .B1(n7962), .B2(n7486), .C1(
        P2_U3151), .C2(n7484), .ZN(P2_U3273) );
  OAI222_X1 U9142 ( .A1(n9616), .A2(n7487), .B1(n7925), .B2(n7486), .C1(
        P1_U3086), .C2(n9050), .ZN(P1_U3333) );
  NAND2_X1 U9143 ( .A1(n7534), .A2(n7488), .ZN(n7489) );
  NAND2_X1 U9144 ( .A1(n7490), .A2(n7489), .ZN(n7598) );
  NAND2_X1 U9145 ( .A1(n7491), .A2(n9705), .ZN(n9023) );
  INV_X1 U9146 ( .A(n7491), .ZN(n9141) );
  NAND2_X1 U9147 ( .A1(n7611), .A2(n9141), .ZN(n8894) );
  NAND2_X1 U9148 ( .A1(n9023), .A2(n8894), .ZN(n8892) );
  NAND2_X1 U9149 ( .A1(n7491), .A2(n7611), .ZN(n7492) );
  OR2_X1 U9150 ( .A1(n7779), .A2(n7548), .ZN(n8895) );
  NAND2_X1 U9151 ( .A1(n7779), .A2(n7548), .ZN(n8883) );
  NAND2_X1 U9152 ( .A1(n8895), .A2(n8883), .ZN(n7496) );
  OAI21_X1 U9153 ( .B1(n7493), .B2(n7496), .A(n7521), .ZN(n9771) );
  INV_X1 U9154 ( .A(n9771), .ZN(n7508) );
  NOR2_X1 U9155 ( .A1(n4419), .A2(n7494), .ZN(n9743) );
  INV_X1 U9156 ( .A(n9743), .ZN(n7507) );
  NAND2_X1 U9157 ( .A1(n7515), .A2(n9024), .ZN(n9067) );
  INV_X1 U9158 ( .A(n8894), .ZN(n7495) );
  NOR2_X1 U9159 ( .A1(n7600), .A2(n7495), .ZN(n7497) );
  INV_X1 U9160 ( .A(n9023), .ZN(n7509) );
  OAI21_X1 U9161 ( .B1(n7497), .B2(n7509), .A(n4952), .ZN(n7539) );
  INV_X1 U9162 ( .A(n7539), .ZN(n7499) );
  NOR3_X1 U9163 ( .A1(n7497), .A2(n7509), .A3(n4952), .ZN(n7498) );
  OAI21_X1 U9164 ( .B1(n7499), .B2(n7498), .A(n9715), .ZN(n7501) );
  INV_X1 U9165 ( .A(n7518), .ZN(n9139) );
  AOI22_X1 U9166 ( .A1(n9461), .A2(n9141), .B1(n9139), .B2(n9460), .ZN(n7500)
         );
  OAI211_X1 U9167 ( .C1(n7508), .C2(n7599), .A(n7501), .B(n7500), .ZN(n9769)
         );
  NAND2_X1 U9168 ( .A1(n9769), .A2(n9471), .ZN(n7506) );
  OAI22_X1 U9169 ( .A1(n9471), .A2(n7502), .B1(n7777), .B2(n9701), .ZN(n7504)
         );
  NAND2_X1 U9170 ( .A1(n7604), .A2(n9768), .ZN(n7545) );
  OAI211_X1 U9171 ( .C1(n7604), .C2(n9768), .A(n9738), .B(n7545), .ZN(n9767)
         );
  NOR2_X1 U9172 ( .A1(n9767), .A2(n9740), .ZN(n7503) );
  AOI211_X1 U9173 ( .C1(n9706), .C2(n7779), .A(n7504), .B(n7503), .ZN(n7505)
         );
  OAI211_X1 U9174 ( .C1(n7508), .C2(n7507), .A(n7506), .B(n7505), .ZN(P1_U3285) );
  NAND2_X1 U9175 ( .A1(n8711), .A2(n8828), .ZN(n9552) );
  INV_X1 U9176 ( .A(n9028), .ZN(n7517) );
  AND2_X1 U9177 ( .A1(n9025), .A2(n5032), .ZN(n7514) );
  OR2_X1 U9178 ( .A1(n8896), .A2(n7509), .ZN(n7511) );
  OR2_X1 U9179 ( .A1(n7627), .A2(n7518), .ZN(n8900) );
  NAND2_X1 U9180 ( .A1(n8900), .A2(n8895), .ZN(n8884) );
  NAND2_X1 U9181 ( .A1(n8884), .A2(n8908), .ZN(n7510) );
  NAND2_X1 U9182 ( .A1(n7511), .A2(n7510), .ZN(n9068) );
  INV_X1 U9183 ( .A(n8884), .ZN(n7513) );
  AND2_X1 U9184 ( .A1(n8894), .A2(n8890), .ZN(n7512) );
  NAND2_X1 U9185 ( .A1(n7513), .A2(n7512), .ZN(n9027) );
  OAI21_X1 U9186 ( .B1(n7517), .B2(n7516), .A(n9554), .ZN(n7520) );
  OAI22_X1 U9187 ( .A1(n7518), .A2(n9393), .B1(n7668), .B2(n9439), .ZN(n7519)
         );
  AOI21_X1 U9188 ( .B1(n7520), .B2(n9715), .A(n7519), .ZN(n9773) );
  INV_X1 U9189 ( .A(n7548), .ZN(n9140) );
  NAND2_X1 U9190 ( .A1(n8900), .A2(n8908), .ZN(n7543) );
  NAND2_X1 U9191 ( .A1(n7544), .A2(n7543), .ZN(n7542) );
  OR2_X1 U9192 ( .A1(n7627), .A2(n9139), .ZN(n7522) );
  OAI21_X1 U9193 ( .B1(n7523), .B2(n9028), .A(n7667), .ZN(n9776) );
  NAND2_X1 U9194 ( .A1(n9776), .A2(n9725), .ZN(n7529) );
  OAI22_X1 U9195 ( .A1(n9471), .A2(n7524), .B1(n8709), .B2(n9701), .ZN(n7527)
         );
  INV_X1 U9196 ( .A(n8711), .ZN(n9774) );
  INV_X1 U9197 ( .A(n7547), .ZN(n7525) );
  INV_X1 U9198 ( .A(n7669), .ZN(n9550) );
  OAI211_X1 U9199 ( .C1(n9774), .C2(n7525), .A(n9550), .B(n9738), .ZN(n9772)
         );
  NOR2_X1 U9200 ( .A1(n9772), .A2(n9740), .ZN(n7526) );
  AOI211_X1 U9201 ( .C1(n9706), .C2(n8711), .A(n7527), .B(n7526), .ZN(n7528)
         );
  OAI211_X1 U9202 ( .C1(n4419), .C2(n9773), .A(n7529), .B(n7528), .ZN(P1_U3283) );
  XNOR2_X1 U9203 ( .A(n7531), .B(n7530), .ZN(n7532) );
  XNOR2_X1 U9204 ( .A(n7533), .B(n7532), .ZN(n7538) );
  OAI22_X1 U9205 ( .A1(n7534), .A2(n9393), .B1(n7548), .B2(n9439), .ZN(n7603)
         );
  AOI22_X1 U9206 ( .A1(n7603), .A2(n8829), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7535) );
  OAI21_X1 U9207 ( .B1(n9702), .B2(n8858), .A(n7535), .ZN(n7536) );
  AOI21_X1 U9208 ( .B1(n9705), .B2(n8864), .A(n7536), .ZN(n7537) );
  OAI21_X1 U9209 ( .B1(n7538), .B2(n8866), .A(n7537), .ZN(P1_U3213) );
  NAND2_X1 U9210 ( .A1(n7539), .A2(n8883), .ZN(n7540) );
  XNOR2_X1 U9211 ( .A(n7540), .B(n7543), .ZN(n7541) );
  NOR2_X1 U9212 ( .A1(n7541), .A2(n9732), .ZN(n7623) );
  INV_X1 U9213 ( .A(n7623), .ZN(n7558) );
  OAI21_X1 U9214 ( .B1(n7544), .B2(n7543), .A(n7542), .ZN(n7625) );
  INV_X1 U9215 ( .A(n7627), .ZN(n8786) );
  NAND2_X1 U9216 ( .A1(n7545), .A2(n7627), .ZN(n7546) );
  NAND3_X1 U9217 ( .A1(n7547), .A2(n9738), .A3(n7546), .ZN(n7552) );
  OR2_X1 U9218 ( .A1(n7548), .A2(n9393), .ZN(n7550) );
  OR2_X1 U9219 ( .A1(n8828), .A2(n9439), .ZN(n7549) );
  NAND2_X1 U9220 ( .A1(n7550), .A2(n7549), .ZN(n8782) );
  INV_X1 U9221 ( .A(n8782), .ZN(n7551) );
  NAND2_X1 U9222 ( .A1(n7552), .A2(n7551), .ZN(n7624) );
  NAND2_X1 U9223 ( .A1(n7624), .A2(n9724), .ZN(n7555) );
  INV_X1 U9224 ( .A(n7553), .ZN(n8783) );
  AOI22_X1 U9225 ( .A1(n4419), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8783), .B2(
        n9736), .ZN(n7554) );
  OAI211_X1 U9226 ( .C1(n8786), .C2(n9741), .A(n7555), .B(n7554), .ZN(n7556)
         );
  AOI21_X1 U9227 ( .B1(n7625), .B2(n9725), .A(n7556), .ZN(n7557) );
  OAI21_X1 U9228 ( .B1(n7558), .B2(n4419), .A(n7557), .ZN(P1_U3284) );
  NOR2_X1 U9229 ( .A1(n9446), .A2(n7560), .ZN(n9150) );
  AOI211_X1 U9230 ( .C1(n9446), .C2(n7560), .A(n9150), .B(n9660), .ZN(n7568)
         );
  OAI21_X1 U9231 ( .B1(n9812), .B2(n7562), .A(n7561), .ZN(n9155) );
  XNOR2_X1 U9232 ( .A(n9155), .B(n9148), .ZN(n7563) );
  NAND2_X1 U9233 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7563), .ZN(n9157) );
  OAI211_X1 U9234 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7563), .A(n9684), .B(
        n9157), .ZN(n7566) );
  NOR2_X1 U9235 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8857), .ZN(n7564) );
  AOI21_X1 U9236 ( .B1(n9673), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n7564), .ZN(
        n7565) );
  OAI211_X1 U9237 ( .C1(n9212), .C2(n9148), .A(n7566), .B(n7565), .ZN(n7567)
         );
  OR2_X1 U9238 ( .A1(n7568), .A2(n7567), .ZN(P1_U3258) );
  XNOR2_X1 U9239 ( .A(n4526), .B(n7576), .ZN(n7685) );
  XNOR2_X1 U9240 ( .A(n7685), .B(n8199), .ZN(n7572) );
  AOI21_X1 U9241 ( .B1(n7572), .B2(n7571), .A(n7686), .ZN(n7582) );
  NOR2_X1 U9242 ( .A1(n8150), .A2(n7573), .ZN(n7580) );
  INV_X1 U9243 ( .A(n8172), .ZN(n8104) );
  INV_X1 U9244 ( .A(n7574), .ZN(n7575) );
  AOI21_X1 U9245 ( .B1(n8177), .B2(n7576), .A(n7575), .ZN(n7577) );
  OAI21_X1 U9246 ( .B1(n8104), .B2(n7578), .A(n7577), .ZN(n7579) );
  AOI211_X1 U9247 ( .C1(n8102), .C2(n8198), .A(n7580), .B(n7579), .ZN(n7581)
         );
  OAI21_X1 U9248 ( .B1(n7582), .B2(n8119), .A(n7581), .ZN(P2_U3153) );
  INV_X1 U9249 ( .A(n8198), .ZN(n7699) );
  XOR2_X1 U9250 ( .A(n7583), .B(n7586), .Z(n7584) );
  OAI222_X1 U9251 ( .A1(n9863), .A2(n8036), .B1(n9865), .B2(n7699), .C1(n9869), 
        .C2(n7584), .ZN(n7615) );
  INV_X1 U9252 ( .A(n7615), .ZN(n7591) );
  XOR2_X1 U9253 ( .A(n7586), .B(n7585), .Z(n7616) );
  INV_X1 U9254 ( .A(n7587), .ZN(n7707) );
  AOI22_X1 U9255 ( .A1(n9874), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n8466), .B2(
        n7707), .ZN(n7588) );
  OAI21_X1 U9256 ( .B1(n7618), .B2(n8534), .A(n7588), .ZN(n7589) );
  AOI21_X1 U9257 ( .B1(n7616), .B2(n8539), .A(n7589), .ZN(n7590) );
  OAI21_X1 U9258 ( .B1(n7591), .B2(n9874), .A(n7590), .ZN(P2_U3224) );
  NAND2_X1 U9259 ( .A1(n7594), .A2(n9608), .ZN(n7592) );
  OAI211_X1 U9260 ( .C1(n7593), .C2(n9616), .A(n7592), .B(n9113), .ZN(P1_U3332) );
  NAND2_X1 U9261 ( .A1(n7594), .A2(n4503), .ZN(n7596) );
  OAI211_X1 U9262 ( .C1(n9986), .C2(n8679), .A(n7596), .B(n7595), .ZN(P2_U3272) );
  OAI21_X1 U9263 ( .B1(n7598), .B2(n8892), .A(n7597), .ZN(n9710) );
  INV_X1 U9264 ( .A(n9710), .ZN(n7607) );
  INV_X1 U9265 ( .A(n7599), .ZN(n9735) );
  NAND2_X1 U9266 ( .A1(n7600), .A2(n8892), .ZN(n7601) );
  AOI21_X1 U9267 ( .B1(n8886), .B2(n7601), .A(n9732), .ZN(n7602) );
  AOI211_X1 U9268 ( .C1(n9735), .C2(n9710), .A(n7603), .B(n7602), .ZN(n9712)
         );
  INV_X1 U9269 ( .A(n7604), .ZN(n7605) );
  OAI211_X1 U9270 ( .C1(n7611), .C2(n7606), .A(n7605), .B(n9738), .ZN(n9708)
         );
  OAI211_X1 U9271 ( .C1(n7607), .C2(n9546), .A(n9712), .B(n9708), .ZN(n7613)
         );
  OAI22_X1 U9272 ( .A1(n9539), .A2(n7611), .B1(n9814), .B2(n6645), .ZN(n7608)
         );
  AOI21_X1 U9273 ( .B1(n7613), .B2(n9814), .A(n7608), .ZN(n7609) );
  INV_X1 U9274 ( .A(n7609), .ZN(P1_U3529) );
  INV_X1 U9275 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7610) );
  OAI22_X1 U9276 ( .A1(n9595), .A2(n7611), .B1(n9788), .B2(n7610), .ZN(n7612)
         );
  AOI21_X1 U9277 ( .B1(n7613), .B2(n9788), .A(n7612), .ZN(n7614) );
  INV_X1 U9278 ( .A(n7614), .ZN(P1_U3474) );
  AOI21_X1 U9279 ( .B1(n7616), .B2(n9920), .A(n7615), .ZN(n7622) );
  INV_X1 U9280 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7617) );
  OAI22_X1 U9281 ( .A1(n7618), .A2(n8667), .B1(n9928), .B2(n7617), .ZN(n7619)
         );
  INV_X1 U9282 ( .A(n7619), .ZN(n7620) );
  OAI21_X1 U9283 ( .B1(n7622), .B2(n9929), .A(n7620), .ZN(P2_U3417) );
  AOI22_X1 U9284 ( .A1(n8607), .A2(n7706), .B1(n9939), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n7621) );
  OAI21_X1 U9285 ( .B1(n7622), .B2(n9939), .A(n7621), .ZN(P2_U3468) );
  AOI211_X1 U9286 ( .C1(n9802), .C2(n7625), .A(n7624), .B(n7623), .ZN(n7630)
         );
  INV_X1 U9287 ( .A(n9539), .ZN(n9560) );
  AOI22_X1 U9288 ( .A1(n9560), .A2(n7627), .B1(n9811), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7626) );
  OAI21_X1 U9289 ( .B1(n7630), .B2(n9811), .A(n7626), .ZN(P1_U3531) );
  INV_X1 U9290 ( .A(n9595), .ZN(n7628) );
  AOI22_X1 U9291 ( .A1(n7628), .A2(n7627), .B1(n9967), .B2(
        P1_REG0_REG_9__SCAN_IN), .ZN(n7629) );
  OAI21_X1 U9292 ( .B1(n7630), .B2(n9967), .A(n7629), .ZN(P1_U3480) );
  NOR2_X1 U9293 ( .A1(n5394), .A2(n7633), .ZN(n7730) );
  AOI21_X1 U9294 ( .B1(n5394), .B2(n7633), .A(n7730), .ZN(n7647) );
  INV_X1 U9295 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10010) );
  NOR2_X1 U9296 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10010), .ZN(n8134) );
  AOI21_X1 U9297 ( .B1(n7635), .B2(n5397), .A(n7712), .ZN(n7636) );
  NOR2_X1 U9298 ( .A1(n9844), .A2(n7636), .ZN(n7637) );
  AOI211_X1 U9299 ( .C1(n7729), .C2(n9819), .A(n8134), .B(n7637), .ZN(n7646)
         );
  MUX2_X1 U9300 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8334), .Z(n7716) );
  XNOR2_X1 U9301 ( .A(n7716), .B(n7729), .ZN(n7643) );
  OR2_X1 U9302 ( .A1(n7639), .A2(n7638), .ZN(n7641) );
  NAND2_X1 U9303 ( .A1(n7641), .A2(n7640), .ZN(n7642) );
  NAND2_X1 U9304 ( .A1(n7643), .A2(n7642), .ZN(n7717) );
  OAI21_X1 U9305 ( .B1(n7643), .B2(n7642), .A(n7717), .ZN(n7644) );
  AOI22_X1 U9306 ( .A1(n9850), .A2(P2_ADDR_REG_11__SCAN_IN), .B1(n9821), .B2(
        n7644), .ZN(n7645) );
  OAI211_X1 U9307 ( .C1(n7647), .C2(n9846), .A(n7646), .B(n7645), .ZN(P2_U3193) );
  INV_X1 U9308 ( .A(n7648), .ZN(n9871) );
  INV_X1 U9309 ( .A(n7651), .ZN(n7649) );
  XNOR2_X1 U9310 ( .A(n7650), .B(n7649), .ZN(n9912) );
  INV_X1 U9311 ( .A(n9912), .ZN(n7656) );
  XNOR2_X1 U9312 ( .A(n7652), .B(n7651), .ZN(n7654) );
  INV_X1 U9313 ( .A(n8197), .ZN(n7817) );
  OAI22_X1 U9314 ( .A1(n7817), .A2(n9865), .B1(n8038), .B2(n9863), .ZN(n7653)
         );
  AOI21_X1 U9315 ( .B1(n7654), .B2(n8494), .A(n7653), .ZN(n7655) );
  OAI21_X1 U9316 ( .B1(n9912), .B2(n9862), .A(n7655), .ZN(n9914) );
  AOI21_X1 U9317 ( .B1(n9871), .B2(n7656), .A(n9914), .ZN(n7659) );
  INV_X1 U9318 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10185) );
  OAI22_X1 U9319 ( .A1(n9872), .A2(n10185), .B1(n7998), .B2(n9860), .ZN(n7657)
         );
  AOI21_X1 U9320 ( .B1(n8524), .B2(n7997), .A(n7657), .ZN(n7658) );
  OAI21_X1 U9321 ( .B1(n7659), .B2(n9874), .A(n7658), .ZN(P2_U3223) );
  OR2_X1 U9322 ( .A1(n4422), .A2(n7668), .ZN(n8912) );
  NAND2_X1 U9323 ( .A1(n4422), .A2(n7668), .ZN(n8910) );
  OR2_X2 U9324 ( .A1(n8738), .A2(n8827), .ZN(n8913) );
  NAND2_X1 U9325 ( .A1(n8738), .A2(n8827), .ZN(n9081) );
  NAND2_X1 U9326 ( .A1(n8913), .A2(n9081), .ZN(n7745) );
  INV_X1 U9327 ( .A(n8910), .ZN(n7660) );
  INV_X1 U9328 ( .A(n7739), .ZN(n7662) );
  INV_X1 U9329 ( .A(n7745), .ZN(n9031) );
  AOI21_X1 U9330 ( .B1(n9556), .B2(n8910), .A(n9031), .ZN(n7661) );
  NOR3_X1 U9331 ( .A1(n7662), .A2(n7661), .A3(n9732), .ZN(n7665) );
  OR2_X1 U9332 ( .A1(n7668), .A2(n9393), .ZN(n7664) );
  OR2_X1 U9333 ( .A1(n8686), .A2(n9439), .ZN(n7663) );
  NAND2_X1 U9334 ( .A1(n7664), .A2(n7663), .ZN(n8733) );
  NOR2_X1 U9335 ( .A1(n7665), .A2(n8733), .ZN(n9779) );
  INV_X1 U9336 ( .A(n8828), .ZN(n9138) );
  OR2_X1 U9337 ( .A1(n8711), .A2(n9138), .ZN(n7666) );
  XNOR2_X1 U9338 ( .A(n7746), .B(n7745), .ZN(n9782) );
  NAND2_X1 U9339 ( .A1(n9782), .A2(n9725), .ZN(n7673) );
  OAI22_X1 U9340 ( .A1(n9471), .A2(n6227), .B1(n8736), .B2(n9701), .ZN(n7671)
         );
  OAI211_X1 U9341 ( .C1(n9548), .C2(n9780), .A(n9738), .B(n7750), .ZN(n9778)
         );
  NOR2_X1 U9342 ( .A1(n9778), .A2(n9740), .ZN(n7670) );
  AOI211_X1 U9343 ( .C1(n9706), .C2(n8738), .A(n7671), .B(n7670), .ZN(n7672)
         );
  OAI211_X1 U9344 ( .C1(n4419), .C2(n9779), .A(n7673), .B(n7672), .ZN(P1_U3281) );
  XNOR2_X1 U9345 ( .A(n7674), .B(n7820), .ZN(n7675) );
  OAI222_X1 U9346 ( .A1(n9863), .A2(n8137), .B1(n9865), .B2(n8036), .C1(n7675), 
        .C2(n9869), .ZN(n9917) );
  INV_X1 U9347 ( .A(n9917), .ZN(n7681) );
  OAI21_X1 U9348 ( .B1(n7677), .B2(n4421), .A(n7676), .ZN(n9919) );
  NOR2_X1 U9349 ( .A1(n8534), .A2(n9916), .ZN(n7679) );
  OAI22_X1 U9350 ( .A1(n9872), .A2(n5394), .B1(n8140), .B2(n9860), .ZN(n7678)
         );
  AOI211_X1 U9351 ( .C1(n9919), .C2(n8539), .A(n7679), .B(n7678), .ZN(n7680)
         );
  OAI21_X1 U9352 ( .B1(n7681), .B2(n9874), .A(n7680), .ZN(P2_U3222) );
  INV_X1 U9353 ( .A(n7682), .ZN(n7770) );
  OAI222_X1 U9354 ( .A1(n7684), .A2(P1_U3086), .B1(n7925), .B2(n7770), .C1(
        n7683), .C2(n9616), .ZN(P1_U3331) );
  INV_X1 U9355 ( .A(n7685), .ZN(n7688) );
  XNOR2_X1 U9356 ( .A(n7847), .B(n9905), .ZN(n7700) );
  XNOR2_X1 U9357 ( .A(n7700), .B(n7699), .ZN(n7689) );
  XNOR2_X1 U9358 ( .A(n7703), .B(n7689), .ZN(n7690) );
  NAND2_X1 U9359 ( .A1(n7690), .A2(n8170), .ZN(n7697) );
  NAND2_X1 U9360 ( .A1(n8172), .A2(n8199), .ZN(n7694) );
  INV_X1 U9361 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7691) );
  NOR2_X1 U9362 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7691), .ZN(n9851) );
  AOI21_X1 U9363 ( .B1(n8177), .B2(n7692), .A(n9851), .ZN(n7693) );
  OAI211_X1 U9364 ( .C1(n7817), .C2(n8175), .A(n7694), .B(n7693), .ZN(n7695)
         );
  INV_X1 U9365 ( .A(n7695), .ZN(n7696) );
  OAI211_X1 U9366 ( .C1(n7698), .C2(n8150), .A(n7697), .B(n7696), .ZN(P2_U3161) );
  NAND2_X1 U9367 ( .A1(n7700), .A2(n7699), .ZN(n7702) );
  INV_X1 U9368 ( .A(n7700), .ZN(n7701) );
  XNOR2_X1 U9369 ( .A(n7847), .B(n7706), .ZN(n7815) );
  XNOR2_X1 U9370 ( .A(n7815), .B(n8197), .ZN(n7818) );
  XNOR2_X1 U9371 ( .A(n7819), .B(n7818), .ZN(n7710) );
  NOR2_X1 U9372 ( .A1(n8175), .A2(n8036), .ZN(n7704) );
  AOI211_X1 U9373 ( .C1(n8172), .C2(n8198), .A(n7705), .B(n7704), .ZN(n7709)
         );
  AOI22_X1 U9374 ( .A1(n8179), .A2(n7707), .B1(n7706), .B2(n8177), .ZN(n7708)
         );
  OAI211_X1 U9375 ( .C1(n7710), .C2(n8119), .A(n7709), .B(n7708), .ZN(P2_U3171) );
  MUX2_X1 U9376 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7714), .S(n7732), .Z(n7715)
         );
  AOI21_X1 U9377 ( .B1(n4495), .B2(n7715), .A(n7789), .ZN(n7738) );
  MUX2_X1 U9378 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8334), .Z(n7796) );
  XNOR2_X1 U9379 ( .A(n7796), .B(n7732), .ZN(n7720) );
  OR2_X1 U9380 ( .A1(n7716), .A2(n7632), .ZN(n7718) );
  NAND2_X1 U9381 ( .A1(n7718), .A2(n7717), .ZN(n7719) );
  NAND2_X1 U9382 ( .A1(n7720), .A2(n7719), .ZN(n7797) );
  OAI21_X1 U9383 ( .B1(n7720), .B2(n7719), .A(n7797), .ZN(n7726) );
  NOR2_X1 U9384 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7721), .ZN(n8041) );
  INV_X1 U9385 ( .A(n8041), .ZN(n7722) );
  OAI21_X1 U9386 ( .B1(n9855), .B2(n7795), .A(n7722), .ZN(n7725) );
  NOR2_X1 U9387 ( .A1(n8341), .A2(n7723), .ZN(n7724) );
  AOI211_X1 U9388 ( .C1(n9821), .C2(n7726), .A(n7725), .B(n7724), .ZN(n7737)
         );
  NOR2_X1 U9389 ( .A1(n7729), .A2(n7728), .ZN(n7731) );
  AOI22_X1 U9390 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7732), .B1(n7795), .B2(
        n7761), .ZN(n7733) );
  NOR2_X1 U9391 ( .A1(n7734), .A2(n7733), .ZN(n7787) );
  AOI21_X1 U9392 ( .B1(n7734), .B2(n7733), .A(n7787), .ZN(n7735) );
  OR2_X1 U9393 ( .A1(n7735), .A2(n9846), .ZN(n7736) );
  OAI211_X1 U9394 ( .C1(n7738), .C2(n9844), .A(n7737), .B(n7736), .ZN(P2_U3194) );
  OR2_X1 U9395 ( .A1(n8807), .A2(n8686), .ZN(n8915) );
  NAND2_X1 U9396 ( .A1(n8807), .A2(n8686), .ZN(n9082) );
  NAND2_X1 U9397 ( .A1(n8915), .A2(n9082), .ZN(n9033) );
  NAND2_X1 U9398 ( .A1(n7740), .A2(n9033), .ZN(n7741) );
  NAND2_X1 U9399 ( .A1(n7909), .A2(n7741), .ZN(n7744) );
  NAND2_X1 U9400 ( .A1(n9437), .A2(n9460), .ZN(n7742) );
  OAI21_X1 U9401 ( .B1(n8827), .B2(n9393), .A(n7742), .ZN(n7743) );
  AOI21_X1 U9402 ( .B1(n7744), .B2(n9715), .A(n7743), .ZN(n9784) );
  NAND2_X1 U9403 ( .A1(n7746), .A2(n7745), .ZN(n7748) );
  INV_X1 U9404 ( .A(n8827), .ZN(n9137) );
  OR2_X1 U9405 ( .A1(n8738), .A2(n9137), .ZN(n7747) );
  XNOR2_X1 U9406 ( .A(n7877), .B(n9033), .ZN(n9786) );
  NAND2_X1 U9407 ( .A1(n9786), .A2(n9725), .ZN(n7755) );
  OAI22_X1 U9408 ( .A1(n9471), .A2(n7749), .B1(n8804), .B2(n9701), .ZN(n7753)
         );
  INV_X1 U9409 ( .A(n7750), .ZN(n7751) );
  OAI211_X1 U9410 ( .C1(n7751), .C2(n4703), .A(n9738), .B(n9466), .ZN(n9783)
         );
  NOR2_X1 U9411 ( .A1(n9783), .A2(n9740), .ZN(n7752) );
  AOI211_X1 U9412 ( .C1(n9706), .C2(n8807), .A(n7753), .B(n7752), .ZN(n7754)
         );
  OAI211_X1 U9413 ( .C1(n4419), .C2(n9784), .A(n7755), .B(n7754), .ZN(P1_U3280) );
  OAI21_X1 U9414 ( .B1(n7757), .B2(n5419), .A(n7756), .ZN(n9923) );
  XNOR2_X1 U9415 ( .A(n7758), .B(n7759), .ZN(n7760) );
  OAI222_X1 U9416 ( .A1(n9863), .A2(n8544), .B1(n9865), .B2(n8038), .C1(n7760), 
        .C2(n9869), .ZN(n9924) );
  NAND2_X1 U9417 ( .A1(n9924), .A2(n9872), .ZN(n7764) );
  OAI22_X1 U9418 ( .A1(n9872), .A2(n7761), .B1(n8042), .B2(n9860), .ZN(n7762)
         );
  AOI21_X1 U9419 ( .B1(n8524), .B2(n9926), .A(n7762), .ZN(n7763) );
  OAI211_X1 U9420 ( .C1(n8552), .C2(n9923), .A(n7764), .B(n7763), .ZN(P2_U3221) );
  INV_X1 U9421 ( .A(n7765), .ZN(n7767) );
  OAI222_X1 U9422 ( .A1(P2_U3151), .A2(n5921), .B1(n7962), .B2(n7767), .C1(
        n7766), .C2(n8679), .ZN(P2_U3270) );
  OAI222_X1 U9423 ( .A1(n7768), .A2(P1_U3086), .B1(n7925), .B2(n7767), .C1(
        n10015), .C2(n9616), .ZN(P1_U3330) );
  OAI222_X1 U9424 ( .A1(P2_U3151), .A2(n5920), .B1(n7962), .B2(n7770), .C1(
        n7769), .C2(n8679), .ZN(P2_U3271) );
  AOI21_X1 U9425 ( .B1(n7773), .B2(n7772), .A(n7771), .ZN(n7781) );
  AOI22_X1 U9426 ( .A1(n8813), .A2(n9141), .B1(n8850), .B2(n9139), .ZN(n7776)
         );
  INV_X1 U9427 ( .A(n7774), .ZN(n7775) );
  OAI211_X1 U9428 ( .C1(n8858), .C2(n7777), .A(n7776), .B(n7775), .ZN(n7778)
         );
  AOI21_X1 U9429 ( .B1(n7779), .B2(n8864), .A(n7778), .ZN(n7780) );
  OAI21_X1 U9430 ( .B1(n7781), .B2(n8866), .A(n7780), .ZN(P1_U3221) );
  INV_X1 U9431 ( .A(n7782), .ZN(n7785) );
  OAI222_X1 U9432 ( .A1(P2_U3151), .A2(n7784), .B1(n7962), .B2(n7785), .C1(
        n7783), .C2(n8679), .ZN(P2_U3269) );
  OAI222_X1 U9433 ( .A1(n7786), .A2(P1_U3086), .B1(n7925), .B2(n7785), .C1(
        n10008), .C2(n9616), .ZN(P1_U3329) );
  AOI21_X1 U9434 ( .B1(n7794), .B2(n7788), .A(n8212), .ZN(n7804) );
  AND2_X1 U9435 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8113) );
  AOI21_X1 U9436 ( .B1(n7790), .B2(n7793), .A(n8206), .ZN(n7791) );
  NOR2_X1 U9437 ( .A1(n9844), .A2(n7791), .ZN(n7792) );
  AOI211_X1 U9438 ( .C1(n8216), .C2(n9819), .A(n8113), .B(n7792), .ZN(n7803)
         );
  MUX2_X1 U9439 ( .A(n7794), .B(n7793), .S(n8334), .Z(n8217) );
  XOR2_X1 U9440 ( .A(n8216), .B(n8217), .Z(n7800) );
  OR2_X1 U9441 ( .A1(n7796), .A2(n7795), .ZN(n7798) );
  NAND2_X1 U9442 ( .A1(n7798), .A2(n7797), .ZN(n7799) );
  NAND2_X1 U9443 ( .A1(n7800), .A2(n7799), .ZN(n8218) );
  OAI21_X1 U9444 ( .B1(n7800), .B2(n7799), .A(n8218), .ZN(n7801) );
  AOI22_X1 U9445 ( .A1(n9850), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(n9821), .B2(
        n7801), .ZN(n7802) );
  OAI211_X1 U9446 ( .C1(n7804), .C2(n9846), .A(n7803), .B(n7802), .ZN(P2_U3195) );
  XNOR2_X1 U9447 ( .A(n7805), .B(n7806), .ZN(n9624) );
  XNOR2_X1 U9448 ( .A(n7807), .B(n7806), .ZN(n7808) );
  OAI222_X1 U9449 ( .A1(n9863), .A2(n8529), .B1(n9865), .B2(n8137), .C1(n7808), 
        .C2(n9869), .ZN(n9626) );
  OAI22_X1 U9450 ( .A1(n9623), .A2(n9858), .B1(n8115), .B2(n9860), .ZN(n7809)
         );
  OAI21_X1 U9451 ( .B1(n9626), .B2(n7809), .A(n9872), .ZN(n7811) );
  NAND2_X1 U9452 ( .A1(n9874), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7810) );
  OAI211_X1 U9453 ( .C1(n8552), .C2(n9624), .A(n7811), .B(n7810), .ZN(P2_U3220) );
  INV_X1 U9454 ( .A(n8675), .ZN(n7812) );
  OAI222_X1 U9455 ( .A1(n9616), .A2(n7894), .B1(P1_U3086), .B2(n6525), .C1(
        n7925), .C2(n7812), .ZN(P1_U3327) );
  XNOR2_X1 U9456 ( .A(n8561), .B(n7847), .ZN(n7866) );
  XNOR2_X1 U9457 ( .A(n7866), .B(n8378), .ZN(n7970) );
  XNOR2_X1 U9458 ( .A(n7813), .B(n4526), .ZN(n7864) );
  INV_X1 U9459 ( .A(n7864), .ZN(n7814) );
  NAND2_X1 U9460 ( .A1(n7814), .A2(n7863), .ZN(n7968) );
  INV_X1 U9461 ( .A(n7815), .ZN(n7816) );
  XNOR2_X1 U9462 ( .A(n4526), .B(n9910), .ZN(n7993) );
  XNOR2_X1 U9463 ( .A(n7847), .B(n7820), .ZN(n8132) );
  OAI21_X1 U9464 ( .B1(n7993), .B2(n8036), .A(n8132), .ZN(n7826) );
  NAND3_X1 U9465 ( .A1(n4526), .A2(n9910), .A3(n8036), .ZN(n7821) );
  OAI211_X1 U9466 ( .C1(n4526), .C2(n8195), .A(n7821), .B(n7820), .ZN(n7824)
         );
  NAND3_X1 U9467 ( .A1(n7069), .A2(n8036), .A3(n7997), .ZN(n7822) );
  OAI211_X1 U9468 ( .C1(n7069), .C2(n8195), .A(n7822), .B(n4421), .ZN(n7823)
         );
  XNOR2_X1 U9469 ( .A(n4526), .B(n9926), .ZN(n7827) );
  XNOR2_X1 U9470 ( .A(n7827), .B(n8194), .ZN(n8039) );
  AOI21_X1 U9471 ( .B1(n7824), .B2(n7823), .A(n8039), .ZN(n7825) );
  XNOR2_X1 U9472 ( .A(n8117), .B(n7069), .ZN(n7828) );
  NAND2_X1 U9473 ( .A1(n7828), .A2(n8544), .ZN(n7831) );
  OAI21_X1 U9474 ( .B1(n7828), .B2(n8544), .A(n7831), .ZN(n8110) );
  NAND2_X1 U9475 ( .A1(n7830), .A2(n7829), .ZN(n8108) );
  NAND2_X1 U9476 ( .A1(n8108), .A2(n7831), .ZN(n7977) );
  XNOR2_X1 U9477 ( .A(n9622), .B(n4526), .ZN(n7832) );
  XNOR2_X1 U9478 ( .A(n7832), .B(n8529), .ZN(n7978) );
  NAND2_X1 U9479 ( .A1(n7977), .A2(n7978), .ZN(n8165) );
  XNOR2_X1 U9480 ( .A(n8533), .B(n7847), .ZN(n7834) );
  XNOR2_X1 U9481 ( .A(n7834), .B(n8191), .ZN(n8166) );
  NOR2_X1 U9482 ( .A1(n7832), .A2(n8192), .ZN(n8167) );
  NOR2_X1 U9483 ( .A1(n8166), .A2(n8167), .ZN(n7833) );
  NAND2_X1 U9484 ( .A1(n8165), .A2(n7833), .ZN(n8169) );
  NAND2_X1 U9485 ( .A1(n7834), .A2(n8191), .ZN(n7835) );
  NAND2_X1 U9486 ( .A1(n8169), .A2(n7835), .ZN(n8064) );
  XNOR2_X1 U9487 ( .A(n8609), .B(n4526), .ZN(n7836) );
  XNOR2_X1 U9488 ( .A(n7836), .B(n8530), .ZN(n8063) );
  NAND2_X1 U9489 ( .A1(n7836), .A2(n8501), .ZN(n7837) );
  XNOR2_X1 U9490 ( .A(n8660), .B(n7069), .ZN(n7839) );
  NAND2_X1 U9491 ( .A1(n7839), .A2(n8514), .ZN(n7840) );
  OAI21_X1 U9492 ( .B1(n7839), .B2(n8514), .A(n7840), .ZN(n8077) );
  XNOR2_X1 U9493 ( .A(n8599), .B(n4526), .ZN(n7841) );
  XNOR2_X1 U9494 ( .A(n7841), .B(n8078), .ZN(n8148) );
  NAND2_X2 U9495 ( .A1(n8147), .A2(n8148), .ZN(n8146) );
  XNOR2_X1 U9496 ( .A(n8477), .B(n4526), .ZN(n7844) );
  XNOR2_X1 U9497 ( .A(n7844), .B(n8484), .ZN(n8016) );
  NOR2_X1 U9498 ( .A1(n7841), .A2(n8498), .ZN(n8017) );
  NOR2_X1 U9499 ( .A1(n8016), .A2(n8017), .ZN(n7842) );
  NAND2_X2 U9500 ( .A1(n8146), .A2(n7842), .ZN(n8098) );
  XNOR2_X1 U9501 ( .A(n8094), .B(n4526), .ZN(n7843) );
  NOR2_X1 U9502 ( .A1(n7843), .A2(n8472), .ZN(n7845) );
  AOI21_X1 U9503 ( .B1(n8472), .B2(n7843), .A(n7845), .ZN(n8096) );
  NAND2_X1 U9504 ( .A1(n7844), .A2(n8484), .ZN(n8097) );
  INV_X1 U9505 ( .A(n7845), .ZN(n7846) );
  XNOR2_X1 U9506 ( .A(n8024), .B(n4526), .ZN(n7848) );
  XNOR2_X1 U9507 ( .A(n7848), .B(n8464), .ZN(n8027) );
  NAND2_X1 U9508 ( .A1(n8026), .A2(n8027), .ZN(n8025) );
  XNOR2_X1 U9509 ( .A(n8646), .B(n7847), .ZN(n7850) );
  XNOR2_X1 U9510 ( .A(n7850), .B(n8189), .ZN(n8121) );
  NOR2_X1 U9511 ( .A1(n7848), .A2(n8190), .ZN(n8122) );
  NOR2_X1 U9512 ( .A1(n8121), .A2(n8122), .ZN(n7849) );
  NAND2_X1 U9513 ( .A1(n8025), .A2(n7849), .ZN(n8124) );
  NAND2_X1 U9514 ( .A1(n7850), .A2(n8189), .ZN(n7851) );
  NAND2_X1 U9515 ( .A1(n8124), .A2(n7851), .ZN(n7853) );
  XNOR2_X1 U9516 ( .A(n8420), .B(n4526), .ZN(n7852) );
  NAND2_X1 U9517 ( .A1(n7986), .A2(n8084), .ZN(n7857) );
  XNOR2_X1 U9518 ( .A(n8398), .B(n4526), .ZN(n7854) );
  NAND2_X1 U9519 ( .A1(n7854), .A2(n8417), .ZN(n8053) );
  INV_X1 U9520 ( .A(n7854), .ZN(n7855) );
  NAND2_X1 U9521 ( .A1(n7855), .A2(n8388), .ZN(n7856) );
  NAND2_X1 U9522 ( .A1(n7857), .A2(n8085), .ZN(n8052) );
  NAND2_X1 U9523 ( .A1(n8052), .A2(n8053), .ZN(n7861) );
  XNOR2_X1 U9524 ( .A(n8051), .B(n7069), .ZN(n7858) );
  NAND2_X1 U9525 ( .A1(n7858), .A2(n8402), .ZN(n7862) );
  INV_X1 U9526 ( .A(n7858), .ZN(n7859) );
  NAND2_X1 U9527 ( .A1(n7859), .A2(n8188), .ZN(n7860) );
  NAND2_X1 U9528 ( .A1(n7861), .A2(n8054), .ZN(n8056) );
  XNOR2_X1 U9529 ( .A(n7864), .B(n7863), .ZN(n8158) );
  XOR2_X1 U9530 ( .A(n4526), .B(n7867), .Z(n7868) );
  AOI22_X1 U9531 ( .A1(n8172), .A2(n8186), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7870) );
  NAND2_X1 U9532 ( .A1(n8179), .A2(n8360), .ZN(n7869) );
  OAI211_X1 U9533 ( .C1(n7871), .C2(n8175), .A(n7870), .B(n7869), .ZN(n7872)
         );
  AOI21_X1 U9534 ( .B1(n7873), .B2(n8177), .A(n7872), .ZN(n7874) );
  OAI21_X1 U9535 ( .B1(n7875), .B2(n8119), .A(n7874), .ZN(P2_U3160) );
  NOR2_X1 U9536 ( .A1(n8807), .A2(n9462), .ZN(n7876) );
  INV_X1 U9537 ( .A(n9452), .ZN(n9642) );
  INV_X1 U9538 ( .A(n9459), .ZN(n8756) );
  NAND2_X1 U9539 ( .A1(n9429), .A2(n9440), .ZN(n9088) );
  NAND2_X1 U9540 ( .A1(n8919), .A2(n9088), .ZN(n9416) );
  NAND2_X1 U9541 ( .A1(n7910), .A2(n9422), .ZN(n7879) );
  INV_X1 U9542 ( .A(n9135), .ZN(n9394) );
  NAND2_X1 U9543 ( .A1(n9524), .A2(n8795), .ZN(n8942) );
  NAND2_X1 U9544 ( .A1(n9521), .A2(n9344), .ZN(n7887) );
  INV_X1 U9545 ( .A(n9344), .ZN(n8947) );
  NAND2_X1 U9546 ( .A1(n9580), .A2(n9256), .ZN(n7892) );
  INV_X1 U9547 ( .A(n9256), .ZN(n9297) );
  NAND2_X1 U9548 ( .A1(n9263), .A2(n9275), .ZN(n7893) );
  NAND2_X1 U9549 ( .A1(n9245), .A2(n9257), .ZN(n8957) );
  NAND2_X1 U9550 ( .A1(n8675), .A2(n8877), .ZN(n7896) );
  OR2_X1 U9551 ( .A1(n8880), .A2(n7894), .ZN(n7895) );
  NOR2_X1 U9552 ( .A1(n9489), .A2(n9240), .ZN(n7897) );
  INV_X1 U9553 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9612) );
  OR2_X1 U9554 ( .A1(n8880), .A2(n9612), .ZN(n7898) );
  INV_X1 U9555 ( .A(n7900), .ZN(n7906) );
  INV_X1 U9556 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7903) );
  NAND2_X1 U9557 ( .A1(n7915), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U9558 ( .A1(n8870), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7901) );
  OAI211_X1 U9559 ( .C1(n8871), .C2(n7903), .A(n7902), .B(n7901), .ZN(n7904)
         );
  AOI21_X1 U9560 ( .B1(n7906), .B2(n6070), .A(n7904), .ZN(n7957) );
  NAND2_X1 U9561 ( .A1(n9483), .A2(n7957), .ZN(n9008) );
  INV_X1 U9562 ( .A(n9429), .ZN(n9636) );
  NAND2_X1 U9563 ( .A1(n9447), .A2(n9636), .ZN(n9425) );
  NOR2_X2 U9564 ( .A1(n9406), .A2(n9542), .ZN(n9395) );
  AND2_X2 U9565 ( .A1(n9395), .A2(n9592), .ZN(n9368) );
  OR2_X2 U9566 ( .A1(n9303), .A2(n9510), .ZN(n9289) );
  AOI211_X1 U9567 ( .C1(n9483), .C2(n7951), .A(n9549), .B(n9231), .ZN(n9482)
         );
  INV_X1 U9568 ( .A(n9483), .ZN(n7908) );
  AOI22_X1 U9569 ( .A1(n7906), .A2(n9736), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n4419), .ZN(n7907) );
  OAI21_X1 U9570 ( .B1(n7908), .B2(n9741), .A(n7907), .ZN(n7922) );
  NAND2_X1 U9571 ( .A1(n9473), .A2(n8861), .ZN(n9084) );
  NAND2_X1 U9572 ( .A1(n8920), .A2(n9084), .ZN(n9457) );
  OR2_X1 U9573 ( .A1(n9452), .A2(n8756), .ZN(n8918) );
  NAND2_X1 U9574 ( .A1(n9452), .A2(n8756), .ZN(n9415) );
  AND2_X1 U9575 ( .A1(n9088), .A2(n9415), .ZN(n9090) );
  NAND2_X1 U9576 ( .A1(n9435), .A2(n9090), .ZN(n9420) );
  NAND2_X1 U9577 ( .A1(n9420), .A2(n8919), .ZN(n9403) );
  OR2_X1 U9578 ( .A1(n7910), .A2(n9392), .ZN(n8927) );
  NAND2_X1 U9579 ( .A1(n7910), .A2(n9392), .ZN(n8933) );
  NAND2_X1 U9580 ( .A1(n9403), .A2(n9402), .ZN(n7911) );
  NAND2_X1 U9581 ( .A1(n7911), .A2(n8927), .ZN(n9389) );
  OR2_X1 U9582 ( .A1(n9542), .A2(n7880), .ZN(n8935) );
  NAND2_X1 U9583 ( .A1(n9542), .A2(n7880), .ZN(n8934) );
  NAND2_X1 U9584 ( .A1(n8935), .A2(n8934), .ZN(n9390) );
  NAND2_X1 U9585 ( .A1(n9387), .A2(n8934), .ZN(n9376) );
  OR2_X1 U9586 ( .A1(n9370), .A2(n9394), .ZN(n8936) );
  NAND2_X1 U9587 ( .A1(n9370), .A2(n9394), .ZN(n9096) );
  XNOR2_X1 U9588 ( .A(n9360), .B(n8930), .ZN(n9351) );
  AND2_X1 U9589 ( .A1(n9588), .A2(n9380), .ZN(n9340) );
  NOR2_X1 U9590 ( .A1(n9339), .A2(n9340), .ZN(n7912) );
  XNOR2_X1 U9591 ( .A(n9521), .B(n9344), .ZN(n9319) );
  OR2_X1 U9592 ( .A1(n9514), .A2(n8771), .ZN(n8949) );
  NAND2_X1 U9593 ( .A1(n9514), .A2(n8771), .ZN(n8981) );
  NAND2_X1 U9594 ( .A1(n8949), .A2(n8981), .ZN(n9308) );
  NOR2_X1 U9595 ( .A1(n9521), .A2(n8947), .ZN(n9309) );
  NOR2_X1 U9596 ( .A1(n9308), .A2(n9309), .ZN(n7913) );
  XNOR2_X1 U9597 ( .A(n9510), .B(n8952), .ZN(n9287) );
  OR2_X1 U9598 ( .A1(n9263), .A2(n8744), .ZN(n8990) );
  NAND2_X1 U9599 ( .A1(n9263), .A2(n8744), .ZN(n8965) );
  NAND2_X1 U9600 ( .A1(n9252), .A2(n8965), .ZN(n9237) );
  NAND2_X1 U9601 ( .A1(n9237), .A2(n9238), .ZN(n9236) );
  INV_X1 U9602 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n7918) );
  NAND2_X1 U9603 ( .A1(n7915), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7917) );
  NAND2_X1 U9604 ( .A1(n8870), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7916) );
  OAI211_X1 U9605 ( .C1(n8871), .C2(n7918), .A(n7917), .B(n7916), .ZN(n9132)
         );
  AND2_X1 U9606 ( .A1(n7919), .A2(P1_B_REG_SCAN_IN), .ZN(n7920) );
  NOR2_X1 U9607 ( .A1(n9439), .A2(n7920), .ZN(n9225) );
  NOR2_X1 U9608 ( .A1(n9485), .A2(n4419), .ZN(n7921) );
  OAI21_X1 U9609 ( .B1(n9487), .B2(n9433), .A(n7923), .ZN(P1_U3356) );
  INV_X1 U9610 ( .A(n8878), .ZN(n7961) );
  OAI222_X1 U9611 ( .A1(n9616), .A2(n8879), .B1(n7925), .B2(n7961), .C1(n7924), 
        .C2(P1_U3086), .ZN(P1_U3325) );
  NAND2_X1 U9612 ( .A1(n9489), .A2(n7926), .ZN(n7929) );
  NAND2_X1 U9613 ( .A1(n9240), .A2(n7927), .ZN(n7928) );
  NAND2_X1 U9614 ( .A1(n7929), .A2(n7928), .ZN(n7930) );
  XNOR2_X1 U9615 ( .A(n7930), .B(n6136), .ZN(n7933) );
  AOI22_X1 U9616 ( .A1(n9489), .A2(n7931), .B1(n7926), .B2(n9240), .ZN(n7932)
         );
  XNOR2_X1 U9617 ( .A(n7933), .B(n7932), .ZN(n7941) );
  INV_X1 U9618 ( .A(n7941), .ZN(n7934) );
  NAND2_X1 U9619 ( .A1(n7934), .A2(n8817), .ZN(n7947) );
  OR2_X1 U9620 ( .A1(n7936), .A2(n7935), .ZN(n7940) );
  NAND4_X1 U9621 ( .A1(n7946), .A2(n8817), .A3(n7941), .A4(n7940), .ZN(n7945)
         );
  NAND2_X1 U9622 ( .A1(n9134), .A2(n8813), .ZN(n7939) );
  INV_X1 U9623 ( .A(n7937), .ZN(n7953) );
  AOI22_X1 U9624 ( .A1(n7953), .A2(n8847), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n7938) );
  OAI211_X1 U9625 ( .C1(n7957), .C2(n8859), .A(n7939), .B(n7938), .ZN(n7943)
         );
  NOR3_X1 U9626 ( .A1(n7941), .A2(n8866), .A3(n7940), .ZN(n7942) );
  AOI211_X1 U9627 ( .C1(n9489), .C2(n8864), .A(n7943), .B(n7942), .ZN(n7944)
         );
  OAI211_X1 U9628 ( .C1(n7947), .C2(n7946), .A(n7945), .B(n7944), .ZN(P1_U3220) );
  INV_X1 U9629 ( .A(n8979), .ZN(n7948) );
  XNOR2_X1 U9630 ( .A(n7950), .B(n7949), .ZN(n9488) );
  INV_X1 U9631 ( .A(n9243), .ZN(n7952) );
  AOI21_X1 U9632 ( .B1(n9489), .B2(n7952), .A(n4710), .ZN(n9490) );
  AOI22_X1 U9633 ( .A1(n7953), .A2(n9736), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n4419), .ZN(n7954) );
  OAI21_X1 U9634 ( .B1(n7955), .B2(n9741), .A(n7954), .ZN(n7959) );
  XOR2_X1 U9635 ( .A(n9044), .B(n7956), .Z(n7958) );
  INV_X1 U9636 ( .A(n7957), .ZN(n9133) );
  INV_X1 U9637 ( .A(n7965), .ZN(n9613) );
  OAI222_X1 U9638 ( .A1(n8679), .A2(n7966), .B1(n7962), .B2(n9613), .C1(n8334), 
        .C2(P2_U3151), .ZN(P2_U3268) );
  OAI222_X1 U9639 ( .A1(n8679), .A2(n7967), .B1(n7962), .B2(n9611), .C1(n5229), 
        .C2(P2_U3151), .ZN(P2_U3266) );
  AND2_X1 U9640 ( .A1(n8156), .A2(n7968), .ZN(n7971) );
  OAI211_X1 U9641 ( .C1(n7971), .C2(n7970), .A(n8170), .B(n7969), .ZN(n7976)
         );
  AOI22_X1 U9642 ( .A1(n8172), .A2(n8389), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7972) );
  OAI21_X1 U9643 ( .B1(n7973), .B2(n8175), .A(n7972), .ZN(n7974) );
  AOI21_X1 U9644 ( .B1(n8373), .B2(n8179), .A(n7974), .ZN(n7975) );
  OAI211_X1 U9645 ( .C1(n5906), .C2(n8164), .A(n7976), .B(n7975), .ZN(P2_U3154) );
  OAI21_X1 U9646 ( .B1(n7978), .B2(n7977), .A(n8165), .ZN(n7979) );
  NAND2_X1 U9647 ( .A1(n7979), .A2(n8170), .ZN(n7985) );
  INV_X1 U9648 ( .A(n8546), .ZN(n7983) );
  INV_X1 U9649 ( .A(n9622), .ZN(n8547) );
  NOR2_X1 U9650 ( .A1(n8547), .A2(n8164), .ZN(n7982) );
  NAND2_X1 U9651 ( .A1(n8172), .A2(n8193), .ZN(n7980) );
  NAND2_X1 U9652 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n8222) );
  OAI211_X1 U9653 ( .C1(n8545), .C2(n8175), .A(n7980), .B(n8222), .ZN(n7981)
         );
  AOI211_X1 U9654 ( .C1(n7983), .C2(n8179), .A(n7982), .B(n7981), .ZN(n7984)
         );
  NAND2_X1 U9655 ( .A1(n7985), .A2(n7984), .ZN(P2_U3155) );
  INV_X1 U9656 ( .A(n7986), .ZN(n8087) );
  AOI21_X1 U9657 ( .B1(n8431), .B2(n7987), .A(n8087), .ZN(n7992) );
  AOI22_X1 U9658 ( .A1(n8102), .A2(n8388), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7989) );
  NAND2_X1 U9659 ( .A1(n8179), .A2(n8421), .ZN(n7988) );
  OAI211_X1 U9660 ( .C1(n8104), .C2(n8451), .A(n7989), .B(n7988), .ZN(n7990)
         );
  AOI21_X1 U9661 ( .B1(n8420), .B2(n8177), .A(n7990), .ZN(n7991) );
  OAI21_X1 U9662 ( .B1(n7992), .B2(n8119), .A(n7991), .ZN(P2_U3156) );
  INV_X1 U9663 ( .A(n7993), .ZN(n7995) );
  XNOR2_X1 U9664 ( .A(n8034), .B(n8196), .ZN(n7994) );
  NOR2_X1 U9665 ( .A1(n7994), .A2(n7995), .ZN(n8035) );
  AOI21_X1 U9666 ( .B1(n7995), .B2(n7994), .A(n8035), .ZN(n8005) );
  AOI21_X1 U9667 ( .B1(n8172), .B2(n8197), .A(n7996), .ZN(n8003) );
  NAND2_X1 U9668 ( .A1(n8177), .A2(n7997), .ZN(n8002) );
  INV_X1 U9669 ( .A(n7998), .ZN(n7999) );
  NAND2_X1 U9670 ( .A1(n8179), .A2(n7999), .ZN(n8001) );
  NAND2_X1 U9671 ( .A1(n8102), .A2(n8195), .ZN(n8000) );
  AND4_X1 U9672 ( .A1(n8003), .A2(n8002), .A3(n8001), .A4(n8000), .ZN(n8004)
         );
  OAI21_X1 U9673 ( .B1(n8005), .B2(n8119), .A(n8004), .ZN(P2_U3157) );
  OAI21_X1 U9674 ( .B1(n8009), .B2(n8008), .A(n8007), .ZN(n8010) );
  NAND3_X1 U9675 ( .A1(n5014), .A2(n8170), .A3(n8010), .ZN(n8015) );
  AOI22_X1 U9676 ( .A1(n8172), .A2(n8204), .B1(n8011), .B2(n8177), .ZN(n8014)
         );
  MUX2_X1 U9677 ( .A(n8150), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n8013) );
  NAND2_X1 U9678 ( .A1(n8102), .A2(n8202), .ZN(n8012) );
  NAND4_X1 U9679 ( .A1(n8015), .A2(n8014), .A3(n8013), .A4(n8012), .ZN(
        P2_U3158) );
  INV_X1 U9680 ( .A(n8477), .ZN(n8598) );
  INV_X1 U9681 ( .A(n8146), .ZN(n8018) );
  OAI21_X1 U9682 ( .B1(n8018), .B2(n8017), .A(n8016), .ZN(n8019) );
  NAND3_X1 U9683 ( .A1(n8019), .A2(n8170), .A3(n8098), .ZN(n8023) );
  NAND2_X1 U9684 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8339) );
  OAI21_X1 U9685 ( .B1(n8175), .B2(n8450), .A(n8339), .ZN(n8021) );
  NOR2_X1 U9686 ( .A1(n8150), .A2(n8474), .ZN(n8020) );
  AOI211_X1 U9687 ( .C1(n8172), .C2(n8498), .A(n8021), .B(n8020), .ZN(n8022)
         );
  OAI211_X1 U9688 ( .C1(n8598), .C2(n8164), .A(n8023), .B(n8022), .ZN(P2_U3159) );
  INV_X1 U9689 ( .A(n8024), .ZN(n8651) );
  OAI21_X1 U9690 ( .B1(n8027), .B2(n8026), .A(n8025), .ZN(n8028) );
  NAND2_X1 U9691 ( .A1(n8028), .A2(n8170), .ZN(n8033) );
  INV_X1 U9692 ( .A(n8029), .ZN(n8452) );
  AOI22_X1 U9693 ( .A1(n8102), .A2(n8189), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8030) );
  OAI21_X1 U9694 ( .B1(n8450), .B2(n8104), .A(n8030), .ZN(n8031) );
  AOI21_X1 U9695 ( .B1(n8452), .B2(n8179), .A(n8031), .ZN(n8032) );
  OAI211_X1 U9696 ( .C1(n8651), .C2(n8164), .A(n8033), .B(n8032), .ZN(P2_U3163) );
  INV_X1 U9697 ( .A(n8034), .ZN(n8037) );
  AOI21_X1 U9698 ( .B1(n8037), .B2(n8036), .A(n8035), .ZN(n8133) );
  NAND2_X1 U9699 ( .A1(n8133), .A2(n8132), .ZN(n8131) );
  OAI21_X1 U9700 ( .B1(n8038), .B2(n8132), .A(n8131), .ZN(n8040) );
  XNOR2_X1 U9701 ( .A(n8040), .B(n8039), .ZN(n8049) );
  AOI21_X1 U9702 ( .B1(n8172), .B2(n8195), .A(n8041), .ZN(n8047) );
  NAND2_X1 U9703 ( .A1(n8177), .A2(n9926), .ZN(n8046) );
  INV_X1 U9704 ( .A(n8042), .ZN(n8043) );
  NAND2_X1 U9705 ( .A1(n8179), .A2(n8043), .ZN(n8045) );
  NAND2_X1 U9706 ( .A1(n8102), .A2(n8193), .ZN(n8044) );
  NAND4_X1 U9707 ( .A1(n8047), .A2(n8046), .A3(n8045), .A4(n8044), .ZN(n8048)
         );
  AOI21_X1 U9708 ( .B1(n8049), .B2(n8170), .A(n8048), .ZN(n8050) );
  INV_X1 U9709 ( .A(n8050), .ZN(P2_U3164) );
  INV_X1 U9710 ( .A(n8051), .ZN(n8635) );
  INV_X1 U9711 ( .A(n8052), .ZN(n8088) );
  INV_X1 U9712 ( .A(n8053), .ZN(n8055) );
  NOR3_X1 U9713 ( .A1(n8088), .A2(n8055), .A3(n8054), .ZN(n8058) );
  INV_X1 U9714 ( .A(n8056), .ZN(n8057) );
  OAI21_X1 U9715 ( .B1(n8058), .B2(n8057), .A(n8170), .ZN(n8062) );
  AOI22_X1 U9716 ( .A1(n8102), .A2(n8389), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8059) );
  OAI21_X1 U9717 ( .B1(n8417), .B2(n8104), .A(n8059), .ZN(n8060) );
  AOI21_X1 U9718 ( .B1(n8393), .B2(n8179), .A(n8060), .ZN(n8061) );
  OAI211_X1 U9719 ( .C1(n8635), .C2(n8164), .A(n8062), .B(n8061), .ZN(P2_U3165) );
  XOR2_X1 U9720 ( .A(n8064), .B(n8063), .Z(n8072) );
  NAND2_X1 U9721 ( .A1(n8609), .A2(n8177), .ZN(n8070) );
  INV_X1 U9722 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8065) );
  NOR2_X1 U9723 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8065), .ZN(n8265) );
  AOI21_X1 U9724 ( .B1(n8172), .B2(n8191), .A(n8265), .ZN(n8069) );
  INV_X1 U9725 ( .A(n8517), .ZN(n8066) );
  NAND2_X1 U9726 ( .A1(n8179), .A2(n8066), .ZN(n8068) );
  NAND2_X1 U9727 ( .A1(n8102), .A2(n8483), .ZN(n8067) );
  NAND4_X1 U9728 ( .A1(n8070), .A2(n8069), .A3(n8068), .A4(n8067), .ZN(n8071)
         );
  AOI21_X1 U9729 ( .B1(n8072), .B2(n8170), .A(n8071), .ZN(n8073) );
  INV_X1 U9730 ( .A(n8073), .ZN(P2_U3166) );
  INV_X1 U9731 ( .A(n8075), .ZN(n8076) );
  AOI21_X1 U9732 ( .B1(n8077), .B2(n8074), .A(n8076), .ZN(n8083) );
  AND2_X1 U9733 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8282) );
  NOR2_X1 U9734 ( .A1(n8175), .A2(n8078), .ZN(n8079) );
  AOI211_X1 U9735 ( .C1(n8172), .C2(n8501), .A(n8282), .B(n8079), .ZN(n8080)
         );
  OAI21_X1 U9736 ( .B1(n8504), .B2(n8150), .A(n8080), .ZN(n8081) );
  AOI21_X1 U9737 ( .B1(n8660), .B2(n8177), .A(n8081), .ZN(n8082) );
  OAI21_X1 U9738 ( .B1(n8083), .B2(n8119), .A(n8082), .ZN(P2_U3168) );
  INV_X1 U9739 ( .A(n8084), .ZN(n8086) );
  NOR3_X1 U9740 ( .A1(n8087), .A2(n8086), .A3(n8085), .ZN(n8089) );
  OAI21_X1 U9741 ( .B1(n8089), .B2(n8088), .A(n8170), .ZN(n8093) );
  AOI22_X1 U9742 ( .A1(n8102), .A2(n8188), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8090) );
  OAI21_X1 U9743 ( .B1(n8401), .B2(n8104), .A(n8090), .ZN(n8091) );
  AOI21_X1 U9744 ( .B1(n8407), .B2(n8179), .A(n8091), .ZN(n8092) );
  OAI211_X1 U9745 ( .C1(n8398), .C2(n8164), .A(n8093), .B(n8092), .ZN(P2_U3169) );
  INV_X1 U9746 ( .A(n8094), .ZN(n8655) );
  INV_X1 U9747 ( .A(n8095), .ZN(n8100) );
  AOI21_X1 U9748 ( .B1(n8098), .B2(n8097), .A(n8096), .ZN(n8099) );
  OAI21_X1 U9749 ( .B1(n8100), .B2(n8099), .A(n8170), .ZN(n8107) );
  INV_X1 U9750 ( .A(n8101), .ZN(n8465) );
  AOI22_X1 U9751 ( .A1(n8102), .A2(n8190), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8103) );
  OAI21_X1 U9752 ( .B1(n8463), .B2(n8104), .A(n8103), .ZN(n8105) );
  AOI21_X1 U9753 ( .B1(n8465), .B2(n8179), .A(n8105), .ZN(n8106) );
  OAI211_X1 U9754 ( .C1(n8655), .C2(n8164), .A(n8107), .B(n8106), .ZN(P2_U3173) );
  INV_X1 U9755 ( .A(n8108), .ZN(n8109) );
  AOI21_X1 U9756 ( .B1(n8111), .B2(n8110), .A(n8109), .ZN(n8120) );
  NOR2_X1 U9757 ( .A1(n8175), .A2(n8529), .ZN(n8112) );
  AOI211_X1 U9758 ( .C1(n8172), .C2(n8194), .A(n8113), .B(n8112), .ZN(n8114)
         );
  OAI21_X1 U9759 ( .B1(n8115), .B2(n8150), .A(n8114), .ZN(n8116) );
  AOI21_X1 U9760 ( .B1(n8117), .B2(n8177), .A(n8116), .ZN(n8118) );
  OAI21_X1 U9761 ( .B1(n8120), .B2(n8119), .A(n8118), .ZN(P2_U3174) );
  INV_X1 U9762 ( .A(n8646), .ZN(n8130) );
  INV_X1 U9763 ( .A(n8025), .ZN(n8123) );
  OAI21_X1 U9764 ( .B1(n8123), .B2(n8122), .A(n8121), .ZN(n8125) );
  NAND3_X1 U9765 ( .A1(n8125), .A2(n8170), .A3(n8124), .ZN(n8129) );
  AOI22_X1 U9766 ( .A1(n8172), .A2(n8190), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8126) );
  OAI21_X1 U9767 ( .B1(n8401), .B2(n8175), .A(n8126), .ZN(n8127) );
  AOI21_X1 U9768 ( .B1(n8435), .B2(n8179), .A(n8127), .ZN(n8128) );
  OAI211_X1 U9769 ( .C1(n8130), .C2(n8164), .A(n8129), .B(n8128), .ZN(P2_U3175) );
  OAI211_X1 U9770 ( .C1(n8133), .C2(n8132), .A(n8131), .B(n8170), .ZN(n8145)
         );
  NAND2_X1 U9771 ( .A1(n8172), .A2(n8196), .ZN(n8136) );
  INV_X1 U9772 ( .A(n8134), .ZN(n8135) );
  OAI211_X1 U9773 ( .C1(n8137), .C2(n8175), .A(n8136), .B(n8135), .ZN(n8138)
         );
  INV_X1 U9774 ( .A(n8138), .ZN(n8144) );
  NAND2_X1 U9775 ( .A1(n8177), .A2(n8139), .ZN(n8143) );
  INV_X1 U9776 ( .A(n8140), .ZN(n8141) );
  NAND2_X1 U9777 ( .A1(n8179), .A2(n8141), .ZN(n8142) );
  NAND4_X1 U9778 ( .A1(n8145), .A2(n8144), .A3(n8143), .A4(n8142), .ZN(
        P2_U3176) );
  INV_X1 U9779 ( .A(n8599), .ZN(n8155) );
  OAI21_X1 U9780 ( .B1(n8148), .B2(n8147), .A(n8146), .ZN(n8149) );
  NAND2_X1 U9781 ( .A1(n8149), .A2(n8170), .ZN(n8154) );
  NAND2_X1 U9782 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8317) );
  OAI21_X1 U9783 ( .B1(n8175), .B2(n8463), .A(n8317), .ZN(n8152) );
  NOR2_X1 U9784 ( .A1(n8150), .A2(n8486), .ZN(n8151) );
  AOI211_X1 U9785 ( .C1(n8172), .C2(n8483), .A(n8152), .B(n8151), .ZN(n8153)
         );
  OAI211_X1 U9786 ( .C1(n8155), .C2(n8164), .A(n8154), .B(n8153), .ZN(P2_U3178) );
  OAI21_X1 U9787 ( .B1(n8158), .B2(n8157), .A(n8156), .ZN(n8159) );
  NAND2_X1 U9788 ( .A1(n8159), .A2(n8170), .ZN(n8163) );
  AOI22_X1 U9789 ( .A1(n8172), .A2(n8188), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8160) );
  OAI21_X1 U9790 ( .B1(n8378), .B2(n8175), .A(n8160), .ZN(n8161) );
  AOI21_X1 U9791 ( .B1(n8381), .B2(n8179), .A(n8161), .ZN(n8162) );
  OAI211_X1 U9792 ( .C1(n8631), .C2(n8164), .A(n8163), .B(n8162), .ZN(P2_U3180) );
  INV_X1 U9793 ( .A(n8165), .ZN(n8168) );
  OAI21_X1 U9794 ( .B1(n8168), .B2(n8167), .A(n8166), .ZN(n8171) );
  NAND3_X1 U9795 ( .A1(n8171), .A2(n8170), .A3(n8169), .ZN(n8183) );
  NAND2_X1 U9796 ( .A1(n8172), .A2(n8192), .ZN(n8174) );
  NOR2_X1 U9797 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5210), .ZN(n8245) );
  INV_X1 U9798 ( .A(n8245), .ZN(n8173) );
  OAI211_X1 U9799 ( .C1(n8530), .C2(n8175), .A(n8174), .B(n8173), .ZN(n8176)
         );
  INV_X1 U9800 ( .A(n8176), .ZN(n8182) );
  NAND2_X1 U9801 ( .A1(n8533), .A2(n8177), .ZN(n8181) );
  INV_X1 U9802 ( .A(n8535), .ZN(n8178) );
  NAND2_X1 U9803 ( .A1(n8179), .A2(n8178), .ZN(n8180) );
  NAND4_X1 U9804 ( .A1(n8183), .A2(n8182), .A3(n8181), .A4(n8180), .ZN(
        P2_U3181) );
  MUX2_X1 U9805 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8184), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9806 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8185), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9807 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8369), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9808 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8186), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9809 ( .A(n8389), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8187), .Z(
        P2_U3517) );
  MUX2_X1 U9810 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8188), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9811 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8388), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9812 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8431), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U9813 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8189), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9814 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8190), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9815 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8472), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9816 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8484), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9817 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8498), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9818 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8483), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9819 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8501), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9820 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8191), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9821 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8192), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9822 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8193), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9823 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8194), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U9824 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8195), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9825 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8196), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U9826 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8197), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U9827 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8198), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U9828 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8199), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U9829 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8200), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U9830 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8201), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U9831 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8202), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U9832 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8203), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U9833 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8204), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U9834 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n5860), .S(P2_U3893), .Z(
        P2_U3492) );
  NOR2_X1 U9835 ( .A1(n8216), .A2(n8205), .ZN(n8207) );
  MUX2_X1 U9836 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8208), .S(n8231), .Z(n8209)
         );
  AOI21_X1 U9837 ( .B1(n4494), .B2(n8209), .A(n8242), .ZN(n8230) );
  NOR2_X1 U9838 ( .A1(n8216), .A2(n8210), .ZN(n8211) );
  INV_X1 U9839 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8213) );
  AOI22_X1 U9840 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8231), .B1(n8243), .B2(
        n8213), .ZN(n8214) );
  AOI21_X1 U9841 ( .B1(n4467), .B2(n8214), .A(n8233), .ZN(n8215) );
  NOR2_X1 U9842 ( .A1(n8215), .A2(n9846), .ZN(n8228) );
  INV_X1 U9843 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8226) );
  NAND2_X1 U9844 ( .A1(n8217), .A2(n8216), .ZN(n8219) );
  NAND2_X1 U9845 ( .A1(n8219), .A2(n8218), .ZN(n8221) );
  MUX2_X1 U9846 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8334), .Z(n8236) );
  XNOR2_X1 U9847 ( .A(n8236), .B(n8231), .ZN(n8220) );
  NAND2_X1 U9848 ( .A1(n8220), .A2(n8221), .ZN(n8237) );
  OAI21_X1 U9849 ( .B1(n8221), .B2(n8220), .A(n8237), .ZN(n8224) );
  OAI21_X1 U9850 ( .B1(n9855), .B2(n8243), .A(n8222), .ZN(n8223) );
  AOI21_X1 U9851 ( .B1(n9821), .B2(n8224), .A(n8223), .ZN(n8225) );
  OAI21_X1 U9852 ( .B1(n8341), .B2(n8226), .A(n8225), .ZN(n8227) );
  NOR2_X1 U9853 ( .A1(n8228), .A2(n8227), .ZN(n8229) );
  OAI21_X1 U9854 ( .B1(n8230), .B2(n9844), .A(n8229), .ZN(P2_U3196) );
  NOR2_X1 U9855 ( .A1(n8231), .A2(n8213), .ZN(n8232) );
  AOI21_X1 U9856 ( .B1(n8235), .B2(n8536), .A(n8255), .ZN(n8253) );
  MUX2_X1 U9857 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8334), .Z(n8268) );
  XNOR2_X1 U9858 ( .A(n8268), .B(n8246), .ZN(n8240) );
  OR2_X1 U9859 ( .A1(n8236), .A2(n8243), .ZN(n8238) );
  NAND2_X1 U9860 ( .A1(n8238), .A2(n8237), .ZN(n8239) );
  NAND2_X1 U9861 ( .A1(n8240), .A2(n8239), .ZN(n8269) );
  OAI21_X1 U9862 ( .B1(n8240), .B2(n8239), .A(n8269), .ZN(n8251) );
  NOR2_X1 U9863 ( .A1(n8341), .A2(n8241), .ZN(n8250) );
  XNOR2_X1 U9864 ( .A(n8258), .B(n8246), .ZN(n8244) );
  AOI21_X1 U9865 ( .B1(n8615), .B2(n8244), .A(n8259), .ZN(n8248) );
  AOI21_X1 U9866 ( .B1(n9819), .B2(n8246), .A(n8245), .ZN(n8247) );
  OAI21_X1 U9867 ( .B1(n8248), .B2(n9844), .A(n8247), .ZN(n8249) );
  AOI211_X1 U9868 ( .C1(n9821), .C2(n8251), .A(n8250), .B(n8249), .ZN(n8252)
         );
  OAI21_X1 U9869 ( .B1(n8253), .B2(n9846), .A(n8252), .ZN(P2_U3197) );
  INV_X1 U9870 ( .A(n8254), .ZN(n8256) );
  AOI22_X1 U9871 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8266), .B1(n8285), .B2(
        n8518), .ZN(n8257) );
  AOI21_X1 U9872 ( .B1(n4469), .B2(n8257), .A(n8277), .ZN(n8276) );
  INV_X1 U9873 ( .A(n8258), .ZN(n8260) );
  XNOR2_X1 U9874 ( .A(n8266), .B(n8261), .ZN(n8262) );
  AOI21_X1 U9875 ( .B1(n4466), .B2(n8262), .A(n8279), .ZN(n8263) );
  NOR2_X1 U9876 ( .A1(n8263), .A2(n9844), .ZN(n8264) );
  AOI211_X1 U9877 ( .C1(n8266), .C2(n9819), .A(n8265), .B(n8264), .ZN(n8275)
         );
  MUX2_X1 U9878 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8334), .Z(n8286) );
  XNOR2_X1 U9879 ( .A(n8286), .B(n8266), .ZN(n8272) );
  OR2_X1 U9880 ( .A1(n8268), .A2(n8267), .ZN(n8270) );
  NAND2_X1 U9881 ( .A1(n8270), .A2(n8269), .ZN(n8271) );
  NAND2_X1 U9882 ( .A1(n8272), .A2(n8271), .ZN(n8287) );
  OAI21_X1 U9883 ( .B1(n8272), .B2(n8271), .A(n8287), .ZN(n8273) );
  AOI22_X1 U9884 ( .A1(n9850), .A2(P2_ADDR_REG_16__SCAN_IN), .B1(n9821), .B2(
        n8273), .ZN(n8274) );
  OAI211_X1 U9885 ( .C1(n8276), .C2(n9846), .A(n8275), .B(n8274), .ZN(P2_U3198) );
  AOI21_X1 U9886 ( .B1(n8505), .B2(n8278), .A(n8296), .ZN(n8294) );
  XNOR2_X1 U9887 ( .A(n8307), .B(n8300), .ZN(n8280) );
  AOI211_X1 U9888 ( .C1(n8307), .C2(n9819), .A(n8282), .B(n8281), .ZN(n8293)
         );
  MUX2_X1 U9889 ( .A(n8505), .B(n8283), .S(n8334), .Z(n8306) );
  XNOR2_X1 U9890 ( .A(n8284), .B(n8306), .ZN(n8290) );
  OR2_X1 U9891 ( .A1(n8286), .A2(n8285), .ZN(n8288) );
  NAND2_X1 U9892 ( .A1(n8288), .A2(n8287), .ZN(n8289) );
  NAND2_X1 U9893 ( .A1(n8290), .A2(n8289), .ZN(n8308) );
  OAI21_X1 U9894 ( .B1(n8290), .B2(n8289), .A(n8308), .ZN(n8291) );
  AOI22_X1 U9895 ( .A1(n9850), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(n9821), .B2(
        n8291), .ZN(n8292) );
  OAI211_X1 U9896 ( .C1(n8294), .C2(n9846), .A(n8293), .B(n8292), .ZN(P2_U3199) );
  NOR2_X1 U9897 ( .A1(n8307), .A2(n8295), .ZN(n8297) );
  NAND2_X1 U9898 ( .A1(n8303), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8324) );
  OAI21_X1 U9899 ( .B1(n8303), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8324), .ZN(
        n8298) );
  AOI21_X1 U9900 ( .B1(n8299), .B2(n8298), .A(n8326), .ZN(n8323) );
  NOR2_X1 U9901 ( .A1(n8307), .A2(n8300), .ZN(n8302) );
  NAND2_X1 U9902 ( .A1(n8303), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8342) );
  OAI21_X1 U9903 ( .B1(n8303), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8342), .ZN(
        n8304) );
  AOI21_X1 U9904 ( .B1(n4463), .B2(n8304), .A(n8344), .ZN(n8305) );
  NOR2_X1 U9905 ( .A1(n8305), .A2(n9844), .ZN(n8321) );
  NAND2_X1 U9906 ( .A1(n8307), .A2(n8306), .ZN(n8309) );
  NAND2_X1 U9907 ( .A1(n8309), .A2(n8308), .ZN(n8311) );
  INV_X1 U9908 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8487) );
  MUX2_X1 U9909 ( .A(n8487), .B(n10233), .S(n8334), .Z(n8310) );
  OR2_X1 U9910 ( .A1(n8311), .A2(n8310), .ZN(n8329) );
  NAND2_X1 U9911 ( .A1(n8311), .A2(n8310), .ZN(n8330) );
  AND2_X1 U9912 ( .A1(n8329), .A2(n8330), .ZN(n8313) );
  INV_X1 U9913 ( .A(n8313), .ZN(n8312) );
  NAND2_X1 U9914 ( .A1(n9821), .A2(n8312), .ZN(n8316) );
  AOI21_X1 U9915 ( .B1(P2_U3893), .B2(n8313), .A(n9819), .ZN(n8315) );
  MUX2_X1 U9916 ( .A(n8316), .B(n8315), .S(n8328), .Z(n8318) );
  OAI211_X1 U9917 ( .C1(n8319), .C2(n8341), .A(n8318), .B(n8317), .ZN(n8320)
         );
  NOR2_X1 U9918 ( .A1(n8321), .A2(n8320), .ZN(n8322) );
  OAI21_X1 U9919 ( .B1(n8323), .B2(n9846), .A(n8322), .ZN(P2_U3200) );
  INV_X1 U9920 ( .A(n8324), .ZN(n8325) );
  MUX2_X1 U9921 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8475), .S(n8333), .Z(n8335)
         );
  XNOR2_X1 U9922 ( .A(n8327), .B(n8335), .ZN(n8350) );
  NAND2_X1 U9923 ( .A1(n8329), .A2(n8328), .ZN(n8331) );
  NAND2_X1 U9924 ( .A1(n8331), .A2(n8330), .ZN(n8337) );
  XNOR2_X1 U9925 ( .A(n8333), .B(n8332), .ZN(n8345) );
  MUX2_X1 U9926 ( .A(n8335), .B(n8345), .S(n8334), .Z(n8336) );
  XNOR2_X1 U9927 ( .A(n8337), .B(n8336), .ZN(n8348) );
  NAND2_X1 U9928 ( .A1(n9819), .A2(n8338), .ZN(n8340) );
  OAI211_X1 U9929 ( .C1(n8341), .C2(n4763), .A(n8340), .B(n8339), .ZN(n8347)
         );
  INV_X1 U9930 ( .A(n8342), .ZN(n8343) );
  OAI21_X1 U9931 ( .B1(n9846), .B2(n8350), .A(n8349), .ZN(P2_U3201) );
  INV_X1 U9932 ( .A(n8555), .ZN(n8621) );
  INV_X1 U9933 ( .A(n8351), .ZN(n8352) );
  OR2_X1 U9934 ( .A1(n8353), .A2(n8352), .ZN(n8619) );
  OAI21_X1 U9935 ( .B1(n9874), .B2(n8619), .A(n8354), .ZN(n8356) );
  AOI21_X1 U9936 ( .B1(n9874), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8356), .ZN(
        n8355) );
  OAI21_X1 U9937 ( .B1(n8621), .B2(n8534), .A(n8355), .ZN(P2_U3202) );
  AOI21_X1 U9938 ( .B1(n9874), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8356), .ZN(
        n8357) );
  OAI21_X1 U9939 ( .B1(n8358), .B2(n8534), .A(n8357), .ZN(P2_U3203) );
  INV_X1 U9940 ( .A(n8359), .ZN(n8366) );
  AOI22_X1 U9941 ( .A1(n9874), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8466), .B2(
        n8360), .ZN(n8361) );
  OAI21_X1 U9942 ( .B1(n8362), .B2(n8534), .A(n8361), .ZN(n8363) );
  AOI21_X1 U9943 ( .B1(n8364), .B2(n8539), .A(n8363), .ZN(n8365) );
  OAI21_X1 U9944 ( .B1(n8366), .B2(n9874), .A(n8365), .ZN(P2_U3205) );
  XNOR2_X1 U9945 ( .A(n8368), .B(n8367), .ZN(n8370) );
  XNOR2_X1 U9946 ( .A(n8372), .B(n8371), .ZN(n8562) );
  AOI22_X1 U9947 ( .A1(n9874), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8466), .B2(
        n8373), .ZN(n8374) );
  OAI21_X1 U9948 ( .B1(n5906), .B2(n8534), .A(n8374), .ZN(n8375) );
  AOI21_X1 U9949 ( .B1(n8562), .B2(n8539), .A(n8375), .ZN(n8376) );
  OAI21_X1 U9950 ( .B1(n8564), .B2(n9874), .A(n8376), .ZN(P2_U3206) );
  INV_X1 U9951 ( .A(n8565), .ZN(n8385) );
  XNOR2_X1 U9952 ( .A(n8380), .B(n8379), .ZN(n8566) );
  AOI22_X1 U9953 ( .A1(n9874), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8466), .B2(
        n8381), .ZN(n8382) );
  OAI21_X1 U9954 ( .B1(n8631), .B2(n8534), .A(n8382), .ZN(n8383) );
  AOI21_X1 U9955 ( .B1(n8566), .B2(n8539), .A(n8383), .ZN(n8384) );
  OAI21_X1 U9956 ( .B1(n8385), .B2(n9874), .A(n8384), .ZN(P2_U3207) );
  NOR2_X1 U9957 ( .A1(n8635), .A2(n9858), .ZN(n8392) );
  OAI21_X1 U9958 ( .B1(n8387), .B2(n8394), .A(n8386), .ZN(n8390) );
  AOI222_X1 U9959 ( .A1(n8494), .A2(n8390), .B1(n8389), .B2(n8499), .C1(n8388), 
        .C2(n8500), .ZN(n8391) );
  INV_X1 U9960 ( .A(n8391), .ZN(n8568) );
  AOI211_X1 U9961 ( .C1(n8466), .C2(n8393), .A(n8392), .B(n8568), .ZN(n8397)
         );
  XNOR2_X1 U9962 ( .A(n8395), .B(n8394), .ZN(n8569) );
  AOI22_X1 U9963 ( .A1(n8569), .A2(n8539), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9874), .ZN(n8396) );
  OAI21_X1 U9964 ( .B1(n8397), .B2(n9874), .A(n8396), .ZN(P2_U3208) );
  NOR2_X1 U9965 ( .A1(n8398), .A2(n9858), .ZN(n8406) );
  XNOR2_X1 U9966 ( .A(n8400), .B(n8411), .ZN(n8404) );
  OAI22_X1 U9967 ( .A1(n8402), .A2(n9863), .B1(n8401), .B2(n9865), .ZN(n8403)
         );
  AOI21_X1 U9968 ( .B1(n8404), .B2(n8494), .A(n8403), .ZN(n8573) );
  INV_X1 U9969 ( .A(n8573), .ZN(n8405) );
  AOI211_X1 U9970 ( .C1(n8466), .C2(n8407), .A(n8406), .B(n8405), .ZN(n8414)
         );
  INV_X1 U9971 ( .A(n8408), .ZN(n8409) );
  OR2_X1 U9972 ( .A1(n8410), .A2(n8409), .ZN(n8412) );
  XNOR2_X1 U9973 ( .A(n8412), .B(n8411), .ZN(n8572) );
  AOI22_X1 U9974 ( .A1(n8572), .A2(n8539), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9874), .ZN(n8413) );
  OAI21_X1 U9975 ( .B1(n8414), .B2(n9874), .A(n8413), .ZN(P2_U3209) );
  XNOR2_X1 U9976 ( .A(n8415), .B(n8418), .ZN(n8416) );
  OAI222_X1 U9977 ( .A1(n9863), .A2(n8417), .B1(n9865), .B2(n8451), .C1(n9869), 
        .C2(n8416), .ZN(n8577) );
  INV_X1 U9978 ( .A(n8577), .ZN(n8425) );
  XNOR2_X1 U9979 ( .A(n8419), .B(n8418), .ZN(n8578) );
  INV_X1 U9980 ( .A(n8420), .ZN(n8643) );
  AOI22_X1 U9981 ( .A1(n9874), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8466), .B2(
        n8421), .ZN(n8422) );
  OAI21_X1 U9982 ( .B1(n8643), .B2(n8534), .A(n8422), .ZN(n8423) );
  AOI21_X1 U9983 ( .B1(n8578), .B2(n8539), .A(n8423), .ZN(n8424) );
  OAI21_X1 U9984 ( .B1(n8425), .B2(n9874), .A(n8424), .ZN(P2_U3210) );
  NAND3_X1 U9985 ( .A1(n8427), .A2(n8429), .A3(n8428), .ZN(n8430) );
  NAND2_X1 U9986 ( .A1(n8426), .A2(n8430), .ZN(n8434) );
  NAND2_X1 U9987 ( .A1(n8431), .A2(n8499), .ZN(n8432) );
  OAI21_X1 U9988 ( .B1(n8464), .B2(n9865), .A(n8432), .ZN(n8433) );
  AOI21_X1 U9989 ( .B1(n8434), .B2(n8494), .A(n8433), .ZN(n8582) );
  INV_X1 U9990 ( .A(n8435), .ZN(n8436) );
  OAI22_X1 U9991 ( .A1(n9872), .A2(n8437), .B1(n8436), .B2(n9860), .ZN(n8438)
         );
  AOI21_X1 U9992 ( .B1(n8646), .B2(n8524), .A(n8438), .ZN(n8442) );
  XNOR2_X1 U9993 ( .A(n8440), .B(n8439), .ZN(n8581) );
  NAND2_X1 U9994 ( .A1(n8581), .A2(n8539), .ZN(n8441) );
  OAI211_X1 U9995 ( .C1(n8582), .C2(n9874), .A(n8442), .B(n8441), .ZN(P2_U3211) );
  XOR2_X1 U9996 ( .A(n8443), .B(n8445), .Z(n8587) );
  INV_X1 U9997 ( .A(n8587), .ZN(n8456) );
  INV_X1 U9998 ( .A(n8445), .ZN(n8447) );
  NAND3_X1 U9999 ( .A1(n8458), .A2(n8447), .A3(n8446), .ZN(n8448) );
  AND2_X1 U10000 ( .A1(n8427), .A2(n8448), .ZN(n8449) );
  OAI222_X1 U10001 ( .A1(n9863), .A2(n8451), .B1(n9865), .B2(n8450), .C1(n9869), .C2(n8449), .ZN(n8586) );
  AOI22_X1 U10002 ( .A1(n9874), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8466), .B2(
        n8452), .ZN(n8453) );
  OAI21_X1 U10003 ( .B1(n8651), .B2(n8534), .A(n8453), .ZN(n8454) );
  AOI21_X1 U10004 ( .B1(n8586), .B2(n9872), .A(n8454), .ZN(n8455) );
  OAI21_X1 U10005 ( .B1(n8552), .B2(n8456), .A(n8455), .ZN(P2_U3212) );
  XOR2_X1 U10006 ( .A(n8461), .B(n8457), .Z(n8591) );
  INV_X1 U10007 ( .A(n8591), .ZN(n8470) );
  INV_X1 U10008 ( .A(n8458), .ZN(n8459) );
  AOI21_X1 U10009 ( .B1(n8461), .B2(n8460), .A(n8459), .ZN(n8462) );
  OAI222_X1 U10010 ( .A1(n9863), .A2(n8464), .B1(n9865), .B2(n8463), .C1(n9869), .C2(n8462), .ZN(n8590) );
  AOI22_X1 U10011 ( .A1(n9874), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8466), .B2(
        n8465), .ZN(n8467) );
  OAI21_X1 U10012 ( .B1(n8655), .B2(n8534), .A(n8467), .ZN(n8468) );
  AOI21_X1 U10013 ( .B1(n8590), .B2(n9872), .A(n8468), .ZN(n8469) );
  OAI21_X1 U10014 ( .B1(n8470), .B2(n8552), .A(n8469), .ZN(P2_U3213) );
  XNOR2_X1 U10015 ( .A(n8471), .B(n8478), .ZN(n8473) );
  AOI222_X1 U10016 ( .A1(n8494), .A2(n8473), .B1(n8472), .B2(n8499), .C1(n8498), .C2(n8500), .ZN(n8597) );
  OAI22_X1 U10017 ( .A1(n9872), .A2(n8475), .B1(n8474), .B2(n9860), .ZN(n8476)
         );
  AOI21_X1 U10018 ( .B1(n8477), .B2(n8524), .A(n8476), .ZN(n8481) );
  OR2_X1 U10019 ( .A1(n8479), .A2(n8478), .ZN(n8595) );
  NAND3_X1 U10020 ( .A1(n8595), .A2(n8594), .A3(n8539), .ZN(n8480) );
  OAI211_X1 U10021 ( .C1(n8597), .C2(n9874), .A(n8481), .B(n8480), .ZN(
        P2_U3214) );
  XNOR2_X1 U10022 ( .A(n8482), .B(n8489), .ZN(n8485) );
  AOI222_X1 U10023 ( .A1(n8494), .A2(n8485), .B1(n8484), .B2(n8499), .C1(n8483), .C2(n8500), .ZN(n8601) );
  OAI22_X1 U10024 ( .A1(n9872), .A2(n8487), .B1(n8486), .B2(n9860), .ZN(n8492)
         );
  OAI21_X1 U10025 ( .B1(n8490), .B2(n8489), .A(n8488), .ZN(n8602) );
  NOR2_X1 U10026 ( .A1(n8602), .A2(n8552), .ZN(n8491) );
  AOI211_X1 U10027 ( .C1(n8524), .C2(n8599), .A(n8492), .B(n8491), .ZN(n8493)
         );
  OAI21_X1 U10028 ( .B1(n9874), .B2(n8601), .A(n8493), .ZN(P2_U3215) );
  OAI211_X1 U10029 ( .C1(n8497), .C2(n8496), .A(n8495), .B(n8494), .ZN(n8503)
         );
  AOI22_X1 U10030 ( .A1(n8501), .A2(n8500), .B1(n8499), .B2(n8498), .ZN(n8502)
         );
  AND2_X1 U10031 ( .A1(n8503), .A2(n8502), .ZN(n8605) );
  OAI22_X1 U10032 ( .A1(n9872), .A2(n8505), .B1(n8504), .B2(n9860), .ZN(n8506)
         );
  AOI21_X1 U10033 ( .B1(n8660), .B2(n8524), .A(n8506), .ZN(n8510) );
  XNOR2_X1 U10034 ( .A(n8508), .B(n8507), .ZN(n8603) );
  NAND2_X1 U10035 ( .A1(n8603), .A2(n8539), .ZN(n8509) );
  OAI211_X1 U10036 ( .C1(n8605), .C2(n9874), .A(n8510), .B(n8509), .ZN(
        P2_U3216) );
  AOI21_X1 U10037 ( .B1(n8512), .B2(n8511), .A(n9869), .ZN(n8516) );
  OAI22_X1 U10038 ( .A1(n8545), .A2(n9865), .B1(n8514), .B2(n9863), .ZN(n8515)
         );
  AOI21_X1 U10039 ( .B1(n8516), .B2(n8513), .A(n8515), .ZN(n8611) );
  OAI22_X1 U10040 ( .A1(n9872), .A2(n8518), .B1(n8517), .B2(n9860), .ZN(n8523)
         );
  INV_X1 U10041 ( .A(n8519), .ZN(n8520) );
  AOI21_X1 U10042 ( .B1(n5890), .B2(n8521), .A(n8520), .ZN(n8612) );
  NOR2_X1 U10043 ( .A1(n8612), .A2(n8552), .ZN(n8522) );
  AOI211_X1 U10044 ( .C1(n8524), .C2(n8609), .A(n8523), .B(n8522), .ZN(n8525)
         );
  OAI21_X1 U10045 ( .B1(n9874), .B2(n8611), .A(n8525), .ZN(P2_U3217) );
  XNOR2_X1 U10046 ( .A(n8527), .B(n8526), .ZN(n8528) );
  OAI222_X1 U10047 ( .A1(n9863), .A2(n8530), .B1(n9865), .B2(n8529), .C1(n9869), .C2(n8528), .ZN(n8613) );
  INV_X1 U10048 ( .A(n8613), .ZN(n8541) );
  XNOR2_X1 U10049 ( .A(n8532), .B(n8531), .ZN(n8614) );
  INV_X1 U10050 ( .A(n8533), .ZN(n8668) );
  NOR2_X1 U10051 ( .A1(n8668), .A2(n8534), .ZN(n8538) );
  OAI22_X1 U10052 ( .A1(n9872), .A2(n8536), .B1(n8535), .B2(n9860), .ZN(n8537)
         );
  AOI211_X1 U10053 ( .C1(n8614), .C2(n8539), .A(n8538), .B(n8537), .ZN(n8540)
         );
  OAI21_X1 U10054 ( .B1(n8541), .B2(n9874), .A(n8540), .ZN(P2_U3218) );
  XOR2_X1 U10055 ( .A(n8551), .B(n8542), .Z(n8543) );
  OAI222_X1 U10056 ( .A1(n9863), .A2(n8545), .B1(n9865), .B2(n8544), .C1(n8543), .C2(n9869), .ZN(n9620) );
  OAI22_X1 U10057 ( .A1(n8547), .A2(n9858), .B1(n8546), .B2(n9860), .ZN(n8548)
         );
  OAI21_X1 U10058 ( .B1(n9620), .B2(n8548), .A(n9872), .ZN(n8554) );
  INV_X1 U10059 ( .A(n8549), .ZN(n9618) );
  NOR2_X1 U10060 ( .A1(n8550), .A2(n8551), .ZN(n9619) );
  OR3_X1 U10061 ( .A1(n9618), .A2(n9619), .A3(n8552), .ZN(n8553) );
  OAI211_X1 U10062 ( .C1(n9872), .C2(n8213), .A(n8554), .B(n8553), .ZN(
        P2_U3219) );
  NAND2_X1 U10063 ( .A1(n8555), .A2(n8607), .ZN(n8557) );
  INV_X1 U10064 ( .A(n8619), .ZN(n8556) );
  NAND2_X1 U10065 ( .A1(n8556), .A2(n9941), .ZN(n8558) );
  OAI211_X1 U10066 ( .C1(n9941), .C2(n5238), .A(n8557), .B(n8558), .ZN(
        P2_U3490) );
  INV_X1 U10067 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U10068 ( .A1(n8622), .A2(n8607), .ZN(n8559) );
  OAI211_X1 U10069 ( .C1(n9941), .C2(n8560), .A(n8559), .B(n8558), .ZN(
        P2_U3489) );
  AOI22_X1 U10070 ( .A1(n8562), .A2(n9920), .B1(n9927), .B2(n8561), .ZN(n8563)
         );
  MUX2_X1 U10071 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8627), .S(n9941), .Z(
        P2_U3486) );
  AOI21_X1 U10072 ( .B1(n8566), .B2(n9920), .A(n8565), .ZN(n8628) );
  MUX2_X1 U10073 ( .A(n10188), .B(n8628), .S(n9941), .Z(n8567) );
  OAI21_X1 U10074 ( .B1(n8631), .B2(n8617), .A(n8567), .ZN(P2_U3485) );
  INV_X1 U10075 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8570) );
  MUX2_X1 U10076 ( .A(n8570), .B(n8632), .S(n9941), .Z(n8571) );
  OAI21_X1 U10077 ( .B1(n8635), .B2(n8617), .A(n8571), .ZN(P2_U3484) );
  NAND2_X1 U10078 ( .A1(n8572), .A2(n9920), .ZN(n8574) );
  NAND2_X1 U10079 ( .A1(n8574), .A2(n8573), .ZN(n8636) );
  MUX2_X1 U10080 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8636), .S(n9941), .Z(n8575) );
  AOI21_X1 U10081 ( .B1(n8607), .B2(n8638), .A(n8575), .ZN(n8576) );
  INV_X1 U10082 ( .A(n8576), .ZN(P2_U3483) );
  INV_X1 U10083 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8579) );
  AOI21_X1 U10084 ( .B1(n9920), .B2(n8578), .A(n8577), .ZN(n8640) );
  MUX2_X1 U10085 ( .A(n8579), .B(n8640), .S(n9941), .Z(n8580) );
  OAI21_X1 U10086 ( .B1(n8643), .B2(n8617), .A(n8580), .ZN(P2_U3482) );
  NAND2_X1 U10087 ( .A1(n8581), .A2(n9920), .ZN(n8583) );
  NAND2_X1 U10088 ( .A1(n8583), .A2(n8582), .ZN(n8644) );
  MUX2_X1 U10089 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8644), .S(n9941), .Z(n8584) );
  AOI21_X1 U10090 ( .B1(n8607), .B2(n8646), .A(n8584), .ZN(n8585) );
  INV_X1 U10091 ( .A(n8585), .ZN(P2_U3481) );
  AOI21_X1 U10092 ( .B1(n8587), .B2(n9920), .A(n8586), .ZN(n8648) );
  MUX2_X1 U10093 ( .A(n8588), .B(n8648), .S(n9941), .Z(n8589) );
  OAI21_X1 U10094 ( .B1(n8651), .B2(n8617), .A(n8589), .ZN(P2_U3480) );
  AOI21_X1 U10095 ( .B1(n9920), .B2(n8591), .A(n8590), .ZN(n8652) );
  MUX2_X1 U10096 ( .A(n8592), .B(n8652), .S(n9941), .Z(n8593) );
  OAI21_X1 U10097 ( .B1(n8655), .B2(n8617), .A(n8593), .ZN(P2_U3479) );
  NAND3_X1 U10098 ( .A1(n8595), .A2(n9920), .A3(n8594), .ZN(n8596) );
  OAI211_X1 U10099 ( .C1(n8598), .C2(n9915), .A(n8597), .B(n8596), .ZN(n8656)
         );
  MUX2_X1 U10100 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8656), .S(n9941), .Z(
        P2_U3478) );
  NAND2_X1 U10101 ( .A1(n8599), .A2(n9927), .ZN(n8600) );
  OAI211_X1 U10102 ( .C1(n9922), .C2(n8602), .A(n8601), .B(n8600), .ZN(n8657)
         );
  MUX2_X1 U10103 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8657), .S(n9941), .Z(
        P2_U3477) );
  NAND2_X1 U10104 ( .A1(n8603), .A2(n9920), .ZN(n8604) );
  NAND2_X1 U10105 ( .A1(n8605), .A2(n8604), .ZN(n8658) );
  MUX2_X1 U10106 ( .A(n8658), .B(P2_REG1_REG_17__SCAN_IN), .S(n9939), .Z(n8606) );
  AOI21_X1 U10107 ( .B1(n8607), .B2(n8660), .A(n8606), .ZN(n8608) );
  INV_X1 U10108 ( .A(n8608), .ZN(P2_U3476) );
  NAND2_X1 U10109 ( .A1(n8609), .A2(n9927), .ZN(n8610) );
  OAI211_X1 U10110 ( .C1(n8612), .C2(n9922), .A(n8611), .B(n8610), .ZN(n8663)
         );
  MUX2_X1 U10111 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8663), .S(n9941), .Z(
        P2_U3475) );
  AOI21_X1 U10112 ( .B1(n9920), .B2(n8614), .A(n8613), .ZN(n8664) );
  MUX2_X1 U10113 ( .A(n8615), .B(n8664), .S(n9941), .Z(n8616) );
  OAI21_X1 U10114 ( .B1(n8668), .B2(n8617), .A(n8616), .ZN(P2_U3474) );
  MUX2_X1 U10115 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n8618), .S(n9941), .Z(
        P2_U3459) );
  NOR2_X1 U10116 ( .A1(n8619), .A2(n9929), .ZN(n8623) );
  AOI21_X1 U10117 ( .B1(P2_REG0_REG_31__SCAN_IN), .B2(n9929), .A(n8623), .ZN(
        n8620) );
  OAI21_X1 U10118 ( .B1(n8621), .B2(n8667), .A(n8620), .ZN(P2_U3458) );
  INV_X1 U10119 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8626) );
  INV_X1 U10120 ( .A(n8667), .ZN(n8661) );
  NAND2_X1 U10121 ( .A1(n8622), .A2(n8661), .ZN(n8625) );
  INV_X1 U10122 ( .A(n8623), .ZN(n8624) );
  OAI211_X1 U10123 ( .C1(n8626), .C2(n9928), .A(n8625), .B(n8624), .ZN(
        P2_U3457) );
  MUX2_X1 U10124 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8627), .S(n9928), .Z(
        P2_U3454) );
  INV_X1 U10125 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8629) );
  MUX2_X1 U10126 ( .A(n8629), .B(n8628), .S(n9928), .Z(n8630) );
  OAI21_X1 U10127 ( .B1(n8631), .B2(n8667), .A(n8630), .ZN(P2_U3453) );
  INV_X1 U10128 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8633) );
  MUX2_X1 U10129 ( .A(n8633), .B(n8632), .S(n9928), .Z(n8634) );
  OAI21_X1 U10130 ( .B1(n8635), .B2(n8667), .A(n8634), .ZN(P2_U3452) );
  MUX2_X1 U10131 ( .A(n8636), .B(P2_REG0_REG_24__SCAN_IN), .S(n9929), .Z(n8637) );
  AOI21_X1 U10132 ( .B1(n8661), .B2(n8638), .A(n8637), .ZN(n8639) );
  INV_X1 U10133 ( .A(n8639), .ZN(P2_U3451) );
  INV_X1 U10134 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8641) );
  MUX2_X1 U10135 ( .A(n8641), .B(n8640), .S(n9928), .Z(n8642) );
  OAI21_X1 U10136 ( .B1(n8643), .B2(n8667), .A(n8642), .ZN(P2_U3450) );
  MUX2_X1 U10137 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8644), .S(n9928), .Z(n8645) );
  AOI21_X1 U10138 ( .B1(n8661), .B2(n8646), .A(n8645), .ZN(n8647) );
  INV_X1 U10139 ( .A(n8647), .ZN(P2_U3449) );
  MUX2_X1 U10140 ( .A(n8649), .B(n8648), .S(n9928), .Z(n8650) );
  OAI21_X1 U10141 ( .B1(n8651), .B2(n8667), .A(n8650), .ZN(P2_U3448) );
  MUX2_X1 U10142 ( .A(n8653), .B(n8652), .S(n9928), .Z(n8654) );
  OAI21_X1 U10143 ( .B1(n8655), .B2(n8667), .A(n8654), .ZN(P2_U3447) );
  MUX2_X1 U10144 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8656), .S(n9928), .Z(
        P2_U3446) );
  MUX2_X1 U10145 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8657), .S(n9928), .Z(
        P2_U3444) );
  MUX2_X1 U10146 ( .A(n8658), .B(P2_REG0_REG_17__SCAN_IN), .S(n9929), .Z(n8659) );
  AOI21_X1 U10147 ( .B1(n8661), .B2(n8660), .A(n8659), .ZN(n8662) );
  INV_X1 U10148 ( .A(n8662), .ZN(P2_U3441) );
  MUX2_X1 U10149 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8663), .S(n9928), .Z(
        P2_U3438) );
  INV_X1 U10150 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8665) );
  MUX2_X1 U10151 ( .A(n8665), .B(n8664), .S(n9928), .Z(n8666) );
  OAI21_X1 U10152 ( .B1(n8668), .B2(n8667), .A(n8666), .ZN(P2_U3435) );
  NAND3_X1 U10153 ( .A1(n8670), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8672) );
  OAI22_X1 U10154 ( .A1(n8669), .A2(n8672), .B1(n8671), .B2(n8679), .ZN(n8673)
         );
  AOI21_X1 U10155 ( .B1(n9609), .B2(n4503), .A(n8673), .ZN(n8674) );
  INV_X1 U10156 ( .A(n8674), .ZN(P2_U3264) );
  NAND2_X1 U10157 ( .A1(n8675), .A2(n4503), .ZN(n8677) );
  OAI211_X1 U10158 ( .C1(n8679), .C2(n8678), .A(n8677), .B(n8676), .ZN(
        P2_U3267) );
  MUX2_X1 U10159 ( .A(n8680), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  XNOR2_X1 U10160 ( .A(n8683), .B(n8682), .ZN(n8684) );
  XNOR2_X1 U10161 ( .A(n8681), .B(n8684), .ZN(n8690) );
  OAI22_X1 U10162 ( .A1(n8858), .A2(n9469), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8685), .ZN(n8688) );
  INV_X1 U10163 ( .A(n8813), .ZN(n8860) );
  OAI22_X1 U10164 ( .A1(n8686), .A2(n8860), .B1(n8859), .B2(n8756), .ZN(n8687)
         );
  AOI211_X1 U10165 ( .C1(n9473), .C2(n8864), .A(n8688), .B(n8687), .ZN(n8689)
         );
  OAI21_X1 U10166 ( .B1(n8690), .B2(n8866), .A(n8689), .ZN(P1_U3215) );
  INV_X1 U10167 ( .A(n8691), .ZN(n8694) );
  INV_X1 U10168 ( .A(n8692), .ZN(n8812) );
  NAND2_X1 U10169 ( .A1(n8811), .A2(n8812), .ZN(n8810) );
  OAI21_X1 U10170 ( .B1(n8694), .B2(n8693), .A(n8810), .ZN(n8698) );
  XNOR2_X1 U10171 ( .A(n8696), .B(n8695), .ZN(n8697) );
  XNOR2_X1 U10172 ( .A(n8698), .B(n8697), .ZN(n8703) );
  OAI22_X1 U10173 ( .A1(n8858), .A2(n9305), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8699), .ZN(n8701) );
  OAI22_X1 U10174 ( .A1(n8952), .A2(n8859), .B1(n8947), .B2(n8860), .ZN(n8700)
         );
  AOI211_X1 U10175 ( .C1(n9514), .C2(n8864), .A(n8701), .B(n8700), .ZN(n8702)
         );
  OAI21_X1 U10176 ( .B1(n8703), .B2(n8866), .A(n8702), .ZN(P1_U3216) );
  XNOR2_X1 U10177 ( .A(n8821), .B(n8822), .ZN(n8706) );
  NOR2_X1 U10178 ( .A1(n8706), .A2(n8705), .ZN(n8820) );
  AOI21_X1 U10179 ( .B1(n8706), .B2(n8705), .A(n8820), .ZN(n8713) );
  AOI22_X1 U10180 ( .A1(n8813), .A2(n9139), .B1(n8850), .B2(n4957), .ZN(n8708)
         );
  NAND2_X1 U10181 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8707) );
  OAI211_X1 U10182 ( .C1(n8858), .C2(n8709), .A(n8708), .B(n8707), .ZN(n8710)
         );
  AOI21_X1 U10183 ( .B1(n8711), .B2(n8864), .A(n8710), .ZN(n8712) );
  OAI21_X1 U10184 ( .B1(n8713), .B2(n8866), .A(n8712), .ZN(P1_U3217) );
  INV_X1 U10185 ( .A(n8714), .ZN(n8718) );
  NAND2_X1 U10186 ( .A1(n5024), .A2(n8717), .ZN(n8716) );
  AOI22_X1 U10187 ( .A1(n8718), .A2(n8717), .B1(n8715), .B2(n8716), .ZN(n8723)
         );
  OAI22_X1 U10188 ( .A1(n8858), .A2(n9371), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8719), .ZN(n8721) );
  OAI22_X1 U10189 ( .A1(n7880), .A2(n8860), .B1(n8859), .B2(n8930), .ZN(n8720)
         );
  AOI211_X1 U10190 ( .C1(n9370), .C2(n8864), .A(n8721), .B(n8720), .ZN(n8722)
         );
  OAI21_X1 U10191 ( .B1(n8723), .B2(n8866), .A(n8722), .ZN(P1_U3219) );
  XOR2_X1 U10192 ( .A(n8725), .B(n8724), .Z(n8730) );
  OAI22_X1 U10193 ( .A1(n8858), .A2(n9335), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8726), .ZN(n8728) );
  OAI22_X1 U10194 ( .A1(n8930), .A2(n8860), .B1(n8859), .B2(n8947), .ZN(n8727)
         );
  AOI211_X1 U10195 ( .C1(n9524), .C2(n8864), .A(n8728), .B(n8727), .ZN(n8729)
         );
  OAI21_X1 U10196 ( .B1(n8730), .B2(n8866), .A(n8729), .ZN(P1_U3223) );
  XOR2_X1 U10197 ( .A(n8732), .B(n8731), .Z(n8740) );
  NAND2_X1 U10198 ( .A1(n8829), .A2(n8733), .ZN(n8734) );
  OAI211_X1 U10199 ( .C1(n8858), .C2(n8736), .A(n8735), .B(n8734), .ZN(n8737)
         );
  AOI21_X1 U10200 ( .B1(n8738), .B2(n8864), .A(n8737), .ZN(n8739) );
  OAI21_X1 U10201 ( .B1(n8740), .B2(n8866), .A(n8739), .ZN(P1_U3224) );
  XOR2_X1 U10202 ( .A(n8742), .B(n8741), .Z(n8748) );
  OAI22_X1 U10203 ( .A1(n9280), .A2(n8858), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8743), .ZN(n8746) );
  OAI22_X1 U10204 ( .A1(n8744), .A2(n8859), .B1(n8952), .B2(n8860), .ZN(n8745)
         );
  AOI211_X1 U10205 ( .C1(n9279), .C2(n8864), .A(n8746), .B(n8745), .ZN(n8747)
         );
  OAI21_X1 U10206 ( .B1(n8748), .B2(n8866), .A(n8747), .ZN(P1_U3225) );
  XNOR2_X1 U10207 ( .A(n8749), .B(n8750), .ZN(n8856) );
  NOR2_X1 U10208 ( .A1(n8856), .A2(n8855), .ZN(n8854) );
  AOI21_X1 U10209 ( .B1(n8750), .B2(n8749), .A(n8854), .ZN(n8754) );
  XNOR2_X1 U10210 ( .A(n8752), .B(n8751), .ZN(n8753) );
  XNOR2_X1 U10211 ( .A(n8754), .B(n8753), .ZN(n8760) );
  OAI22_X1 U10212 ( .A1(n8858), .A2(n9426), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8755), .ZN(n8758) );
  OAI22_X1 U10213 ( .A1(n8756), .A2(n8860), .B1(n8859), .B2(n9392), .ZN(n8757)
         );
  AOI211_X1 U10214 ( .C1(n9429), .C2(n8864), .A(n8758), .B(n8757), .ZN(n8759)
         );
  OAI21_X1 U10215 ( .B1(n8760), .B2(n8866), .A(n8759), .ZN(P1_U3226) );
  OAI211_X1 U10216 ( .C1(n8763), .C2(n8762), .A(n8761), .B(n8817), .ZN(n8768)
         );
  AND2_X1 U10217 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9173) );
  OR2_X1 U10218 ( .A1(n9440), .A2(n9393), .ZN(n8765) );
  NAND2_X1 U10219 ( .A1(n9379), .A2(n9460), .ZN(n8764) );
  AND2_X1 U10220 ( .A1(n8765), .A2(n8764), .ZN(n9404) );
  NOR2_X1 U10221 ( .A1(n8797), .A2(n9404), .ZN(n8766) );
  AOI211_X1 U10222 ( .C1(n8847), .C2(n9408), .A(n9173), .B(n8766), .ZN(n8767)
         );
  OAI211_X1 U10223 ( .C1(n9631), .C2(n8853), .A(n8768), .B(n8767), .ZN(
        P1_U3228) );
  XOR2_X1 U10224 ( .A(n8770), .B(n8769), .Z(n8775) );
  OAI22_X1 U10225 ( .A1(n9291), .A2(n8858), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10044), .ZN(n8773) );
  OAI22_X1 U10226 ( .A1(n9256), .A2(n8859), .B1(n8771), .B2(n8860), .ZN(n8772)
         );
  AOI211_X1 U10227 ( .C1(n9510), .C2(n8864), .A(n8773), .B(n8772), .ZN(n8774)
         );
  OAI21_X1 U10228 ( .B1(n8775), .B2(n8866), .A(n8774), .ZN(P1_U3229) );
  INV_X1 U10229 ( .A(n8776), .ZN(n8778) );
  NAND2_X1 U10230 ( .A1(n8778), .A2(n8777), .ZN(n8779) );
  XNOR2_X1 U10231 ( .A(n8780), .B(n8779), .ZN(n8788) );
  AOI21_X1 U10232 ( .B1(n8829), .B2(n8782), .A(n8781), .ZN(n8785) );
  NAND2_X1 U10233 ( .A1(n8847), .A2(n8783), .ZN(n8784) );
  OAI211_X1 U10234 ( .C1(n8786), .C2(n8853), .A(n8785), .B(n8784), .ZN(n8787)
         );
  AOI21_X1 U10235 ( .B1(n8788), .B2(n8817), .A(n8787), .ZN(n8789) );
  INV_X1 U10236 ( .A(n8789), .ZN(P1_U3231) );
  OAI21_X1 U10237 ( .B1(n8792), .B2(n8791), .A(n8790), .ZN(n8793) );
  NAND2_X1 U10238 ( .A1(n8793), .A2(n8817), .ZN(n8800) );
  INV_X1 U10239 ( .A(n8794), .ZN(n9361) );
  OAI22_X1 U10240 ( .A1(n8795), .A2(n9439), .B1(n9394), .B2(n9393), .ZN(n8796)
         );
  INV_X1 U10241 ( .A(n8796), .ZN(n9355) );
  OAI22_X1 U10242 ( .A1(n9355), .A2(n8797), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10016), .ZN(n8798) );
  AOI21_X1 U10243 ( .B1(n9361), .B2(n8847), .A(n8798), .ZN(n8799) );
  OAI211_X1 U10244 ( .C1(n9588), .C2(n8853), .A(n8800), .B(n8799), .ZN(
        P1_U3233) );
  XOR2_X1 U10245 ( .A(n8802), .B(n8801), .Z(n8809) );
  OAI22_X1 U10246 ( .A1(n8858), .A2(n8804), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8803), .ZN(n8806) );
  OAI22_X1 U10247 ( .A1(n8827), .A2(n8860), .B1(n8859), .B2(n8861), .ZN(n8805)
         );
  AOI211_X1 U10248 ( .C1(n8807), .C2(n8864), .A(n8806), .B(n8805), .ZN(n8808)
         );
  OAI21_X1 U10249 ( .B1(n8809), .B2(n8866), .A(n8808), .ZN(P1_U3234) );
  OAI21_X1 U10250 ( .B1(n8812), .B2(n8811), .A(n8810), .ZN(n8818) );
  AOI22_X1 U10251 ( .A1(n8847), .A2(n9327), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n8815) );
  AOI22_X1 U10252 ( .A1(n9322), .A2(n8850), .B1(n8813), .B2(n9321), .ZN(n8814)
         );
  OAI211_X1 U10253 ( .C1(n9330), .C2(n8853), .A(n8815), .B(n8814), .ZN(n8816)
         );
  AOI21_X1 U10254 ( .B1(n8818), .B2(n8817), .A(n8816), .ZN(n8819) );
  INV_X1 U10255 ( .A(n8819), .ZN(P1_U3235) );
  AOI21_X1 U10256 ( .B1(n8822), .B2(n8821), .A(n8820), .ZN(n8826) );
  XNOR2_X1 U10257 ( .A(n8824), .B(n8823), .ZN(n8825) );
  XNOR2_X1 U10258 ( .A(n8826), .B(n8825), .ZN(n8833) );
  OAI22_X1 U10259 ( .A1(n8828), .A2(n9393), .B1(n8827), .B2(n9439), .ZN(n9557)
         );
  AOI22_X1 U10260 ( .A1(n9557), .A2(n8829), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n8830) );
  OAI21_X1 U10261 ( .B1(n9692), .B2(n8858), .A(n8830), .ZN(n8831) );
  AOI21_X1 U10262 ( .B1(n4422), .B2(n8864), .A(n8831), .ZN(n8832) );
  OAI21_X1 U10263 ( .B1(n8833), .B2(n8866), .A(n8832), .ZN(P1_U3236) );
  XOR2_X1 U10264 ( .A(n8835), .B(n8834), .Z(n8836) );
  XNOR2_X1 U10265 ( .A(n8837), .B(n8836), .ZN(n8843) );
  INV_X1 U10266 ( .A(n9396), .ZN(n8839) );
  OAI22_X1 U10267 ( .A1(n8858), .A2(n8839), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8838), .ZN(n8841) );
  OAI22_X1 U10268 ( .A1(n9392), .A2(n8860), .B1(n8859), .B2(n9394), .ZN(n8840)
         );
  AOI211_X1 U10269 ( .C1(n9542), .C2(n8864), .A(n8841), .B(n8840), .ZN(n8842)
         );
  OAI21_X1 U10270 ( .B1(n8843), .B2(n8866), .A(n8842), .ZN(P1_U3238) );
  AOI22_X1 U10271 ( .A1(n9264), .A2(n8847), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n8848) );
  OAI21_X1 U10272 ( .B1(n9256), .B2(n8860), .A(n8848), .ZN(n8849) );
  AOI21_X1 U10273 ( .B1(n9134), .B2(n8850), .A(n8849), .ZN(n8851) );
  OAI211_X1 U10274 ( .C1(n9576), .C2(n8853), .A(n8852), .B(n8851), .ZN(
        P1_U3240) );
  AOI21_X1 U10275 ( .B1(n8856), .B2(n8855), .A(n8854), .ZN(n8867) );
  OAI22_X1 U10276 ( .A1(n8858), .A2(n9445), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8857), .ZN(n8863) );
  OAI22_X1 U10277 ( .A1(n8861), .A2(n8860), .B1(n8859), .B2(n9440), .ZN(n8862)
         );
  AOI211_X1 U10278 ( .C1(n9452), .C2(n8864), .A(n8863), .B(n8862), .ZN(n8865)
         );
  OAI21_X1 U10279 ( .B1(n8867), .B2(n8866), .A(n8865), .ZN(P1_U3241) );
  NAND2_X1 U10280 ( .A1(n4539), .A2(n9050), .ZN(n8970) );
  INV_X1 U10281 ( .A(n8970), .ZN(n8976) );
  NAND2_X1 U10282 ( .A1(n9609), .A2(n8877), .ZN(n8869) );
  OR2_X1 U10283 ( .A1(n8880), .A2(n9604), .ZN(n8868) );
  NAND2_X1 U10284 ( .A1(n8870), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8876) );
  INV_X1 U10285 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9478) );
  OR2_X1 U10286 ( .A1(n8871), .A2(n9478), .ZN(n8875) );
  INV_X1 U10287 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8872) );
  OR2_X1 U10288 ( .A1(n8873), .A2(n8872), .ZN(n8874) );
  AND3_X1 U10289 ( .A1(n8876), .A2(n8875), .A3(n8874), .ZN(n9227) );
  NAND2_X1 U10290 ( .A1(n8878), .A2(n8877), .ZN(n8882) );
  OR2_X1 U10291 ( .A1(n8880), .A2(n8879), .ZN(n8881) );
  INV_X1 U10292 ( .A(n9132), .ZN(n9007) );
  AND2_X1 U10293 ( .A1(n8883), .A2(n9023), .ZN(n8885) );
  INV_X1 U10294 ( .A(n8887), .ZN(n9071) );
  OAI211_X1 U10295 ( .C1(n8889), .C2(n9071), .A(n9024), .B(n8888), .ZN(n8891)
         );
  NAND2_X1 U10296 ( .A1(n8891), .A2(n8890), .ZN(n8893) );
  NAND2_X1 U10297 ( .A1(n8893), .A2(n4949), .ZN(n8898) );
  AND2_X1 U10298 ( .A1(n8895), .A2(n8894), .ZN(n8897) );
  AOI21_X1 U10299 ( .B1(n8898), .B2(n8897), .A(n8896), .ZN(n8899) );
  INV_X1 U10300 ( .A(n8900), .ZN(n8901) );
  OAI21_X1 U10301 ( .B1(n8907), .B2(n8901), .A(n9552), .ZN(n8902) );
  NAND2_X1 U10302 ( .A1(n8903), .A2(n8919), .ZN(n8904) );
  INV_X1 U10303 ( .A(n8919), .ZN(n9421) );
  OR2_X1 U10304 ( .A1(n9090), .A2(n9421), .ZN(n8905) );
  NAND3_X1 U10305 ( .A1(n8904), .A2(n8976), .A3(n8905), .ZN(n8925) );
  INV_X1 U10306 ( .A(n8905), .ZN(n8906) );
  NAND2_X1 U10307 ( .A1(n8906), .A2(n8970), .ZN(n8924) );
  INV_X1 U10308 ( .A(n8907), .ZN(n8909) );
  NAND2_X1 U10309 ( .A1(n8909), .A2(n8908), .ZN(n8911) );
  NAND2_X1 U10310 ( .A1(n8910), .A2(n9552), .ZN(n9075) );
  AOI21_X1 U10311 ( .B1(n8911), .B2(n9073), .A(n9075), .ZN(n8914) );
  NAND2_X1 U10312 ( .A1(n8913), .A2(n8912), .ZN(n9078) );
  OAI21_X1 U10313 ( .B1(n8914), .B2(n9078), .A(n9081), .ZN(n8916) );
  NAND2_X1 U10314 ( .A1(n8916), .A2(n8915), .ZN(n8917) );
  INV_X1 U10315 ( .A(n9457), .ZN(n9455) );
  NAND3_X1 U10316 ( .A1(n8917), .A2(n9455), .A3(n9082), .ZN(n8921) );
  AND2_X1 U10317 ( .A1(n8919), .A2(n8918), .ZN(n9087) );
  NAND4_X1 U10318 ( .A1(n8921), .A2(n9087), .A3(n8920), .A4(n8970), .ZN(n8923)
         );
  NAND4_X1 U10319 ( .A1(n9088), .A2(n9642), .A3(n8976), .A4(n9459), .ZN(n8922)
         );
  NAND4_X1 U10320 ( .A1(n8925), .A2(n8924), .A3(n8923), .A4(n8922), .ZN(n8926)
         );
  NAND2_X1 U10321 ( .A1(n8926), .A2(n9402), .ZN(n8937) );
  AND2_X1 U10322 ( .A1(n8935), .A2(n8927), .ZN(n9095) );
  NAND2_X1 U10323 ( .A1(n8937), .A2(n9095), .ZN(n8928) );
  NAND3_X1 U10324 ( .A1(n8928), .A2(n9096), .A3(n8934), .ZN(n8929) );
  INV_X1 U10325 ( .A(n9340), .ZN(n8939) );
  NAND3_X1 U10326 ( .A1(n8929), .A2(n8936), .A3(n8939), .ZN(n8931) );
  NAND2_X1 U10327 ( .A1(n9360), .A2(n8930), .ZN(n8938) );
  AND2_X1 U10328 ( .A1(n8942), .A2(n8938), .ZN(n8994) );
  NAND2_X1 U10329 ( .A1(n8931), .A2(n8994), .ZN(n8932) );
  NAND2_X1 U10330 ( .A1(n8932), .A2(n8995), .ZN(n8945) );
  AND2_X1 U10331 ( .A1(n8934), .A2(n8933), .ZN(n9092) );
  NAND2_X1 U10332 ( .A1(n8936), .A2(n8935), .ZN(n9097) );
  AOI21_X1 U10333 ( .B1(n8937), .B2(n9092), .A(n9097), .ZN(n8941) );
  NAND2_X1 U10334 ( .A1(n8938), .A2(n9096), .ZN(n8940) );
  AND2_X1 U10335 ( .A1(n8995), .A2(n8939), .ZN(n8988) );
  OAI21_X1 U10336 ( .B1(n8941), .B2(n8940), .A(n8988), .ZN(n8943) );
  NAND2_X1 U10337 ( .A1(n8943), .A2(n8942), .ZN(n8944) );
  INV_X1 U10338 ( .A(n9309), .ZN(n8946) );
  NAND2_X1 U10339 ( .A1(n8946), .A2(n8949), .ZN(n8982) );
  NAND2_X1 U10340 ( .A1(n9521), .A2(n8947), .ZN(n8948) );
  NAND2_X1 U10341 ( .A1(n8981), .A2(n8948), .ZN(n8993) );
  MUX2_X1 U10342 ( .A(n8982), .B(n8993), .S(n8970), .Z(n8951) );
  INV_X1 U10343 ( .A(n9287), .ZN(n9295) );
  MUX2_X1 U10344 ( .A(n8981), .B(n8949), .S(n8970), .Z(n8950) );
  NAND2_X1 U10345 ( .A1(n9510), .A2(n8952), .ZN(n8998) );
  MUX2_X1 U10346 ( .A(n8983), .B(n8998), .S(n8970), .Z(n8953) );
  INV_X1 U10347 ( .A(n9000), .ZN(n8954) );
  INV_X1 U10348 ( .A(n8965), .ZN(n9099) );
  AOI211_X1 U10349 ( .C1(n8987), .C2(n8963), .A(n8954), .B(n9099), .ZN(n8956)
         );
  INV_X1 U10350 ( .A(n8990), .ZN(n8955) );
  NOR2_X1 U10351 ( .A1(n8956), .A2(n8955), .ZN(n8961) );
  INV_X1 U10352 ( .A(n8957), .ZN(n8958) );
  NOR2_X1 U10353 ( .A1(n8959), .A2(n8958), .ZN(n8962) );
  NAND2_X1 U10354 ( .A1(n8962), .A2(n8970), .ZN(n8960) );
  INV_X1 U10355 ( .A(n8962), .ZN(n9005) );
  NAND3_X1 U10356 ( .A1(n9005), .A2(n8976), .A3(n8979), .ZN(n8969) );
  NAND2_X1 U10357 ( .A1(n8963), .A2(n9000), .ZN(n8964) );
  NAND3_X1 U10358 ( .A1(n8964), .A2(n8990), .A3(n8987), .ZN(n8966) );
  NAND2_X1 U10359 ( .A1(n8966), .A2(n8965), .ZN(n8967) );
  NAND4_X1 U10360 ( .A1(n8979), .A2(n8967), .A3(n8976), .A4(n8991), .ZN(n8968)
         );
  INV_X1 U10361 ( .A(n9227), .ZN(n9131) );
  AOI21_X1 U10362 ( .B1(n8976), .B2(n9053), .A(n9051), .ZN(n9130) );
  NOR2_X1 U10363 ( .A1(n9113), .A2(n4550), .ZN(n9123) );
  INV_X1 U10364 ( .A(n8977), .ZN(n8978) );
  OAI211_X1 U10365 ( .C1(n4728), .C2(n7035), .A(n9123), .B(n8978), .ZN(n9129)
         );
  AND2_X1 U10366 ( .A1(n8980), .A2(n8979), .ZN(n9057) );
  NAND2_X1 U10367 ( .A1(n8982), .A2(n8981), .ZN(n8984) );
  NAND2_X1 U10368 ( .A1(n8984), .A2(n8983), .ZN(n8985) );
  NAND2_X1 U10369 ( .A1(n8985), .A2(n8998), .ZN(n8986) );
  NAND2_X1 U10370 ( .A1(n8987), .A2(n8986), .ZN(n8992) );
  INV_X1 U10371 ( .A(n8988), .ZN(n8989) );
  NOR2_X1 U10372 ( .A1(n8992), .A2(n8989), .ZN(n9101) );
  AOI21_X1 U10373 ( .B1(n9101), .B2(n9352), .A(n9099), .ZN(n9006) );
  NAND2_X1 U10374 ( .A1(n8991), .A2(n8990), .ZN(n9102) );
  NAND2_X1 U10375 ( .A1(n8992), .A2(n9000), .ZN(n9002) );
  INV_X1 U10376 ( .A(n8993), .ZN(n8999) );
  INV_X1 U10377 ( .A(n8994), .ZN(n8996) );
  NAND2_X1 U10378 ( .A1(n8996), .A2(n8995), .ZN(n8997) );
  NAND4_X1 U10379 ( .A1(n9000), .A2(n8999), .A3(n8998), .A4(n8997), .ZN(n9001)
         );
  NAND2_X1 U10380 ( .A1(n9002), .A2(n9001), .ZN(n9003) );
  NOR2_X1 U10381 ( .A1(n9102), .A2(n9003), .ZN(n9004) );
  NOR2_X1 U10382 ( .A1(n9005), .A2(n9004), .ZN(n9058) );
  OAI21_X1 U10383 ( .B1(n9006), .B2(n9102), .A(n9058), .ZN(n9009) );
  NAND2_X1 U10384 ( .A1(n9223), .A2(n9007), .ZN(n9047) );
  NAND2_X1 U10385 ( .A1(n9047), .A2(n9008), .ZN(n9111) );
  AOI21_X1 U10386 ( .B1(n9057), .B2(n9009), .A(n9111), .ZN(n9010) );
  AOI21_X1 U10387 ( .B1(n4562), .B2(n9131), .A(n9010), .ZN(n9011) );
  AOI211_X1 U10388 ( .C1(n9227), .C2(n9223), .A(n9012), .B(n9011), .ZN(n9014)
         );
  NOR2_X1 U10389 ( .A1(n9014), .A2(n9013), .ZN(n9049) );
  INV_X1 U10390 ( .A(n9238), .ZN(n9043) );
  INV_X1 U10391 ( .A(n9319), .ZN(n9040) );
  INV_X1 U10392 ( .A(n9390), .ZN(n9037) );
  NOR2_X1 U10393 ( .A1(n9720), .A2(n4420), .ZN(n9019) );
  INV_X1 U10394 ( .A(n9015), .ZN(n9017) );
  NAND4_X1 U10395 ( .A1(n9019), .A2(n9018), .A3(n9017), .A4(n9016), .ZN(n9022)
         );
  NOR3_X1 U10396 ( .A1(n9022), .A2(n9021), .A3(n9020), .ZN(n9026) );
  NAND4_X1 U10397 ( .A1(n9026), .A2(n9025), .A3(n9024), .A4(n9023), .ZN(n9029)
         );
  NOR3_X1 U10398 ( .A1(n9029), .A2(n9028), .A3(n9027), .ZN(n9030) );
  NAND3_X1 U10399 ( .A1(n9031), .A2(n9551), .A3(n9030), .ZN(n9032) );
  NOR2_X1 U10400 ( .A1(n9033), .A2(n9032), .ZN(n9034) );
  NAND3_X1 U10401 ( .A1(n9443), .A2(n9455), .A3(n9034), .ZN(n9035) );
  NOR2_X1 U10402 ( .A1(n9416), .A2(n9035), .ZN(n9036) );
  NAND4_X1 U10403 ( .A1(n9377), .A2(n9037), .A3(n9402), .A4(n9036), .ZN(n9038)
         );
  OR3_X1 U10404 ( .A1(n9339), .A2(n9351), .A3(n9038), .ZN(n9039) );
  NOR3_X1 U10405 ( .A1(n9308), .A2(n9040), .A3(n9039), .ZN(n9041) );
  NAND4_X1 U10406 ( .A1(n9254), .A2(n4880), .A3(n9041), .A4(n9295), .ZN(n9042)
         );
  OR3_X1 U10407 ( .A1(n9044), .A2(n9043), .A3(n9042), .ZN(n9045) );
  NOR2_X1 U10408 ( .A1(n9046), .A2(n9045), .ZN(n9048) );
  INV_X1 U10409 ( .A(n9053), .ZN(n9109) );
  OAI21_X1 U10410 ( .B1(n9049), .B2(n4436), .A(n9109), .ZN(n9055) );
  INV_X1 U10411 ( .A(n9057), .ZN(n9107) );
  INV_X1 U10412 ( .A(n9058), .ZN(n9105) );
  INV_X1 U10413 ( .A(n9059), .ZN(n9060) );
  AND2_X1 U10414 ( .A1(n9061), .A2(n9060), .ZN(n9066) );
  AOI21_X1 U10415 ( .B1(n9749), .B2(n6964), .A(n9062), .ZN(n9065) );
  NAND4_X1 U10416 ( .A1(n9066), .A2(n9065), .A3(n9064), .A4(n9063), .ZN(n9070)
         );
  INV_X1 U10417 ( .A(n9067), .ZN(n9069) );
  OAI211_X1 U10418 ( .C1(n9071), .C2(n9070), .A(n9069), .B(n9068), .ZN(n9074)
         );
  NAND3_X1 U10419 ( .A1(n9074), .A2(n9073), .A3(n9072), .ZN(n9077) );
  INV_X1 U10420 ( .A(n9075), .ZN(n9076) );
  NAND2_X1 U10421 ( .A1(n9077), .A2(n9076), .ZN(n9080) );
  INV_X1 U10422 ( .A(n9078), .ZN(n9079) );
  NAND2_X1 U10423 ( .A1(n9080), .A2(n9079), .ZN(n9083) );
  NAND3_X1 U10424 ( .A1(n9083), .A2(n9082), .A3(n9081), .ZN(n9086) );
  INV_X1 U10425 ( .A(n9084), .ZN(n9085) );
  AOI21_X1 U10426 ( .B1(n9086), .B2(n4490), .A(n9085), .ZN(n9091) );
  INV_X1 U10427 ( .A(n9087), .ZN(n9089) );
  AOI22_X1 U10428 ( .A1(n9091), .A2(n9090), .B1(n9089), .B2(n9088), .ZN(n9094)
         );
  INV_X1 U10429 ( .A(n9092), .ZN(n9093) );
  AOI21_X1 U10430 ( .B1(n9095), .B2(n9094), .A(n9093), .ZN(n9098) );
  OAI21_X1 U10431 ( .B1(n9098), .B2(n9097), .A(n9096), .ZN(n9100) );
  AOI21_X1 U10432 ( .B1(n9101), .B2(n9100), .A(n9099), .ZN(n9103) );
  NOR2_X1 U10433 ( .A1(n9103), .A2(n9102), .ZN(n9104) );
  NOR2_X1 U10434 ( .A1(n9105), .A2(n9104), .ZN(n9106) );
  NOR2_X1 U10435 ( .A1(n9107), .A2(n9106), .ZN(n9110) );
  OAI211_X1 U10436 ( .C1(n9111), .C2(n9110), .A(n9109), .B(n9108), .ZN(n9112)
         );
  NAND2_X1 U10437 ( .A1(n9112), .A2(n4728), .ZN(n9114) );
  AOI21_X1 U10438 ( .B1(n9114), .B2(n6000), .A(n9113), .ZN(n9118) );
  INV_X1 U10439 ( .A(n9114), .ZN(n9116) );
  NAND2_X1 U10440 ( .A1(n9116), .A2(n6754), .ZN(n9117) );
  INV_X1 U10441 ( .A(n9120), .ZN(n9599) );
  NAND3_X1 U10442 ( .A1(n9122), .A2(n9599), .A3(n9121), .ZN(n9126) );
  INV_X1 U10443 ( .A(n9123), .ZN(n9124) );
  OAI211_X1 U10444 ( .C1(n9126), .C2(n9125), .A(P1_B_REG_SCAN_IN), .B(n9124), 
        .ZN(n9127) );
  OAI211_X1 U10445 ( .C1(n9130), .C2(n9129), .A(n9128), .B(n9127), .ZN(
        P1_U3242) );
  MUX2_X1 U10446 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9131), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10447 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9132), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10448 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9133), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10449 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9240), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10450 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9134), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10451 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9275), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10452 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9297), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10453 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9312), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10454 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9322), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10455 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9344), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10456 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9321), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10457 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9380), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10458 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9135), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10459 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9379), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10460 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9422), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10461 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9136), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10462 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9459), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10463 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9437), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10464 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9462), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10465 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9137), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10466 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n4957), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10467 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9138), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10468 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9139), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10469 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9140), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10470 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9141), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10471 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9142), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10472 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9143), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10473 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9144), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10474 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9145), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10475 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9146), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10476 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6964), .S(n9147), .Z(
        P1_U3555) );
  NOR2_X1 U10477 ( .A1(n9149), .A2(n9148), .ZN(n9151) );
  NOR2_X1 U10478 ( .A1(n9151), .A2(n9150), .ZN(n9154) );
  NAND2_X1 U10479 ( .A1(n9170), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9152) );
  OAI21_X1 U10480 ( .B1(n9170), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9152), .ZN(
        n9153) );
  NOR2_X1 U10481 ( .A1(n9154), .A2(n9153), .ZN(n9169) );
  AOI211_X1 U10482 ( .C1(n9154), .C2(n9153), .A(n9169), .B(n9660), .ZN(n9168)
         );
  NAND2_X1 U10483 ( .A1(n9156), .A2(n9155), .ZN(n9158) );
  NAND2_X1 U10484 ( .A1(n9158), .A2(n9157), .ZN(n9162) );
  NOR2_X1 U10485 ( .A1(n9170), .A2(n9159), .ZN(n9160) );
  AOI21_X1 U10486 ( .B1(n9170), .B2(n9159), .A(n9160), .ZN(n9161) );
  NOR2_X1 U10487 ( .A1(n9161), .A2(n9162), .ZN(n9176) );
  AOI21_X1 U10488 ( .B1(n9162), .B2(n9161), .A(n9176), .ZN(n9166) );
  AND2_X1 U10489 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9163) );
  AOI21_X1 U10490 ( .B1(n9673), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n9163), .ZN(
        n9165) );
  NAND2_X1 U10491 ( .A1(n9677), .A2(n9170), .ZN(n9164) );
  OAI211_X1 U10492 ( .C1(n9166), .C2(n9213), .A(n9165), .B(n9164), .ZN(n9167)
         );
  OR2_X1 U10493 ( .A1(n9168), .A2(n9167), .ZN(P1_U3259) );
  AOI21_X1 U10494 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9170), .A(n9169), .ZN(
        n9172) );
  MUX2_X1 U10495 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n9192), .S(n9188), .Z(n9171) );
  NAND2_X1 U10496 ( .A1(n9172), .A2(n9171), .ZN(n9195) );
  OAI21_X1 U10497 ( .B1(n9172), .B2(n9171), .A(n9195), .ZN(n9185) );
  AOI21_X1 U10498 ( .B1(n9673), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n9173), .ZN(
        n9183) );
  NAND2_X1 U10499 ( .A1(n9188), .A2(n9175), .ZN(n9174) );
  OAI21_X1 U10500 ( .B1(n9188), .B2(n9175), .A(n9174), .ZN(n9180) );
  AOI21_X1 U10501 ( .B1(n9177), .B2(n9159), .A(n9176), .ZN(n9178) );
  INV_X1 U10502 ( .A(n9178), .ZN(n9179) );
  NAND2_X1 U10503 ( .A1(n9180), .A2(n9179), .ZN(n9187) );
  OAI21_X1 U10504 ( .B1(n9180), .B2(n9179), .A(n9187), .ZN(n9181) );
  NAND2_X1 U10505 ( .A1(n9684), .A2(n9181), .ZN(n9182) );
  OAI211_X1 U10506 ( .C1(n9212), .C2(n9193), .A(n9183), .B(n9182), .ZN(n9184)
         );
  AOI21_X1 U10507 ( .B1(n9185), .B2(n9682), .A(n9184), .ZN(n9186) );
  INV_X1 U10508 ( .A(n9186), .ZN(P1_U3260) );
  INV_X1 U10509 ( .A(n9210), .ZN(n9205) );
  XNOR2_X1 U10510 ( .A(n9210), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9190) );
  OAI21_X1 U10511 ( .B1(n9188), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9187), .ZN(
        n9189) );
  NOR2_X1 U10512 ( .A1(n9189), .A2(n9190), .ZN(n9209) );
  AOI211_X1 U10513 ( .C1(n9190), .C2(n9189), .A(n9209), .B(n9213), .ZN(n9191)
         );
  INV_X1 U10514 ( .A(n9191), .ZN(n9204) );
  AND2_X1 U10515 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9202) );
  NAND2_X1 U10516 ( .A1(n9193), .A2(n9192), .ZN(n9194) );
  NAND2_X1 U10517 ( .A1(n9195), .A2(n9194), .ZN(n9200) );
  INV_X1 U10518 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9196) );
  OR2_X1 U10519 ( .A1(n9210), .A2(n9196), .ZN(n9198) );
  NAND2_X1 U10520 ( .A1(n9210), .A2(n9196), .ZN(n9197) );
  AND2_X1 U10521 ( .A1(n9198), .A2(n9197), .ZN(n9199) );
  NOR2_X1 U10522 ( .A1(n9200), .A2(n9199), .ZN(n9207) );
  AOI211_X1 U10523 ( .C1(n9200), .C2(n9199), .A(n9207), .B(n9660), .ZN(n9201)
         );
  AOI211_X1 U10524 ( .C1(n9673), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9202), .B(
        n9201), .ZN(n9203) );
  OAI211_X1 U10525 ( .C1(n9212), .C2(n9205), .A(n9204), .B(n9203), .ZN(
        P1_U3261) );
  AND2_X1 U10526 ( .A1(n9210), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9206) );
  OR2_X1 U10527 ( .A1(n9207), .A2(n9206), .ZN(n9208) );
  XNOR2_X1 U10528 ( .A(n9208), .B(n9372), .ZN(n9217) );
  INV_X1 U10529 ( .A(n9217), .ZN(n9215) );
  AOI21_X1 U10530 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9210), .A(n9209), .ZN(
        n9211) );
  XNOR2_X1 U10531 ( .A(n9211), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9216) );
  OAI21_X1 U10532 ( .B1(n9216), .B2(n9213), .A(n9212), .ZN(n9214) );
  AOI21_X1 U10533 ( .B1(n9215), .B2(n9682), .A(n9214), .ZN(n9219) );
  AOI22_X1 U10534 ( .A1(n9217), .A2(n9682), .B1(n9684), .B2(n9216), .ZN(n9218)
         );
  MUX2_X1 U10535 ( .A(n9219), .B(n9218), .S(n7035), .Z(n9221) );
  NAND2_X1 U10536 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9220) );
  OAI211_X1 U10537 ( .C1(n4764), .C2(n9222), .A(n9221), .B(n9220), .ZN(
        P1_U3262) );
  NAND2_X1 U10538 ( .A1(n8974), .A2(n9231), .ZN(n9230) );
  INV_X1 U10539 ( .A(n9225), .ZN(n9226) );
  OR2_X1 U10540 ( .A1(n9227), .A2(n9226), .ZN(n9479) );
  NOR2_X1 U10541 ( .A1(n4419), .A2(n9479), .ZN(n9233) );
  NOR2_X1 U10542 ( .A1(n9565), .A2(n9741), .ZN(n9228) );
  AOI211_X1 U10543 ( .C1(n4419), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9233), .B(
        n9228), .ZN(n9229) );
  OAI21_X1 U10544 ( .B1(n9477), .B2(n9740), .A(n9229), .ZN(P1_U3263) );
  OAI211_X1 U10545 ( .C1(n8974), .C2(n9231), .A(n9738), .B(n9230), .ZN(n9480)
         );
  NOR2_X1 U10546 ( .A1(n8974), .A2(n9741), .ZN(n9232) );
  AOI211_X1 U10547 ( .C1(n4419), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9233), .B(
        n9232), .ZN(n9234) );
  OAI21_X1 U10548 ( .B1(n9480), .B2(n9740), .A(n9234), .ZN(P1_U3264) );
  XNOR2_X1 U10549 ( .A(n9235), .B(n9238), .ZN(n9497) );
  INV_X1 U10550 ( .A(n9497), .ZN(n9251) );
  OAI21_X1 U10551 ( .B1(n9238), .B2(n9237), .A(n9236), .ZN(n9239) );
  NAND2_X1 U10552 ( .A1(n9239), .A2(n9715), .ZN(n9242) );
  AOI22_X1 U10553 ( .A1(n9240), .A2(n9460), .B1(n9461), .B2(n9275), .ZN(n9241)
         );
  NAND2_X1 U10554 ( .A1(n9242), .A2(n9241), .ZN(n9495) );
  INV_X1 U10555 ( .A(n9261), .ZN(n9244) );
  AOI211_X1 U10556 ( .C1(n9245), .C2(n9244), .A(n9549), .B(n9243), .ZN(n9496)
         );
  NAND2_X1 U10557 ( .A1(n9496), .A2(n9724), .ZN(n9248) );
  AOI22_X1 U10558 ( .A1(n9246), .A2(n9736), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n4419), .ZN(n9247) );
  OAI211_X1 U10559 ( .C1(n9573), .C2(n9741), .A(n9248), .B(n9247), .ZN(n9249)
         );
  AOI21_X1 U10560 ( .B1(n9495), .B2(n9471), .A(n9249), .ZN(n9250) );
  OAI21_X1 U10561 ( .B1(n9251), .B2(n9433), .A(n9250), .ZN(P1_U3266) );
  INV_X1 U10562 ( .A(n9502), .ZN(n9269) );
  OAI21_X1 U10563 ( .B1(n9254), .B2(n9253), .A(n9252), .ZN(n9255) );
  NAND2_X1 U10564 ( .A1(n9255), .A2(n9715), .ZN(n9260) );
  OAI22_X1 U10565 ( .A1(n9257), .A2(n9439), .B1(n9256), .B2(n9393), .ZN(n9258)
         );
  INV_X1 U10566 ( .A(n9258), .ZN(n9259) );
  NAND2_X1 U10567 ( .A1(n9260), .A2(n9259), .ZN(n9500) );
  INV_X1 U10568 ( .A(n9278), .ZN(n9262) );
  AOI211_X1 U10569 ( .C1(n9263), .C2(n9262), .A(n9549), .B(n9261), .ZN(n9501)
         );
  NAND2_X1 U10570 ( .A1(n9501), .A2(n9724), .ZN(n9266) );
  AOI22_X1 U10571 ( .A1(n9264), .A2(n9736), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n4419), .ZN(n9265) );
  OAI211_X1 U10572 ( .C1(n9576), .C2(n9741), .A(n9266), .B(n9265), .ZN(n9267)
         );
  AOI21_X1 U10573 ( .B1(n9500), .B2(n9471), .A(n9267), .ZN(n9268) );
  OAI21_X1 U10574 ( .B1(n9269), .B2(n9433), .A(n9268), .ZN(P1_U3267) );
  XNOR2_X1 U10575 ( .A(n4478), .B(n4880), .ZN(n9506) );
  INV_X1 U10576 ( .A(n9506), .ZN(n9286) );
  NAND2_X1 U10577 ( .A1(n9271), .A2(n9270), .ZN(n9272) );
  NAND2_X1 U10578 ( .A1(n9273), .A2(n9272), .ZN(n9274) );
  NAND2_X1 U10579 ( .A1(n9274), .A2(n9715), .ZN(n9277) );
  AOI22_X1 U10580 ( .A1(n9275), .A2(n9460), .B1(n9461), .B2(n9312), .ZN(n9276)
         );
  NAND2_X1 U10581 ( .A1(n9277), .A2(n9276), .ZN(n9504) );
  AOI211_X1 U10582 ( .C1(n9279), .C2(n9289), .A(n9549), .B(n9278), .ZN(n9505)
         );
  NAND2_X1 U10583 ( .A1(n9505), .A2(n9724), .ZN(n9283) );
  INV_X1 U10584 ( .A(n9280), .ZN(n9281) );
  AOI22_X1 U10585 ( .A1(n9281), .A2(n9736), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n4419), .ZN(n9282) );
  OAI211_X1 U10586 ( .C1(n9580), .C2(n9741), .A(n9283), .B(n9282), .ZN(n9284)
         );
  AOI21_X1 U10587 ( .B1(n9504), .B2(n9471), .A(n9284), .ZN(n9285) );
  OAI21_X1 U10588 ( .B1(n9286), .B2(n9433), .A(n9285), .ZN(P1_U3268) );
  XNOR2_X1 U10589 ( .A(n9288), .B(n9287), .ZN(n9513) );
  INV_X1 U10590 ( .A(n9289), .ZN(n9290) );
  AOI211_X1 U10591 ( .C1(n9510), .C2(n9303), .A(n9549), .B(n9290), .ZN(n9509)
         );
  INV_X1 U10592 ( .A(n9291), .ZN(n9292) );
  AOI22_X1 U10593 ( .A1(n9292), .A2(n9736), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n4419), .ZN(n9293) );
  OAI21_X1 U10594 ( .B1(n9294), .B2(n9741), .A(n9293), .ZN(n9300) );
  XNOR2_X1 U10595 ( .A(n9296), .B(n9295), .ZN(n9298) );
  AOI222_X1 U10596 ( .A1(n9715), .A2(n9298), .B1(n9297), .B2(n9460), .C1(n9322), .C2(n9461), .ZN(n9512) );
  NOR2_X1 U10597 ( .A1(n9512), .A2(n4419), .ZN(n9299) );
  AOI211_X1 U10598 ( .C1(n9509), .C2(n9724), .A(n9300), .B(n9299), .ZN(n9301)
         );
  OAI21_X1 U10599 ( .B1(n9513), .B2(n9433), .A(n9301), .ZN(P1_U3269) );
  XNOR2_X1 U10600 ( .A(n9302), .B(n9308), .ZN(n9518) );
  INV_X1 U10601 ( .A(n9303), .ZN(n9304) );
  AOI21_X1 U10602 ( .B1(n9514), .B2(n9325), .A(n9304), .ZN(n9515) );
  INV_X1 U10603 ( .A(n9305), .ZN(n9306) );
  AOI22_X1 U10604 ( .A1(n9306), .A2(n9736), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n4419), .ZN(n9307) );
  OAI21_X1 U10605 ( .B1(n4705), .B2(n9741), .A(n9307), .ZN(n9315) );
  OAI21_X1 U10606 ( .B1(n4505), .B2(n9309), .A(n9308), .ZN(n9311) );
  NAND2_X1 U10607 ( .A1(n9311), .A2(n9310), .ZN(n9313) );
  AOI222_X1 U10608 ( .A1(n9715), .A2(n9313), .B1(n9312), .B2(n9460), .C1(n9344), .C2(n9461), .ZN(n9517) );
  NOR2_X1 U10609 ( .A1(n9517), .A2(n4419), .ZN(n9314) );
  AOI211_X1 U10610 ( .C1(n9515), .C2(n9348), .A(n9315), .B(n9314), .ZN(n9316)
         );
  OAI21_X1 U10611 ( .B1(n9518), .B2(n9433), .A(n9316), .ZN(P1_U3270) );
  XNOR2_X1 U10612 ( .A(n9317), .B(n9319), .ZN(n9523) );
  OAI211_X1 U10613 ( .C1(n9320), .C2(n9319), .A(n9318), .B(n9715), .ZN(n9324)
         );
  AOI22_X1 U10614 ( .A1(n9322), .A2(n9460), .B1(n9461), .B2(n9321), .ZN(n9323)
         );
  NAND2_X1 U10615 ( .A1(n9324), .A2(n9323), .ZN(n9519) );
  INV_X1 U10616 ( .A(n9325), .ZN(n9326) );
  AOI211_X1 U10617 ( .C1(n9521), .C2(n4709), .A(n9549), .B(n9326), .ZN(n9520)
         );
  NAND2_X1 U10618 ( .A1(n9520), .A2(n9724), .ZN(n9329) );
  AOI22_X1 U10619 ( .A1(n9327), .A2(n9736), .B1(n4419), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9328) );
  OAI211_X1 U10620 ( .C1(n9330), .C2(n9741), .A(n9329), .B(n9328), .ZN(n9331)
         );
  AOI21_X1 U10621 ( .B1(n9471), .B2(n9519), .A(n9331), .ZN(n9332) );
  OAI21_X1 U10622 ( .B1(n9523), .B2(n9433), .A(n9332), .ZN(P1_U3271) );
  XNOR2_X1 U10623 ( .A(n9333), .B(n9339), .ZN(n9528) );
  AOI21_X1 U10624 ( .B1(n9524), .B2(n9357), .A(n9334), .ZN(n9525) );
  INV_X1 U10625 ( .A(n9524), .ZN(n9338) );
  INV_X1 U10626 ( .A(n9335), .ZN(n9336) );
  AOI22_X1 U10627 ( .A1(n4419), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9336), .B2(
        n9736), .ZN(n9337) );
  OAI21_X1 U10628 ( .B1(n9338), .B2(n9741), .A(n9337), .ZN(n9347) );
  INV_X1 U10629 ( .A(n9353), .ZN(n9341) );
  OAI21_X1 U10630 ( .B1(n9341), .B2(n9340), .A(n9339), .ZN(n9343) );
  NAND2_X1 U10631 ( .A1(n9343), .A2(n9342), .ZN(n9345) );
  AOI222_X1 U10632 ( .A1(n9715), .A2(n9345), .B1(n9344), .B2(n9460), .C1(n9380), .C2(n9461), .ZN(n9527) );
  NOR2_X1 U10633 ( .A1(n9527), .A2(n4419), .ZN(n9346) );
  AOI211_X1 U10634 ( .C1(n9525), .C2(n9348), .A(n9347), .B(n9346), .ZN(n9349)
         );
  OAI21_X1 U10635 ( .B1(n9528), .B2(n9433), .A(n9349), .ZN(P1_U3272) );
  XOR2_X1 U10636 ( .A(n9351), .B(n9350), .Z(n9531) );
  INV_X1 U10637 ( .A(n9531), .ZN(n9366) );
  AOI21_X1 U10638 ( .B1(n9352), .B2(n9351), .A(n9732), .ZN(n9354) );
  NAND2_X1 U10639 ( .A1(n9354), .A2(n9353), .ZN(n9356) );
  NAND2_X1 U10640 ( .A1(n9356), .A2(n9355), .ZN(n9529) );
  INV_X1 U10641 ( .A(n9368), .ZN(n9359) );
  INV_X1 U10642 ( .A(n9357), .ZN(n9358) );
  AOI211_X1 U10643 ( .C1(n9360), .C2(n9359), .A(n9549), .B(n9358), .ZN(n9530)
         );
  NAND2_X1 U10644 ( .A1(n9530), .A2(n9724), .ZN(n9363) );
  AOI22_X1 U10645 ( .A1(n4419), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9361), .B2(
        n9736), .ZN(n9362) );
  OAI211_X1 U10646 ( .C1(n9588), .C2(n9741), .A(n9363), .B(n9362), .ZN(n9364)
         );
  AOI21_X1 U10647 ( .B1(n9471), .B2(n9529), .A(n9364), .ZN(n9365) );
  OAI21_X1 U10648 ( .B1(n9366), .B2(n9433), .A(n9365), .ZN(P1_U3273) );
  XNOR2_X1 U10649 ( .A(n9367), .B(n9377), .ZN(n9536) );
  INV_X1 U10650 ( .A(n9536), .ZN(n9385) );
  INV_X1 U10651 ( .A(n9395), .ZN(n9369) );
  AOI211_X1 U10652 ( .C1(n9370), .C2(n9369), .A(n9549), .B(n9368), .ZN(n9535)
         );
  NOR2_X1 U10653 ( .A1(n9592), .A2(n9741), .ZN(n9374) );
  OAI22_X1 U10654 ( .A1(n9471), .A2(n9372), .B1(n9371), .B2(n9701), .ZN(n9373)
         );
  AOI211_X1 U10655 ( .C1(n9535), .C2(n9724), .A(n9374), .B(n9373), .ZN(n9384)
         );
  OAI21_X1 U10656 ( .B1(n9377), .B2(n9376), .A(n9375), .ZN(n9378) );
  NAND2_X1 U10657 ( .A1(n9378), .A2(n9715), .ZN(n9382) );
  AOI22_X1 U10658 ( .A1(n9380), .A2(n9460), .B1(n9461), .B2(n9379), .ZN(n9381)
         );
  NAND2_X1 U10659 ( .A1(n9382), .A2(n9381), .ZN(n9534) );
  NAND2_X1 U10660 ( .A1(n9534), .A2(n9471), .ZN(n9383) );
  OAI211_X1 U10661 ( .C1(n9385), .C2(n9433), .A(n9384), .B(n9383), .ZN(
        P1_U3274) );
  XNOR2_X1 U10662 ( .A(n9386), .B(n9390), .ZN(n9545) );
  INV_X1 U10663 ( .A(n9387), .ZN(n9388) );
  AOI21_X1 U10664 ( .B1(n9390), .B2(n9389), .A(n9388), .ZN(n9391) );
  OAI222_X1 U10665 ( .A1(n9439), .A2(n9394), .B1(n9393), .B2(n9392), .C1(n9732), .C2(n9391), .ZN(n9540) );
  AOI211_X1 U10666 ( .C1(n9542), .C2(n9406), .A(n9549), .B(n9395), .ZN(n9541)
         );
  NAND2_X1 U10667 ( .A1(n9541), .A2(n9724), .ZN(n9398) );
  AOI22_X1 U10668 ( .A1(n4419), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9396), .B2(
        n9736), .ZN(n9397) );
  OAI211_X1 U10669 ( .C1(n7881), .C2(n9741), .A(n9398), .B(n9397), .ZN(n9399)
         );
  AOI21_X1 U10670 ( .B1(n9540), .B2(n9471), .A(n9399), .ZN(n9400) );
  OAI21_X1 U10671 ( .B1(n9545), .B2(n9433), .A(n9400), .ZN(P1_U3275) );
  XOR2_X1 U10672 ( .A(n9402), .B(n9401), .Z(n9634) );
  INV_X1 U10673 ( .A(n9634), .ZN(n9413) );
  XNOR2_X1 U10674 ( .A(n9403), .B(n9402), .ZN(n9405) );
  OAI21_X1 U10675 ( .B1(n9405), .B2(n9732), .A(n9404), .ZN(n9633) );
  INV_X1 U10676 ( .A(n9425), .ZN(n9407) );
  OAI211_X1 U10677 ( .C1(n9407), .C2(n9631), .A(n9406), .B(n9738), .ZN(n9630)
         );
  NOR2_X1 U10678 ( .A1(n9630), .A2(n9740), .ZN(n9411) );
  AOI22_X1 U10679 ( .A1(n4419), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9408), .B2(
        n9736), .ZN(n9409) );
  OAI21_X1 U10680 ( .B1(n9631), .B2(n9741), .A(n9409), .ZN(n9410) );
  AOI211_X1 U10681 ( .C1(n9633), .C2(n9471), .A(n9411), .B(n9410), .ZN(n9412)
         );
  OAI21_X1 U10682 ( .B1(n9413), .B2(n9433), .A(n9412), .ZN(P1_U3276) );
  XOR2_X1 U10683 ( .A(n9414), .B(n9416), .Z(n9639) );
  INV_X1 U10684 ( .A(n9639), .ZN(n9434) );
  INV_X1 U10685 ( .A(n9435), .ZN(n9418) );
  INV_X1 U10686 ( .A(n9415), .ZN(n9417) );
  OAI21_X1 U10687 ( .B1(n9418), .B2(n9417), .A(n9416), .ZN(n9419) );
  OAI211_X1 U10688 ( .C1(n9421), .C2(n9420), .A(n9419), .B(n9715), .ZN(n9424)
         );
  AOI22_X1 U10689 ( .A1(n9461), .A2(n9459), .B1(n9422), .B2(n9460), .ZN(n9423)
         );
  NAND2_X1 U10690 ( .A1(n9424), .A2(n9423), .ZN(n9638) );
  OAI211_X1 U10691 ( .C1(n9447), .C2(n9636), .A(n9425), .B(n9738), .ZN(n9635)
         );
  OAI22_X1 U10692 ( .A1(n9471), .A2(n9427), .B1(n9426), .B2(n9701), .ZN(n9428)
         );
  AOI21_X1 U10693 ( .B1(n9429), .B2(n9706), .A(n9428), .ZN(n9430) );
  OAI21_X1 U10694 ( .B1(n9635), .B2(n9740), .A(n9430), .ZN(n9431) );
  AOI21_X1 U10695 ( .B1(n9638), .B2(n9471), .A(n9431), .ZN(n9432) );
  OAI21_X1 U10696 ( .B1(n9434), .B2(n9433), .A(n9432), .ZN(P1_U3277) );
  OAI21_X1 U10697 ( .B1(n9443), .B2(n9436), .A(n9435), .ZN(n9442) );
  NAND2_X1 U10698 ( .A1(n9437), .A2(n9461), .ZN(n9438) );
  OAI21_X1 U10699 ( .B1(n9440), .B2(n9439), .A(n9438), .ZN(n9441) );
  AOI21_X1 U10700 ( .B1(n9442), .B2(n9715), .A(n9441), .ZN(n9641) );
  XNOR2_X1 U10701 ( .A(n9444), .B(n9443), .ZN(n9644) );
  NAND2_X1 U10702 ( .A1(n9644), .A2(n9725), .ZN(n9454) );
  OAI22_X1 U10703 ( .A1(n9471), .A2(n9446), .B1(n9445), .B2(n9701), .ZN(n9451)
         );
  INV_X1 U10704 ( .A(n9467), .ZN(n9449) );
  INV_X1 U10705 ( .A(n9447), .ZN(n9448) );
  OAI211_X1 U10706 ( .C1(n9642), .C2(n9449), .A(n9448), .B(n9738), .ZN(n9640)
         );
  NOR2_X1 U10707 ( .A1(n9640), .A2(n9740), .ZN(n9450) );
  AOI211_X1 U10708 ( .C1(n9706), .C2(n9452), .A(n9451), .B(n9450), .ZN(n9453)
         );
  OAI211_X1 U10709 ( .C1(n4419), .C2(n9641), .A(n9454), .B(n9453), .ZN(
        P1_U3278) );
  XNOR2_X1 U10710 ( .A(n9456), .B(n9455), .ZN(n9793) );
  XNOR2_X1 U10711 ( .A(n9458), .B(n9457), .ZN(n9464) );
  AOI22_X1 U10712 ( .A1(n9462), .A2(n9461), .B1(n9460), .B2(n9459), .ZN(n9463)
         );
  OAI21_X1 U10713 ( .B1(n9464), .B2(n9732), .A(n9463), .ZN(n9465) );
  AOI21_X1 U10714 ( .B1(n9793), .B2(n9735), .A(n9465), .ZN(n9795) );
  AOI21_X1 U10715 ( .B1(n9466), .B2(n9473), .A(n9549), .ZN(n9468) );
  NAND2_X1 U10716 ( .A1(n9468), .A2(n9467), .ZN(n9789) );
  OAI22_X1 U10717 ( .A1(n9471), .A2(n9470), .B1(n9469), .B2(n9701), .ZN(n9472)
         );
  AOI21_X1 U10718 ( .B1(n9473), .B2(n9706), .A(n9472), .ZN(n9474) );
  OAI21_X1 U10719 ( .B1(n9789), .B2(n9740), .A(n9474), .ZN(n9475) );
  AOI21_X1 U10720 ( .B1(n9793), .B2(n9743), .A(n9475), .ZN(n9476) );
  OAI21_X1 U10721 ( .B1(n9795), .B2(n4419), .A(n9476), .ZN(P1_U3279) );
  AND2_X1 U10722 ( .A1(n9480), .A2(n9479), .ZN(n9566) );
  MUX2_X1 U10723 ( .A(n7918), .B(n9566), .S(n9814), .Z(n9481) );
  OAI21_X1 U10724 ( .B1(n8974), .B2(n9539), .A(n9481), .ZN(P1_U3552) );
  AOI21_X1 U10725 ( .B1(n9629), .B2(n9483), .A(n9482), .ZN(n9484) );
  AND2_X1 U10726 ( .A1(n9485), .A2(n9484), .ZN(n9486) );
  OAI21_X1 U10727 ( .B1(n9487), .B2(n9544), .A(n9486), .ZN(n9569) );
  MUX2_X1 U10728 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9569), .S(n9814), .Z(
        P1_U3551) );
  AOI22_X1 U10729 ( .A1(n9490), .A2(n9738), .B1(n9629), .B2(n9489), .ZN(n9491)
         );
  NAND2_X1 U10730 ( .A1(n9494), .A2(n9493), .ZN(n9570) );
  MUX2_X1 U10731 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9570), .S(n9814), .Z(
        P1_U3550) );
  INV_X1 U10732 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9498) );
  MUX2_X1 U10733 ( .A(n9498), .B(n9571), .S(n9814), .Z(n9499) );
  OAI21_X1 U10734 ( .B1(n9573), .B2(n9539), .A(n9499), .ZN(P1_U3549) );
  MUX2_X1 U10735 ( .A(n10059), .B(n9574), .S(n9814), .Z(n9503) );
  OAI21_X1 U10736 ( .B1(n9576), .B2(n9539), .A(n9503), .ZN(P1_U3548) );
  MUX2_X1 U10737 ( .A(n9507), .B(n9577), .S(n9814), .Z(n9508) );
  OAI21_X1 U10738 ( .B1(n9580), .B2(n9539), .A(n9508), .ZN(P1_U3547) );
  AOI21_X1 U10739 ( .B1(n9629), .B2(n9510), .A(n9509), .ZN(n9511) );
  OAI211_X1 U10740 ( .C1(n9513), .C2(n9544), .A(n9512), .B(n9511), .ZN(n9581)
         );
  MUX2_X1 U10741 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9581), .S(n9814), .Z(
        P1_U3546) );
  AOI22_X1 U10742 ( .A1(n9515), .A2(n9738), .B1(n9629), .B2(n9514), .ZN(n9516)
         );
  OAI211_X1 U10743 ( .C1(n9518), .C2(n9544), .A(n9517), .B(n9516), .ZN(n9582)
         );
  MUX2_X1 U10744 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9582), .S(n9814), .Z(
        P1_U3545) );
  AOI211_X1 U10745 ( .C1(n9629), .C2(n9521), .A(n9520), .B(n9519), .ZN(n9522)
         );
  OAI21_X1 U10746 ( .B1(n9523), .B2(n9544), .A(n9522), .ZN(n9583) );
  MUX2_X1 U10747 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9583), .S(n9814), .Z(
        P1_U3544) );
  AOI22_X1 U10748 ( .A1(n9525), .A2(n9738), .B1(n9629), .B2(n9524), .ZN(n9526)
         );
  OAI211_X1 U10749 ( .C1(n9528), .C2(n9544), .A(n9527), .B(n9526), .ZN(n9584)
         );
  MUX2_X1 U10750 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9584), .S(n9814), .Z(
        P1_U3543) );
  INV_X1 U10751 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9532) );
  AOI211_X1 U10752 ( .C1(n9531), .C2(n9802), .A(n9530), .B(n9529), .ZN(n9585)
         );
  MUX2_X1 U10753 ( .A(n9532), .B(n9585), .S(n9814), .Z(n9533) );
  OAI21_X1 U10754 ( .B1(n9588), .B2(n9539), .A(n9533), .ZN(P1_U3542) );
  AOI211_X1 U10755 ( .C1(n9536), .C2(n9802), .A(n9535), .B(n9534), .ZN(n9589)
         );
  MUX2_X1 U10756 ( .A(n9537), .B(n9589), .S(n9814), .Z(n9538) );
  OAI21_X1 U10757 ( .B1(n9592), .B2(n9539), .A(n9538), .ZN(P1_U3541) );
  AOI211_X1 U10758 ( .C1(n9629), .C2(n9542), .A(n9541), .B(n9540), .ZN(n9543)
         );
  OAI21_X1 U10759 ( .B1(n9545), .B2(n9544), .A(n9543), .ZN(n9593) );
  MUX2_X1 U10760 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9593), .S(n9814), .Z(
        P1_U3540) );
  INV_X1 U10761 ( .A(n9546), .ZN(n9792) );
  XOR2_X1 U10762 ( .A(n9551), .B(n9547), .Z(n9698) );
  AOI211_X1 U10763 ( .C1(n4422), .C2(n9550), .A(n9549), .B(n9548), .ZN(n9691)
         );
  INV_X1 U10764 ( .A(n9551), .ZN(n9553) );
  NAND3_X1 U10765 ( .A1(n9554), .A2(n9553), .A3(n9552), .ZN(n9555) );
  AOI21_X1 U10766 ( .B1(n9556), .B2(n9555), .A(n9732), .ZN(n9558) );
  AOI211_X1 U10767 ( .C1(n9698), .C2(n9735), .A(n9558), .B(n9557), .ZN(n9700)
         );
  INV_X1 U10768 ( .A(n9700), .ZN(n9559) );
  AOI211_X1 U10769 ( .C1(n9792), .C2(n9698), .A(n9691), .B(n9559), .ZN(n9598)
         );
  AOI22_X1 U10770 ( .A1(n4422), .A2(n9560), .B1(n9811), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n9561) );
  OAI21_X1 U10771 ( .B1(n9598), .B2(n9811), .A(n9561), .ZN(P1_U3533) );
  INV_X1 U10772 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9563) );
  MUX2_X1 U10773 ( .A(n9563), .B(n9562), .S(n9788), .Z(n9564) );
  OAI21_X1 U10774 ( .B1(n9565), .B2(n9595), .A(n9564), .ZN(P1_U3521) );
  INV_X1 U10775 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9567) );
  MUX2_X1 U10776 ( .A(n9567), .B(n9566), .S(n9788), .Z(n9568) );
  OAI21_X1 U10777 ( .B1(n8974), .B2(n9595), .A(n9568), .ZN(P1_U3520) );
  MUX2_X1 U10778 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9569), .S(n9788), .Z(
        P1_U3519) );
  MUX2_X1 U10779 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9570), .S(n9788), .Z(
        P1_U3518) );
  MUX2_X1 U10780 ( .A(n10035), .B(n9571), .S(n9788), .Z(n9572) );
  OAI21_X1 U10781 ( .B1(n9573), .B2(n9595), .A(n9572), .ZN(P1_U3517) );
  MUX2_X1 U10782 ( .A(n9997), .B(n9574), .S(n9788), .Z(n9575) );
  OAI21_X1 U10783 ( .B1(n9576), .B2(n9595), .A(n9575), .ZN(P1_U3516) );
  INV_X1 U10784 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9578) );
  MUX2_X1 U10785 ( .A(n9578), .B(n9577), .S(n9788), .Z(n9579) );
  OAI21_X1 U10786 ( .B1(n9580), .B2(n9595), .A(n9579), .ZN(P1_U3515) );
  MUX2_X1 U10787 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9581), .S(n9788), .Z(
        P1_U3514) );
  MUX2_X1 U10788 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9582), .S(n9788), .Z(
        P1_U3513) );
  MUX2_X1 U10789 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9583), .S(n9788), .Z(
        P1_U3512) );
  MUX2_X1 U10790 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9584), .S(n9788), .Z(
        P1_U3511) );
  INV_X1 U10791 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9586) );
  MUX2_X1 U10792 ( .A(n9586), .B(n9585), .S(n9788), .Z(n9587) );
  OAI21_X1 U10793 ( .B1(n9588), .B2(n9595), .A(n9587), .ZN(P1_U3510) );
  MUX2_X1 U10794 ( .A(n9590), .B(n9589), .S(n9788), .Z(n9591) );
  OAI21_X1 U10795 ( .B1(n9592), .B2(n9595), .A(n9591), .ZN(P1_U3509) );
  MUX2_X1 U10796 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9593), .S(n9788), .Z(
        P1_U3507) );
  INV_X1 U10797 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9594) );
  OAI22_X1 U10798 ( .A1(n9696), .A2(n9595), .B1(n9788), .B2(n9594), .ZN(n9596)
         );
  INV_X1 U10799 ( .A(n9596), .ZN(n9597) );
  OAI21_X1 U10800 ( .B1(n9598), .B2(n9967), .A(n9597), .ZN(P1_U3486) );
  AND2_X1 U10801 ( .A1(n9600), .A2(n9599), .ZN(n9747) );
  MUX2_X1 U10802 ( .A(P1_D_REG_1__SCAN_IN), .B(n9601), .S(n9747), .Z(P1_U3440)
         );
  MUX2_X1 U10803 ( .A(P1_D_REG_0__SCAN_IN), .B(n9602), .S(n9747), .Z(P1_U3439)
         );
  NAND3_X1 U10804 ( .A1(n9603), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n9605) );
  OAI22_X1 U10805 ( .A1(n9606), .A2(n9605), .B1(n9604), .B2(n9616), .ZN(n9607)
         );
  AOI21_X1 U10806 ( .B1(n9609), .B2(n9608), .A(n9607), .ZN(n9610) );
  INV_X1 U10807 ( .A(n9610), .ZN(P1_U3324) );
  OAI222_X1 U10808 ( .A1(n9616), .A2(n9612), .B1(P1_U3086), .B2(n6011), .C1(
        n7925), .C2(n9611), .ZN(P1_U3326) );
  MUX2_X1 U10809 ( .A(n9617), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR3_X1 U10810 ( .A1(n9619), .A2(n9618), .A3(n9922), .ZN(n9621) );
  AOI211_X1 U10811 ( .C1(n9927), .C2(n9622), .A(n9621), .B(n9620), .ZN(n9627)
         );
  AOI22_X1 U10812 ( .A1(n9941), .A2(n9627), .B1(n8208), .B2(n9939), .ZN(
        P2_U3473) );
  OAI22_X1 U10813 ( .A1(n9624), .A2(n9922), .B1(n9623), .B2(n9915), .ZN(n9625)
         );
  NOR2_X1 U10814 ( .A1(n9626), .A2(n9625), .ZN(n9628) );
  AOI22_X1 U10815 ( .A1(n9941), .A2(n9628), .B1(n7793), .B2(n9939), .ZN(
        P2_U3472) );
  AOI22_X1 U10816 ( .A1(n9929), .A2(n5441), .B1(n9627), .B2(n9928), .ZN(
        P2_U3432) );
  INV_X1 U10817 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9976) );
  AOI22_X1 U10818 ( .A1(n9929), .A2(n9976), .B1(n9628), .B2(n9928), .ZN(
        P2_U3429) );
  INV_X1 U10819 ( .A(n9629), .ZN(n9799) );
  OAI21_X1 U10820 ( .B1(n9631), .B2(n9799), .A(n9630), .ZN(n9632) );
  AOI211_X1 U10821 ( .C1(n9634), .C2(n9802), .A(n9633), .B(n9632), .ZN(n9645)
         );
  AOI22_X1 U10822 ( .A1(n9814), .A2(n9645), .B1(n9175), .B2(n9811), .ZN(
        P1_U3539) );
  OAI21_X1 U10823 ( .B1(n9636), .B2(n9799), .A(n9635), .ZN(n9637) );
  AOI211_X1 U10824 ( .C1(n9639), .C2(n9802), .A(n9638), .B(n9637), .ZN(n9647)
         );
  AOI22_X1 U10825 ( .A1(n9814), .A2(n9647), .B1(n9159), .B2(n9811), .ZN(
        P1_U3538) );
  OAI211_X1 U10826 ( .C1(n9642), .C2(n9799), .A(n9641), .B(n9640), .ZN(n9643)
         );
  AOI21_X1 U10827 ( .B1(n9644), .B2(n9802), .A(n9643), .ZN(n9649) );
  AOI22_X1 U10828 ( .A1(n9814), .A2(n9649), .B1(n6290), .B2(n9811), .ZN(
        P1_U3537) );
  AOI22_X1 U10829 ( .A1(n9788), .A2(n9645), .B1(n6315), .B2(n9967), .ZN(
        P1_U3504) );
  INV_X1 U10830 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9646) );
  AOI22_X1 U10831 ( .A1(n9788), .A2(n9647), .B1(n9646), .B2(n9967), .ZN(
        P1_U3501) );
  INV_X1 U10832 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9648) );
  AOI22_X1 U10833 ( .A1(n9788), .A2(n9649), .B1(n9648), .B2(n9967), .ZN(
        P1_U3498) );
  XNOR2_X1 U10834 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10835 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10836 ( .A(n9650), .ZN(n9652) );
  NAND2_X1 U10837 ( .A1(n9651), .A2(n6013), .ZN(n9653) );
  NAND2_X1 U10838 ( .A1(n9652), .A2(n9653), .ZN(n9654) );
  MUX2_X1 U10839 ( .A(n9654), .B(n9653), .S(n9666), .Z(n9656) );
  NAND2_X1 U10840 ( .A1(n9656), .A2(n9655), .ZN(n9658) );
  AOI22_X1 U10841 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9673), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9657) );
  OAI21_X1 U10842 ( .B1(n9659), .B2(n9658), .A(n9657), .ZN(P1_U3243) );
  AOI22_X1 U10843 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n9673), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9672) );
  AOI211_X1 U10844 ( .C1(n9663), .C2(n9662), .A(n9661), .B(n9660), .ZN(n9664)
         );
  AOI21_X1 U10845 ( .B1(n9677), .B2(n9665), .A(n9664), .ZN(n9671) );
  NOR2_X1 U10846 ( .A1(n9666), .A2(n6013), .ZN(n9669) );
  OAI211_X1 U10847 ( .C1(n9669), .C2(n9668), .A(n9684), .B(n9667), .ZN(n9670)
         );
  NAND3_X1 U10848 ( .A1(n9672), .A2(n9671), .A3(n9670), .ZN(P1_U3244) );
  AOI22_X1 U10849 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(n9673), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9690) );
  INV_X1 U10850 ( .A(n9674), .ZN(n9675) );
  AOI21_X1 U10851 ( .B1(n9677), .B2(n9676), .A(n9675), .ZN(n9689) );
  AOI21_X1 U10852 ( .B1(n9680), .B2(n9679), .A(n9678), .ZN(n9681) );
  NAND2_X1 U10853 ( .A1(n9682), .A2(n9681), .ZN(n9688) );
  OAI211_X1 U10854 ( .C1(n9686), .C2(n9685), .A(n9684), .B(n9683), .ZN(n9687)
         );
  NAND4_X1 U10855 ( .A1(n9690), .A2(n9689), .A3(n9688), .A4(n9687), .ZN(
        P1_U3245) );
  NAND2_X1 U10856 ( .A1(n9691), .A2(n9724), .ZN(n9695) );
  INV_X1 U10857 ( .A(n9692), .ZN(n9693) );
  AOI22_X1 U10858 ( .A1(n4419), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9693), .B2(
        n9736), .ZN(n9694) );
  OAI211_X1 U10859 ( .C1(n9696), .C2(n9741), .A(n9695), .B(n9694), .ZN(n9697)
         );
  AOI21_X1 U10860 ( .B1(n9698), .B2(n9743), .A(n9697), .ZN(n9699) );
  OAI21_X1 U10861 ( .B1(n4419), .B2(n9700), .A(n9699), .ZN(P1_U3282) );
  OAI22_X1 U10862 ( .A1(n9471), .A2(n9703), .B1(n9702), .B2(n9701), .ZN(n9704)
         );
  AOI21_X1 U10863 ( .B1(n9706), .B2(n9705), .A(n9704), .ZN(n9707) );
  OAI21_X1 U10864 ( .B1(n9708), .B2(n9740), .A(n9707), .ZN(n9709) );
  AOI21_X1 U10865 ( .B1(n9710), .B2(n9743), .A(n9709), .ZN(n9711) );
  OAI21_X1 U10866 ( .B1(n4419), .B2(n9712), .A(n9711), .ZN(P1_U3286) );
  XOR2_X1 U10867 ( .A(n9720), .B(n9713), .Z(n9716) );
  AOI21_X1 U10868 ( .B1(n9716), .B2(n9715), .A(n9714), .ZN(n9757) );
  AOI22_X1 U10869 ( .A1(n4419), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9736), .ZN(n9717) );
  OAI21_X1 U10870 ( .B1(n9741), .B2(n9756), .A(n9717), .ZN(n9718) );
  INV_X1 U10871 ( .A(n9718), .ZN(n9727) );
  XNOR2_X1 U10872 ( .A(n9719), .B(n9720), .ZN(n9760) );
  INV_X1 U10873 ( .A(n9737), .ZN(n9722) );
  OAI211_X1 U10874 ( .C1(n9722), .C2(n9756), .A(n9738), .B(n9721), .ZN(n9755)
         );
  INV_X1 U10875 ( .A(n9755), .ZN(n9723) );
  AOI22_X1 U10876 ( .A1(n9760), .A2(n9725), .B1(n9724), .B2(n9723), .ZN(n9726)
         );
  OAI211_X1 U10877 ( .C1(n4419), .C2(n9757), .A(n9727), .B(n9726), .ZN(
        P1_U3291) );
  XNOR2_X1 U10878 ( .A(n9730), .B(n9728), .ZN(n9753) );
  XNOR2_X1 U10879 ( .A(n9730), .B(n9729), .ZN(n9733) );
  OAI21_X1 U10880 ( .B1(n9733), .B2(n9732), .A(n9731), .ZN(n9734) );
  AOI21_X1 U10881 ( .B1(n9735), .B2(n9753), .A(n9734), .ZN(n9750) );
  AOI22_X1 U10882 ( .A1(n9736), .A2(P1_REG3_REG_1__SCAN_IN), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(n4419), .ZN(n9745) );
  OAI211_X1 U10883 ( .C1(n9739), .C2(n9749), .A(n9738), .B(n9737), .ZN(n9748)
         );
  OAI22_X1 U10884 ( .A1(n9749), .A2(n9741), .B1(n9740), .B2(n9748), .ZN(n9742)
         );
  AOI21_X1 U10885 ( .B1(n9743), .B2(n9753), .A(n9742), .ZN(n9744) );
  OAI211_X1 U10886 ( .C1(n4419), .C2(n9750), .A(n9745), .B(n9744), .ZN(
        P1_U3292) );
  AND2_X1 U10887 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9746), .ZN(P1_U3294) );
  AND2_X1 U10888 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9746), .ZN(P1_U3295) );
  AND2_X1 U10889 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9746), .ZN(P1_U3296) );
  AND2_X1 U10890 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9746), .ZN(P1_U3297) );
  AND2_X1 U10891 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9746), .ZN(P1_U3298) );
  AND2_X1 U10892 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9746), .ZN(P1_U3299) );
  INV_X1 U10893 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10265) );
  NOR2_X1 U10894 ( .A1(n9747), .A2(n10265), .ZN(P1_U3300) );
  AND2_X1 U10895 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9746), .ZN(P1_U3301) );
  NOR2_X1 U10896 ( .A1(n9747), .A2(n10078), .ZN(P1_U3302) );
  AND2_X1 U10897 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9746), .ZN(P1_U3303) );
  AND2_X1 U10898 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9746), .ZN(P1_U3304) );
  NOR2_X1 U10899 ( .A1(n9747), .A2(n10173), .ZN(P1_U3305) );
  AND2_X1 U10900 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9746), .ZN(P1_U3306) );
  INV_X1 U10901 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10257) );
  NOR2_X1 U10902 ( .A1(n9747), .A2(n10257), .ZN(P1_U3307) );
  AND2_X1 U10903 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9746), .ZN(P1_U3308) );
  INV_X1 U10904 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10194) );
  NOR2_X1 U10905 ( .A1(n9747), .A2(n10194), .ZN(P1_U3309) );
  AND2_X1 U10906 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9746), .ZN(P1_U3310) );
  AND2_X1 U10907 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9746), .ZN(P1_U3311) );
  AND2_X1 U10908 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9746), .ZN(P1_U3312) );
  INV_X1 U10909 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10196) );
  NOR2_X1 U10910 ( .A1(n9747), .A2(n10196), .ZN(P1_U3313) );
  NOR2_X1 U10911 ( .A1(n9747), .A2(n10160), .ZN(P1_U3314) );
  AND2_X1 U10912 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9746), .ZN(P1_U3315) );
  AND2_X1 U10913 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9746), .ZN(P1_U3316) );
  AND2_X1 U10914 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9746), .ZN(P1_U3317) );
  AND2_X1 U10915 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9746), .ZN(P1_U3318) );
  AND2_X1 U10916 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9746), .ZN(P1_U3319) );
  AND2_X1 U10917 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9746), .ZN(P1_U3320) );
  NOR2_X1 U10918 ( .A1(n9747), .A2(n10056), .ZN(P1_U3321) );
  AND2_X1 U10919 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9746), .ZN(P1_U3322) );
  INV_X1 U10920 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10195) );
  NOR2_X1 U10921 ( .A1(n9747), .A2(n10195), .ZN(P1_U3323) );
  OAI21_X1 U10922 ( .B1(n9749), .B2(n9799), .A(n9748), .ZN(n9752) );
  INV_X1 U10923 ( .A(n9750), .ZN(n9751) );
  AOI211_X1 U10924 ( .C1(n9792), .C2(n9753), .A(n9752), .B(n9751), .ZN(n9796)
         );
  INV_X1 U10925 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9754) );
  AOI22_X1 U10926 ( .A1(n9788), .A2(n9796), .B1(n9754), .B2(n9967), .ZN(
        P1_U3456) );
  OAI21_X1 U10927 ( .B1(n9756), .B2(n9799), .A(n9755), .ZN(n9759) );
  INV_X1 U10928 ( .A(n9757), .ZN(n9758) );
  AOI211_X1 U10929 ( .C1(n9802), .C2(n9760), .A(n9759), .B(n9758), .ZN(n9797)
         );
  AOI22_X1 U10930 ( .A1(n9788), .A2(n9797), .B1(n6042), .B2(n9967), .ZN(
        P1_U3459) );
  OAI21_X1 U10931 ( .B1(n9762), .B2(n9799), .A(n9761), .ZN(n9765) );
  INV_X1 U10932 ( .A(n9763), .ZN(n9764) );
  AOI211_X1 U10933 ( .C1(n9766), .C2(n9802), .A(n9765), .B(n9764), .ZN(n9806)
         );
  INV_X1 U10934 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U10935 ( .A1(n9788), .A2(n9806), .B1(n10184), .B2(n9967), .ZN(
        P1_U3465) );
  OAI21_X1 U10936 ( .B1(n9768), .B2(n9799), .A(n9767), .ZN(n9770) );
  AOI211_X1 U10937 ( .C1(n9792), .C2(n9771), .A(n9770), .B(n9769), .ZN(n9807)
         );
  INV_X1 U10938 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10256) );
  AOI22_X1 U10939 ( .A1(n9788), .A2(n9807), .B1(n10256), .B2(n9967), .ZN(
        P1_U3477) );
  OAI211_X1 U10940 ( .C1(n9774), .C2(n9799), .A(n9773), .B(n9772), .ZN(n9775)
         );
  AOI21_X1 U10941 ( .B1(n9776), .B2(n9802), .A(n9775), .ZN(n9808) );
  INV_X1 U10942 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9777) );
  AOI22_X1 U10943 ( .A1(n9788), .A2(n9808), .B1(n9777), .B2(n9967), .ZN(
        P1_U3483) );
  OAI211_X1 U10944 ( .C1(n9780), .C2(n9799), .A(n9779), .B(n9778), .ZN(n9781)
         );
  AOI21_X1 U10945 ( .B1(n9782), .B2(n9802), .A(n9781), .ZN(n9809) );
  INV_X1 U10946 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9970) );
  AOI22_X1 U10947 ( .A1(n9788), .A2(n9809), .B1(n9970), .B2(n9967), .ZN(
        P1_U3489) );
  OAI211_X1 U10948 ( .C1(n4703), .C2(n9799), .A(n9784), .B(n9783), .ZN(n9785)
         );
  AOI21_X1 U10949 ( .B1(n9786), .B2(n9802), .A(n9785), .ZN(n9810) );
  INV_X1 U10950 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9787) );
  AOI22_X1 U10951 ( .A1(n9788), .A2(n9810), .B1(n9787), .B2(n9967), .ZN(
        P1_U3492) );
  OAI21_X1 U10952 ( .B1(n9790), .B2(n9799), .A(n9789), .ZN(n9791) );
  AOI21_X1 U10953 ( .B1(n9793), .B2(n9792), .A(n9791), .ZN(n9794) );
  AND2_X1 U10954 ( .A1(n9795), .A2(n9794), .ZN(n9813) );
  AOI22_X1 U10955 ( .A1(n9788), .A2(n9813), .B1(n6259), .B2(n9967), .ZN(
        P1_U3495) );
  AOI22_X1 U10956 ( .A1(n9814), .A2(n9796), .B1(n6640), .B2(n9811), .ZN(
        P1_U3523) );
  AOI22_X1 U10957 ( .A1(n9814), .A2(n9797), .B1(n6639), .B2(n9811), .ZN(
        P1_U3524) );
  OAI21_X1 U10958 ( .B1(n9800), .B2(n9799), .A(n9798), .ZN(n9801) );
  AOI21_X1 U10959 ( .B1(n9803), .B2(n9802), .A(n9801), .ZN(n9805) );
  AND2_X1 U10960 ( .A1(n9805), .A2(n9804), .ZN(n9966) );
  AOI22_X1 U10961 ( .A1(n9814), .A2(n9966), .B1(n6638), .B2(n9811), .ZN(
        P1_U3525) );
  AOI22_X1 U10962 ( .A1(n9814), .A2(n9806), .B1(n6068), .B2(n9811), .ZN(
        P1_U3526) );
  AOI22_X1 U10963 ( .A1(n9814), .A2(n9807), .B1(n6674), .B2(n9811), .ZN(
        P1_U3530) );
  AOI22_X1 U10964 ( .A1(n9814), .A2(n9808), .B1(n6739), .B2(n9811), .ZN(
        P1_U3532) );
  AOI22_X1 U10965 ( .A1(n9814), .A2(n9809), .B1(n6222), .B2(n9811), .ZN(
        P1_U3534) );
  AOI22_X1 U10966 ( .A1(n9814), .A2(n9810), .B1(n6955), .B2(n9811), .ZN(
        P1_U3535) );
  AOI22_X1 U10967 ( .A1(n9814), .A2(n9813), .B1(n9812), .B2(n9811), .ZN(
        P1_U3536) );
  AOI21_X1 U10968 ( .B1(n9817), .B2(n9816), .A(n9815), .ZN(n9826) );
  NAND2_X1 U10969 ( .A1(n9819), .A2(n9818), .ZN(n9825) );
  OAI211_X1 U10970 ( .C1(n9823), .C2(n9822), .A(n9821), .B(n9820), .ZN(n9824)
         );
  OAI211_X1 U10971 ( .C1(n9826), .C2(n9846), .A(n9825), .B(n9824), .ZN(n9827)
         );
  AOI21_X1 U10972 ( .B1(n9850), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n9827), .ZN(
        n9834) );
  INV_X1 U10973 ( .A(n9828), .ZN(n9832) );
  AND2_X1 U10974 ( .A1(n9829), .A2(n7125), .ZN(n9831) );
  OAI21_X1 U10975 ( .B1(n9832), .B2(n9831), .A(n9830), .ZN(n9833) );
  OAI211_X1 U10976 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7015), .A(n9834), .B(
        n9833), .ZN(P2_U3183) );
  XOR2_X1 U10977 ( .A(n9836), .B(n9835), .Z(n9838) );
  NOR2_X1 U10978 ( .A1(n9838), .A2(n9837), .ZN(n9849) );
  AOI21_X1 U10979 ( .B1(n9841), .B2(n9840), .A(n9839), .ZN(n9847) );
  AOI21_X1 U10980 ( .B1(n4501), .B2(n9843), .A(n9842), .ZN(n9845) );
  OAI22_X1 U10981 ( .A1(n9847), .A2(n9846), .B1(n9845), .B2(n9844), .ZN(n9848)
         );
  AOI211_X1 U10982 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n9850), .A(n9849), .B(
        n9848), .ZN(n9853) );
  INV_X1 U10983 ( .A(n9851), .ZN(n9852) );
  OAI211_X1 U10984 ( .C1(n9855), .C2(n9854), .A(n9853), .B(n9852), .ZN(
        P2_U3190) );
  OAI21_X1 U10985 ( .B1(n9857), .B2(n5655), .A(n9856), .ZN(n9885) );
  OAI22_X1 U10986 ( .A1(n9860), .A2(n9859), .B1(n9882), .B2(n9858), .ZN(n9870)
         );
  XNOR2_X1 U10987 ( .A(n9861), .B(n5655), .ZN(n9868) );
  INV_X1 U10988 ( .A(n9862), .ZN(n9880) );
  OAI22_X1 U10989 ( .A1(n4640), .A2(n9865), .B1(n9864), .B2(n9863), .ZN(n9866)
         );
  AOI21_X1 U10990 ( .B1(n9885), .B2(n9880), .A(n9866), .ZN(n9867) );
  OAI21_X1 U10991 ( .B1(n9869), .B2(n9868), .A(n9867), .ZN(n9883) );
  AOI211_X1 U10992 ( .C1(n9871), .C2(n9885), .A(n9870), .B(n9883), .ZN(n9873)
         );
  AOI22_X1 U10993 ( .A1(n9874), .A2(n5263), .B1(n9873), .B2(n9872), .ZN(
        P2_U3231) );
  INV_X1 U10994 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9881) );
  INV_X1 U10995 ( .A(n9911), .ZN(n9886) );
  NAND2_X1 U10996 ( .A1(n9879), .A2(n9886), .ZN(n9875) );
  OAI21_X1 U10997 ( .B1(n9876), .B2(n9915), .A(n9875), .ZN(n9877) );
  AOI211_X1 U10998 ( .C1(n9880), .C2(n9879), .A(n9878), .B(n9877), .ZN(n9930)
         );
  AOI22_X1 U10999 ( .A1(n9929), .A2(n9881), .B1(n9930), .B2(n9928), .ZN(
        P2_U3393) );
  INV_X1 U11000 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9887) );
  NOR2_X1 U11001 ( .A1(n9882), .A2(n9915), .ZN(n9884) );
  AOI211_X1 U11002 ( .C1(n9886), .C2(n9885), .A(n9884), .B(n9883), .ZN(n9931)
         );
  AOI22_X1 U11003 ( .A1(n9929), .A2(n9887), .B1(n9931), .B2(n9928), .ZN(
        P2_U3396) );
  INV_X1 U11004 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9984) );
  NOR2_X1 U11005 ( .A1(n9888), .A2(n9915), .ZN(n9890) );
  AOI211_X1 U11006 ( .C1(n9920), .C2(n9891), .A(n9890), .B(n9889), .ZN(n9932)
         );
  AOI22_X1 U11007 ( .A1(n9929), .A2(n9984), .B1(n9932), .B2(n9928), .ZN(
        P2_U3399) );
  NOR2_X1 U11008 ( .A1(n9892), .A2(n9915), .ZN(n9894) );
  AOI211_X1 U11009 ( .C1(n9920), .C2(n9895), .A(n9894), .B(n9893), .ZN(n9933)
         );
  AOI22_X1 U11010 ( .A1(n9929), .A2(n5292), .B1(n9933), .B2(n9928), .ZN(
        P2_U3402) );
  NOR2_X1 U11011 ( .A1(n9896), .A2(n9915), .ZN(n9898) );
  AOI211_X1 U11012 ( .C1(n9920), .C2(n9899), .A(n9898), .B(n9897), .ZN(n9934)
         );
  AOI22_X1 U11013 ( .A1(n9929), .A2(n5320), .B1(n9934), .B2(n9928), .ZN(
        P2_U3408) );
  INV_X1 U11014 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9904) );
  OAI22_X1 U11015 ( .A1(n9901), .A2(n9911), .B1(n9900), .B2(n9915), .ZN(n9902)
         );
  NOR2_X1 U11016 ( .A1(n9903), .A2(n9902), .ZN(n9935) );
  AOI22_X1 U11017 ( .A1(n9929), .A2(n9904), .B1(n9935), .B2(n9928), .ZN(
        P2_U3411) );
  OAI22_X1 U11018 ( .A1(n9906), .A2(n9922), .B1(n9905), .B2(n9915), .ZN(n9907)
         );
  INV_X1 U11019 ( .A(n9907), .ZN(n9909) );
  AND2_X1 U11020 ( .A1(n9909), .A2(n9908), .ZN(n9936) );
  AOI22_X1 U11021 ( .A1(n9929), .A2(n5349), .B1(n9936), .B2(n9928), .ZN(
        P2_U3414) );
  OAI22_X1 U11022 ( .A1(n9912), .A2(n9911), .B1(n9910), .B2(n9915), .ZN(n9913)
         );
  NOR2_X1 U11023 ( .A1(n9914), .A2(n9913), .ZN(n9937) );
  AOI22_X1 U11024 ( .A1(n9929), .A2(n5378), .B1(n9937), .B2(n9928), .ZN(
        P2_U3420) );
  INV_X1 U11025 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9921) );
  NOR2_X1 U11026 ( .A1(n9916), .A2(n9915), .ZN(n9918) );
  AOI211_X1 U11027 ( .C1(n9920), .C2(n9919), .A(n9918), .B(n9917), .ZN(n9938)
         );
  AOI22_X1 U11028 ( .A1(n9929), .A2(n9921), .B1(n9938), .B2(n9928), .ZN(
        P2_U3423) );
  INV_X1 U11029 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10175) );
  NOR2_X1 U11030 ( .A1(n9923), .A2(n9922), .ZN(n9925) );
  AOI211_X1 U11031 ( .C1(n9927), .C2(n9926), .A(n9925), .B(n9924), .ZN(n9940)
         );
  AOI22_X1 U11032 ( .A1(n9929), .A2(n10175), .B1(n9940), .B2(n9928), .ZN(
        P2_U3426) );
  AOI22_X1 U11033 ( .A1(n9941), .A2(n9930), .B1(n7125), .B2(n9939), .ZN(
        P2_U3460) );
  AOI22_X1 U11034 ( .A1(n9941), .A2(n9931), .B1(n5264), .B2(n9939), .ZN(
        P2_U3461) );
  AOI22_X1 U11035 ( .A1(n9941), .A2(n9932), .B1(n5277), .B2(n9939), .ZN(
        P2_U3462) );
  AOI22_X1 U11036 ( .A1(n9941), .A2(n9933), .B1(n5294), .B2(n9939), .ZN(
        P2_U3463) );
  AOI22_X1 U11037 ( .A1(n9941), .A2(n9934), .B1(n7248), .B2(n9939), .ZN(
        P2_U3465) );
  AOI22_X1 U11038 ( .A1(n9941), .A2(n9935), .B1(n5337), .B2(n9939), .ZN(
        P2_U3466) );
  AOI22_X1 U11039 ( .A1(n9941), .A2(n9936), .B1(n7368), .B2(n9939), .ZN(
        P2_U3467) );
  AOI22_X1 U11040 ( .A1(n9941), .A2(n9937), .B1(n7451), .B2(n9939), .ZN(
        P2_U3469) );
  AOI22_X1 U11041 ( .A1(n9941), .A2(n9938), .B1(n5397), .B2(n9939), .ZN(
        P2_U3470) );
  AOI22_X1 U11042 ( .A1(n9941), .A2(n9940), .B1(n7714), .B2(n9939), .ZN(
        P2_U3471) );
  NOR2_X1 U11043 ( .A1(n9943), .A2(n9942), .ZN(n9944) );
  XOR2_X1 U11044 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9944), .Z(ADD_1068_U5) );
  AOI21_X1 U11045 ( .B1(n9946), .B2(n10013), .A(n9945), .ZN(ADD_1068_U46) );
  OAI21_X1 U11046 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9948), .A(n9947), .ZN(
        n9949) );
  XNOR2_X1 U11047 ( .A(n9949), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  XNOR2_X1 U11048 ( .A(n9951), .B(n9950), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11049 ( .A(n9953), .B(n9952), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11050 ( .A(n9955), .B(n9954), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11051 ( .A(n9957), .B(n9956), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11052 ( .A(n9959), .B(n9958), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11053 ( .A(n9961), .B(n9960), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11054 ( .A(n9963), .B(n9962), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11055 ( .A(n9965), .B(n9964), .ZN(ADD_1068_U63) );
  INV_X1 U11056 ( .A(n9966), .ZN(n9968) );
  AOI22_X1 U11057 ( .A1(n9788), .A2(n9968), .B1(P1_REG0_REG_3__SCAN_IN), .B2(
        n9967), .ZN(n10281) );
  AOI22_X1 U11058 ( .A1(n9971), .A2(keyinput50), .B1(keyinput64), .B2(n9970), 
        .ZN(n9969) );
  OAI221_X1 U11059 ( .B1(n9971), .B2(keyinput50), .C1(n9970), .C2(keyinput64), 
        .A(n9969), .ZN(n9982) );
  AOI22_X1 U11060 ( .A1(n9973), .A2(keyinput114), .B1(keyinput51), .B2(n7471), 
        .ZN(n9972) );
  OAI221_X1 U11061 ( .B1(n9973), .B2(keyinput114), .C1(n7471), .C2(keyinput51), 
        .A(n9972), .ZN(n9981) );
  AOI22_X1 U11062 ( .A1(n9976), .A2(keyinput6), .B1(n9975), .B2(keyinput54), 
        .ZN(n9974) );
  OAI221_X1 U11063 ( .B1(n9976), .B2(keyinput6), .C1(n9975), .C2(keyinput54), 
        .A(n9974), .ZN(n9980) );
  XNOR2_X1 U11064 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput66), .ZN(n9978) );
  XNOR2_X1 U11065 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput11), .ZN(n9977) );
  NAND2_X1 U11066 ( .A1(n9978), .A2(n9977), .ZN(n9979) );
  NOR4_X1 U11067 ( .A1(n9982), .A2(n9981), .A3(n9980), .A4(n9979), .ZN(n10279)
         );
  AOI22_X1 U11068 ( .A1(n9984), .A2(keyinput125), .B1(keyinput47), .B2(n6217), 
        .ZN(n9983) );
  OAI221_X1 U11069 ( .B1(n9984), .B2(keyinput125), .C1(n6217), .C2(keyinput47), 
        .A(n9983), .ZN(n9994) );
  AOI22_X1 U11070 ( .A1(n9986), .A2(keyinput92), .B1(keyinput127), .B2(n5349), 
        .ZN(n9985) );
  OAI221_X1 U11071 ( .B1(n9986), .B2(keyinput92), .C1(n5349), .C2(keyinput127), 
        .A(n9985), .ZN(n9993) );
  AOI22_X1 U11072 ( .A1(n9988), .A2(keyinput82), .B1(n5378), .B2(keyinput41), 
        .ZN(n9987) );
  OAI221_X1 U11073 ( .B1(n9988), .B2(keyinput82), .C1(n5378), .C2(keyinput41), 
        .A(n9987), .ZN(n9992) );
  XNOR2_X1 U11074 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput17), .ZN(n9990) );
  XNOR2_X1 U11075 ( .A(P1_REG3_REG_26__SCAN_IN), .B(keyinput49), .ZN(n9989) );
  NAND2_X1 U11076 ( .A1(n9990), .A2(n9989), .ZN(n9991) );
  NOR4_X1 U11077 ( .A1(n9994), .A2(n9993), .A3(n9992), .A4(n9991), .ZN(n10278)
         );
  AOI22_X1 U11078 ( .A1(n9997), .A2(keyinput73), .B1(keyinput106), .B2(n9996), 
        .ZN(n9995) );
  OAI221_X1 U11079 ( .B1(n9997), .B2(keyinput73), .C1(n9996), .C2(keyinput106), 
        .A(n9995), .ZN(n10090) );
  AOI22_X1 U11080 ( .A1(n9999), .A2(keyinput75), .B1(keyinput90), .B2(n8685), 
        .ZN(n9998) );
  OAI221_X1 U11081 ( .B1(n9999), .B2(keyinput75), .C1(n8685), .C2(keyinput90), 
        .A(n9998), .ZN(n10089) );
  INV_X1 U11082 ( .A(keyinput9), .ZN(n10023) );
  XNOR2_X1 U11083 ( .A(n10000), .B(keyinput76), .ZN(n10005) );
  XNOR2_X1 U11084 ( .A(n10001), .B(keyinput15), .ZN(n10004) );
  INV_X1 U11085 ( .A(keyinput119), .ZN(n10002) );
  MUX2_X1 U11086 ( .A(keyinput119), .B(n10002), .S(P2_DATAO_REG_15__SCAN_IN), 
        .Z(n10003) );
  NOR3_X1 U11087 ( .A1(n10005), .A2(n10004), .A3(n10003), .ZN(n10022) );
  INV_X1 U11088 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10007) );
  AOI22_X1 U11089 ( .A1(n10008), .A2(keyinput109), .B1(keyinput4), .B2(n10007), 
        .ZN(n10006) );
  OAI221_X1 U11090 ( .B1(n10008), .B2(keyinput109), .C1(n10007), .C2(keyinput4), .A(n10006), .ZN(n10020) );
  AOI22_X1 U11091 ( .A1(n10010), .A2(keyinput28), .B1(keyinput63), .B2(n6633), 
        .ZN(n10009) );
  OAI221_X1 U11092 ( .B1(n10010), .B2(keyinput28), .C1(n6633), .C2(keyinput63), 
        .A(n10009), .ZN(n10019) );
  AOI22_X1 U11093 ( .A1(n10013), .A2(keyinput126), .B1(n10012), .B2(keyinput34), .ZN(n10011) );
  OAI221_X1 U11094 ( .B1(n10013), .B2(keyinput126), .C1(n10012), .C2(
        keyinput34), .A(n10011), .ZN(n10018) );
  AOI22_X1 U11095 ( .A1(n10016), .A2(keyinput118), .B1(n10015), .B2(keyinput61), .ZN(n10014) );
  OAI221_X1 U11096 ( .B1(n10016), .B2(keyinput118), .C1(n10015), .C2(
        keyinput61), .A(n10014), .ZN(n10017) );
  NOR4_X1 U11097 ( .A1(n10020), .A2(n10019), .A3(n10018), .A4(n10017), .ZN(
        n10021) );
  OAI211_X1 U11098 ( .C1(P1_REG3_REG_25__SCAN_IN), .C2(n10023), .A(n10022), 
        .B(n10021), .ZN(n10088) );
  INV_X1 U11099 ( .A(P2_B_REG_SCAN_IN), .ZN(n10026) );
  AOI22_X1 U11100 ( .A1(n10026), .A2(keyinput24), .B1(keyinput36), .B2(n10025), 
        .ZN(n10024) );
  OAI221_X1 U11101 ( .B1(n10026), .B2(keyinput24), .C1(n10025), .C2(keyinput36), .A(n10024), .ZN(n10031) );
  XNOR2_X1 U11102 ( .A(n10027), .B(keyinput97), .ZN(n10030) );
  XNOR2_X1 U11103 ( .A(n10028), .B(keyinput67), .ZN(n10029) );
  OR3_X1 U11104 ( .A1(n10031), .A2(n10030), .A3(n10029), .ZN(n10039) );
  AOI22_X1 U11105 ( .A1(n10033), .A2(keyinput14), .B1(keyinput96), .B2(n9427), 
        .ZN(n10032) );
  OAI221_X1 U11106 ( .B1(n10033), .B2(keyinput14), .C1(n9427), .C2(keyinput96), 
        .A(n10032), .ZN(n10038) );
  INV_X1 U11107 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n10036) );
  AOI22_X1 U11108 ( .A1(n10036), .A2(keyinput13), .B1(keyinput68), .B2(n10035), 
        .ZN(n10034) );
  OAI221_X1 U11109 ( .B1(n10036), .B2(keyinput13), .C1(n10035), .C2(keyinput68), .A(n10034), .ZN(n10037) );
  NOR3_X1 U11110 ( .A1(n10039), .A2(n10038), .A3(n10037), .ZN(n10086) );
  AOI22_X1 U11111 ( .A1(n10042), .A2(keyinput101), .B1(keyinput78), .B2(n10041), .ZN(n10040) );
  OAI221_X1 U11112 ( .B1(n10042), .B2(keyinput101), .C1(n10041), .C2(
        keyinput78), .A(n10040), .ZN(n10053) );
  AOI22_X1 U11113 ( .A1(n10045), .A2(keyinput33), .B1(n10044), .B2(keyinput30), 
        .ZN(n10043) );
  OAI221_X1 U11114 ( .B1(n10045), .B2(keyinput33), .C1(n10044), .C2(keyinput30), .A(n10043), .ZN(n10052) );
  INV_X1 U11115 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10046) );
  XOR2_X1 U11116 ( .A(n10046), .B(keyinput107), .Z(n10050) );
  XNOR2_X1 U11117 ( .A(keyinput46), .B(P1_REG0_REG_9__SCAN_IN), .ZN(n10049) );
  XNOR2_X1 U11118 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput25), .ZN(n10048) );
  XNOR2_X1 U11119 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput77), .ZN(n10047) );
  NAND4_X1 U11120 ( .A1(n10050), .A2(n10049), .A3(n10048), .A4(n10047), .ZN(
        n10051) );
  NOR3_X1 U11121 ( .A1(n10053), .A2(n10052), .A3(n10051), .ZN(n10085) );
  INV_X1 U11122 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n10055) );
  AOI22_X1 U11123 ( .A1(n10056), .A2(keyinput38), .B1(keyinput22), .B2(n10055), 
        .ZN(n10054) );
  OAI221_X1 U11124 ( .B1(n10056), .B2(keyinput38), .C1(n10055), .C2(keyinput22), .A(n10054), .ZN(n10066) );
  AOI22_X1 U11125 ( .A1(n8518), .A2(keyinput1), .B1(n5043), .B2(keyinput98), 
        .ZN(n10057) );
  OAI221_X1 U11126 ( .B1(n8518), .B2(keyinput1), .C1(n5043), .C2(keyinput98), 
        .A(n10057), .ZN(n10065) );
  AOI22_X1 U11127 ( .A1(n10060), .A2(keyinput93), .B1(keyinput88), .B2(n10059), 
        .ZN(n10058) );
  OAI221_X1 U11128 ( .B1(n10060), .B2(keyinput93), .C1(n10059), .C2(keyinput88), .A(n10058), .ZN(n10064) );
  XNOR2_X1 U11129 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput89), .ZN(n10062) );
  XNOR2_X1 U11130 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput56), .ZN(n10061)
         );
  NAND2_X1 U11131 ( .A1(n10062), .A2(n10061), .ZN(n10063) );
  NOR4_X1 U11132 ( .A1(n10066), .A2(n10065), .A3(n10064), .A4(n10063), .ZN(
        n10084) );
  AOI22_X1 U11133 ( .A1(n10069), .A2(keyinput104), .B1(keyinput60), .B2(n10068), .ZN(n10067) );
  OAI221_X1 U11134 ( .B1(n10069), .B2(keyinput104), .C1(n10068), .C2(
        keyinput60), .A(n10067), .ZN(n10070) );
  INV_X1 U11135 ( .A(n10070), .ZN(n10082) );
  AOI22_X1 U11136 ( .A1(n9703), .A2(keyinput111), .B1(n10072), .B2(keyinput45), 
        .ZN(n10071) );
  OAI221_X1 U11137 ( .B1(n9703), .B2(keyinput111), .C1(n10072), .C2(keyinput45), .A(n10071), .ZN(n10073) );
  INV_X1 U11138 ( .A(n10073), .ZN(n10081) );
  XNOR2_X1 U11139 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput40), .ZN(n10076) );
  XNOR2_X1 U11140 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput53), .ZN(n10075) );
  XNOR2_X1 U11141 ( .A(keyinput74), .B(P1_REG0_REG_15__SCAN_IN), .ZN(n10074)
         );
  AND3_X1 U11142 ( .A1(n10076), .A2(n10075), .A3(n10074), .ZN(n10080) );
  INV_X1 U11143 ( .A(keyinput72), .ZN(n10077) );
  XNOR2_X1 U11144 ( .A(n10078), .B(n10077), .ZN(n10079) );
  AND4_X1 U11145 ( .A1(n10082), .A2(n10081), .A3(n10080), .A4(n10079), .ZN(
        n10083) );
  NAND4_X1 U11146 ( .A1(n10086), .A2(n10085), .A3(n10084), .A4(n10083), .ZN(
        n10087) );
  NOR4_X1 U11147 ( .A1(n10090), .A2(n10089), .A3(n10088), .A4(n10087), .ZN(
        n10277) );
  INV_X1 U11148 ( .A(keyinput15), .ZN(n10093) );
  INV_X1 U11149 ( .A(keyinput90), .ZN(n10091) );
  NAND4_X1 U11150 ( .A1(keyinput76), .A2(keyinput119), .A3(keyinput73), .A4(
        n10091), .ZN(n10092) );
  NOR4_X1 U11151 ( .A1(keyinput108), .A2(keyinput75), .A3(n10093), .A4(n10092), 
        .ZN(n10106) );
  NOR4_X1 U11152 ( .A1(keyinput63), .A2(keyinput109), .A3(keyinput61), .A4(
        keyinput126), .ZN(n10105) );
  NAND2_X1 U11153 ( .A1(keyinput4), .A2(keyinput28), .ZN(n10094) );
  NOR3_X1 U11154 ( .A1(keyinput106), .A2(keyinput118), .A3(n10094), .ZN(n10104) );
  INV_X1 U11155 ( .A(keyinput82), .ZN(n10095) );
  NAND4_X1 U11156 ( .A1(keyinput125), .A2(keyinput127), .A3(keyinput47), .A4(
        n10095), .ZN(n10102) );
  NOR2_X1 U11157 ( .A1(keyinput34), .A2(keyinput17), .ZN(n10096) );
  NAND3_X1 U11158 ( .A1(keyinput49), .A2(keyinput92), .A3(n10096), .ZN(n10101)
         );
  NOR2_X1 U11159 ( .A1(keyinput50), .A2(keyinput114), .ZN(n10097) );
  NAND3_X1 U11160 ( .A1(keyinput11), .A2(keyinput64), .A3(n10097), .ZN(n10100)
         );
  NOR3_X1 U11161 ( .A1(keyinput41), .A2(keyinput66), .A3(keyinput6), .ZN(
        n10098) );
  NAND2_X1 U11162 ( .A1(keyinput54), .A2(n10098), .ZN(n10099) );
  NOR4_X1 U11163 ( .A1(n10102), .A2(n10101), .A3(n10100), .A4(n10099), .ZN(
        n10103) );
  NAND4_X1 U11164 ( .A1(n10106), .A2(n10105), .A3(n10104), .A4(n10103), .ZN(
        n10157) );
  NAND2_X1 U11165 ( .A1(keyinput35), .A2(keyinput79), .ZN(n10107) );
  NOR3_X1 U11166 ( .A1(keyinput27), .A2(keyinput110), .A3(n10107), .ZN(n10155)
         );
  NAND2_X1 U11167 ( .A1(keyinput21), .A2(keyinput58), .ZN(n10108) );
  NOR3_X1 U11168 ( .A1(keyinput43), .A2(keyinput48), .A3(n10108), .ZN(n10154)
         );
  NAND4_X1 U11169 ( .A1(keyinput123), .A2(keyinput26), .A3(keyinput70), .A4(
        keyinput71), .ZN(n10119) );
  INV_X1 U11170 ( .A(keyinput23), .ZN(n10109) );
  NAND4_X1 U11171 ( .A1(keyinput122), .A2(keyinput120), .A3(keyinput65), .A4(
        n10109), .ZN(n10118) );
  NAND2_X1 U11172 ( .A1(keyinput86), .A2(keyinput16), .ZN(n10110) );
  NOR3_X1 U11173 ( .A1(keyinput52), .A2(keyinput91), .A3(n10110), .ZN(n10116)
         );
  INV_X1 U11174 ( .A(keyinput29), .ZN(n10111) );
  NOR4_X1 U11175 ( .A1(keyinput12), .A2(keyinput3), .A3(keyinput87), .A4(
        n10111), .ZN(n10115) );
  NAND2_X1 U11176 ( .A1(keyinput32), .A2(keyinput113), .ZN(n10112) );
  NOR3_X1 U11177 ( .A1(keyinput18), .A2(keyinput81), .A3(n10112), .ZN(n10114)
         );
  NOR4_X1 U11178 ( .A1(keyinput31), .A2(keyinput0), .A3(keyinput94), .A4(
        keyinput59), .ZN(n10113) );
  NAND4_X1 U11179 ( .A1(n10116), .A2(n10115), .A3(n10114), .A4(n10113), .ZN(
        n10117) );
  NOR3_X1 U11180 ( .A1(n10119), .A2(n10118), .A3(n10117), .ZN(n10153) );
  NAND2_X1 U11181 ( .A1(keyinput72), .A2(keyinput111), .ZN(n10120) );
  NOR3_X1 U11182 ( .A1(keyinput74), .A2(keyinput45), .A3(n10120), .ZN(n10126)
         );
  INV_X1 U11183 ( .A(keyinput104), .ZN(n10121) );
  NOR4_X1 U11184 ( .A1(keyinput68), .A2(keyinput60), .A3(keyinput40), .A4(
        n10121), .ZN(n10125) );
  NOR4_X1 U11185 ( .A1(keyinput22), .A2(keyinput1), .A3(keyinput88), .A4(
        keyinput56), .ZN(n10124) );
  NAND3_X1 U11186 ( .A1(keyinput93), .A2(keyinput98), .A3(keyinput53), .ZN(
        n10122) );
  NOR2_X1 U11187 ( .A1(keyinput38), .A2(n10122), .ZN(n10123) );
  NAND4_X1 U11188 ( .A1(n10126), .A2(n10125), .A3(n10124), .A4(n10123), .ZN(
        n10151) );
  INV_X1 U11189 ( .A(keyinput107), .ZN(n10127) );
  NOR4_X1 U11190 ( .A1(keyinput46), .A2(keyinput77), .A3(keyinput101), .A4(
        n10127), .ZN(n10133) );
  NOR4_X1 U11191 ( .A1(keyinput51), .A2(keyinput33), .A3(keyinput30), .A4(
        keyinput25), .ZN(n10132) );
  NAND2_X1 U11192 ( .A1(keyinput36), .A2(keyinput24), .ZN(n10128) );
  NOR3_X1 U11193 ( .A1(keyinput97), .A2(keyinput13), .A3(n10128), .ZN(n10131)
         );
  NAND2_X1 U11194 ( .A1(keyinput96), .A2(keyinput78), .ZN(n10129) );
  NOR3_X1 U11195 ( .A1(keyinput14), .A2(keyinput67), .A3(n10129), .ZN(n10130)
         );
  NAND4_X1 U11196 ( .A1(n10133), .A2(n10132), .A3(n10131), .A4(n10130), .ZN(
        n10150) );
  NOR2_X1 U11197 ( .A1(keyinput116), .A2(keyinput85), .ZN(n10134) );
  NAND3_X1 U11198 ( .A1(keyinput2), .A2(keyinput57), .A3(n10134), .ZN(n10140)
         );
  INV_X1 U11199 ( .A(keyinput8), .ZN(n10135) );
  NAND4_X1 U11200 ( .A1(keyinput69), .A2(keyinput80), .A3(keyinput99), .A4(
        n10135), .ZN(n10139) );
  NAND4_X1 U11201 ( .A1(keyinput44), .A2(keyinput20), .A3(keyinput19), .A4(
        keyinput7), .ZN(n10138) );
  NOR2_X1 U11202 ( .A1(keyinput124), .A2(keyinput117), .ZN(n10136) );
  NAND3_X1 U11203 ( .A1(keyinput100), .A2(keyinput95), .A3(n10136), .ZN(n10137) );
  OR4_X1 U11204 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(
        n10149) );
  NAND2_X1 U11205 ( .A1(keyinput105), .A2(keyinput62), .ZN(n10141) );
  NOR3_X1 U11206 ( .A1(keyinput83), .A2(keyinput102), .A3(n10141), .ZN(n10147)
         );
  INV_X1 U11207 ( .A(keyinput103), .ZN(n10142) );
  NOR4_X1 U11208 ( .A1(keyinput89), .A2(keyinput39), .A3(keyinput121), .A4(
        n10142), .ZN(n10146) );
  NAND2_X1 U11209 ( .A1(keyinput37), .A2(keyinput5), .ZN(n10143) );
  NOR3_X1 U11210 ( .A1(keyinput84), .A2(keyinput55), .A3(n10143), .ZN(n10145)
         );
  NOR4_X1 U11211 ( .A1(keyinput42), .A2(keyinput112), .A3(keyinput10), .A4(
        keyinput115), .ZN(n10144) );
  NAND4_X1 U11212 ( .A1(n10147), .A2(n10146), .A3(n10145), .A4(n10144), .ZN(
        n10148) );
  NOR4_X1 U11213 ( .A1(n10151), .A2(n10150), .A3(n10149), .A4(n10148), .ZN(
        n10152) );
  NAND4_X1 U11214 ( .A1(n10155), .A2(n10154), .A3(n10153), .A4(n10152), .ZN(
        n10156) );
  OAI21_X1 U11215 ( .B1(n10157), .B2(n10156), .A(keyinput9), .ZN(n10275) );
  AOI22_X1 U11216 ( .A1(n10160), .A2(keyinput105), .B1(n10159), .B2(keyinput69), .ZN(n10158) );
  OAI221_X1 U11217 ( .B1(n10160), .B2(keyinput105), .C1(n10159), .C2(
        keyinput69), .A(n10158), .ZN(n10169) );
  AOI22_X1 U11218 ( .A1(n6009), .A2(keyinput62), .B1(n5264), .B2(keyinput102), 
        .ZN(n10161) );
  OAI221_X1 U11219 ( .B1(n6009), .B2(keyinput62), .C1(n5264), .C2(keyinput102), 
        .A(n10161), .ZN(n10168) );
  AOI22_X1 U11220 ( .A1(n6168), .A2(keyinput121), .B1(n10163), .B2(keyinput83), 
        .ZN(n10162) );
  OAI221_X1 U11221 ( .B1(n6168), .B2(keyinput121), .C1(n10163), .C2(keyinput83), .A(n10162), .ZN(n10167) );
  XNOR2_X1 U11222 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput39), .ZN(n10165)
         );
  XNOR2_X1 U11223 ( .A(P1_REG3_REG_15__SCAN_IN), .B(keyinput103), .ZN(n10164)
         );
  NAND2_X1 U11224 ( .A1(n10165), .A2(n10164), .ZN(n10166) );
  NOR4_X1 U11225 ( .A1(n10169), .A2(n10168), .A3(n10167), .A4(n10166), .ZN(
        n10215) );
  AOI22_X1 U11226 ( .A1(n10171), .A2(keyinput8), .B1(n5210), .B2(keyinput80), 
        .ZN(n10170) );
  OAI221_X1 U11227 ( .B1(n10171), .B2(keyinput8), .C1(n5210), .C2(keyinput80), 
        .A(n10170), .ZN(n10182) );
  AOI22_X1 U11228 ( .A1(n10173), .A2(keyinput99), .B1(keyinput116), .B2(n8872), 
        .ZN(n10172) );
  OAI221_X1 U11229 ( .B1(n10173), .B2(keyinput99), .C1(n8872), .C2(keyinput116), .A(n10172), .ZN(n10181) );
  AOI22_X1 U11230 ( .A1(n10175), .A2(keyinput2), .B1(keyinput85), .B2(P1_U3086), .ZN(n10174) );
  OAI221_X1 U11231 ( .B1(n10175), .B2(keyinput2), .C1(P1_U3086), .C2(
        keyinput85), .A(n10174), .ZN(n10180) );
  INV_X1 U11232 ( .A(keyinput124), .ZN(n10177) );
  AOI22_X1 U11233 ( .A1(n10178), .A2(keyinput57), .B1(P2_WR_REG_SCAN_IN), .B2(
        n10177), .ZN(n10176) );
  OAI221_X1 U11234 ( .B1(n10178), .B2(keyinput57), .C1(n10177), .C2(
        P2_WR_REG_SCAN_IN), .A(n10176), .ZN(n10179) );
  NOR4_X1 U11235 ( .A1(n10182), .A2(n10181), .A3(n10180), .A4(n10179), .ZN(
        n10214) );
  AOI22_X1 U11236 ( .A1(n10185), .A2(keyinput20), .B1(keyinput95), .B2(n10184), 
        .ZN(n10183) );
  OAI221_X1 U11237 ( .B1(n10185), .B2(keyinput20), .C1(n10184), .C2(keyinput95), .A(n10183), .ZN(n10192) );
  AOI22_X1 U11238 ( .A1(n10188), .A2(keyinput7), .B1(n10187), .B2(keyinput42), 
        .ZN(n10186) );
  OAI221_X1 U11239 ( .B1(n10188), .B2(keyinput7), .C1(n10187), .C2(keyinput42), 
        .A(n10186), .ZN(n10191) );
  XNOR2_X1 U11240 ( .A(n10189), .B(keyinput100), .ZN(n10190) );
  OR3_X1 U11241 ( .A1(n10192), .A2(n10191), .A3(n10190), .ZN(n10199) );
  AOI22_X1 U11242 ( .A1(n10195), .A2(keyinput117), .B1(keyinput19), .B2(n10194), .ZN(n10193) );
  OAI221_X1 U11243 ( .B1(n10195), .B2(keyinput117), .C1(n10194), .C2(
        keyinput19), .A(n10193), .ZN(n10198) );
  XNOR2_X1 U11244 ( .A(n10196), .B(keyinput44), .ZN(n10197) );
  NOR3_X1 U11245 ( .A1(n10199), .A2(n10198), .A3(n10197), .ZN(n10213) );
  AOI22_X1 U11246 ( .A1(n10201), .A2(keyinput37), .B1(keyinput58), .B2(n8226), 
        .ZN(n10200) );
  OAI221_X1 U11247 ( .B1(n10201), .B2(keyinput37), .C1(n8226), .C2(keyinput58), 
        .A(n10200), .ZN(n10211) );
  AOI22_X1 U11248 ( .A1(n10203), .A2(keyinput115), .B1(keyinput84), .B2(n6290), 
        .ZN(n10202) );
  OAI221_X1 U11249 ( .B1(n10203), .B2(keyinput115), .C1(n6290), .C2(keyinput84), .A(n10202), .ZN(n10210) );
  INV_X1 U11250 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10205) );
  AOI22_X1 U11251 ( .A1(n10205), .A2(keyinput112), .B1(keyinput10), .B2(n5995), 
        .ZN(n10204) );
  OAI221_X1 U11252 ( .B1(n10205), .B2(keyinput112), .C1(n5995), .C2(keyinput10), .A(n10204), .ZN(n10209) );
  XNOR2_X1 U11253 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput5), .ZN(n10207) );
  XNOR2_X1 U11254 ( .A(P1_REG3_REG_2__SCAN_IN), .B(keyinput55), .ZN(n10206) );
  NAND2_X1 U11255 ( .A1(n10207), .A2(n10206), .ZN(n10208) );
  NOR4_X1 U11256 ( .A1(n10211), .A2(n10210), .A3(n10209), .A4(n10208), .ZN(
        n10212) );
  NAND4_X1 U11257 ( .A1(n10215), .A2(n10214), .A3(n10213), .A4(n10212), .ZN(
        n10274) );
  AOI22_X1 U11258 ( .A1(n5985), .A2(keyinput110), .B1(keyinput120), .B2(n10217), .ZN(n10216) );
  OAI221_X1 U11259 ( .B1(n5985), .B2(keyinput110), .C1(n10217), .C2(
        keyinput120), .A(n10216), .ZN(n10228) );
  AOI22_X1 U11260 ( .A1(n10219), .A2(keyinput79), .B1(keyinput35), .B2(n5009), 
        .ZN(n10218) );
  OAI221_X1 U11261 ( .B1(n10219), .B2(keyinput79), .C1(n5009), .C2(keyinput35), 
        .A(n10218), .ZN(n10227) );
  INV_X1 U11262 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10222) );
  AOI22_X1 U11263 ( .A1(n10222), .A2(keyinput48), .B1(keyinput27), .B2(n10221), 
        .ZN(n10220) );
  OAI221_X1 U11264 ( .B1(n10222), .B2(keyinput48), .C1(n10221), .C2(keyinput27), .A(n10220), .ZN(n10226) );
  XOR2_X1 U11265 ( .A(n6520), .B(keyinput21), .Z(n10224) );
  XNOR2_X1 U11266 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput43), .ZN(n10223) );
  NAND2_X1 U11267 ( .A1(n10224), .A2(n10223), .ZN(n10225) );
  NOR4_X1 U11268 ( .A1(n10228), .A2(n10227), .A3(n10226), .A4(n10225), .ZN(
        n10272) );
  INV_X1 U11269 ( .A(SI_18_), .ZN(n10230) );
  AOI22_X1 U11270 ( .A1(n10230), .A2(keyinput122), .B1(keyinput23), .B2(n6227), 
        .ZN(n10229) );
  OAI221_X1 U11271 ( .B1(n10230), .B2(keyinput122), .C1(n6227), .C2(keyinput23), .A(n10229), .ZN(n10241) );
  AOI22_X1 U11272 ( .A1(n10233), .A2(keyinput65), .B1(n10232), .B2(keyinput123), .ZN(n10231) );
  OAI221_X1 U11273 ( .B1(n10233), .B2(keyinput65), .C1(n10232), .C2(
        keyinput123), .A(n10231), .ZN(n10240) );
  XOR2_X1 U11274 ( .A(n10234), .B(keyinput70), .Z(n10238) );
  XOR2_X1 U11275 ( .A(n9603), .B(keyinput71), .Z(n10237) );
  XNOR2_X1 U11276 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput26), .ZN(n10236) );
  XNOR2_X1 U11277 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput12), .ZN(n10235) );
  NAND4_X1 U11278 ( .A1(n10238), .A2(n10237), .A3(n10236), .A4(n10235), .ZN(
        n10239) );
  NOR3_X1 U11279 ( .A1(n10241), .A2(n10240), .A3(n10239), .ZN(n10271) );
  AOI22_X1 U11280 ( .A1(n5509), .A2(keyinput29), .B1(keyinput3), .B2(n10243), 
        .ZN(n10242) );
  OAI221_X1 U11281 ( .B1(n5509), .B2(keyinput29), .C1(n10243), .C2(keyinput3), 
        .A(n10242), .ZN(n10253) );
  AOI22_X1 U11282 ( .A1(n10246), .A2(keyinput87), .B1(n10245), .B2(keyinput52), 
        .ZN(n10244) );
  OAI221_X1 U11283 ( .B1(n10246), .B2(keyinput87), .C1(n10245), .C2(keyinput52), .A(n10244), .ZN(n10252) );
  XOR2_X1 U11284 ( .A(n6165), .B(keyinput31), .Z(n10250) );
  XNOR2_X1 U11285 ( .A(keyinput16), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n10249)
         );
  XNOR2_X1 U11286 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput91), .ZN(n10248) );
  XNOR2_X1 U11287 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput86), .ZN(n10247) );
  NAND4_X1 U11288 ( .A1(n10250), .A2(n10249), .A3(n10248), .A4(n10247), .ZN(
        n10251) );
  NOR3_X1 U11289 ( .A1(n10253), .A2(n10252), .A3(n10251), .ZN(n10270) );
  INV_X1 U11290 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U11291 ( .A1(n10256), .A2(keyinput108), .B1(n10255), .B2(keyinput59), .ZN(n10254) );
  OAI221_X1 U11292 ( .B1(n10256), .B2(keyinput108), .C1(n10255), .C2(
        keyinput59), .A(n10254), .ZN(n10260) );
  XNOR2_X1 U11293 ( .A(n10257), .B(keyinput0), .ZN(n10259) );
  XNOR2_X1 U11294 ( .A(n5003), .B(keyinput113), .ZN(n10258) );
  OR3_X1 U11295 ( .A1(n10260), .A2(n10259), .A3(n10258), .ZN(n10268) );
  AOI22_X1 U11296 ( .A1(n10263), .A2(keyinput81), .B1(keyinput94), .B2(n10262), 
        .ZN(n10261) );
  OAI221_X1 U11297 ( .B1(n10263), .B2(keyinput81), .C1(n10262), .C2(keyinput94), .A(n10261), .ZN(n10267) );
  AOI22_X1 U11298 ( .A1(n10265), .A2(keyinput18), .B1(n5292), .B2(keyinput32), 
        .ZN(n10264) );
  OAI221_X1 U11299 ( .B1(n10265), .B2(keyinput18), .C1(n5292), .C2(keyinput32), 
        .A(n10264), .ZN(n10266) );
  NOR3_X1 U11300 ( .A1(n10268), .A2(n10267), .A3(n10266), .ZN(n10269) );
  NAND4_X1 U11301 ( .A1(n10272), .A2(n10271), .A3(n10270), .A4(n10269), .ZN(
        n10273) );
  AOI211_X1 U11302 ( .C1(P1_REG3_REG_25__SCAN_IN), .C2(n10275), .A(n10274), 
        .B(n10273), .ZN(n10276) );
  NAND4_X1 U11303 ( .A1(n10279), .A2(n10278), .A3(n10277), .A4(n10276), .ZN(
        n10280) );
  XOR2_X1 U11304 ( .A(n10281), .B(n10280), .Z(P1_U3462) );
  XNOR2_X1 U11305 ( .A(n10283), .B(n10282), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11306 ( .A(n10285), .B(n10284), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11307 ( .A(n10287), .B(n10286), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11308 ( .A(n10289), .B(n10288), .ZN(ADD_1068_U48) );
  XNOR2_X1 U11309 ( .A(n10291), .B(n10290), .ZN(ADD_1068_U50) );
  XOR2_X1 U11310 ( .A(n10293), .B(n10292), .Z(ADD_1068_U54) );
  XOR2_X1 U11311 ( .A(n10295), .B(n10294), .Z(ADD_1068_U53) );
  XNOR2_X1 U11312 ( .A(n10297), .B(n10296), .ZN(ADD_1068_U52) );
  INV_X2 U5196 ( .A(n5288), .ZN(n5610) );
  BUF_X2 U6127 ( .A(n7847), .Z(n4526) );
  CLKBUF_X1 U4951 ( .A(n8704), .Z(n8821) );
  XNOR2_X1 U5116 ( .A(n5403), .B(n5402), .ZN(n6611) );
  XNOR2_X1 U5713 ( .A(n5846), .B(n5845), .ZN(n5921) );
endmodule

