

module b14_C_AntiSAT_k_128_9 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590;

  NOR2_X1 U2294 ( .A1(n2751), .A2(n4580), .ZN(n3606) );
  AND2_X1 U2295 ( .A1(n2059), .A2(n2274), .ZN(n2273) );
  INV_X1 U2296 ( .A(n2841), .ZN(n3225) );
  INV_X1 U2297 ( .A(n3226), .ZN(n3210) );
  OAI21_X1 U2298 ( .B1(n2918), .B2(n2917), .A(n2916), .ZN(n3250) );
  INV_X2 U2299 ( .A(n3198), .ZN(n3223) );
  INV_X2 U2300 ( .A(n2827), .ZN(n2841) );
  NOR2_X1 U2301 ( .A1(n2775), .A2(n2774), .ZN(n2780) );
  NAND2_X2 U2302 ( .A1(n3612), .A2(n4301), .ZN(n3613) );
  OAI21_X2 U2303 ( .B1(n3314), .B2(n3150), .A(n3149), .ZN(n3377) );
  NAND2_X2 U2304 ( .A1(n3144), .A2(n3143), .ZN(n3314) );
  NOR3_X2 U2305 ( .A1(n3911), .A2(n3146), .A3(n2115), .ZN(n2113) );
  OAI21_X2 U2306 ( .B1(n4498), .B2(n4174), .A(n4373), .ZN(n3619) );
  AOI21_X2 U2307 ( .B1(n4243), .B2(n3607), .A(n3606), .ZN(n4261) );
  OAI22_X2 U2308 ( .A1(n2877), .A2(n2876), .B1(n2875), .B2(n2874), .ZN(n2918)
         );
  OAI21_X2 U2309 ( .B1(n2239), .B2(n2780), .A(n2238), .ZN(n2877) );
  AND2_X2 U2310 ( .A1(n2785), .A2(STATE_REG_SCAN_IN), .ZN(n3403) );
  NAND4_X2 U2311 ( .A1(n2341), .A2(n2340), .A3(n2339), .A4(n2338), .ZN(n3919)
         );
  AND4_X1 U2312 ( .A1(n2354), .A2(n2353), .A3(n2352), .A4(n2351), .ZN(n2829)
         );
  INV_X2 U2313 ( .A(n2323), .ZN(n2708) );
  INV_X4 U2314 ( .A(n3222), .ZN(n2709) );
  INV_X4 U2315 ( .A(n4569), .ZN(n4548) );
  AND2_X4 U2316 ( .A1(n2673), .A2(n4235), .ZN(n2333) );
  OR2_X2 U2317 ( .A1(n2647), .A2(n3104), .ZN(n2783) );
  XNOR2_X1 U2318 ( .A(n2627), .B(n2626), .ZN(n3104) );
  NAND3_X2 U2319 ( .A1(n2313), .A2(n2312), .A3(n2311), .ZN(n2052) );
  AND2_X1 U2320 ( .A1(n2273), .A2(n2078), .ZN(n2111) );
  NAND2_X1 U2321 ( .A1(n3583), .A2(n3582), .ZN(n3581) );
  NAND2_X1 U2322 ( .A1(IR_REG_31__SCAN_IN), .A2(n2227), .ZN(n2330) );
  AND2_X1 U2323 ( .A1(n2277), .A2(n2190), .ZN(n2056) );
  AND4_X1 U2324 ( .A1(n2292), .A2(n2165), .A3(n2164), .A4(n2163), .ZN(n2059)
         );
  AND2_X1 U2325 ( .A1(n2582), .A2(n2293), .ZN(n2275) );
  NOR2_X1 U2326 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2289)
         );
  NOR2_X1 U2327 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2290)
         );
  INV_X1 U2328 ( .A(IR_REG_21__SCAN_IN), .ZN(n2582) );
  INV_X1 U2329 ( .A(IR_REG_3__SCAN_IN), .ZN(n2343) );
  INV_X1 U2330 ( .A(IR_REG_0__SCAN_IN), .ZN(n2228) );
  INV_X1 U2331 ( .A(IR_REG_1__SCAN_IN), .ZN(n2191) );
  NOR2_X1 U2332 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2288)
         );
  AOI21_X2 U2333 ( .B1(n4167), .B2(n4494), .A(n4394), .ZN(n4405) );
  NAND3_X2 U2334 ( .A1(n2313), .A2(n2312), .A3(n2311), .ZN(n2053) );
  NAND3_X1 U2335 ( .A1(n2313), .A2(n2312), .A3(n2311), .ZN(n2346) );
  AND2_X2 U2336 ( .A1(n2304), .A2(n2303), .ZN(n2337) );
  NOR2_X2 U2337 ( .A1(n4273), .A2(n4272), .ZN(n4271) );
  AOI21_X2 U2338 ( .B1(n4515), .B2(REG1_REG_5__SCAN_IN), .A(n4259), .ZN(n3608)
         );
  NAND2_X1 U2339 ( .A1(n3538), .A2(n3532), .ZN(n2187) );
  NAND2_X1 U2340 ( .A1(n2186), .A2(n3538), .ZN(n2185) );
  INV_X1 U2341 ( .A(n3535), .ZN(n2186) );
  AND2_X1 U2342 ( .A1(n3504), .A2(n3718), .ZN(n3538) );
  NAND2_X1 U2343 ( .A1(n2215), .A2(n2214), .ZN(n2213) );
  NAND2_X1 U2344 ( .A1(n3649), .A2(REG2_REG_15__SCAN_IN), .ZN(n2214) );
  NOR2_X1 U2345 ( .A1(n2161), .A2(n2159), .ZN(n2158) );
  INV_X1 U2346 ( .A(n2160), .ZN(n2159) );
  NOR2_X1 U2347 ( .A1(n2145), .A2(n2473), .ZN(n2143) );
  INV_X1 U2348 ( .A(n3429), .ZN(n2197) );
  INV_X1 U2349 ( .A(n2331), .ZN(n2815) );
  INV_X1 U2350 ( .A(IR_REG_17__SCAN_IN), .ZN(n2274) );
  NAND2_X1 U2351 ( .A1(n2705), .A2(n2596), .ZN(n4473) );
  INV_X1 U2352 ( .A(n2242), .ZN(n2241) );
  OAI21_X1 U2353 ( .B1(n2243), .B2(n3373), .A(n3159), .ZN(n2242) );
  OR2_X1 U2354 ( .A1(n3158), .A2(n3157), .ZN(n3159) );
  AND2_X1 U2355 ( .A1(n2570), .A2(n2569), .ZN(n3389) );
  NAND2_X1 U2356 ( .A1(n2333), .A2(REG3_REG_1__SCAN_IN), .ZN(n2307) );
  NAND2_X1 U2357 ( .A1(n2097), .A2(n2096), .ZN(n3579) );
  NAND2_X1 U2358 ( .A1(n2315), .A2(REG2_REG_1__SCAN_IN), .ZN(n2096) );
  OR2_X1 U2359 ( .A1(n2315), .A2(REG2_REG_1__SCAN_IN), .ZN(n2097) );
  NAND2_X1 U2360 ( .A1(n4306), .A2(n4305), .ZN(n4304) );
  NAND2_X1 U2361 ( .A1(n4324), .A2(n4325), .ZN(n4323) );
  XNOR2_X1 U2362 ( .A(n3643), .B(n4504), .ZN(n4336) );
  NAND2_X1 U2363 ( .A1(n4336), .A2(REG2_REG_12__SCAN_IN), .ZN(n4335) );
  INV_X1 U2364 ( .A(IR_REG_19__SCAN_IN), .ZN(n2584) );
  INV_X1 U2365 ( .A(n2130), .ZN(n3701) );
  AOI21_X1 U2366 ( .B1(n2127), .B2(n2125), .A(n2082), .ZN(n2124) );
  NAND2_X1 U2367 ( .A1(n2127), .A2(n2549), .ZN(n2126) );
  NOR2_X1 U2368 ( .A1(n2132), .A2(n2129), .ZN(n2128) );
  NOR2_X1 U2369 ( .A1(n2064), .A2(n2525), .ZN(n2129) );
  NAND2_X1 U2370 ( .A1(n2134), .A2(n2133), .ZN(n2132) );
  INV_X1 U2371 ( .A(n2541), .ZN(n2133) );
  AOI22_X1 U2372 ( .A1(n3805), .A2(n2513), .B1(n3817), .B2(n3795), .ZN(n3787)
         );
  NAND2_X1 U2373 ( .A1(n2231), .A2(n3125), .ZN(n2230) );
  NAND2_X1 U2374 ( .A1(n2232), .A2(n2236), .ZN(n2231) );
  INV_X1 U2375 ( .A(n3042), .ZN(n2235) );
  NAND2_X1 U2376 ( .A1(n3384), .A2(n3383), .ZN(n2253) );
  INV_X1 U2377 ( .A(n3191), .ZN(n2258) );
  OR2_X1 U2378 ( .A1(n3287), .A2(n2087), .ZN(n2256) );
  INV_X1 U2379 ( .A(n3182), .ZN(n2259) );
  AND2_X1 U2380 ( .A1(n3153), .A2(n3152), .ZN(n3154) );
  NOR2_X1 U2381 ( .A1(n2496), .A2(n3378), .ZN(n2504) );
  NAND2_X1 U2382 ( .A1(n2783), .A2(n2804), .ZN(n2827) );
  NAND2_X1 U2383 ( .A1(n3596), .A2(n2220), .ZN(n2219) );
  NAND2_X1 U2384 ( .A1(n4245), .A2(REG2_REG_2__SCAN_IN), .ZN(n2220) );
  OAI21_X1 U2385 ( .B1(n3998), .B2(n4512), .A(n4286), .ZN(n3637) );
  NAND2_X1 U2386 ( .A1(n2182), .A2(n2185), .ZN(n3704) );
  NOR2_X1 U2387 ( .A1(n3420), .A2(n2207), .ZN(n2206) );
  AND2_X1 U2388 ( .A1(n2443), .A2(REG3_REG_13__SCAN_IN), .ZN(n2453) );
  NAND2_X1 U2389 ( .A1(n4410), .A2(n3425), .ZN(n2198) );
  OR2_X1 U2390 ( .A1(n2969), .A2(n3347), .ZN(n2410) );
  AND2_X1 U2391 ( .A1(n2154), .A2(n2284), .ZN(n2151) );
  OAI21_X1 U2392 ( .B1(n2811), .B2(n2348), .A(n2347), .ZN(n2851) );
  NAND2_X1 U2393 ( .A1(n2600), .A2(n3515), .ZN(n2814) );
  NAND2_X1 U2394 ( .A1(n2323), .A2(n2710), .ZN(n3437) );
  INV_X1 U2395 ( .A(n4460), .ZN(n4474) );
  AOI21_X1 U2396 ( .B1(n2204), .B2(IR_REG_31__SCAN_IN), .A(n2076), .ZN(n2203)
         );
  NAND2_X1 U2397 ( .A1(n3267), .A2(n3182), .ZN(n3270) );
  INV_X1 U2398 ( .A(n2271), .ZN(n2267) );
  AND2_X1 U2399 ( .A1(n2270), .A2(n3343), .ZN(n2269) );
  NAND2_X1 U2400 ( .A1(n2272), .A2(n2271), .ZN(n2270) );
  INV_X1 U2401 ( .A(n3709), .ZN(n3298) );
  OR2_X1 U2402 ( .A1(n3332), .A2(n3333), .ZN(n2835) );
  OR2_X1 U2403 ( .A1(n2965), .A2(n2966), .ZN(n2271) );
  NAND2_X1 U2404 ( .A1(n3354), .A2(n3355), .ZN(n3353) );
  AND2_X1 U2405 ( .A1(n3017), .A2(n3016), .ZN(n3019) );
  XNOR2_X1 U2406 ( .A(n2707), .B(n3223), .ZN(n2757) );
  OAI22_X1 U2407 ( .A1(n2708), .A2(n2827), .B1(n2710), .B2(n3222), .ZN(n2707)
         );
  INV_X1 U2408 ( .A(n2333), .ZN(n2595) );
  NAND2_X1 U2410 ( .A1(n3579), .A2(n2692), .ZN(n3593) );
  XNOR2_X1 U2411 ( .A(n2219), .B(n2218), .ZN(n2695) );
  NAND2_X1 U2412 ( .A1(n2695), .A2(REG2_REG_3__SCAN_IN), .ZN(n2746) );
  NOR2_X1 U2413 ( .A1(n2749), .A2(n2071), .ZN(n3605) );
  NAND2_X1 U2414 ( .A1(n4292), .A2(REG2_REG_8__SCAN_IN), .ZN(n4291) );
  NAND2_X1 U2415 ( .A1(n4304), .A2(n3639), .ZN(n3640) );
  NAND2_X1 U2416 ( .A1(n4323), .A2(n2081), .ZN(n3643) );
  NAND2_X1 U2417 ( .A1(n4329), .A2(n2278), .ZN(n3615) );
  OAI21_X1 U2418 ( .B1(n4347), .B2(n2088), .A(n2221), .ZN(n3646) );
  NAND2_X1 U2419 ( .A1(n4356), .A2(n4344), .ZN(n2221) );
  NAND2_X1 U2420 ( .A1(n4380), .A2(n3652), .ZN(n4388) );
  INV_X1 U2421 ( .A(n2213), .ZN(n3651) );
  OR2_X1 U2422 ( .A1(n2571), .A2(n3230), .ZN(n3118) );
  NAND2_X1 U2423 ( .A1(n2180), .A2(n2178), .ZN(n3668) );
  NAND2_X1 U2424 ( .A1(n2179), .A2(n3665), .ZN(n2178) );
  INV_X1 U2425 ( .A(n2181), .ZN(n2179) );
  NAND2_X1 U2426 ( .A1(n2177), .A2(n2181), .ZN(n3666) );
  NAND2_X1 U2427 ( .A1(n3774), .A2(n2058), .ZN(n2177) );
  AND2_X1 U2428 ( .A1(n2562), .A2(n2554), .ZN(n2160) );
  OR2_X1 U2429 ( .A1(n3694), .A2(n3712), .ZN(n2554) );
  NOR2_X1 U2430 ( .A1(n2055), .A2(n3685), .ZN(n3684) );
  AOI21_X1 U2431 ( .B1(n2128), .B2(n2064), .A(n2542), .ZN(n2127) );
  NAND2_X1 U2432 ( .A1(n2184), .A2(n3535), .ZN(n3719) );
  OR2_X1 U2433 ( .A1(n3774), .A2(n2618), .ZN(n2184) );
  AOI21_X1 U2434 ( .B1(n3787), .B2(n3508), .A(n3510), .ZN(n3772) );
  AND2_X1 U2435 ( .A1(n3851), .A2(n3841), .ZN(n2503) );
  AOI21_X1 U2436 ( .B1(n2143), .B2(n2140), .A(n2085), .ZN(n2139) );
  INV_X1 U2437 ( .A(n2147), .ZN(n2140) );
  INV_X1 U2438 ( .A(n2143), .ZN(n2141) );
  NOR2_X1 U2439 ( .A1(n3899), .A2(n2148), .ZN(n2147) );
  INV_X1 U2440 ( .A(n2452), .ZN(n2148) );
  OAI22_X1 U2441 ( .A1(n3899), .A2(n2146), .B1(n3566), .B2(n3910), .ZN(n2145)
         );
  INV_X1 U2442 ( .A(n2451), .ZN(n2146) );
  NAND2_X1 U2443 ( .A1(n2607), .A2(n3432), .ZN(n3898) );
  AOI21_X1 U2444 ( .B1(n2195), .B2(n2194), .A(n2193), .ZN(n2192) );
  INV_X1 U2445 ( .A(n3425), .ZN(n2194) );
  AND2_X1 U2446 ( .A1(n3877), .A2(n3421), .ZN(n3899) );
  AOI21_X1 U2447 ( .B1(n2991), .B2(n2442), .A(n2441), .ZN(n3003) );
  MUX2_X1 U2448 ( .A(n4501), .B(DATAI_13_), .S(n2052), .Z(n3070) );
  OR2_X1 U2449 ( .A1(n2412), .A2(n2981), .ZN(n2431) );
  NAND2_X1 U2450 ( .A1(n2605), .A2(n3455), .ZN(n2937) );
  INV_X1 U2451 ( .A(n4446), .ZN(n3881) );
  AND2_X1 U2452 ( .A1(n4445), .A2(n2324), .ZN(n3918) );
  NOR2_X1 U2453 ( .A1(n3944), .A2(n4569), .ZN(n2102) );
  NOR2_X1 U2454 ( .A1(n3944), .A2(n2104), .ZN(n2103) );
  INV_X1 U2455 ( .A(n2106), .ZN(n2104) );
  NOR2_X1 U2456 ( .A1(n3944), .A2(n3410), .ZN(n2100) );
  AND2_X1 U2457 ( .A1(n3684), .A2(n3676), .ZN(n3674) );
  NAND2_X1 U2458 ( .A1(n3674), .A2(n3231), .ZN(n3110) );
  NOR2_X2 U2459 ( .A1(n4473), .A2(n4241), .ZN(n4569) );
  XNOR2_X1 U2460 ( .A(n2302), .B(n2667), .ZN(n2303) );
  NAND2_X1 U2461 ( .A1(n2670), .A2(IR_REG_31__SCAN_IN), .ZN(n2302) );
  XNOR2_X1 U2462 ( .A(n2299), .B(n2298), .ZN(n2304) );
  NOR2_X1 U2463 ( .A1(n2590), .A2(n2297), .ZN(n2299) );
  AND2_X1 U2464 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .ZN(n2297)
         );
  INV_X1 U2465 ( .A(n2295), .ZN(n2166) );
  NOR2_X1 U2466 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2629)
         );
  NAND2_X1 U2467 ( .A1(n2625), .A2(IR_REG_31__SCAN_IN), .ZN(n2649) );
  MUX2_X1 U2468 ( .A(IR_REG_31__SCAN_IN), .B(n2579), .S(IR_REG_22__SCAN_IN), 
        .Z(n2580) );
  XNOR2_X1 U2469 ( .A(n2583), .B(n2582), .ZN(n2596) );
  XNOR2_X1 U2470 ( .A(n2588), .B(n2587), .ZN(n2652) );
  OR2_X1 U2471 ( .A1(n3142), .A2(n3141), .ZN(n3143) );
  NOR2_X1 U2472 ( .A1(n2700), .A2(n4578), .ZN(n2749) );
  XNOR2_X1 U2473 ( .A(n3605), .B(n3628), .ZN(n2751) );
  NAND2_X1 U2474 ( .A1(n4330), .A2(n4331), .ZN(n4329) );
  XNOR2_X1 U2475 ( .A(n3615), .B(n4504), .ZN(n4341) );
  NAND2_X1 U2476 ( .A1(n4352), .A2(n4353), .ZN(n4351) );
  XNOR2_X1 U2477 ( .A(n2585), .B(n2584), .ZN(n3659) );
  NAND2_X1 U2478 ( .A1(n3110), .A2(n3115), .ZN(n2107) );
  NOR2_X1 U2479 ( .A1(n2623), .A2(n2210), .ZN(n3237) );
  NAND2_X1 U2480 ( .A1(n2212), .A2(n2211), .ZN(n2210) );
  INV_X1 U2481 ( .A(n2624), .ZN(n2212) );
  NAND2_X1 U2482 ( .A1(n2797), .A2(n4482), .ZN(n4477) );
  AND2_X1 U2483 ( .A1(n2998), .A2(n2996), .ZN(n3428) );
  NOR2_X1 U2484 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2291)
         );
  INV_X1 U2485 ( .A(n2804), .ZN(n2706) );
  NAND2_X1 U2486 ( .A1(n3279), .A2(n2244), .ZN(n2243) );
  NAND2_X1 U2487 ( .A1(n3654), .A2(REG2_REG_18__SCAN_IN), .ZN(n2225) );
  NAND2_X1 U2488 ( .A1(n2062), .A2(n2188), .ZN(n2181) );
  NAND2_X1 U2489 ( .A1(n2185), .A2(n2187), .ZN(n2183) );
  NOR2_X1 U2490 ( .A1(n2128), .A2(n2131), .ZN(n2125) );
  AND2_X1 U2491 ( .A1(n2504), .A2(REG3_REG_19__SCAN_IN), .ZN(n2514) );
  INV_X1 U2492 ( .A(n3428), .ZN(n2193) );
  NOR2_X1 U2493 ( .A1(n2431), .A2(n2428), .ZN(n2443) );
  AND2_X1 U2494 ( .A1(n2657), .A2(n2645), .ZN(n2715) );
  NAND2_X1 U2495 ( .A1(n2121), .A2(n3728), .ZN(n2120) );
  NOR2_X1 U2496 ( .A1(n3272), .A2(n3767), .ZN(n2121) );
  AND2_X1 U2497 ( .A1(n2052), .A2(DATAI_21_), .ZN(n3171) );
  AND2_X1 U2498 ( .A1(n2053), .A2(DATAI_20_), .ZN(n3163) );
  NAND2_X1 U2499 ( .A1(n2116), .A2(n3870), .ZN(n2115) );
  INV_X1 U2500 ( .A(n2117), .ZN(n2116) );
  NAND2_X1 U2501 ( .A1(n3889), .A2(n3082), .ZN(n2117) );
  INV_X1 U2502 ( .A(IR_REG_18__SCAN_IN), .ZN(n2190) );
  INV_X1 U2503 ( .A(IR_REG_20__SCAN_IN), .ZN(n2587) );
  INV_X1 U2504 ( .A(IR_REG_16__SCAN_IN), .ZN(n2163) );
  INV_X1 U2505 ( .A(IR_REG_13__SCAN_IN), .ZN(n2292) );
  INV_X1 U2506 ( .A(IR_REG_6__SCAN_IN), .ZN(n2404) );
  INV_X1 U2507 ( .A(IR_REG_7__SCAN_IN), .ZN(n2403) );
  INV_X1 U2508 ( .A(IR_REG_2__SCAN_IN), .ZN(n2285) );
  NAND2_X1 U2509 ( .A1(n2237), .A2(n3044), .ZN(n2236) );
  INV_X1 U2510 ( .A(n3078), .ZN(n2237) );
  INV_X1 U2511 ( .A(n2233), .ZN(n2232) );
  OAI21_X1 U2512 ( .B1(n3078), .B2(n2234), .A(n3077), .ZN(n2233) );
  NAND2_X1 U2513 ( .A1(n3044), .A2(n2235), .ZN(n2234) );
  NOR2_X1 U2514 ( .A1(n3260), .A2(n2255), .ZN(n2254) );
  INV_X1 U2515 ( .A(n2252), .ZN(n2251) );
  OAI22_X1 U2516 ( .A1(n3260), .A2(n2253), .B1(n3220), .B2(n3221), .ZN(n2252)
         );
  OAI21_X1 U2517 ( .B1(n3229), .B2(n2251), .A(n2248), .ZN(n2247) );
  OAI21_X1 U2518 ( .B1(n3229), .B2(n2254), .A(n2251), .ZN(n2248) );
  AND2_X1 U2519 ( .A1(n2061), .A2(n2316), .ZN(n2710) );
  NAND2_X1 U2520 ( .A1(n2053), .A2(DATAI_1_), .ZN(n2316) );
  AND2_X1 U2521 ( .A1(n2346), .A2(DATAI_25_), .ZN(n3200) );
  AOI21_X1 U2522 ( .B1(n3182), .B2(n2261), .A(n2258), .ZN(n2257) );
  AND2_X1 U2523 ( .A1(n2965), .A2(n2966), .ZN(n2272) );
  NAND2_X1 U2524 ( .A1(n2968), .A2(n2271), .ZN(n2265) );
  AOI21_X1 U2525 ( .B1(n2711), .B2(REG1_REG_0__SCAN_IN), .A(n2713), .ZN(n2712)
         );
  NAND2_X1 U2526 ( .A1(n2264), .A2(n2260), .ZN(n3267) );
  NAND2_X1 U2527 ( .A1(n3285), .A2(n3284), .ZN(n2263) );
  NAND2_X1 U2528 ( .A1(n3041), .A2(n3042), .ZN(n3040) );
  NAND2_X1 U2529 ( .A1(n2309), .A2(IR_REG_27__SCAN_IN), .ZN(n2312) );
  OR2_X1 U2530 ( .A1(n2309), .A2(IR_REG_28__SCAN_IN), .ZN(n2313) );
  OR2_X1 U2531 ( .A1(n2484), .A2(n2483), .ZN(n2496) );
  INV_X1 U2532 ( .A(n4490), .ZN(n2731) );
  NAND2_X1 U2533 ( .A1(n2217), .A2(REG2_REG_1__SCAN_IN), .ZN(n3592) );
  INV_X1 U2534 ( .A(n2219), .ZN(n2747) );
  INV_X1 U2535 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4098) );
  NAND2_X1 U2536 ( .A1(n2168), .A2(n2167), .ZN(n3610) );
  OR2_X1 U2537 ( .A1(n4283), .A2(n4584), .ZN(n2167) );
  NAND2_X1 U2538 ( .A1(n2169), .A2(n4280), .ZN(n2168) );
  NAND2_X1 U2539 ( .A1(n4283), .A2(n4584), .ZN(n2169) );
  NAND2_X1 U2540 ( .A1(n4291), .A2(n3638), .ZN(n4306) );
  NAND2_X1 U2541 ( .A1(n4315), .A2(n3641), .ZN(n4324) );
  XNOR2_X1 U2542 ( .A(n3646), .B(n4367), .ZN(n4358) );
  NAND2_X1 U2543 ( .A1(n4351), .A2(n2093), .ZN(n3617) );
  OR2_X1 U2544 ( .A1(n4370), .A2(n4369), .ZN(n2215) );
  XNOR2_X1 U2545 ( .A(n2213), .B(n4496), .ZN(n4381) );
  INV_X1 U2546 ( .A(n4393), .ZN(n2176) );
  OR2_X1 U2547 ( .A1(n3653), .A2(REG2_REG_17__SCAN_IN), .ZN(n2226) );
  NAND2_X1 U2548 ( .A1(n4388), .A2(n4390), .ZN(n4389) );
  INV_X1 U2549 ( .A(n2225), .ZN(n2222) );
  INV_X1 U2550 ( .A(n2226), .ZN(n2224) );
  NOR2_X1 U2551 ( .A1(n2578), .A2(n3115), .ZN(n2106) );
  OAI21_X1 U2552 ( .B1(n2054), .B2(n2066), .A(n2162), .ZN(n2157) );
  AND2_X1 U2553 ( .A1(n3112), .A2(n3408), .ZN(n3501) );
  NAND2_X1 U2554 ( .A1(n3411), .A2(n4447), .ZN(n2211) );
  AND2_X1 U2555 ( .A1(n2053), .A2(DATAI_26_), .ZN(n3685) );
  AND2_X1 U2556 ( .A1(n2053), .A2(DATAI_22_), .ZN(n3767) );
  NAND2_X1 U2557 ( .A1(n2616), .A2(n3470), .ZN(n3774) );
  NAND2_X1 U2558 ( .A1(n2208), .A2(n2065), .ZN(n2616) );
  NAND2_X1 U2559 ( .A1(n2208), .A2(n2206), .ZN(n3790) );
  INV_X1 U2560 ( .A(n3834), .ZN(n3841) );
  NAND2_X1 U2561 ( .A1(n2493), .A2(n3146), .ZN(n2494) );
  AOI21_X1 U2562 ( .B1(n2138), .B2(n2136), .A(n2135), .ZN(n3848) );
  NOR2_X1 U2563 ( .A1(n2141), .A2(n2137), .ZN(n2136) );
  OAI21_X1 U2564 ( .B1(n2139), .B2(n2137), .A(n2084), .ZN(n2135) );
  INV_X1 U2565 ( .A(n3003), .ZN(n2138) );
  AND4_X1 U2566 ( .A1(n2501), .A2(n2500), .A3(n2499), .A4(n2498), .ZN(n3851)
         );
  NAND2_X1 U2567 ( .A1(n2208), .A2(n3419), .ZN(n3849) );
  AND4_X1 U2568 ( .A1(n2477), .A2(n2476), .A3(n2475), .A4(n2474), .ZN(n3882)
         );
  AND4_X1 U2569 ( .A1(n2460), .A2(n2459), .A3(n2458), .A4(n2457), .ZN(n3880)
         );
  AND2_X1 U2570 ( .A1(n4240), .A2(n2652), .ZN(n2804) );
  NAND2_X1 U2571 ( .A1(n3898), .A2(n3899), .ZN(n3897) );
  OR2_X1 U2572 ( .A1(n3004), .A2(n3070), .ZN(n3911) );
  NAND2_X1 U2573 ( .A1(n2198), .A2(n2195), .ZN(n2997) );
  NAND2_X1 U2574 ( .A1(n2198), .A2(n3427), .ZN(n2987) );
  OAI21_X1 U2575 ( .B1(n3052), .B2(n2419), .A(n2420), .ZN(n4415) );
  NAND2_X1 U2576 ( .A1(n3053), .A2(n3424), .ZN(n2606) );
  OAI21_X1 U2577 ( .B1(n2937), .B2(n2935), .A(n3459), .ZN(n3053) );
  INV_X1 U2578 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2981) );
  OR2_X1 U2579 ( .A1(n2396), .A2(n3346), .ZN(n2412) );
  OAI21_X1 U2580 ( .B1(n2947), .B2(n2395), .A(n2394), .ZN(n2936) );
  INV_X1 U2581 ( .A(n2941), .ZN(n3347) );
  OAI21_X1 U2582 ( .B1(n2903), .B2(n2604), .A(n3456), .ZN(n2948) );
  INV_X1 U2583 ( .A(n3571), .ZN(n2928) );
  INV_X1 U2584 ( .A(n2920), .ZN(n3253) );
  NAND2_X1 U2585 ( .A1(n2201), .A2(n3452), .ZN(n2903) );
  NAND2_X1 U2586 ( .A1(n2863), .A2(n3448), .ZN(n2201) );
  AOI21_X1 U2587 ( .B1(n2151), .B2(n2368), .A(n2070), .ZN(n2149) );
  OAI21_X1 U2588 ( .B1(n2852), .B2(n2601), .A(n3450), .ZN(n2799) );
  INV_X1 U2589 ( .A(n2853), .ZN(n3336) );
  NAND2_X1 U2590 ( .A1(n2850), .A2(n3336), .ZN(n2849) );
  NAND2_X1 U2591 ( .A1(n2814), .A2(n3445), .ZN(n2852) );
  NOR2_X1 U2592 ( .A1(n4528), .A2(n3443), .ZN(n2850) );
  NAND2_X1 U2593 ( .A1(n3917), .A2(n2332), .ZN(n2811) );
  NAND2_X1 U2594 ( .A1(n3918), .A2(n2598), .ZN(n3917) );
  NAND3_X1 U2595 ( .A1(n2199), .A2(n2597), .A3(n3437), .ZN(n4455) );
  INV_X1 U2596 ( .A(n3577), .ZN(n4450) );
  NAND2_X1 U2597 ( .A1(n4236), .A2(n2718), .ZN(n4449) );
  NAND2_X1 U2598 ( .A1(n4452), .A2(n4443), .ZN(n4445) );
  NAND2_X1 U2599 ( .A1(n2597), .A2(n3437), .ZN(n4452) );
  INV_X1 U2600 ( .A(n2108), .ZN(n3939) );
  NOR2_X1 U2601 ( .A1(n3779), .A2(n2119), .ZN(n3748) );
  INV_X1 U2602 ( .A(n2121), .ZN(n2119) );
  OR2_X1 U2603 ( .A1(n3798), .A2(n3171), .ZN(n3779) );
  INV_X1 U2604 ( .A(n3171), .ZN(n3780) );
  NAND2_X1 U2605 ( .A1(n3821), .A2(n3799), .ZN(n3798) );
  INV_X1 U2606 ( .A(n3163), .ZN(n3799) );
  MUX2_X1 U2607 ( .A(n3659), .B(n4067), .S(n2052), .Z(n3823) );
  NOR2_X1 U2608 ( .A1(n3856), .A2(n3834), .ZN(n3839) );
  AND2_X1 U2609 ( .A1(n3839), .A2(n3823), .ZN(n3821) );
  INV_X1 U2610 ( .A(n2480), .ZN(n3870) );
  NOR2_X1 U2611 ( .A1(n3911), .A2(n3910), .ZN(n3909) );
  NOR2_X1 U2612 ( .A1(n3911), .A2(n2117), .ZN(n3887) );
  NOR2_X1 U2613 ( .A1(n4423), .A2(n4424), .ZN(n4422) );
  NAND2_X1 U2614 ( .A1(n4422), .A2(n3027), .ZN(n3004) );
  NAND2_X1 U2615 ( .A1(n2099), .A2(n2098), .ZN(n4423) );
  INV_X1 U2616 ( .A(n2949), .ZN(n2956) );
  AND2_X1 U2617 ( .A1(n2907), .A2(n3253), .ZN(n2957) );
  NAND2_X1 U2618 ( .A1(n2957), .A2(n2956), .ZN(n2955) );
  OR2_X1 U2619 ( .A1(n2849), .A2(n2842), .ZN(n2867) );
  NOR2_X1 U2620 ( .A1(n2867), .A2(n2881), .ZN(n2907) );
  NAND2_X1 U2621 ( .A1(n2110), .A2(IR_REG_31__SCAN_IN), .ZN(n2309) );
  NAND4_X1 U2622 ( .A1(n2111), .A2(n2056), .A3(n2189), .A4(n2205), .ZN(n2110)
         );
  AND2_X1 U2623 ( .A1(n2478), .A2(n2472), .ZN(n3649) );
  OR2_X1 U2624 ( .A1(n2425), .A2(IR_REG_10__SCAN_IN), .ZN(n2426) );
  AOI21_X1 U2625 ( .B1(n2269), .B2(n2267), .A(n2075), .ZN(n2266) );
  INV_X1 U2626 ( .A(n2269), .ZN(n2268) );
  NOR2_X1 U2627 ( .A1(n2780), .A2(n2779), .ZN(n3334) );
  MUX2_X1 U2628 ( .A(n4244), .B(DATAI_3_), .S(n2052), .Z(n3443) );
  NAND2_X1 U2629 ( .A1(n2247), .A2(n2249), .ZN(n2246) );
  NAND2_X1 U2630 ( .A1(n2250), .A2(n2251), .ZN(n2249) );
  INV_X1 U2631 ( .A(n3229), .ZN(n2250) );
  AND2_X1 U2632 ( .A1(n3118), .A2(n2572), .ZN(n3238) );
  INV_X1 U2633 ( .A(n3570), .ZN(n2969) );
  AND4_X1 U2634 ( .A1(n2380), .A2(n2379), .A3(n2378), .A4(n2377), .ZN(n2951)
         );
  INV_X1 U2635 ( .A(n2710), .ZN(n4459) );
  AND4_X1 U2636 ( .A1(n2424), .A2(n2423), .A3(n2422), .A4(n2421), .ZN(n3056)
         );
  INV_X1 U2637 ( .A(n3200), .ZN(n3712) );
  NAND2_X1 U2638 ( .A1(n2835), .A2(n2067), .ZN(n2238) );
  NAND2_X1 U2639 ( .A1(n2240), .A2(n2067), .ZN(n2239) );
  INV_X1 U2640 ( .A(n3187), .ZN(n3728) );
  NAND2_X1 U2641 ( .A1(n2322), .A2(n2321), .ZN(n4460) );
  NAND2_X1 U2642 ( .A1(n2346), .A2(DATAI_0_), .ZN(n2321) );
  OR2_X1 U2643 ( .A1(n2052), .A2(n2228), .ZN(n2322) );
  AND2_X1 U2644 ( .A1(n2723), .A2(n2722), .ZN(n3344) );
  AND4_X1 U2645 ( .A1(n2511), .A2(n2510), .A3(n2509), .A4(n2508), .ZN(n3833)
         );
  NAND2_X1 U2646 ( .A1(n2264), .A2(n2263), .ZN(n3365) );
  AND4_X1 U2647 ( .A1(n2436), .A2(n2435), .A3(n2434), .A4(n2433), .ZN(n4414)
         );
  OR2_X1 U2648 ( .A1(n2726), .A2(n4458), .ZN(n3273) );
  INV_X1 U2649 ( .A(n3273), .ZN(n3401) );
  INV_X1 U2650 ( .A(n3388), .ZN(n3398) );
  INV_X1 U2651 ( .A(n3387), .ZN(n3399) );
  OAI211_X1 U2652 ( .C1(n2361), .C2(n3687), .A(n2561), .B(n2560), .ZN(n3709)
         );
  OR2_X1 U2653 ( .A1(n3686), .A2(n2595), .ZN(n2561) );
  OAI211_X1 U2654 ( .C1(n3297), .C2(n2595), .A(n2553), .B(n2552), .ZN(n3724)
         );
  OR2_X1 U2655 ( .A1(n3326), .A2(n2595), .ZN(n2547) );
  AND4_X1 U2656 ( .A1(n2524), .A2(n2523), .A3(n2522), .A4(n2521), .ZN(n3793)
         );
  NAND4_X1 U2657 ( .A1(n2520), .A2(n2519), .A3(n2518), .A4(n2517), .ZN(n3818)
         );
  INV_X1 U2658 ( .A(n3833), .ZN(n3795) );
  INV_X1 U2659 ( .A(n3882), .ZN(n3853) );
  INV_X1 U2660 ( .A(n4414), .ZN(n3568) );
  INV_X1 U2661 ( .A(n3056), .ZN(n3569) );
  INV_X1 U2662 ( .A(n2951), .ZN(n3572) );
  INV_X1 U2663 ( .A(n2829), .ZN(n3575) );
  NAND2_X1 U2664 ( .A1(n2335), .A2(REG1_REG_1__SCAN_IN), .ZN(n2308) );
  NAND2_X1 U2665 ( .A1(n2336), .A2(REG2_REG_1__SCAN_IN), .ZN(n2306) );
  NAND2_X1 U2666 ( .A1(n2200), .A2(n2057), .ZN(n3577) );
  AND2_X1 U2667 ( .A1(n2319), .A2(n2320), .ZN(n2200) );
  NAND2_X1 U2668 ( .A1(n2217), .A2(REG1_REG_1__SCAN_IN), .ZN(n2698) );
  XNOR2_X1 U2669 ( .A(n2750), .B(n4244), .ZN(n2700) );
  NOR2_X1 U2670 ( .A1(n4261), .A2(n4260), .ZN(n4259) );
  XNOR2_X1 U2671 ( .A(n3610), .B(n4510), .ZN(n4297) );
  NAND2_X1 U2672 ( .A1(n4297), .A2(REG1_REG_8__SCAN_IN), .ZN(n4296) );
  NAND2_X1 U2673 ( .A1(n4313), .A2(n3614), .ZN(n4330) );
  NAND2_X1 U2674 ( .A1(n4335), .A2(n3645), .ZN(n4347) );
  NAND2_X1 U2675 ( .A1(n4340), .A2(n3616), .ZN(n4352) );
  XNOR2_X1 U2676 ( .A(n3617), .B(n4367), .ZN(n4364) );
  INV_X1 U2677 ( .A(n2215), .ZN(n4368) );
  XNOR2_X1 U2678 ( .A(n3619), .B(n3650), .ZN(n4384) );
  INV_X1 U2679 ( .A(n2175), .ZN(n4385) );
  OR2_X1 U2680 ( .A1(n4384), .A2(REG1_REG_16__SCAN_IN), .ZN(n2175) );
  INV_X1 U2681 ( .A(n3620), .ZN(n2174) );
  NAND2_X1 U2682 ( .A1(n2171), .A2(n2170), .ZN(n4394) );
  NAND2_X1 U2683 ( .A1(n3620), .A2(n2176), .ZN(n2170) );
  OR2_X1 U2684 ( .A1(n4384), .A2(n2172), .ZN(n2171) );
  NAND2_X1 U2685 ( .A1(n2176), .A2(n2173), .ZN(n2172) );
  NAND2_X1 U2686 ( .A1(n4389), .A2(n2226), .ZN(n4398) );
  OR2_X1 U2687 ( .A1(n4258), .A2(n4237), .ZN(n4270) );
  NAND2_X1 U2688 ( .A1(n2223), .A2(n2095), .ZN(n3656) );
  AOI21_X1 U2689 ( .B1(n2555), .B2(n2160), .A(n2054), .ZN(n3664) );
  NAND2_X1 U2690 ( .A1(n3772), .A2(n2128), .ZN(n2123) );
  OR2_X1 U2691 ( .A1(n4466), .A2(n4242), .ZN(n3844) );
  OAI21_X1 U2692 ( .B1(n3003), .B2(n2141), .A(n2139), .ZN(n3863) );
  NAND2_X1 U2693 ( .A1(n2144), .A2(n2142), .ZN(n3876) );
  INV_X1 U2694 ( .A(n2145), .ZN(n2142) );
  NAND2_X1 U2695 ( .A1(n3003), .A2(n2147), .ZN(n2144) );
  AOI21_X1 U2696 ( .B1(n3003), .B2(n2452), .A(n2451), .ZN(n3904) );
  NAND2_X1 U2697 ( .A1(n2153), .A2(n2154), .ZN(n2862) );
  OR2_X1 U2698 ( .A1(n2803), .A2(n2368), .ZN(n2153) );
  INV_X1 U2699 ( .A(n3914), .ZN(n4468) );
  NAND2_X1 U2700 ( .A1(n2725), .A2(n2727), .ZN(n4482) );
  NAND2_X1 U2701 ( .A1(n2105), .A2(n2101), .ZN(n3946) );
  NAND2_X1 U2702 ( .A1(n3110), .A2(n2100), .ZN(n2105) );
  INV_X2 U2703 ( .A(n4570), .ZN(n4572) );
  INV_X1 U2704 ( .A(n2741), .ZN(n4236) );
  NAND2_X1 U2705 ( .A1(n2633), .A2(IR_REG_31__SCAN_IN), .ZN(n2634) );
  XNOR2_X1 U2706 ( .A(n2631), .B(n2294), .ZN(n4238) );
  NAND2_X1 U2707 ( .A1(n2651), .A2(IR_REG_31__SCAN_IN), .ZN(n2627) );
  INV_X1 U2708 ( .A(n2596), .ZN(n4240) );
  INV_X1 U2709 ( .A(n2652), .ZN(n4241) );
  AND2_X1 U2710 ( .A1(n2409), .A2(n2425), .ZN(n4300) );
  NAND2_X1 U2711 ( .A1(n3584), .A2(n2217), .ZN(n3585) );
  AND2_X1 U2712 ( .A1(n2107), .A2(n2108), .ZN(n3945) );
  OAI21_X1 U2713 ( .B1(n2664), .B2(n4587), .A(n2092), .ZN(n2661) );
  MUX2_X1 U2714 ( .A(REG0_REG_28__SCAN_IN), .B(n2664), .S(n4572), .Z(n2665) );
  NAND2_X1 U2715 ( .A1(U3149), .A2(DATAI_1_), .ZN(n2216) );
  AND2_X1 U2716 ( .A1(n3298), .A2(n3693), .ZN(n2054) );
  OR3_X1 U2717 ( .A1(n3779), .A2(n2120), .A3(n3200), .ZN(n2055) );
  NAND2_X1 U2718 ( .A1(n2708), .A2(n4459), .ZN(n2597) );
  NAND2_X1 U2719 ( .A1(n2287), .A2(n2277), .ZN(n2366) );
  INV_X2 U2720 ( .A(n2361), .ZN(n2350) );
  AND2_X1 U2721 ( .A1(n2318), .A2(n2317), .ZN(n2057) );
  AND2_X1 U2722 ( .A1(n2188), .A2(n2185), .ZN(n2058) );
  AND4_X1 U2723 ( .A1(n2289), .A2(n2290), .A3(n2291), .A4(n2288), .ZN(n2060)
         );
  OR2_X1 U2724 ( .A1(n2053), .A2(n2315), .ZN(n2061) );
  NAND2_X1 U2725 ( .A1(n3473), .A2(n2183), .ZN(n2062) );
  INV_X1 U2726 ( .A(IR_REG_31__SCAN_IN), .ZN(n2628) );
  AND2_X1 U2727 ( .A1(n4389), .A2(n2091), .ZN(n2063) );
  NOR2_X1 U2728 ( .A1(n3793), .A2(n3780), .ZN(n2064) );
  INV_X1 U2729 ( .A(n3486), .ZN(n2137) );
  INV_X1 U2730 ( .A(n3054), .ZN(n2098) );
  AND2_X1 U2731 ( .A1(n2206), .A2(n2209), .ZN(n2065) );
  AND2_X1 U2732 ( .A1(n3389), .A2(n3676), .ZN(n2066) );
  INV_X1 U2733 ( .A(n3900), .ZN(n3309) );
  INV_X2 U2734 ( .A(n4587), .ZN(n4590) );
  NAND2_X1 U2735 ( .A1(n2837), .A2(n2836), .ZN(n2067) );
  AOI21_X1 U2736 ( .B1(n3772), .B2(n2525), .A(n2064), .ZN(n3734) );
  AND2_X1 U2737 ( .A1(n2584), .A2(n2587), .ZN(n2068) );
  AND2_X1 U2738 ( .A1(n2123), .A2(n2127), .ZN(n2069) );
  AND2_X1 U2739 ( .A1(n2355), .A2(n2345), .ZN(n4244) );
  INV_X1 U2740 ( .A(n4244), .ZN(n2218) );
  AND2_X1 U2741 ( .A1(n3573), .A2(n2881), .ZN(n2070) );
  OAI21_X1 U2742 ( .B1(n3377), .B2(n2243), .A(n2241), .ZN(n3354) );
  AND2_X1 U2743 ( .A1(n2750), .A2(n4244), .ZN(n2071) );
  NAND4_X1 U2744 ( .A1(n2308), .A2(n2307), .A3(n2306), .A4(n2305), .ZN(n2323)
         );
  INV_X1 U2745 ( .A(n2205), .ZN(n2204) );
  NOR2_X1 U2746 ( .A1(n2295), .A2(IR_REG_26__SCAN_IN), .ZN(n2205) );
  INV_X1 U2747 ( .A(n2335), .ZN(n2359) );
  AND2_X1 U2748 ( .A1(n2673), .A2(n2303), .ZN(n2335) );
  AND3_X1 U2749 ( .A1(n2319), .A2(n2320), .A3(n4460), .ZN(n2072) );
  AND2_X1 U2750 ( .A1(n2175), .A2(n2174), .ZN(n2073) );
  NAND2_X1 U2751 ( .A1(n2581), .A2(n2582), .ZN(n2074) );
  INV_X1 U2752 ( .A(n2112), .ZN(n2581) );
  NAND2_X1 U2753 ( .A1(n2980), .A2(n2979), .ZN(n2075) );
  AND2_X1 U2754 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2076)
         );
  AND2_X1 U2755 ( .A1(n2058), .A2(n3665), .ZN(n2077) );
  AND2_X1 U2756 ( .A1(n2068), .A2(n2275), .ZN(n2078) );
  AND2_X1 U2757 ( .A1(n2166), .A2(n2275), .ZN(n2079) );
  AND3_X1 U2758 ( .A1(n2060), .A2(n2287), .A3(n2277), .ZN(n2080) );
  NAND2_X1 U2759 ( .A1(n3040), .A2(n3044), .ZN(n3079) );
  INV_X1 U2760 ( .A(n2842), .ZN(n2155) );
  AND2_X1 U2761 ( .A1(n2080), .A2(n2292), .ZN(n2461) );
  INV_X1 U2762 ( .A(n2336), .ZN(n2361) );
  AOI21_X1 U2763 ( .B1(n4415), .B2(n4416), .A(n2427), .ZN(n2991) );
  OAI21_X1 U2764 ( .B1(n2936), .B2(n2411), .A(n2410), .ZN(n3052) );
  INV_X1 U2765 ( .A(n3418), .ZN(n2188) );
  INV_X1 U2766 ( .A(n3383), .ZN(n2255) );
  INV_X1 U2767 ( .A(n3136), .ZN(n3889) );
  INV_X1 U2768 ( .A(n4280), .ZN(n4512) );
  OR2_X1 U2769 ( .A1(n4334), .A2(n3642), .ZN(n2081) );
  INV_X1 U2770 ( .A(n2122), .ZN(n4146) );
  NOR2_X1 U2771 ( .A1(n3779), .A2(n3767), .ZN(n2122) );
  INV_X1 U2772 ( .A(n3760), .ZN(n2134) );
  INV_X1 U2773 ( .A(n2118), .ZN(n3727) );
  NOR2_X1 U2774 ( .A1(n3779), .A2(n2120), .ZN(n2118) );
  AND2_X1 U2775 ( .A1(n3818), .A2(n3799), .ZN(n3533) );
  INV_X1 U2776 ( .A(n3533), .ZN(n2209) );
  INV_X1 U2777 ( .A(n2261), .ZN(n2260) );
  NAND2_X1 U2778 ( .A1(n2262), .A2(n2263), .ZN(n2261) );
  INV_X1 U2779 ( .A(n2549), .ZN(n2131) );
  AND2_X1 U2780 ( .A1(n3707), .A2(n3728), .ZN(n2082) );
  AND2_X1 U2781 ( .A1(n3741), .A2(n3739), .ZN(n3532) );
  NAND2_X1 U2782 ( .A1(n3229), .A2(n2254), .ZN(n2083) );
  NAND2_X1 U2783 ( .A1(n3853), .A2(n2480), .ZN(n2084) );
  NAND2_X1 U2784 ( .A1(n2072), .A2(n2057), .ZN(n4451) );
  INV_X1 U2785 ( .A(n4451), .ZN(n2199) );
  INV_X1 U2786 ( .A(n2162), .ZN(n2161) );
  AND2_X1 U2787 ( .A1(n3900), .A2(n3136), .ZN(n2085) );
  AND2_X1 U2788 ( .A1(n2247), .A2(n2083), .ZN(n2086) );
  OR2_X1 U2789 ( .A1(n2259), .A2(n3174), .ZN(n2087) );
  INV_X1 U2790 ( .A(n2196), .ZN(n2195) );
  NAND2_X1 U2791 ( .A1(n2197), .A2(n3427), .ZN(n2196) );
  INV_X1 U2792 ( .A(n2598), .ZN(n3490) );
  NAND2_X1 U2793 ( .A1(n3439), .A2(n3440), .ZN(n2598) );
  NAND2_X1 U2794 ( .A1(n2265), .A2(n2269), .ZN(n2978) );
  NOR2_X1 U2795 ( .A1(n2955), .A2(n2941), .ZN(n2099) );
  XNOR2_X1 U2796 ( .A(n2634), .B(IR_REG_26__SCAN_IN), .ZN(n2646) );
  INV_X1 U2797 ( .A(IR_REG_15__SCAN_IN), .ZN(n2165) );
  AND2_X1 U2798 ( .A1(n4501), .A2(REG2_REG_13__SCAN_IN), .ZN(n2088) );
  INV_X1 U2799 ( .A(n3419), .ZN(n2207) );
  NAND2_X1 U2800 ( .A1(n2080), .A2(n2059), .ZN(n2490) );
  INV_X1 U2801 ( .A(IR_REG_14__SCAN_IN), .ZN(n2164) );
  INV_X1 U2802 ( .A(n2114), .ZN(n3869) );
  NOR2_X1 U2803 ( .A1(n3911), .A2(n2115), .ZN(n2114) );
  NAND2_X1 U2804 ( .A1(n2273), .A2(n2080), .ZN(n2089) );
  OR2_X1 U2805 ( .A1(n3334), .A2(n2835), .ZN(n2090) );
  NOR2_X1 U2806 ( .A1(n4399), .A2(n2224), .ZN(n2091) );
  INV_X1 U2807 ( .A(n2109), .ZN(n3926) );
  NAND2_X1 U2808 ( .A1(n4474), .A2(n2710), .ZN(n2109) );
  OR2_X1 U2809 ( .A1(n4590), .A2(REG1_REG_28__SCAN_IN), .ZN(n2092) );
  INV_X1 U2810 ( .A(n2578), .ZN(n3231) );
  OR2_X1 U2811 ( .A1(n4356), .A2(n4042), .ZN(n2093) );
  AND2_X1 U2812 ( .A1(n4390), .A2(n2225), .ZN(n2094) );
  OR2_X1 U2813 ( .A1(n2091), .A2(n2222), .ZN(n2095) );
  INV_X1 U2814 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2173) );
  XNOR2_X2 U2815 ( .A(n2191), .B(n2314), .ZN(n2315) );
  NAND2_X1 U2816 ( .A1(n2693), .A2(n2694), .ZN(n3596) );
  NOR2_X1 U2817 ( .A1(n4357), .A2(n3647), .ZN(n4370) );
  NAND2_X1 U2818 ( .A1(n3674), .A2(n2106), .ZN(n2108) );
  AOI21_X1 U2819 ( .B1(n3674), .B2(n2103), .A(n2102), .ZN(n2101) );
  NAND3_X1 U2820 ( .A1(n2111), .A2(n2056), .A3(n2189), .ZN(n2625) );
  NAND4_X1 U2821 ( .A1(n2189), .A2(n2056), .A3(n2273), .A4(n2068), .ZN(n2112)
         );
  INV_X1 U2822 ( .A(n2113), .ZN(n3856) );
  OAI21_X1 U2823 ( .B1(n3772), .B2(n2126), .A(n2124), .ZN(n2130) );
  INV_X1 U2824 ( .A(n3574), .ZN(n2152) );
  NAND2_X1 U2825 ( .A1(n2150), .A2(n2149), .ZN(n2912) );
  NAND2_X1 U2826 ( .A1(n2803), .A2(n2151), .ZN(n2150) );
  NAND2_X1 U2827 ( .A1(n2152), .A2(n2155), .ZN(n2154) );
  NAND2_X1 U2828 ( .A1(n2555), .A2(n2158), .ZN(n2156) );
  NAND2_X1 U2829 ( .A1(n2156), .A2(n2157), .ZN(n3108) );
  NAND2_X1 U2830 ( .A1(n2555), .A2(n2554), .ZN(n3683) );
  NAND2_X1 U2831 ( .A1(n3696), .A2(n3669), .ZN(n2162) );
  NAND2_X1 U2832 ( .A1(n2581), .A2(n2079), .ZN(n2633) );
  INV_X1 U2833 ( .A(n2633), .ZN(n2301) );
  NOR2_X2 U2834 ( .A1(n4271), .A2(n3609), .ZN(n4283) );
  NAND2_X1 U2835 ( .A1(n2301), .A2(n2276), .ZN(n2670) );
  NAND2_X1 U2836 ( .A1(n3774), .A2(n2077), .ZN(n2180) );
  OR2_X1 U2837 ( .A1(n3774), .A2(n2187), .ZN(n2182) );
  NAND3_X1 U2838 ( .A1(n2273), .A2(n2189), .A3(n2056), .ZN(n2512) );
  AND2_X2 U2839 ( .A1(n2060), .A2(n2287), .ZN(n2189) );
  NAND2_X1 U2840 ( .A1(n2228), .A2(n2191), .ZN(n2227) );
  NAND3_X1 U2841 ( .A1(n2228), .A2(n2285), .A3(n2191), .ZN(n2342) );
  OAI21_X1 U2842 ( .B1(n4410), .B2(n2196), .A(n2192), .ZN(n2607) );
  INV_X1 U2843 ( .A(n2625), .ZN(n2202) );
  OAI21_X1 U2844 ( .B1(n2202), .B2(n2628), .A(n2203), .ZN(n2590) );
  NAND2_X1 U2845 ( .A1(n3864), .A2(n2137), .ZN(n2208) );
  XNOR2_X1 U2846 ( .A(n3108), .B(n3501), .ZN(n3244) );
  OAI21_X1 U2847 ( .B1(n3244), .B2(n4557), .A(n3237), .ZN(n2664) );
  OAI21_X1 U2848 ( .B1(n2315), .B2(U3149), .A(n2216), .ZN(U3351) );
  MUX2_X1 U2849 ( .A(n4575), .B(REG1_REG_1__SCAN_IN), .S(n2315), .Z(n3583) );
  INV_X1 U2850 ( .A(n2315), .ZN(n2217) );
  NAND2_X1 U2851 ( .A1(n4388), .A2(n2094), .ZN(n2223) );
  OAI21_X1 U2852 ( .B1(n3041), .B2(n2236), .A(n2232), .ZN(n3124) );
  INV_X1 U2853 ( .A(n2229), .ZN(n3123) );
  AOI21_X1 U2854 ( .B1(n3041), .B2(n2232), .A(n2230), .ZN(n2229) );
  INV_X1 U2855 ( .A(n2779), .ZN(n2240) );
  OAI21_X1 U2856 ( .B1(n3377), .B2(n3375), .A(n3373), .ZN(n3278) );
  NAND2_X1 U2857 ( .A1(n3375), .A2(n3373), .ZN(n2244) );
  NAND2_X1 U2858 ( .A1(n3386), .A2(n2086), .ZN(n2245) );
  OAI211_X1 U2859 ( .C1(n3386), .C2(n2246), .A(n2245), .B(n3344), .ZN(n3236)
         );
  OAI21_X1 U2860 ( .B1(n3386), .B2(n3384), .A(n3383), .ZN(n3259) );
  OR2_X1 U2861 ( .A1(n3287), .A2(n3174), .ZN(n2264) );
  NAND2_X1 U2862 ( .A1(n2256), .A2(n2257), .ZN(n3194) );
  INV_X1 U2863 ( .A(n3366), .ZN(n2262) );
  OAI21_X1 U2864 ( .B1(n2968), .B2(n2268), .A(n2266), .ZN(n3014) );
  OAI21_X1 U2865 ( .B1(n2968), .B2(n2272), .A(n2271), .ZN(n2279) );
  OAI21_X1 U2866 ( .B1(n3108), .B2(n3501), .A(n3107), .ZN(n3109) );
  AND2_X1 U2867 ( .A1(n3304), .A2(n3308), .ZN(n3140) );
  INV_X1 U2868 ( .A(n2303), .ZN(n4235) );
  OR2_X1 U2869 ( .A1(n2783), .A2(n4490), .ZN(n3576) );
  AND2_X1 U2870 ( .A1(n2783), .A2(n2731), .ZN(n2725) );
  NAND2_X1 U2871 ( .A1(n3251), .A2(n2927), .ZN(n2968) );
  NAND2_X1 U2872 ( .A1(n3132), .A2(n3133), .ZN(n3304) );
  NAND2_X1 U2873 ( .A1(n3353), .A2(n3357), .ZN(n3287) );
  AND4_X1 U2874 ( .A1(n2296), .A2(n2310), .A3(n2300), .A4(n2298), .ZN(n2276)
         );
  AND2_X1 U2875 ( .A1(n2343), .A2(n2286), .ZN(n2277) );
  OAI22_X1 U2876 ( .A1(n2708), .A2(n3226), .B1(n2827), .B2(n2710), .ZN(n2756)
         );
  OR2_X1 U2877 ( .A1(n4334), .A2(n4588), .ZN(n2278) );
  OR2_X1 U2878 ( .A1(n2493), .A2(n3146), .ZN(n2280) );
  OR2_X1 U2879 ( .A1(n3240), .A2(n4231), .ZN(n2281) );
  OR2_X1 U2880 ( .A1(n3240), .A2(n4176), .ZN(n2282) );
  INV_X1 U2881 ( .A(IR_REG_27__SCAN_IN), .ZN(n2310) );
  OR2_X1 U2882 ( .A1(n3724), .A2(n3200), .ZN(n2283) );
  INV_X1 U2883 ( .A(IR_REG_26__SCAN_IN), .ZN(n2296) );
  NAND2_X1 U2884 ( .A1(n3270), .A2(n3189), .ZN(n3323) );
  OR2_X1 U2886 ( .A1(n3573), .A2(n2881), .ZN(n2284) );
  INV_X1 U2887 ( .A(n3865), .ZN(n2493) );
  INV_X1 U2888 ( .A(IR_REG_4__SCAN_IN), .ZN(n2286) );
  AND2_X1 U2889 ( .A1(n3191), .A2(n3192), .ZN(n3189) );
  OR2_X1 U2890 ( .A1(n3788), .A2(n2615), .ZN(n3529) );
  INV_X1 U2891 ( .A(IR_REG_25__SCAN_IN), .ZN(n2294) );
  INV_X1 U2892 ( .A(n3133), .ZN(n3134) );
  INV_X1 U2893 ( .A(IR_REG_29__SCAN_IN), .ZN(n2298) );
  INV_X1 U2894 ( .A(IR_REG_22__SCAN_IN), .ZN(n2293) );
  AND2_X1 U2895 ( .A1(n2453), .A2(REG3_REG_14__SCAN_IN), .ZN(n2463) );
  OR2_X1 U2896 ( .A1(n2545), .A2(n3327), .ZN(n2550) );
  NAND2_X1 U2897 ( .A1(n2335), .A2(REG1_REG_2__SCAN_IN), .ZN(n2327) );
  INV_X1 U2898 ( .A(n4472), .ZN(n4447) );
  OR2_X1 U2899 ( .A1(n3671), .A2(n3231), .ZN(n3107) );
  INV_X1 U2900 ( .A(n4449), .ZN(n4411) );
  NAND2_X1 U2901 ( .A1(n3446), .A2(n3450), .ZN(n3489) );
  NOR2_X1 U2902 ( .A1(n2375), .A2(n4098), .ZN(n2386) );
  INV_X1 U2903 ( .A(n3745), .ZN(n3707) );
  AND3_X1 U2904 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2369) );
  NAND2_X1 U2905 ( .A1(n2514), .A2(REG3_REG_20__SCAN_IN), .ZN(n2534) );
  OR2_X1 U2906 ( .A1(n2534), .A2(n2526), .ZN(n2535) );
  INV_X1 U2907 ( .A(n3685), .ZN(n3693) );
  NAND2_X1 U2908 ( .A1(n2463), .A2(REG3_REG_15__SCAN_IN), .ZN(n2484) );
  OR2_X1 U2909 ( .A1(n2550), .A2(n3299), .ZN(n2557) );
  INV_X1 U2910 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3346) );
  OR2_X1 U2911 ( .A1(n4258), .A2(n3557), .ZN(n4397) );
  AND2_X1 U2912 ( .A1(n3111), .A2(n3477), .ZN(n3665) );
  AND2_X1 U2913 ( .A1(n3741), .A2(n2617), .ZN(n3760) );
  INV_X1 U2914 ( .A(n4463), .ZN(n3892) );
  INV_X1 U2915 ( .A(n3927), .ZN(n2762) );
  OR2_X1 U2916 ( .A1(n2676), .A2(D_REG_0__SCAN_IN), .ZN(n2660) );
  AND2_X1 U2917 ( .A1(n2052), .A2(DATAI_24_), .ZN(n3187) );
  INV_X1 U2918 ( .A(n3857), .ZN(n3146) );
  INV_X1 U2919 ( .A(n4469), .ZN(n4453) );
  INV_X1 U2920 ( .A(n2715), .ZN(n2795) );
  AND2_X1 U2921 ( .A1(n2635), .A2(n2646), .ZN(n2657) );
  AND2_X1 U2922 ( .A1(n2053), .A2(DATAI_23_), .ZN(n3272) );
  AND2_X1 U2923 ( .A1(n2577), .A2(n2576), .ZN(n3671) );
  AND4_X1 U2924 ( .A1(n2540), .A2(n2539), .A3(n2538), .A4(n2537), .ZN(n3775)
         );
  AND4_X1 U2925 ( .A1(n2489), .A2(n2488), .A3(n2487), .A4(n2486), .ZN(n3865)
         );
  INV_X1 U2926 ( .A(n4270), .ZN(n4404) );
  INV_X1 U2927 ( .A(n4397), .ZN(n4345) );
  OR2_X1 U2928 ( .A1(n4466), .A2(n2805), .ZN(n3914) );
  NAND2_X1 U2929 ( .A1(n2660), .A2(n2659), .ZN(n2793) );
  INV_X1 U2930 ( .A(n2657), .ZN(n2676) );
  NAND2_X1 U2931 ( .A1(n2782), .A2(STATE_REG_SCAN_IN), .ZN(n4490) );
  OR2_X1 U2932 ( .A1(n2408), .A2(IR_REG_9__SCAN_IN), .ZN(n2425) );
  AND2_X1 U2933 ( .A1(n2392), .A2(n2383), .ZN(n4280) );
  AND2_X1 U2934 ( .A1(n2690), .A2(n2681), .ZN(n4402) );
  INV_X1 U2935 ( .A(n3344), .ZN(n3406) );
  INV_X1 U2936 ( .A(n3389), .ZN(n3696) );
  INV_X1 U2937 ( .A(n3775), .ZN(n3564) );
  INV_X1 U2938 ( .A(n3880), .ZN(n3566) );
  INV_X1 U2939 ( .A(n4505), .ZN(n4334) );
  OR2_X1 U2940 ( .A1(n4258), .A2(n4236), .ZN(n4409) );
  AND2_X1 U2941 ( .A1(n3914), .A2(n2806), .ZN(n3896) );
  NAND2_X1 U2943 ( .A1(n4590), .A2(n4569), .ZN(n4176) );
  OR2_X1 U2944 ( .A1(n2663), .A2(n2793), .ZN(n4587) );
  NAND2_X1 U2945 ( .A1(n4572), .A2(n4569), .ZN(n4231) );
  OR2_X1 U2946 ( .A1(n2663), .A2(n2662), .ZN(n4570) );
  NAND2_X1 U2947 ( .A1(n2676), .A2(n2725), .ZN(n4489) );
  INV_X1 U2948 ( .A(n3653), .ZN(n4494) );
  INV_X1 U2949 ( .A(n2342), .ZN(n2287) );
  NAND2_X1 U2950 ( .A1(n2629), .A2(n2294), .ZN(n2295) );
  INV_X1 U2951 ( .A(n2304), .ZN(n2673) );
  INV_X1 U2952 ( .A(IR_REG_28__SCAN_IN), .ZN(n2300) );
  INV_X1 U2953 ( .A(IR_REG_30__SCAN_IN), .ZN(n2667) );
  AND2_X2 U2954 ( .A1(n2304), .A2(n4235), .ZN(n2336) );
  NAND2_X1 U2955 ( .A1(n2337), .A2(REG0_REG_1__SCAN_IN), .ZN(n2305) );
  NAND2_X1 U2956 ( .A1(n2310), .A2(IR_REG_28__SCAN_IN), .ZN(n2311) );
  NAND2_X1 U2957 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2314)
         );
  NAND2_X1 U2958 ( .A1(n2333), .A2(REG3_REG_0__SCAN_IN), .ZN(n2320) );
  NAND2_X1 U2959 ( .A1(n2335), .A2(REG1_REG_0__SCAN_IN), .ZN(n2319) );
  NAND2_X1 U2960 ( .A1(n2336), .A2(REG2_REG_0__SCAN_IN), .ZN(n2318) );
  NAND2_X1 U2961 ( .A1(n2337), .A2(REG0_REG_0__SCAN_IN), .ZN(n2317) );
  AND2_X1 U2962 ( .A1(n3577), .A2(n4460), .ZN(n4443) );
  NAND2_X1 U2963 ( .A1(n2323), .A2(n4459), .ZN(n2324) );
  NAND2_X1 U2964 ( .A1(n2336), .A2(REG2_REG_2__SCAN_IN), .ZN(n2329) );
  NAND2_X1 U2965 ( .A1(n2333), .A2(REG3_REG_2__SCAN_IN), .ZN(n2326) );
  NAND2_X1 U2966 ( .A1(n2337), .A2(REG0_REG_2__SCAN_IN), .ZN(n2325) );
  AND3_X1 U2967 ( .A1(n2327), .A2(n2326), .A3(n2325), .ZN(n2328) );
  NAND2_X1 U2968 ( .A1(n2329), .A2(n2328), .ZN(n2331) );
  XNOR2_X2 U2969 ( .A(n2330), .B(IR_REG_2__SCAN_IN), .ZN(n4245) );
  MUX2_X1 U2970 ( .A(n4245), .B(DATAI_2_), .S(n2052), .Z(n3927) );
  NAND2_X1 U2971 ( .A1(n2815), .A2(n3927), .ZN(n3439) );
  NAND2_X1 U2972 ( .A1(n2331), .A2(n2762), .ZN(n3440) );
  NAND2_X1 U2973 ( .A1(n2815), .A2(n2762), .ZN(n2332) );
  INV_X1 U2974 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2334) );
  NAND2_X1 U2975 ( .A1(n2333), .A2(n2334), .ZN(n2341) );
  NAND2_X1 U2976 ( .A1(n2335), .A2(REG1_REG_3__SCAN_IN), .ZN(n2340) );
  NAND2_X1 U2977 ( .A1(n2350), .A2(REG2_REG_3__SCAN_IN), .ZN(n2339) );
  NAND2_X1 U2978 ( .A1(n2337), .A2(REG0_REG_3__SCAN_IN), .ZN(n2338) );
  NAND2_X1 U2979 ( .A1(n2342), .A2(IR_REG_31__SCAN_IN), .ZN(n2344) );
  NAND2_X1 U2980 ( .A1(n2344), .A2(n2343), .ZN(n2355) );
  OR2_X1 U2981 ( .A1(n2344), .A2(n2343), .ZN(n2345) );
  NOR2_X1 U2982 ( .A1(n3919), .A2(n3443), .ZN(n2348) );
  NAND2_X1 U2983 ( .A1(n3919), .A2(n3443), .ZN(n2347) );
  NAND2_X1 U2984 ( .A1(n2337), .A2(REG0_REG_4__SCAN_IN), .ZN(n2354) );
  NAND2_X1 U2985 ( .A1(n2335), .A2(REG1_REG_4__SCAN_IN), .ZN(n2353) );
  INV_X1 U2986 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2349) );
  XNOR2_X1 U2987 ( .A(n2349), .B(REG3_REG_3__SCAN_IN), .ZN(n3339) );
  NAND2_X1 U2988 ( .A1(n2333), .A2(n3339), .ZN(n2352) );
  NAND2_X1 U2989 ( .A1(n2350), .A2(REG2_REG_4__SCAN_IN), .ZN(n2351) );
  NAND2_X1 U2990 ( .A1(n2355), .A2(IR_REG_31__SCAN_IN), .ZN(n2356) );
  XNOR2_X1 U2991 ( .A(n2356), .B(IR_REG_4__SCAN_IN), .ZN(n4243) );
  MUX2_X1 U2992 ( .A(n4243), .B(DATAI_4_), .S(n2053), .Z(n2853) );
  NAND2_X1 U2993 ( .A1(n2829), .A2(n2853), .ZN(n3446) );
  NAND2_X1 U2994 ( .A1(n3575), .A2(n3336), .ZN(n3450) );
  NAND2_X1 U2995 ( .A1(n2851), .A2(n3489), .ZN(n2358) );
  NAND2_X1 U2996 ( .A1(n3575), .A2(n2853), .ZN(n2357) );
  NAND2_X1 U2997 ( .A1(n2358), .A2(n2357), .ZN(n2803) );
  NAND2_X1 U2998 ( .A1(n2337), .A2(REG0_REG_5__SCAN_IN), .ZN(n2365) );
  INV_X2 U2999 ( .A(n2359), .ZN(n2559) );
  NAND2_X1 U3000 ( .A1(n2559), .A2(REG1_REG_5__SCAN_IN), .ZN(n2364) );
  AOI21_X1 U3001 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2360) );
  NOR2_X1 U3002 ( .A1(n2360), .A2(n2369), .ZN(n2845) );
  NAND2_X1 U3003 ( .A1(n2333), .A2(n2845), .ZN(n2363) );
  NAND2_X1 U3004 ( .A1(n2350), .A2(REG2_REG_5__SCAN_IN), .ZN(n2362) );
  NAND4_X1 U3005 ( .A1(n2365), .A2(n2364), .A3(n2363), .A4(n2362), .ZN(n3574)
         );
  NAND2_X1 U3006 ( .A1(n2366), .A2(IR_REG_31__SCAN_IN), .ZN(n2367) );
  XNOR2_X1 U3007 ( .A(n2367), .B(IR_REG_5__SCAN_IN), .ZN(n4515) );
  MUX2_X1 U3008 ( .A(n4515), .B(DATAI_5_), .S(n2052), .Z(n2842) );
  AND2_X1 U3009 ( .A1(n3574), .A2(n2842), .ZN(n2368) );
  NAND2_X1 U3010 ( .A1(n2337), .A2(REG0_REG_6__SCAN_IN), .ZN(n2373) );
  NAND2_X1 U3011 ( .A1(n2559), .A2(REG1_REG_6__SCAN_IN), .ZN(n2372) );
  NAND2_X1 U3012 ( .A1(n2369), .A2(REG3_REG_6__SCAN_IN), .ZN(n2375) );
  OAI21_X1 U3013 ( .B1(n2369), .B2(REG3_REG_6__SCAN_IN), .A(n2375), .ZN(n2868)
         );
  INV_X1 U3014 ( .A(n2868), .ZN(n2889) );
  NAND2_X1 U3015 ( .A1(n2333), .A2(n2889), .ZN(n2371) );
  NAND2_X1 U3016 ( .A1(n2350), .A2(REG2_REG_6__SCAN_IN), .ZN(n2370) );
  NAND4_X1 U3017 ( .A1(n2373), .A2(n2372), .A3(n2371), .A4(n2370), .ZN(n3573)
         );
  NOR2_X1 U3018 ( .A1(n2366), .A2(IR_REG_5__SCAN_IN), .ZN(n2406) );
  OR2_X1 U3019 ( .A1(n2406), .A2(n2628), .ZN(n2374) );
  XNOR2_X1 U3020 ( .A(n2374), .B(IR_REG_6__SCAN_IN), .ZN(n3634) );
  MUX2_X1 U3021 ( .A(n3634), .B(DATAI_6_), .S(n2053), .Z(n2881) );
  NAND2_X1 U3022 ( .A1(n2337), .A2(REG0_REG_7__SCAN_IN), .ZN(n2380) );
  NAND2_X1 U3023 ( .A1(n2559), .A2(REG1_REG_7__SCAN_IN), .ZN(n2379) );
  AND2_X1 U3024 ( .A1(n2375), .A2(n4098), .ZN(n2376) );
  NOR2_X1 U3025 ( .A1(n2386), .A2(n2376), .ZN(n3255) );
  NAND2_X1 U3026 ( .A1(n2333), .A2(n3255), .ZN(n2378) );
  NAND2_X1 U3027 ( .A1(n2350), .A2(REG2_REG_7__SCAN_IN), .ZN(n2377) );
  NAND2_X1 U3028 ( .A1(n2406), .A2(n2404), .ZN(n2381) );
  NAND2_X1 U3029 ( .A1(n2381), .A2(IR_REG_31__SCAN_IN), .ZN(n2382) );
  NAND2_X1 U3030 ( .A1(n2382), .A2(n2403), .ZN(n2392) );
  OR2_X1 U3031 ( .A1(n2382), .A2(n2403), .ZN(n2383) );
  MUX2_X1 U3032 ( .A(n4280), .B(DATAI_7_), .S(n2052), .Z(n2920) );
  NAND2_X1 U3033 ( .A1(n2951), .A2(n2920), .ZN(n2603) );
  NAND2_X1 U3034 ( .A1(n3572), .A2(n3253), .ZN(n3456) );
  NAND2_X1 U3035 ( .A1(n2603), .A2(n3456), .ZN(n3491) );
  NAND2_X1 U3036 ( .A1(n2912), .A2(n3491), .ZN(n2385) );
  NAND2_X1 U3037 ( .A1(n3572), .A2(n2920), .ZN(n2384) );
  NAND2_X1 U3038 ( .A1(n2385), .A2(n2384), .ZN(n2947) );
  NAND2_X1 U3039 ( .A1(n2337), .A2(REG0_REG_8__SCAN_IN), .ZN(n2391) );
  NAND2_X1 U3040 ( .A1(n2559), .A2(REG1_REG_8__SCAN_IN), .ZN(n2390) );
  NAND2_X1 U3041 ( .A1(n2386), .A2(REG3_REG_8__SCAN_IN), .ZN(n2396) );
  OR2_X1 U3042 ( .A1(n2386), .A2(REG3_REG_8__SCAN_IN), .ZN(n2387) );
  AND2_X1 U3043 ( .A1(n2396), .A2(n2387), .ZN(n4435) );
  NAND2_X1 U3044 ( .A1(n2333), .A2(n4435), .ZN(n2389) );
  NAND2_X1 U3045 ( .A1(n2350), .A2(REG2_REG_8__SCAN_IN), .ZN(n2388) );
  NAND4_X1 U3046 ( .A1(n2391), .A2(n2390), .A3(n2389), .A4(n2388), .ZN(n3571)
         );
  NAND2_X1 U3047 ( .A1(n2392), .A2(IR_REG_31__SCAN_IN), .ZN(n2393) );
  XNOR2_X1 U3048 ( .A(n2393), .B(IR_REG_8__SCAN_IN), .ZN(n3636) );
  MUX2_X1 U3049 ( .A(n3636), .B(DATAI_8_), .S(n2053), .Z(n2949) );
  AND2_X1 U3050 ( .A1(n3571), .A2(n2949), .ZN(n2395) );
  NAND2_X1 U3051 ( .A1(n2928), .A2(n2956), .ZN(n2394) );
  NAND2_X1 U3052 ( .A1(n2337), .A2(REG0_REG_9__SCAN_IN), .ZN(n2401) );
  NAND2_X1 U3053 ( .A1(n2559), .A2(REG1_REG_9__SCAN_IN), .ZN(n2400) );
  NAND2_X1 U3054 ( .A1(n2396), .A2(n3346), .ZN(n2397) );
  AND2_X1 U3055 ( .A1(n2412), .A2(n2397), .ZN(n3349) );
  NAND2_X1 U3056 ( .A1(n2333), .A2(n3349), .ZN(n2399) );
  NAND2_X1 U3057 ( .A1(n2350), .A2(REG2_REG_9__SCAN_IN), .ZN(n2398) );
  NAND4_X1 U3058 ( .A1(n2401), .A2(n2400), .A3(n2399), .A4(n2398), .ZN(n3570)
         );
  INV_X1 U3059 ( .A(IR_REG_8__SCAN_IN), .ZN(n2402) );
  AND3_X1 U3060 ( .A1(n2404), .A2(n2403), .A3(n2402), .ZN(n2405) );
  NAND2_X1 U3061 ( .A1(n2406), .A2(n2405), .ZN(n2408) );
  NAND2_X1 U3062 ( .A1(n2408), .A2(IR_REG_31__SCAN_IN), .ZN(n2407) );
  MUX2_X1 U3063 ( .A(IR_REG_31__SCAN_IN), .B(n2407), .S(IR_REG_9__SCAN_IN), 
        .Z(n2409) );
  MUX2_X1 U3064 ( .A(n4300), .B(DATAI_9_), .S(n2052), .Z(n2941) );
  NOR2_X1 U3065 ( .A1(n3570), .A2(n2941), .ZN(n2411) );
  NAND2_X1 U3066 ( .A1(n2412), .A2(n2981), .ZN(n2413) );
  AND2_X1 U3067 ( .A1(n2431), .A2(n2413), .ZN(n4428) );
  NAND2_X1 U3068 ( .A1(n2333), .A2(n4428), .ZN(n2417) );
  NAND2_X1 U3069 ( .A1(n2559), .A2(REG1_REG_10__SCAN_IN), .ZN(n2416) );
  NAND2_X1 U3070 ( .A1(n2350), .A2(REG2_REG_10__SCAN_IN), .ZN(n2415) );
  NAND2_X1 U3071 ( .A1(n3412), .A2(REG0_REG_10__SCAN_IN), .ZN(n2414) );
  NAND4_X1 U3072 ( .A1(n2417), .A2(n2416), .A3(n2415), .A4(n2414), .ZN(n4412)
         );
  NAND2_X1 U3073 ( .A1(n2425), .A2(IR_REG_31__SCAN_IN), .ZN(n2418) );
  XNOR2_X1 U3074 ( .A(n2418), .B(IR_REG_10__SCAN_IN), .ZN(n4507) );
  MUX2_X1 U3075 ( .A(n4507), .B(DATAI_10_), .S(n2052), .Z(n3054) );
  AND2_X1 U3076 ( .A1(n4412), .A2(n3054), .ZN(n2419) );
  INV_X1 U3077 ( .A(n4412), .ZN(n3046) );
  NAND2_X1 U3078 ( .A1(n3046), .A2(n2098), .ZN(n2420) );
  NAND2_X1 U3079 ( .A1(n2337), .A2(REG0_REG_11__SCAN_IN), .ZN(n2424) );
  NAND2_X1 U3080 ( .A1(n2559), .A2(REG1_REG_11__SCAN_IN), .ZN(n2423) );
  XNOR2_X1 U3081 ( .A(n2431), .B(REG3_REG_11__SCAN_IN), .ZN(n4421) );
  NAND2_X1 U3082 ( .A1(n2333), .A2(n4421), .ZN(n2422) );
  NAND2_X1 U3083 ( .A1(n2350), .A2(REG2_REG_11__SCAN_IN), .ZN(n2421) );
  NAND2_X1 U3084 ( .A1(n2426), .A2(IR_REG_31__SCAN_IN), .ZN(n2438) );
  XNOR2_X1 U3085 ( .A(n2438), .B(IR_REG_11__SCAN_IN), .ZN(n4505) );
  MUX2_X1 U3086 ( .A(n4505), .B(DATAI_11_), .S(n2053), .Z(n4424) );
  NAND2_X1 U3087 ( .A1(n3056), .A2(n4424), .ZN(n3427) );
  INV_X1 U3088 ( .A(n4424), .ZN(n3048) );
  NAND2_X1 U3089 ( .A1(n3569), .A2(n3048), .ZN(n3425) );
  NAND2_X1 U3090 ( .A1(n3427), .A2(n3425), .ZN(n4416) );
  NOR2_X1 U3091 ( .A1(n3569), .A2(n4424), .ZN(n2427) );
  NAND2_X1 U3092 ( .A1(n2337), .A2(REG0_REG_12__SCAN_IN), .ZN(n2436) );
  NAND2_X1 U3093 ( .A1(n2559), .A2(REG1_REG_12__SCAN_IN), .ZN(n2435) );
  NAND2_X1 U3094 ( .A1(REG3_REG_12__SCAN_IN), .A2(REG3_REG_11__SCAN_IN), .ZN(
        n2428) );
  INV_X1 U3095 ( .A(n2443), .ZN(n2444) );
  INV_X1 U3096 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2430) );
  INV_X1 U3097 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2429) );
  OAI21_X1 U3098 ( .B1(n2431), .B2(n2430), .A(n2429), .ZN(n2432) );
  AND2_X1 U3099 ( .A1(n2444), .A2(n2432), .ZN(n3030) );
  NAND2_X1 U3100 ( .A1(n2333), .A2(n3030), .ZN(n2434) );
  NAND2_X1 U3101 ( .A1(n2350), .A2(REG2_REG_12__SCAN_IN), .ZN(n2433) );
  INV_X1 U3102 ( .A(IR_REG_11__SCAN_IN), .ZN(n2437) );
  NAND2_X1 U3103 ( .A1(n2438), .A2(n2437), .ZN(n2439) );
  NAND2_X1 U3104 ( .A1(n2439), .A2(IR_REG_31__SCAN_IN), .ZN(n2440) );
  XNOR2_X1 U3105 ( .A(n2440), .B(IR_REG_12__SCAN_IN), .ZN(n3644) );
  INV_X1 U3106 ( .A(n3644), .ZN(n4504) );
  INV_X1 U3107 ( .A(DATAI_12_), .ZN(n4503) );
  MUX2_X1 U3108 ( .A(n4504), .B(n4503), .S(n2053), .Z(n3027) );
  NAND2_X1 U3109 ( .A1(n4414), .A2(n3027), .ZN(n2442) );
  INV_X1 U3110 ( .A(n3027), .ZN(n3023) );
  AND2_X1 U3111 ( .A1(n3568), .A2(n3023), .ZN(n2441) );
  NAND2_X1 U3112 ( .A1(n2337), .A2(REG0_REG_13__SCAN_IN), .ZN(n2449) );
  NAND2_X1 U3113 ( .A1(n2559), .A2(REG1_REG_13__SCAN_IN), .ZN(n2448) );
  INV_X1 U3114 ( .A(n2453), .ZN(n2455) );
  INV_X1 U3115 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3097) );
  NAND2_X1 U3116 ( .A1(n2444), .A2(n3097), .ZN(n2445) );
  AND2_X1 U3117 ( .A1(n2455), .A2(n2445), .ZN(n3100) );
  NAND2_X1 U3118 ( .A1(n2333), .A2(n3100), .ZN(n2447) );
  NAND2_X1 U3119 ( .A1(n2350), .A2(REG2_REG_13__SCAN_IN), .ZN(n2446) );
  NAND4_X1 U3120 ( .A1(n2449), .A2(n2448), .A3(n2447), .A4(n2446), .ZN(n3567)
         );
  OR2_X1 U3121 ( .A1(n2080), .A2(n2628), .ZN(n2450) );
  XNOR2_X1 U3122 ( .A(n2450), .B(IR_REG_13__SCAN_IN), .ZN(n4501) );
  NAND2_X1 U3123 ( .A1(n3567), .A2(n3070), .ZN(n2452) );
  NOR2_X1 U3124 ( .A1(n3567), .A2(n3070), .ZN(n2451) );
  NAND2_X1 U3125 ( .A1(n3412), .A2(REG0_REG_14__SCAN_IN), .ZN(n2460) );
  NAND2_X1 U3126 ( .A1(n2559), .A2(REG1_REG_14__SCAN_IN), .ZN(n2459) );
  INV_X1 U3127 ( .A(n2463), .ZN(n2464) );
  INV_X1 U3128 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2454) );
  NAND2_X1 U3129 ( .A1(n2455), .A2(n2454), .ZN(n2456) );
  AND2_X1 U3130 ( .A1(n2464), .A2(n2456), .ZN(n3908) );
  NAND2_X1 U3131 ( .A1(n2333), .A2(n3908), .ZN(n2458) );
  NAND2_X1 U3132 ( .A1(n2350), .A2(REG2_REG_14__SCAN_IN), .ZN(n2457) );
  OR2_X1 U3133 ( .A1(n2461), .A2(n2628), .ZN(n2462) );
  XNOR2_X1 U3134 ( .A(n2462), .B(IR_REG_14__SCAN_IN), .ZN(n4499) );
  MUX2_X1 U3135 ( .A(n4499), .B(DATAI_14_), .S(n2052), .Z(n3910) );
  NAND2_X1 U3136 ( .A1(n3880), .A2(n3910), .ZN(n3877) );
  INV_X1 U3137 ( .A(n3910), .ZN(n3082) );
  NAND2_X1 U3138 ( .A1(n3566), .A2(n3082), .ZN(n3421) );
  NAND2_X1 U3139 ( .A1(n3412), .A2(REG0_REG_15__SCAN_IN), .ZN(n2469) );
  NAND2_X1 U3140 ( .A1(n2559), .A2(REG1_REG_15__SCAN_IN), .ZN(n2468) );
  INV_X1 U3141 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3400) );
  NAND2_X1 U3142 ( .A1(n2464), .A2(n3400), .ZN(n2465) );
  AND2_X1 U3143 ( .A1(n2484), .A2(n2465), .ZN(n3890) );
  NAND2_X1 U3144 ( .A1(n2333), .A2(n3890), .ZN(n2467) );
  NAND2_X1 U3145 ( .A1(n2350), .A2(REG2_REG_15__SCAN_IN), .ZN(n2466) );
  NAND4_X1 U3146 ( .A1(n2469), .A2(n2468), .A3(n2467), .A4(n2466), .ZN(n3900)
         );
  NAND2_X1 U3147 ( .A1(n2461), .A2(n2164), .ZN(n2470) );
  NAND2_X1 U31480 ( .A1(n2470), .A2(IR_REG_31__SCAN_IN), .ZN(n2471) );
  NAND2_X1 U31490 ( .A1(n2471), .A2(n2165), .ZN(n2478) );
  OR2_X1 U3150 ( .A1(n2471), .A2(n2165), .ZN(n2472) );
  MUX2_X1 U3151 ( .A(n3649), .B(DATAI_15_), .S(n2053), .Z(n3136) );
  NOR2_X1 U3152 ( .A1(n3900), .A2(n3136), .ZN(n2473) );
  NAND2_X1 U3153 ( .A1(n3412), .A2(REG0_REG_16__SCAN_IN), .ZN(n2477) );
  NAND2_X1 U3154 ( .A1(n2559), .A2(REG1_REG_16__SCAN_IN), .ZN(n2476) );
  XNOR2_X1 U3155 ( .A(n2484), .B(REG3_REG_16__SCAN_IN), .ZN(n3871) );
  NAND2_X1 U3156 ( .A1(n2333), .A2(n3871), .ZN(n2475) );
  NAND2_X1 U3157 ( .A1(n2350), .A2(REG2_REG_16__SCAN_IN), .ZN(n2474) );
  NAND2_X1 U3158 ( .A1(n2478), .A2(IR_REG_31__SCAN_IN), .ZN(n2479) );
  XNOR2_X1 U3159 ( .A(n2479), .B(IR_REG_16__SCAN_IN), .ZN(n3650) );
  MUX2_X1 U3160 ( .A(n3650), .B(DATAI_16_), .S(n2052), .Z(n2480) );
  NAND2_X1 U3161 ( .A1(n3882), .A2(n2480), .ZN(n3526) );
  NAND2_X1 U3162 ( .A1(n3853), .A2(n3870), .ZN(n3419) );
  NAND2_X1 U3163 ( .A1(n3526), .A2(n3419), .ZN(n3486) );
  NAND2_X1 U3164 ( .A1(n3412), .A2(REG0_REG_17__SCAN_IN), .ZN(n2489) );
  NAND2_X1 U3165 ( .A1(n2559), .A2(REG1_REG_17__SCAN_IN), .ZN(n2488) );
  INV_X1 U3166 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2482) );
  INV_X1 U3167 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2481) );
  OAI21_X1 U3168 ( .B1(n2484), .B2(n2482), .A(n2481), .ZN(n2485) );
  NAND2_X1 U3169 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .ZN(
        n2483) );
  AND2_X1 U3170 ( .A1(n2485), .A2(n2496), .ZN(n3858) );
  NAND2_X1 U3171 ( .A1(n2333), .A2(n3858), .ZN(n2487) );
  NAND2_X1 U3172 ( .A1(n2336), .A2(REG2_REG_17__SCAN_IN), .ZN(n2486) );
  NAND2_X1 U3173 ( .A1(n2490), .A2(IR_REG_31__SCAN_IN), .ZN(n2491) );
  XNOR2_X1 U3174 ( .A(n2491), .B(IR_REG_17__SCAN_IN), .ZN(n3653) );
  INV_X1 U3175 ( .A(DATAI_17_), .ZN(n2492) );
  MUX2_X1 U3176 ( .A(n4494), .B(n2492), .S(n2346), .Z(n3857) );
  NAND2_X1 U3177 ( .A1(n3848), .A2(n2494), .ZN(n2495) );
  NAND2_X1 U3178 ( .A1(n2495), .A2(n2280), .ZN(n3829) );
  NAND2_X1 U3179 ( .A1(n3412), .A2(REG0_REG_18__SCAN_IN), .ZN(n2501) );
  NAND2_X1 U3180 ( .A1(n2559), .A2(REG1_REG_18__SCAN_IN), .ZN(n2500) );
  INV_X1 U3181 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3378) );
  INV_X1 U3182 ( .A(n2504), .ZN(n2506) );
  NAND2_X1 U3183 ( .A1(n2496), .A2(n3378), .ZN(n2497) );
  AND2_X1 U3184 ( .A1(n2506), .A2(n2497), .ZN(n3842) );
  NAND2_X1 U3185 ( .A1(n2333), .A2(n3842), .ZN(n2499) );
  NAND2_X1 U3186 ( .A1(n2336), .A2(REG2_REG_18__SCAN_IN), .ZN(n2498) );
  NAND2_X1 U3187 ( .A1(n2089), .A2(IR_REG_31__SCAN_IN), .ZN(n2502) );
  XNOR2_X1 U3188 ( .A(n2502), .B(IR_REG_18__SCAN_IN), .ZN(n3654) );
  MUX2_X1 U3189 ( .A(n3654), .B(DATAI_18_), .S(n2053), .Z(n3834) );
  NAND2_X1 U3190 ( .A1(n3851), .A2(n3834), .ZN(n3811) );
  INV_X1 U3191 ( .A(n3851), .ZN(n3565) );
  NAND2_X1 U3192 ( .A1(n3565), .A2(n3841), .ZN(n3812) );
  NAND2_X1 U3193 ( .A1(n3811), .A2(n3812), .ZN(n3830) );
  AOI21_X1 U3194 ( .B1(n3829), .B2(n3830), .A(n2503), .ZN(n3805) );
  NAND2_X1 U3195 ( .A1(n3412), .A2(REG0_REG_19__SCAN_IN), .ZN(n2511) );
  NAND2_X1 U3196 ( .A1(n2559), .A2(REG1_REG_19__SCAN_IN), .ZN(n2510) );
  INV_X1 U3197 ( .A(n2514), .ZN(n2515) );
  INV_X1 U3198 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2505) );
  NAND2_X1 U3199 ( .A1(n2506), .A2(n2505), .ZN(n2507) );
  AND2_X1 U3200 ( .A1(n2515), .A2(n2507), .ZN(n3824) );
  NAND2_X1 U3201 ( .A1(n2333), .A2(n3824), .ZN(n2509) );
  NAND2_X1 U3202 ( .A1(n2336), .A2(REG2_REG_19__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U3203 ( .A1(n2512), .A2(IR_REG_31__SCAN_IN), .ZN(n2585) );
  INV_X1 U3204 ( .A(DATAI_19_), .ZN(n4067) );
  NAND2_X1 U3205 ( .A1(n3833), .A2(n3823), .ZN(n2513) );
  INV_X1 U3206 ( .A(n3823), .ZN(n3817) );
  NAND2_X1 U3207 ( .A1(n3412), .A2(REG0_REG_20__SCAN_IN), .ZN(n2520) );
  NAND2_X1 U3208 ( .A1(n2559), .A2(REG1_REG_20__SCAN_IN), .ZN(n2519) );
  INV_X1 U3209 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3359) );
  NAND2_X1 U32100 ( .A1(n2515), .A2(n3359), .ZN(n2516) );
  AND2_X1 U32110 ( .A1(n2534), .A2(n2516), .ZN(n3800) );
  NAND2_X1 U32120 ( .A1(n2333), .A2(n3800), .ZN(n2518) );
  NAND2_X1 U32130 ( .A1(n2336), .A2(REG2_REG_20__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U32140 ( .A1(n3818), .A2(n3163), .ZN(n3508) );
  NOR2_X1 U32150 ( .A1(n3818), .A2(n3163), .ZN(n3510) );
  XNOR2_X1 U32160 ( .A(n2534), .B(REG3_REG_21__SCAN_IN), .ZN(n3782) );
  NAND2_X1 U32170 ( .A1(n2333), .A2(n3782), .ZN(n2524) );
  NAND2_X1 U32180 ( .A1(n2559), .A2(REG1_REG_21__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U32190 ( .A1(n2336), .A2(REG2_REG_21__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U32200 ( .A1(n3412), .A2(REG0_REG_21__SCAN_IN), .ZN(n2521) );
  NAND2_X1 U32210 ( .A1(n3793), .A2(n3780), .ZN(n2525) );
  NAND2_X1 U32220 ( .A1(n3412), .A2(REG0_REG_23__SCAN_IN), .ZN(n2533) );
  NAND2_X1 U32230 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2526) );
  INV_X1 U32240 ( .A(n2535), .ZN(n2527) );
  NAND2_X1 U32250 ( .A1(n2527), .A2(REG3_REG_23__SCAN_IN), .ZN(n2545) );
  INV_X1 U32260 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2528) );
  NAND2_X1 U32270 ( .A1(n2535), .A2(n2528), .ZN(n2529) );
  AND2_X1 U32280 ( .A1(n2545), .A2(n2529), .ZN(n3751) );
  NAND2_X1 U32290 ( .A1(n3751), .A2(n2333), .ZN(n2532) );
  NAND2_X1 U32300 ( .A1(n2559), .A2(REG1_REG_23__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U32310 ( .A1(n2350), .A2(REG2_REG_23__SCAN_IN), .ZN(n2530) );
  NAND4_X1 U32320 ( .A1(n2533), .A2(n2532), .A3(n2531), .A4(n2530), .ZN(n3761)
         );
  NOR2_X1 U32330 ( .A1(n3761), .A2(n3272), .ZN(n2541) );
  NAND2_X1 U32340 ( .A1(n3412), .A2(REG0_REG_22__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U32350 ( .A1(n2559), .A2(REG1_REG_22__SCAN_IN), .ZN(n2539) );
  INV_X1 U32360 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3288) );
  INV_X1 U32370 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3367) );
  OAI21_X1 U32380 ( .B1(n2534), .B2(n3288), .A(n3367), .ZN(n2536) );
  AND2_X1 U32390 ( .A1(n2536), .A2(n2535), .ZN(n3766) );
  NAND2_X1 U32400 ( .A1(n2333), .A2(n3766), .ZN(n2538) );
  NAND2_X1 U32410 ( .A1(n2350), .A2(REG2_REG_22__SCAN_IN), .ZN(n2537) );
  NAND2_X1 U32420 ( .A1(n3775), .A2(n3767), .ZN(n3741) );
  INV_X1 U32430 ( .A(n3767), .ZN(n3368) );
  NAND2_X1 U32440 ( .A1(n3564), .A2(n3368), .ZN(n2617) );
  NAND2_X1 U32450 ( .A1(n3564), .A2(n3767), .ZN(n3735) );
  INV_X1 U32460 ( .A(n3761), .ZN(n3722) );
  INV_X1 U32470 ( .A(n3272), .ZN(n3750) );
  OAI22_X1 U32480 ( .A1(n2541), .A2(n3735), .B1(n3722), .B2(n3750), .ZN(n2542)
         );
  INV_X1 U32490 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4095) );
  NAND2_X1 U32500 ( .A1(n3412), .A2(REG0_REG_24__SCAN_IN), .ZN(n2544) );
  NAND2_X1 U32510 ( .A1(n2559), .A2(REG1_REG_24__SCAN_IN), .ZN(n2543) );
  AND2_X1 U32520 ( .A1(n2544), .A2(n2543), .ZN(n2548) );
  INV_X1 U32530 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3327) );
  NAND2_X1 U32540 ( .A1(n2545), .A2(n3327), .ZN(n2546) );
  NAND2_X1 U32550 ( .A1(n2550), .A2(n2546), .ZN(n3326) );
  OAI211_X1 U32560 ( .C1(n2361), .C2(n4095), .A(n2548), .B(n2547), .ZN(n3745)
         );
  NAND2_X1 U32570 ( .A1(n3745), .A2(n3187), .ZN(n2549) );
  INV_X1 U32580 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3299) );
  NAND2_X1 U32590 ( .A1(n2550), .A2(n3299), .ZN(n2551) );
  NAND2_X1 U32600 ( .A1(n2557), .A2(n2551), .ZN(n3297) );
  AOI22_X1 U32610 ( .A1(n2336), .A2(REG2_REG_25__SCAN_IN), .B1(n2559), .B2(
        REG1_REG_25__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U32620 ( .A1(n3412), .A2(REG0_REG_25__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U32630 ( .A1(n3701), .A2(n2283), .ZN(n2555) );
  INV_X1 U32640 ( .A(n3724), .ZN(n3694) );
  INV_X1 U32650 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3687) );
  INV_X1 U32660 ( .A(n2557), .ZN(n2556) );
  NAND2_X1 U32670 ( .A1(n2556), .A2(REG3_REG_26__SCAN_IN), .ZN(n2564) );
  INV_X1 U32680 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3390) );
  NAND2_X1 U32690 ( .A1(n2557), .A2(n3390), .ZN(n2558) );
  NAND2_X1 U32700 ( .A1(n2564), .A2(n2558), .ZN(n3686) );
  AOI22_X1 U32710 ( .A1(n3412), .A2(REG0_REG_26__SCAN_IN), .B1(n2559), .B2(
        REG1_REG_26__SCAN_IN), .ZN(n2560) );
  NAND2_X1 U32720 ( .A1(n3709), .A2(n3685), .ZN(n2562) );
  INV_X1 U32730 ( .A(n2564), .ZN(n2563) );
  NAND2_X1 U32740 ( .A1(n2563), .A2(REG3_REG_27__SCAN_IN), .ZN(n2571) );
  INV_X1 U32750 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3262) );
  NAND2_X1 U32760 ( .A1(n2564), .A2(n3262), .ZN(n2565) );
  NAND2_X1 U32770 ( .A1(n2571), .A2(n2565), .ZN(n3261) );
  OR2_X1 U32780 ( .A1(n3261), .A2(n2595), .ZN(n2570) );
  INV_X1 U32790 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4061) );
  NAND2_X1 U32800 ( .A1(n2336), .A2(REG2_REG_27__SCAN_IN), .ZN(n2567) );
  NAND2_X1 U32810 ( .A1(n3412), .A2(REG0_REG_27__SCAN_IN), .ZN(n2566) );
  OAI211_X1 U32820 ( .C1(n4061), .C2(n2359), .A(n2567), .B(n2566), .ZN(n2568)
         );
  INV_X1 U32830 ( .A(n2568), .ZN(n2569) );
  NAND2_X1 U32840 ( .A1(n2346), .A2(DATAI_27_), .ZN(n3676) );
  INV_X1 U32850 ( .A(n3676), .ZN(n3669) );
  INV_X1 U32860 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3230) );
  NAND2_X1 U32870 ( .A1(n2571), .A2(n3230), .ZN(n2572) );
  NAND2_X1 U32880 ( .A1(n3238), .A2(n2333), .ZN(n2577) );
  INV_X1 U32890 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4115) );
  NAND2_X1 U32900 ( .A1(n3412), .A2(REG0_REG_28__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U32910 ( .A1(n2336), .A2(REG2_REG_28__SCAN_IN), .ZN(n2573) );
  OAI211_X1 U32920 ( .C1(n2359), .C2(n4115), .A(n2574), .B(n2573), .ZN(n2575)
         );
  INV_X1 U32930 ( .A(n2575), .ZN(n2576) );
  AND2_X1 U32940 ( .A1(n2346), .A2(DATAI_28_), .ZN(n2578) );
  NAND2_X1 U32950 ( .A1(n3671), .A2(n2578), .ZN(n3112) );
  INV_X1 U32960 ( .A(n3671), .ZN(n3563) );
  NAND2_X1 U32970 ( .A1(n3563), .A2(n3231), .ZN(n3408) );
  NAND2_X1 U32980 ( .A1(n2074), .A2(IR_REG_31__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U32990 ( .A1(n2580), .A2(n2625), .ZN(n2705) );
  NAND2_X1 U33000 ( .A1(n2112), .A2(IR_REG_31__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U33010 ( .A1(n2585), .A2(n2584), .ZN(n2586) );
  NAND2_X1 U33020 ( .A1(n2586), .A2(IR_REG_31__SCAN_IN), .ZN(n2588) );
  XNOR2_X1 U33030 ( .A(n2705), .B(n2804), .ZN(n2589) );
  NAND2_X1 U33040 ( .A1(n2589), .A2(n3659), .ZN(n4417) );
  INV_X1 U33050 ( .A(n3659), .ZN(n4242) );
  AND2_X1 U33060 ( .A1(n2652), .A2(n4242), .ZN(n4475) );
  NAND2_X1 U33070 ( .A1(n2705), .A2(n4475), .ZN(n4563) );
  NAND2_X1 U33080 ( .A1(n4417), .A2(n4563), .ZN(n4554) );
  INV_X1 U33090 ( .A(n4554), .ZN(n4557) );
  XNOR2_X1 U33100 ( .A(n2590), .B(IR_REG_28__SCAN_IN), .ZN(n2741) );
  NOR2_X1 U33110 ( .A1(n2705), .A2(n2596), .ZN(n2718) );
  NAND2_X1 U33120 ( .A1(n2741), .A2(n2718), .ZN(n4472) );
  INV_X1 U33130 ( .A(REG1_REG_29__SCAN_IN), .ZN(n4003) );
  NAND2_X1 U33140 ( .A1(n2336), .A2(REG2_REG_29__SCAN_IN), .ZN(n2592) );
  NAND2_X1 U33150 ( .A1(n3412), .A2(REG0_REG_29__SCAN_IN), .ZN(n2591) );
  OAI211_X1 U33160 ( .C1(n2359), .C2(n4003), .A(n2592), .B(n2591), .ZN(n2593)
         );
  INV_X1 U33170 ( .A(n2593), .ZN(n2594) );
  OAI21_X1 U33180 ( .B1(n3118), .B2(n2595), .A(n2594), .ZN(n3411) );
  NOR2_X2 U33190 ( .A1(n4473), .A2(n2652), .ZN(n4446) );
  OAI22_X1 U33200 ( .A1(n3389), .A2(n4449), .B1(n3881), .B2(n3231), .ZN(n2624)
         );
  NAND2_X1 U33210 ( .A1(n4455), .A2(n2597), .ZN(n2599) );
  NAND2_X1 U33220 ( .A1(n2599), .A2(n3490), .ZN(n3922) );
  NAND2_X1 U33230 ( .A1(n3922), .A2(n3439), .ZN(n2600) );
  XNOR2_X1 U33240 ( .A(n3919), .B(n3443), .ZN(n3515) );
  INV_X1 U33250 ( .A(n3919), .ZN(n3442) );
  NAND2_X1 U33260 ( .A1(n3442), .A2(n3443), .ZN(n3445) );
  INV_X1 U33270 ( .A(n3446), .ZN(n2601) );
  AND2_X1 U33280 ( .A1(n3574), .A2(n2155), .ZN(n2798) );
  NAND2_X1 U33290 ( .A1(n2152), .A2(n2842), .ZN(n3435) );
  OAI21_X1 U33300 ( .B1(n2799), .B2(n2798), .A(n3435), .ZN(n2863) );
  INV_X1 U33310 ( .A(n2881), .ZN(n2887) );
  NAND2_X1 U33320 ( .A1(n3573), .A2(n2887), .ZN(n3448) );
  INV_X1 U33330 ( .A(n3573), .ZN(n2602) );
  NAND2_X1 U33340 ( .A1(n2602), .A2(n2881), .ZN(n3452) );
  INV_X1 U33350 ( .A(n2603), .ZN(n2604) );
  NAND2_X1 U33360 ( .A1(n2928), .A2(n2949), .ZN(n3458) );
  NAND2_X1 U33370 ( .A1(n2948), .A2(n3458), .ZN(n2605) );
  NAND2_X1 U33380 ( .A1(n3571), .A2(n2956), .ZN(n3455) );
  AND2_X1 U33390 ( .A1(n3570), .A2(n3347), .ZN(n2935) );
  NAND2_X1 U33400 ( .A1(n2969), .A2(n2941), .ZN(n3459) );
  NAND2_X1 U33410 ( .A1(n4412), .A2(n2098), .ZN(n3424) );
  NAND2_X1 U33420 ( .A1(n3046), .A2(n3054), .ZN(n3423) );
  NAND2_X1 U33430 ( .A1(n2606), .A2(n3423), .ZN(n4410) );
  NOR2_X1 U33440 ( .A1(n3568), .A2(n3027), .ZN(n3429) );
  INV_X1 U33450 ( .A(n3070), .ZN(n3098) );
  NAND2_X1 U33460 ( .A1(n3567), .A2(n3098), .ZN(n2998) );
  NAND2_X1 U33470 ( .A1(n3568), .A2(n3027), .ZN(n2996) );
  INV_X1 U33480 ( .A(n3567), .ZN(n3902) );
  NAND2_X1 U33490 ( .A1(n3902), .A2(n3070), .ZN(n3432) );
  NAND2_X1 U33500 ( .A1(n3309), .A2(n3136), .ZN(n3523) );
  NAND2_X1 U33510 ( .A1(n3900), .A2(n3889), .ZN(n3422) );
  NAND2_X1 U33520 ( .A1(n3523), .A2(n3422), .ZN(n3879) );
  INV_X1 U3353 ( .A(n3877), .ZN(n3525) );
  NOR2_X1 U33540 ( .A1(n3879), .A2(n3525), .ZN(n2608) );
  NAND2_X1 U3355 ( .A1(n3897), .A2(n2608), .ZN(n2609) );
  NAND2_X1 U3356 ( .A1(n2609), .A2(n3422), .ZN(n3864) );
  NAND2_X1 U3357 ( .A1(n3795), .A2(n3823), .ZN(n2610) );
  AND2_X1 U3358 ( .A1(n3812), .A2(n2610), .ZN(n2611) );
  NAND2_X1 U3359 ( .A1(n2493), .A2(n3857), .ZN(n3807) );
  NAND2_X1 U3360 ( .A1(n2611), .A2(n3807), .ZN(n3420) );
  NAND2_X1 U3361 ( .A1(n3865), .A2(n3146), .ZN(n3809) );
  NAND2_X1 U3362 ( .A1(n3811), .A2(n3809), .ZN(n2612) );
  NAND2_X1 U3363 ( .A1(n2612), .A2(n2611), .ZN(n2614) );
  NAND2_X1 U3364 ( .A1(n3833), .A2(n3817), .ZN(n2613) );
  NAND2_X1 U3365 ( .A1(n2614), .A2(n2613), .ZN(n3788) );
  NOR2_X1 U3366 ( .A1(n3818), .A2(n3799), .ZN(n2615) );
  NAND2_X1 U3367 ( .A1(n3529), .A2(n2209), .ZN(n3470) );
  NAND2_X1 U3368 ( .A1(n3793), .A2(n3171), .ZN(n3739) );
  INV_X1 U3369 ( .A(n3532), .ZN(n2618) );
  NOR2_X1 U3370 ( .A1(n3793), .A2(n3171), .ZN(n3737) );
  NAND2_X1 U3371 ( .A1(n3761), .A2(n3750), .ZN(n3505) );
  NAND2_X1 U3372 ( .A1(n2617), .A2(n3505), .ZN(n3475) );
  AOI21_X1 U3373 ( .B1(n3737), .B2(n3741), .A(n3475), .ZN(n3535) );
  NAND2_X1 U3374 ( .A1(n3707), .A2(n3187), .ZN(n3504) );
  NAND2_X1 U3375 ( .A1(n3722), .A2(n3272), .ZN(n3718) );
  NAND2_X1 U3376 ( .A1(n3298), .A2(n3685), .ZN(n3497) );
  OR2_X1 U3377 ( .A1(n3724), .A2(n3712), .ZN(n3689) );
  NAND2_X1 U3378 ( .A1(n3497), .A2(n3689), .ZN(n3541) );
  INV_X1 U3379 ( .A(n3541), .ZN(n3473) );
  NAND2_X1 U3380 ( .A1(n3724), .A2(n3712), .ZN(n3511) );
  NAND2_X1 U3381 ( .A1(n3745), .A2(n3728), .ZN(n3702) );
  AND2_X1 U3382 ( .A1(n3511), .A2(n3702), .ZN(n3537) );
  NAND2_X1 U3383 ( .A1(n3709), .A2(n3693), .ZN(n3521) );
  OAI21_X1 U3384 ( .B1(n3541), .B2(n3537), .A(n3521), .ZN(n3418) );
  NAND2_X1 U3385 ( .A1(n3389), .A2(n3669), .ZN(n3111) );
  NAND2_X1 U3386 ( .A1(n3696), .A2(n3676), .ZN(n3477) );
  INV_X1 U3387 ( .A(n3111), .ZN(n2619) );
  NOR2_X1 U3388 ( .A1(n3668), .A2(n2619), .ZN(n2620) );
  XNOR2_X1 U3389 ( .A(n2620), .B(n3501), .ZN(n2622) );
  NAND2_X1 U3390 ( .A1(n4240), .A2(n4241), .ZN(n2621) );
  OAI21_X2 U3391 ( .B1(n2705), .B2(n3659), .A(n2621), .ZN(n4469) );
  NOR2_X1 U3392 ( .A1(n2622), .A2(n4453), .ZN(n2623) );
  INV_X1 U3393 ( .A(IR_REG_23__SCAN_IN), .ZN(n2648) );
  NAND2_X1 U3394 ( .A1(n2649), .A2(n2648), .ZN(n2651) );
  INV_X1 U3395 ( .A(IR_REG_24__SCAN_IN), .ZN(n2626) );
  OR2_X1 U3396 ( .A1(n2629), .A2(n2628), .ZN(n2630) );
  NAND2_X1 U3397 ( .A1(n2649), .A2(n2630), .ZN(n2631) );
  INV_X1 U3398 ( .A(n4238), .ZN(n2653) );
  NAND2_X1 U3399 ( .A1(n3104), .A2(n2653), .ZN(n2632) );
  MUX2_X1 U3400 ( .A(n3104), .B(n2632), .S(B_REG_SCAN_IN), .Z(n2635) );
  NOR4_X1 U3401 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2644) );
  NOR4_X1 U3402 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2643) );
  INV_X1 U3403 ( .A(D_REG_18__SCAN_IN), .ZN(n4486) );
  INV_X1 U3404 ( .A(D_REG_3__SCAN_IN), .ZN(n4487) );
  INV_X1 U3405 ( .A(D_REG_22__SCAN_IN), .ZN(n4484) );
  INV_X1 U3406 ( .A(D_REG_21__SCAN_IN), .ZN(n4485) );
  NAND4_X1 U3407 ( .A1(n4486), .A2(n4487), .A3(n4484), .A4(n4485), .ZN(n2641)
         );
  NOR4_X1 U3408 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2639) );
  NOR4_X1 U3409 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2638) );
  NOR4_X1 U3410 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2637) );
  NOR4_X1 U3411 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2636) );
  NAND4_X1 U3412 ( .A1(n2639), .A2(n2638), .A3(n2637), .A4(n2636), .ZN(n2640)
         );
  NOR4_X1 U3413 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(n2641), 
        .A4(n2640), .ZN(n2642) );
  NAND3_X1 U3414 ( .A1(n2644), .A2(n2643), .A3(n2642), .ZN(n2645) );
  NAND2_X1 U3415 ( .A1(n2646), .A2(n4238), .ZN(n2647) );
  OR2_X1 U3416 ( .A1(n2649), .A2(n2648), .ZN(n2650) );
  NAND2_X1 U3417 ( .A1(n2651), .A2(n2650), .ZN(n2782) );
  NAND2_X1 U3418 ( .A1(n2652), .A2(n3659), .ZN(n2717) );
  NAND2_X1 U3419 ( .A1(n2718), .A2(n2717), .ZN(n2781) );
  NAND2_X1 U3420 ( .A1(n2725), .A2(n2781), .ZN(n2729) );
  NOR2_X1 U3421 ( .A1(n4563), .A2(n4240), .ZN(n2727) );
  NOR2_X1 U3422 ( .A1(n2729), .A2(n2727), .ZN(n2656) );
  INV_X1 U3423 ( .A(D_REG_1__SCAN_IN), .ZN(n2678) );
  NAND2_X1 U3424 ( .A1(n2657), .A2(n2678), .ZN(n2655) );
  INV_X1 U3425 ( .A(n2646), .ZN(n2658) );
  NAND2_X1 U3426 ( .A1(n2658), .A2(n2653), .ZN(n2654) );
  NAND2_X1 U3427 ( .A1(n2655), .A2(n2654), .ZN(n2792) );
  NAND3_X1 U3428 ( .A1(n2795), .A2(n2656), .A3(n2792), .ZN(n2663) );
  NAND2_X1 U3429 ( .A1(n3104), .A2(n2658), .ZN(n2659) );
  NAND2_X1 U3430 ( .A1(n3926), .A2(n2762), .ZN(n4528) );
  OAI21_X1 U3431 ( .B1(n3674), .B2(n3231), .A(n3110), .ZN(n3240) );
  NAND2_X1 U3432 ( .A1(n2661), .A2(n2282), .ZN(U3546) );
  INV_X1 U3433 ( .A(n2793), .ZN(n2662) );
  INV_X1 U3434 ( .A(n2665), .ZN(n2666) );
  NAND2_X1 U3435 ( .A1(n2666), .A2(n2281), .ZN(U3514) );
  INV_X2 U3436 ( .A(n3576), .ZN(U4043) );
  INV_X2 U3437 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND3_X1 U3438 ( .A1(n2667), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n2669) );
  INV_X1 U3439 ( .A(DATAI_31_), .ZN(n2668) );
  OAI22_X1 U3440 ( .A1(n2670), .A2(n2669), .B1(STATE_REG_SCAN_IN), .B2(n2668), 
        .ZN(U3321) );
  INV_X1 U3441 ( .A(DATAI_24_), .ZN(n2671) );
  MUX2_X1 U3442 ( .A(n2671), .B(n3104), .S(STATE_REG_SCAN_IN), .Z(n2672) );
  INV_X1 U3443 ( .A(n2672), .ZN(U3328) );
  INV_X1 U3444 ( .A(DATAI_29_), .ZN(n2675) );
  NAND2_X1 U3445 ( .A1(n2673), .A2(STATE_REG_SCAN_IN), .ZN(n2674) );
  OAI21_X1 U3446 ( .B1(STATE_REG_SCAN_IN), .B2(n2675), .A(n2674), .ZN(U3323)
         );
  NOR3_X1 U3447 ( .A1(n4238), .A2(n2646), .A3(n4490), .ZN(n2677) );
  AOI21_X1 U3448 ( .B1(n4489), .B2(n2678), .A(n2677), .ZN(U3459) );
  INV_X1 U3449 ( .A(n2725), .ZN(n2724) );
  INV_X1 U3450 ( .A(n2782), .ZN(n2679) );
  NAND2_X1 U3451 ( .A1(n2679), .A2(STATE_REG_SCAN_IN), .ZN(n3561) );
  NAND2_X1 U3452 ( .A1(n2724), .A2(n3561), .ZN(n2690) );
  NAND2_X1 U3453 ( .A1(n2718), .A2(n2782), .ZN(n2680) );
  AND2_X1 U3454 ( .A1(n2053), .A2(n2680), .ZN(n2689) );
  INV_X1 U3455 ( .A(n2689), .ZN(n2681) );
  NOR2_X1 U3456 ( .A1(n4402), .A2(U4043), .ZN(U3148) );
  NAND2_X1 U3457 ( .A1(n3576), .A2(DATAO_REG_21__SCAN_IN), .ZN(n2682) );
  OAI21_X1 U34580 ( .B1(n3793), .B2(n3576), .A(n2682), .ZN(U3571) );
  INV_X1 U34590 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4057) );
  NAND2_X1 U3460 ( .A1(n2559), .A2(REG1_REG_30__SCAN_IN), .ZN(n2685) );
  NAND2_X1 U3461 ( .A1(n2336), .A2(REG2_REG_30__SCAN_IN), .ZN(n2684) );
  NAND2_X1 U3462 ( .A1(n2337), .A2(REG0_REG_30__SCAN_IN), .ZN(n2683) );
  NAND3_X1 U3463 ( .A1(n2685), .A2(n2684), .A3(n2683), .ZN(n3478) );
  NAND2_X1 U3464 ( .A1(n3478), .A2(U4043), .ZN(n2686) );
  OAI21_X1 U3465 ( .B1(U4043), .B2(n4057), .A(n2686), .ZN(U3580) );
  INV_X1 U3466 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4062) );
  NAND2_X1 U34670 ( .A1(n3818), .A2(U4043), .ZN(n2687) );
  OAI21_X1 U3468 ( .B1(n4062), .B2(U4043), .A(n2687), .ZN(U3570) );
  INV_X1 U34690 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4039) );
  NAND2_X1 U3470 ( .A1(n3761), .A2(U4043), .ZN(n2688) );
  OAI21_X1 U34710 ( .B1(U4043), .B2(n4039), .A(n2688), .ZN(U3573) );
  NAND2_X1 U3472 ( .A1(n2690), .A2(n2689), .ZN(n4258) );
  INV_X1 U34730 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3925) );
  MUX2_X1 U3474 ( .A(REG2_REG_2__SCAN_IN), .B(n3925), .S(n4245), .Z(n2694) );
  INV_X1 U34750 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2691) );
  AND2_X1 U3476 ( .A1(REG2_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2692)
         );
  NAND2_X1 U34770 ( .A1(n3593), .A2(n3592), .ZN(n2693) );
  XNOR2_X1 U3478 ( .A(n2309), .B(IR_REG_27__SCAN_IN), .ZN(n4237) );
  INV_X1 U34790 ( .A(n4237), .ZN(n4254) );
  OR2_X1 U3480 ( .A1(n4254), .A2(n2741), .ZN(n3557) );
  OAI211_X1 U34810 ( .C1(REG2_REG_3__SCAN_IN), .C2(n2695), .A(n4345), .B(n2746), .ZN(n2697) );
  NOR2_X1 U3482 ( .A1(STATE_REG_SCAN_IN), .A2(n2334), .ZN(n2788) );
  AOI21_X1 U34830 ( .B1(n4402), .B2(ADDR_REG_3__SCAN_IN), .A(n2788), .ZN(n2696) );
  OAI211_X1 U3484 ( .C1(n4409), .C2(n2218), .A(n2697), .B(n2696), .ZN(n2702)
         );
  INV_X1 U34850 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4578) );
  INV_X1 U3486 ( .A(n4245), .ZN(n3590) );
  INV_X1 U34870 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2699) );
  MUX2_X1 U3488 ( .A(REG1_REG_2__SCAN_IN), .B(n2699), .S(n4245), .Z(n3599) );
  INV_X1 U34890 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4575) );
  AND2_X1 U3490 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3582)
         );
  NAND2_X1 U34910 ( .A1(n3581), .A2(n2698), .ZN(n3598) );
  NAND2_X1 U3492 ( .A1(n3599), .A2(n3598), .ZN(n3597) );
  OAI21_X1 U34930 ( .B1(n3590), .B2(n2699), .A(n3597), .ZN(n2750) );
  AOI211_X1 U3494 ( .C1(n4578), .C2(n2700), .A(n2749), .B(n4270), .ZN(n2701)
         );
  OR2_X1 U34950 ( .A1(n2702), .A2(n2701), .ZN(U3243) );
  INV_X1 U3496 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n2704) );
  NAND2_X1 U34970 ( .A1(n3411), .A2(U4043), .ZN(n2703) );
  OAI21_X1 U3498 ( .B1(U4043), .B2(n2704), .A(n2703), .ZN(U3579) );
  NAND2_X4 U34990 ( .A1(n2783), .A2(n2706), .ZN(n3222) );
  INV_X1 U3500 ( .A(n2705), .ZN(n4239) );
  NAND2_X1 U35010 ( .A1(n4239), .A2(n3659), .ZN(n2730) );
  AND2_X2 U3502 ( .A1(n2730), .A2(n2706), .ZN(n3198) );
  NAND2_X4 U35030 ( .A1(n2709), .A2(n4548), .ZN(n3226) );
  XNOR2_X1 U3504 ( .A(n2757), .B(n2756), .ZN(n2760) );
  OAI222_X1 U35050 ( .A1(n4474), .A2(n2827), .B1(n3226), .B2(n4450), .C1(n2783), .C2(n2228), .ZN(n2739) );
  INV_X1 U35060 ( .A(n2783), .ZN(n2711) );
  NOR2_X1 U35070 ( .A1(n4474), .A2(n3222), .ZN(n2713) );
  OAI21_X1 U35080 ( .B1(n4450), .B2(n2827), .A(n2712), .ZN(n2738) );
  INV_X1 U35090 ( .A(n2713), .ZN(n2714) );
  AOI22_X1 U35100 ( .A1(n2739), .A2(n2738), .B1(n3198), .B2(n2714), .ZN(n2761)
         );
  XNOR2_X1 U35110 ( .A(n2760), .B(n2761), .ZN(n2737) );
  OR2_X1 U35120 ( .A1(n2715), .A2(n2792), .ZN(n2716) );
  NOR2_X1 U35130 ( .A1(n2793), .A2(n2716), .ZN(n2723) );
  INV_X1 U35140 ( .A(n2717), .ZN(n2720) );
  INV_X1 U35150 ( .A(n2718), .ZN(n2719) );
  OAI211_X1 U35160 ( .C1(n2720), .C2(n4473), .A(n2725), .B(n2719), .ZN(n2721)
         );
  INV_X1 U35170 ( .A(n2721), .ZN(n2722) );
  INV_X1 U35180 ( .A(n2723), .ZN(n2733) );
  NOR3_X1 U35190 ( .A1(n2733), .A2(n2724), .A3(n3881), .ZN(n2726) );
  INV_X2 U35200 ( .A(n4482), .ZN(n4458) );
  INV_X1 U35210 ( .A(n2727), .ZN(n2728) );
  NAND2_X1 U35220 ( .A1(n2733), .A2(n2728), .ZN(n2784) );
  INV_X1 U35230 ( .A(n2729), .ZN(n2794) );
  NAND2_X1 U35240 ( .A1(n2784), .A2(n2794), .ZN(n3246) );
  AOI22_X1 U35250 ( .A1(n3273), .A2(n4459), .B1(REG3_REG_1__SCAN_IN), .B2(
        n3246), .ZN(n2736) );
  INV_X1 U35260 ( .A(n2730), .ZN(n2732) );
  NAND3_X1 U35270 ( .A1(n2841), .A2(n2732), .A3(n2731), .ZN(n3558) );
  NOR2_X1 U35280 ( .A1(n2733), .A2(n3558), .ZN(n2734) );
  NAND2_X1 U35290 ( .A1(n2734), .A2(n4236), .ZN(n3387) );
  NAND2_X1 U35300 ( .A1(n2734), .A2(n2741), .ZN(n3388) );
  AOI22_X1 U35310 ( .A1(n3399), .A2(n3577), .B1(n3398), .B2(n2331), .ZN(n2735)
         );
  OAI211_X1 U35320 ( .C1(n2737), .C2(n3406), .A(n2736), .B(n2735), .ZN(U3219)
         );
  XOR2_X1 U35330 ( .A(n2739), .B(n2738), .Z(n3245) );
  NOR3_X1 U35340 ( .A1(n3245), .A2(n2741), .A3(n4237), .ZN(n2745) );
  NAND2_X1 U35350 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(
        n3578) );
  INV_X1 U35360 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2740) );
  AND2_X1 U35370 ( .A1(n4237), .A2(n2740), .ZN(n2742) );
  OR2_X1 U35380 ( .A1(n2742), .A2(n2741), .ZN(n4253) );
  NAND2_X1 U35390 ( .A1(n4253), .A2(n2228), .ZN(n2743) );
  OAI211_X1 U35400 ( .C1(n3578), .C2(n3557), .A(U4043), .B(n2743), .ZN(n2744)
         );
  OR2_X1 U35410 ( .A1(n2745), .A2(n2744), .ZN(n3603) );
  INV_X1 U35420 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3630) );
  OAI21_X1 U35430 ( .B1(n2747), .B2(n2218), .A(n2746), .ZN(n3627) );
  XNOR2_X1 U35440 ( .A(n3627), .B(n4243), .ZN(n3631) );
  XOR2_X1 U35450 ( .A(n3630), .B(n3631), .Z(n2754) );
  INV_X1 U35460 ( .A(n4243), .ZN(n3628) );
  AND2_X1 U35470 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3338) );
  AOI21_X1 U35480 ( .B1(n4402), .B2(ADDR_REG_4__SCAN_IN), .A(n3338), .ZN(n2748) );
  OAI21_X1 U35490 ( .B1(n4409), .B2(n3628), .A(n2748), .ZN(n2753) );
  INV_X1 U35500 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4580) );
  AOI211_X1 U35510 ( .C1(n4580), .C2(n2751), .A(n4270), .B(n3606), .ZN(n2752)
         );
  AOI211_X1 U35520 ( .C1(n4345), .C2(n2754), .A(n2753), .B(n2752), .ZN(n2755)
         );
  NAND2_X1 U35530 ( .A1(n3603), .A2(n2755), .ZN(U3244) );
  INV_X1 U35540 ( .A(n2756), .ZN(n2759) );
  INV_X1 U35550 ( .A(n2757), .ZN(n2758) );
  OAI22_X1 U35560 ( .A1(n2761), .A2(n2760), .B1(n2759), .B2(n2758), .ZN(n2769)
         );
  OAI22_X1 U35570 ( .A1(n2815), .A2(n2827), .B1(n3222), .B2(n2762), .ZN(n2763)
         );
  XNOR2_X1 U35580 ( .A(n2763), .B(n3198), .ZN(n2767) );
  OR2_X1 U35590 ( .A1(n2815), .A2(n3226), .ZN(n2765) );
  NAND2_X1 U35600 ( .A1(n3927), .A2(n2841), .ZN(n2764) );
  AND2_X1 U35610 ( .A1(n2765), .A2(n2764), .ZN(n2766) );
  NAND2_X1 U35620 ( .A1(n2767), .A2(n2766), .ZN(n2773) );
  OAI21_X1 U35630 ( .B1(n2767), .B2(n2766), .A(n2773), .ZN(n2768) );
  NOR2_X1 U35640 ( .A1(n2769), .A2(n2768), .ZN(n2775) );
  AOI21_X1 U35650 ( .B1(n2769), .B2(n2768), .A(n2775), .ZN(n2772) );
  AOI22_X1 U35660 ( .A1(n3273), .A2(n3927), .B1(REG3_REG_2__SCAN_IN), .B2(
        n3246), .ZN(n2771) );
  AOI22_X1 U35670 ( .A1(n3398), .A2(n3919), .B1(n3399), .B2(n2323), .ZN(n2770)
         );
  OAI211_X1 U35680 ( .C1(n2772), .C2(n3406), .A(n2771), .B(n2770), .ZN(U3234)
         );
  INV_X1 U35690 ( .A(n2773), .ZN(n2774) );
  AOI22_X1 U35700 ( .A1(n3919), .A2(n3210), .B1(n2841), .B2(n3443), .ZN(n2832)
         );
  NAND2_X1 U35710 ( .A1(n3919), .A2(n2841), .ZN(n2777) );
  NAND2_X1 U35720 ( .A1(n3443), .A2(n2709), .ZN(n2776) );
  NAND2_X1 U35730 ( .A1(n2777), .A2(n2776), .ZN(n2778) );
  XNOR2_X1 U35740 ( .A(n2778), .B(n3223), .ZN(n2834) );
  XOR2_X1 U35750 ( .A(n2832), .B(n2834), .Z(n2779) );
  AOI21_X1 U35760 ( .B1(n2780), .B2(n2779), .A(n3334), .ZN(n2791) );
  AOI22_X1 U35770 ( .A1(n3399), .A2(n2331), .B1(n3398), .B2(n3575), .ZN(n2790)
         );
  NAND4_X1 U35780 ( .A1(n2784), .A2(n2783), .A3(n2782), .A4(n2781), .ZN(n2785)
         );
  INV_X1 U35790 ( .A(n3403), .ZN(n2786) );
  NOR2_X1 U35800 ( .A1(n2786), .A2(REG3_REG_3__SCAN_IN), .ZN(n2787) );
  AOI211_X1 U35810 ( .C1(n3443), .C2(n3273), .A(n2788), .B(n2787), .ZN(n2789)
         );
  OAI211_X1 U3582 ( .C1(n2791), .C2(n3406), .A(n2790), .B(n2789), .ZN(U3215)
         );
  INV_X1 U3583 ( .A(n2792), .ZN(n2796) );
  NAND4_X1 U3584 ( .A1(n2796), .A2(n2795), .A3(n2794), .A4(n2793), .ZN(n2797)
         );
  INV_X1 U3585 ( .A(n2798), .ZN(n3449) );
  NAND2_X1 U3586 ( .A1(n3449), .A2(n3435), .ZN(n3506) );
  XNOR2_X1 U3587 ( .A(n2799), .B(n3506), .ZN(n2802) );
  AOI22_X1 U3588 ( .A1(n3573), .A2(n4447), .B1(n4446), .B2(n2842), .ZN(n2800)
         );
  OAI21_X1 U3589 ( .B1(n2829), .B2(n4449), .A(n2800), .ZN(n2801) );
  AOI21_X1 U3590 ( .B1(n2802), .B2(n4469), .A(n2801), .ZN(n4546) );
  XOR2_X1 U3591 ( .A(n3506), .B(n2803), .Z(n4550) );
  NAND2_X1 U3592 ( .A1(n2804), .A2(n4242), .ZN(n2805) );
  OR2_X1 U3593 ( .A1(n4466), .A2(n4417), .ZN(n2806) );
  INV_X1 U3594 ( .A(n3896), .ZN(n3008) );
  NOR2_X2 U3595 ( .A1(n3844), .A2(n4548), .ZN(n4463) );
  NAND2_X1 U3596 ( .A1(n2849), .A2(n2842), .ZN(n2807) );
  NAND2_X1 U3597 ( .A1(n2867), .A2(n2807), .ZN(n4547) );
  AOI22_X1 U3598 ( .A1(n4466), .A2(REG2_REG_5__SCAN_IN), .B1(n2845), .B2(n4458), .ZN(n2808) );
  OAI21_X1 U3599 ( .B1(n3892), .B2(n4547), .A(n2808), .ZN(n2809) );
  AOI21_X1 U3600 ( .B1(n4550), .B2(n3008), .A(n2809), .ZN(n2810) );
  OAI21_X1 U3601 ( .B1(n4466), .B2(n4546), .A(n2810), .ZN(U3285) );
  INV_X1 U3602 ( .A(n3515), .ZN(n2812) );
  XNOR2_X1 U3603 ( .A(n2811), .B(n2812), .ZN(n4536) );
  INV_X1 U3604 ( .A(n4417), .ZN(n4470) );
  NAND2_X1 U3605 ( .A1(n4536), .A2(n4470), .ZN(n2821) );
  NAND3_X1 U3606 ( .A1(n3922), .A2(n3439), .A3(n2812), .ZN(n2813) );
  NAND2_X1 U3607 ( .A1(n2814), .A2(n2813), .ZN(n2819) );
  OR2_X1 U3608 ( .A1(n2815), .A2(n4449), .ZN(n2817) );
  NAND2_X1 U3609 ( .A1(n3443), .A2(n4446), .ZN(n2816) );
  OAI211_X1 U3610 ( .C1(n2829), .C2(n4472), .A(n2817), .B(n2816), .ZN(n2818)
         );
  AOI21_X1 U3611 ( .B1(n2819), .B2(n4469), .A(n2818), .ZN(n2820) );
  AND2_X1 U3612 ( .A1(n2821), .A2(n2820), .ZN(n4538) );
  AND2_X1 U3613 ( .A1(n4528), .A2(n3443), .ZN(n2822) );
  NOR2_X1 U3614 ( .A1(n2850), .A2(n2822), .ZN(n4535) );
  INV_X1 U3615 ( .A(n4535), .ZN(n2824) );
  AOI22_X1 U3616 ( .A1(n4466), .A2(REG2_REG_3__SCAN_IN), .B1(n4458), .B2(n2334), .ZN(n2823) );
  OAI21_X1 U3617 ( .B1(n3892), .B2(n2824), .A(n2823), .ZN(n2825) );
  AOI21_X1 U3618 ( .B1(n4536), .B2(n4468), .A(n2825), .ZN(n2826) );
  OAI21_X1 U3619 ( .B1(n4538), .B2(n4466), .A(n2826), .ZN(U3287) );
  OAI22_X1 U3620 ( .A1(n2829), .A2(n2827), .B1(n3222), .B2(n3336), .ZN(n2828)
         );
  XNOR2_X1 U3621 ( .A(n2828), .B(n3223), .ZN(n2837) );
  OR2_X1 U3622 ( .A1(n2829), .A2(n3226), .ZN(n2831) );
  NAND2_X1 U3623 ( .A1(n2853), .A2(n2841), .ZN(n2830) );
  NAND2_X1 U3624 ( .A1(n2831), .A2(n2830), .ZN(n2836) );
  XNOR2_X1 U3625 ( .A(n2837), .B(n2836), .ZN(n3332) );
  INV_X1 U3626 ( .A(n2832), .ZN(n2833) );
  NOR2_X1 U3627 ( .A1(n2834), .A2(n2833), .ZN(n3333) );
  NAND2_X1 U3628 ( .A1(n3574), .A2(n2841), .ZN(n2839) );
  NAND2_X1 U3629 ( .A1(n2842), .A2(n2709), .ZN(n2838) );
  NAND2_X1 U3630 ( .A1(n2839), .A2(n2838), .ZN(n2840) );
  XNOR2_X1 U3631 ( .A(n2840), .B(n3198), .ZN(n2874) );
  AOI22_X1 U3632 ( .A1(n3574), .A2(n3210), .B1(n2841), .B2(n2842), .ZN(n2875)
         );
  XNOR2_X1 U3633 ( .A(n2874), .B(n2875), .ZN(n2876) );
  XNOR2_X1 U3634 ( .A(n2877), .B(n2876), .ZN(n2848) );
  AOI22_X1 U3635 ( .A1(n3399), .A2(n3575), .B1(n3398), .B2(n3573), .ZN(n2847)
         );
  INV_X1 U3636 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2843) );
  NOR2_X1 U3637 ( .A1(STATE_REG_SCAN_IN), .A2(n2843), .ZN(n4262) );
  NOR2_X1 U3638 ( .A1(n3401), .A2(n2155), .ZN(n2844) );
  AOI211_X1 U3639 ( .C1(n3403), .C2(n2845), .A(n4262), .B(n2844), .ZN(n2846)
         );
  OAI211_X1 U3640 ( .C1(n2848), .C2(n3406), .A(n2847), .B(n2846), .ZN(U3224)
         );
  OAI211_X1 U3641 ( .C1(n2850), .C2(n3336), .A(n2849), .B(n4569), .ZN(n4540)
         );
  NOR2_X1 U3642 ( .A1(n4540), .A2(n4242), .ZN(n2858) );
  XNOR2_X1 U3643 ( .A(n2851), .B(n3489), .ZN(n2859) );
  XOR2_X1 U3644 ( .A(n3489), .B(n2852), .Z(n2856) );
  AOI22_X1 U3645 ( .A1(n3574), .A2(n4447), .B1(n2853), .B2(n4446), .ZN(n2854)
         );
  OAI21_X1 U3646 ( .B1(n3442), .B2(n4449), .A(n2854), .ZN(n2855) );
  AOI21_X1 U3647 ( .B1(n2856), .B2(n4469), .A(n2855), .ZN(n2857) );
  OAI21_X1 U3648 ( .B1(n4417), .B2(n2859), .A(n2857), .ZN(n4541) );
  AOI211_X1 U3649 ( .C1(n4458), .C2(n3339), .A(n2858), .B(n4541), .ZN(n2861)
         );
  INV_X1 U3650 ( .A(n2859), .ZN(n4544) );
  AOI22_X1 U3651 ( .A1(n4544), .A2(n4468), .B1(REG2_REG_4__SCAN_IN), .B2(n4466), .ZN(n2860) );
  OAI21_X1 U3652 ( .B1(n2861), .B2(n4466), .A(n2860), .ZN(U3286) );
  NAND2_X1 U3653 ( .A1(n3452), .A2(n3448), .ZN(n3488) );
  XNOR2_X1 U3654 ( .A(n2862), .B(n3488), .ZN(n2894) );
  INV_X1 U3655 ( .A(n2894), .ZN(n2873) );
  XNOR2_X1 U3656 ( .A(n2863), .B(n3488), .ZN(n2866) );
  OAI22_X1 U3657 ( .A1(n2951), .A2(n4472), .B1(n3881), .B2(n2887), .ZN(n2864)
         );
  AOI21_X1 U3658 ( .B1(n4411), .B2(n3574), .A(n2864), .ZN(n2865) );
  OAI21_X1 U3659 ( .B1(n2866), .B2(n4453), .A(n2865), .ZN(n2893) );
  NAND2_X1 U3660 ( .A1(n2893), .A2(n4477), .ZN(n2872) );
  AOI21_X1 U3661 ( .B1(n2881), .B2(n2867), .A(n2907), .ZN(n2900) );
  INV_X1 U3662 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2869) );
  OAI22_X1 U3663 ( .A1(n4477), .A2(n2869), .B1(n2868), .B2(n4482), .ZN(n2870)
         );
  AOI21_X1 U3664 ( .B1(n2900), .B2(n4463), .A(n2870), .ZN(n2871) );
  OAI211_X1 U3665 ( .C1(n3896), .C2(n2873), .A(n2872), .B(n2871), .ZN(U3284)
         );
  NAND2_X1 U3666 ( .A1(n3573), .A2(n2841), .ZN(n2879) );
  NAND2_X1 U3667 ( .A1(n2881), .A2(n2709), .ZN(n2878) );
  NAND2_X1 U3668 ( .A1(n2879), .A2(n2878), .ZN(n2880) );
  XNOR2_X1 U3669 ( .A(n2880), .B(n3198), .ZN(n2883) );
  AOI22_X1 U3670 ( .A1(n3573), .A2(n3210), .B1(n2841), .B2(n2881), .ZN(n2882)
         );
  NOR2_X1 U3671 ( .A1(n2883), .A2(n2882), .ZN(n2917) );
  NAND2_X1 U3672 ( .A1(n2883), .A2(n2882), .ZN(n2916) );
  INV_X1 U3673 ( .A(n2916), .ZN(n2884) );
  NOR2_X1 U3674 ( .A1(n2917), .A2(n2884), .ZN(n2885) );
  XNOR2_X1 U3675 ( .A(n2918), .B(n2885), .ZN(n2892) );
  AOI22_X1 U3676 ( .A1(n3399), .A2(n3574), .B1(n3398), .B2(n3572), .ZN(n2891)
         );
  INV_X1 U3677 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2886) );
  NOR2_X1 U3678 ( .A1(STATE_REG_SCAN_IN), .A2(n2886), .ZN(n4274) );
  NOR2_X1 U3679 ( .A1(n3401), .A2(n2887), .ZN(n2888) );
  AOI211_X1 U3680 ( .C1(n3403), .C2(n2889), .A(n4274), .B(n2888), .ZN(n2890)
         );
  OAI211_X1 U3681 ( .C1(n2892), .C2(n3406), .A(n2891), .B(n2890), .ZN(U3236)
         );
  AOI21_X1 U3682 ( .B1(n4554), .B2(n2894), .A(n2893), .ZN(n2902) );
  INV_X1 U3683 ( .A(n4176), .ZN(n2895) );
  AOI22_X1 U3684 ( .A1(n2900), .A2(n2895), .B1(n4587), .B2(REG1_REG_6__SCAN_IN), .ZN(n2896) );
  OAI21_X1 U3685 ( .B1(n2902), .B2(n4587), .A(n2896), .ZN(U3524) );
  INV_X1 U3686 ( .A(n4231), .ZN(n2899) );
  INV_X1 U3687 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2897) );
  NOR2_X1 U3688 ( .A1(n4572), .A2(n2897), .ZN(n2898) );
  AOI21_X1 U3689 ( .B1(n2900), .B2(n2899), .A(n2898), .ZN(n2901) );
  OAI21_X1 U3690 ( .B1(n2902), .B2(n4570), .A(n2901), .ZN(U3479) );
  XNOR2_X1 U3691 ( .A(n2903), .B(n3491), .ZN(n2906) );
  OAI22_X1 U3692 ( .A1(n2928), .A2(n4472), .B1(n3881), .B2(n3253), .ZN(n2904)
         );
  AOI21_X1 U3693 ( .B1(n4411), .B2(n3573), .A(n2904), .ZN(n2905) );
  OAI21_X1 U3694 ( .B1(n2906), .B2(n4453), .A(n2905), .ZN(n4552) );
  INV_X1 U3695 ( .A(n4552), .ZN(n2915) );
  INV_X1 U3696 ( .A(n2907), .ZN(n2908) );
  AOI211_X1 U3697 ( .C1(n2920), .C2(n2908), .A(n4548), .B(n2957), .ZN(n4553)
         );
  INV_X1 U3698 ( .A(n3844), .ZN(n2911) );
  INV_X1 U3699 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3998) );
  INV_X1 U3700 ( .A(n3255), .ZN(n2909) );
  OAI22_X1 U3701 ( .A1(n4477), .A2(n3998), .B1(n2909), .B2(n4482), .ZN(n2910)
         );
  AOI21_X1 U3702 ( .B1(n4553), .B2(n2911), .A(n2910), .ZN(n2914) );
  XOR2_X1 U3703 ( .A(n2912), .B(n3491), .Z(n4555) );
  NAND2_X1 U3704 ( .A1(n4555), .A2(n3008), .ZN(n2913) );
  OAI211_X1 U3705 ( .C1(n2915), .C2(n4466), .A(n2914), .B(n2913), .ZN(U3283)
         );
  INV_X1 U3706 ( .A(n3250), .ZN(n2924) );
  OAI22_X1 U3707 ( .A1(n2951), .A2(n3225), .B1(n3222), .B2(n3253), .ZN(n2919)
         );
  XNOR2_X1 U3708 ( .A(n2919), .B(n3223), .ZN(n2925) );
  OR2_X1 U3709 ( .A1(n2951), .A2(n3226), .ZN(n2922) );
  NAND2_X1 U3710 ( .A1(n2920), .A2(n2841), .ZN(n2921) );
  NAND2_X1 U3711 ( .A1(n2922), .A2(n2921), .ZN(n2926) );
  XNOR2_X1 U3712 ( .A(n2925), .B(n2926), .ZN(n3249) );
  INV_X1 U3713 ( .A(n3249), .ZN(n2923) );
  NAND2_X1 U3714 ( .A1(n2924), .A2(n2923), .ZN(n3251) );
  NAND2_X1 U3715 ( .A1(n2925), .A2(n2926), .ZN(n2927) );
  OAI22_X1 U3716 ( .A1(n2928), .A2(n3225), .B1(n3222), .B2(n2956), .ZN(n2929)
         );
  XNOR2_X1 U3717 ( .A(n2929), .B(n3223), .ZN(n2965) );
  AOI22_X1 U3718 ( .A1(n3571), .A2(n3210), .B1(n2841), .B2(n2949), .ZN(n2967)
         );
  XNOR2_X1 U3719 ( .A(n2965), .B(n2967), .ZN(n2930) );
  XNOR2_X1 U3720 ( .A(n2968), .B(n2930), .ZN(n2934) );
  OAI22_X1 U3721 ( .A1(n2951), .A2(n3387), .B1(n3388), .B2(n2969), .ZN(n2932)
         );
  NAND2_X1 U3722 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4293) );
  OAI21_X1 U3723 ( .B1(n3401), .B2(n2956), .A(n4293), .ZN(n2931) );
  AOI211_X1 U3724 ( .C1(n4435), .C2(n3403), .A(n2932), .B(n2931), .ZN(n2933)
         );
  OAI21_X1 U3725 ( .B1(n2934), .B2(n3406), .A(n2933), .ZN(U3218) );
  INV_X1 U3726 ( .A(n2935), .ZN(n3464) );
  NAND2_X1 U3727 ( .A1(n3464), .A2(n3459), .ZN(n3507) );
  XOR2_X1 U3728 ( .A(n3507), .B(n2936), .Z(n4558) );
  XOR2_X1 U3729 ( .A(n3507), .B(n2937), .Z(n2940) );
  OAI22_X1 U3730 ( .A1(n3046), .A2(n4472), .B1(n3881), .B2(n3347), .ZN(n2938)
         );
  AOI21_X1 U3731 ( .B1(n4411), .B2(n3571), .A(n2938), .ZN(n2939) );
  OAI21_X1 U3732 ( .B1(n2940), .B2(n4453), .A(n2939), .ZN(n4560) );
  NAND2_X1 U3733 ( .A1(n4560), .A2(n4477), .ZN(n2946) );
  AOI21_X1 U3734 ( .B1(n2941), .B2(n2955), .A(n2099), .ZN(n4561) );
  INV_X1 U3735 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2943) );
  INV_X1 U3736 ( .A(n3349), .ZN(n2942) );
  OAI22_X1 U3737 ( .A1(n4477), .A2(n2943), .B1(n2942), .B2(n4482), .ZN(n2944)
         );
  AOI21_X1 U3738 ( .B1(n4561), .B2(n4463), .A(n2944), .ZN(n2945) );
  OAI211_X1 U3739 ( .C1(n3896), .C2(n4558), .A(n2946), .B(n2945), .ZN(U3281)
         );
  NAND2_X1 U3740 ( .A1(n3458), .A2(n3455), .ZN(n3487) );
  XNOR2_X1 U3741 ( .A(n2947), .B(n3487), .ZN(n4436) );
  XNOR2_X1 U3742 ( .A(n2948), .B(n3487), .ZN(n2954) );
  AOI22_X1 U3743 ( .A1(n3570), .A2(n4447), .B1(n4446), .B2(n2949), .ZN(n2950)
         );
  OAI21_X1 U3744 ( .B1(n2951), .B2(n4449), .A(n2950), .ZN(n2953) );
  NOR2_X1 U3745 ( .A1(n4436), .A2(n4417), .ZN(n2952) );
  AOI211_X1 U3746 ( .C1(n4469), .C2(n2954), .A(n2953), .B(n2952), .ZN(n4442)
         );
  OAI21_X1 U3747 ( .B1(n4563), .B2(n4436), .A(n4442), .ZN(n2963) );
  OAI21_X1 U3748 ( .B1(n2957), .B2(n2956), .A(n2955), .ZN(n4437) );
  INV_X1 U3749 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2958) );
  OAI22_X1 U3750 ( .A1(n4437), .A2(n4231), .B1(n4572), .B2(n2958), .ZN(n2959)
         );
  AOI21_X1 U3751 ( .B1(n2963), .B2(n4572), .A(n2959), .ZN(n2960) );
  INV_X1 U3752 ( .A(n2960), .ZN(U3483) );
  INV_X1 U3753 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2961) );
  OAI22_X1 U3754 ( .A1(n4437), .A2(n4176), .B1(n4590), .B2(n2961), .ZN(n2962)
         );
  AOI21_X1 U3755 ( .B1(n2963), .B2(n4590), .A(n2962), .ZN(n2964) );
  INV_X1 U3756 ( .A(n2964), .ZN(U3526) );
  INV_X1 U3757 ( .A(n2967), .ZN(n2966) );
  OAI22_X1 U3758 ( .A1(n2969), .A2(n3226), .B1(n3225), .B2(n3347), .ZN(n2972)
         );
  OAI22_X1 U3759 ( .A1(n2969), .A2(n3225), .B1(n3222), .B2(n3347), .ZN(n2970)
         );
  XNOR2_X1 U3760 ( .A(n2970), .B(n3223), .ZN(n2971) );
  XOR2_X1 U3761 ( .A(n2972), .B(n2971), .Z(n3343) );
  INV_X1 U3762 ( .A(n2971), .ZN(n2974) );
  INV_X1 U3763 ( .A(n2972), .ZN(n2973) );
  NAND2_X1 U3764 ( .A1(n2974), .A2(n2973), .ZN(n2980) );
  NAND2_X1 U3765 ( .A1(n4412), .A2(n2841), .ZN(n2976) );
  NAND2_X1 U3766 ( .A1(n3054), .A2(n2709), .ZN(n2975) );
  NAND2_X1 U3767 ( .A1(n2976), .A2(n2975), .ZN(n2977) );
  XNOR2_X1 U3768 ( .A(n2977), .B(n3223), .ZN(n3010) );
  AOI22_X1 U3769 ( .A1(n4412), .A2(n3210), .B1(n2841), .B2(n3054), .ZN(n3011)
         );
  XNOR2_X1 U3770 ( .A(n3010), .B(n3011), .ZN(n2979) );
  NAND2_X1 U3771 ( .A1(n3014), .A2(n3344), .ZN(n2986) );
  AOI21_X1 U3772 ( .B1(n2978), .B2(n2980), .A(n2979), .ZN(n2985) );
  AOI22_X1 U3773 ( .A1(n3399), .A2(n3570), .B1(n3398), .B2(n3569), .ZN(n2984)
         );
  NOR2_X1 U3774 ( .A1(STATE_REG_SCAN_IN), .A2(n2981), .ZN(n4321) );
  NOR2_X1 U3775 ( .A1(n3401), .A2(n2098), .ZN(n2982) );
  AOI211_X1 U3776 ( .C1(n3403), .C2(n4428), .A(n4321), .B(n2982), .ZN(n2983)
         );
  OAI211_X1 U3777 ( .C1(n2986), .C2(n2985), .A(n2984), .B(n2983), .ZN(U3214)
         );
  XNOR2_X1 U3778 ( .A(n4414), .B(n3023), .ZN(n3519) );
  XNOR2_X1 U3779 ( .A(n2987), .B(n3519), .ZN(n2990) );
  OAI22_X1 U3780 ( .A1(n3902), .A2(n4472), .B1(n3881), .B2(n3027), .ZN(n2988)
         );
  AOI21_X1 U3781 ( .B1(n4411), .B2(n3569), .A(n2988), .ZN(n2989) );
  OAI21_X1 U3782 ( .B1(n2990), .B2(n4453), .A(n2989), .ZN(n3033) );
  INV_X1 U3783 ( .A(n3033), .ZN(n2995) );
  XOR2_X1 U3784 ( .A(n3519), .B(n2991), .Z(n3034) );
  OAI21_X1 U3785 ( .B1(n4422), .B2(n3027), .A(n3004), .ZN(n3039) );
  AOI22_X1 U3786 ( .A1(n4466), .A2(REG2_REG_12__SCAN_IN), .B1(n3030), .B2(
        n4458), .ZN(n2992) );
  OAI21_X1 U3787 ( .B1(n3039), .B2(n3892), .A(n2992), .ZN(n2993) );
  AOI21_X1 U3788 ( .B1(n3034), .B2(n3008), .A(n2993), .ZN(n2994) );
  OAI21_X1 U3789 ( .B1(n4466), .B2(n2995), .A(n2994), .ZN(U3278) );
  NAND2_X1 U3790 ( .A1(n2997), .A2(n2996), .ZN(n2999) );
  NAND2_X1 U3791 ( .A1(n3432), .A2(n2998), .ZN(n3483) );
  XNOR2_X1 U3792 ( .A(n2999), .B(n3483), .ZN(n3002) );
  AOI22_X1 U3793 ( .A1(n3566), .A2(n4447), .B1(n4446), .B2(n3070), .ZN(n3000)
         );
  OAI21_X1 U3794 ( .B1(n4414), .B2(n4449), .A(n3000), .ZN(n3001) );
  AOI21_X1 U3795 ( .B1(n3002), .B2(n4469), .A(n3001), .ZN(n4183) );
  XNOR2_X1 U3796 ( .A(n3003), .B(n3483), .ZN(n4182) );
  NAND2_X1 U3797 ( .A1(n3004), .A2(n3070), .ZN(n3005) );
  NAND2_X1 U3798 ( .A1(n3911), .A2(n3005), .ZN(n4185) );
  AOI22_X1 U3799 ( .A1(n4466), .A2(REG2_REG_13__SCAN_IN), .B1(n3100), .B2(
        n4458), .ZN(n3006) );
  OAI21_X1 U3800 ( .B1(n4185), .B2(n3892), .A(n3006), .ZN(n3007) );
  AOI21_X1 U3801 ( .B1(n4182), .B2(n3008), .A(n3007), .ZN(n3009) );
  OAI21_X1 U3802 ( .B1(n4466), .B2(n4183), .A(n3009), .ZN(U3277) );
  INV_X1 U3803 ( .A(n3010), .ZN(n3012) );
  OR2_X1 U3804 ( .A1(n3012), .A2(n3011), .ZN(n3013) );
  NAND2_X1 U3805 ( .A1(n3014), .A2(n3013), .ZN(n3041) );
  OAI22_X1 U3806 ( .A1(n3056), .A2(n3225), .B1(n3222), .B2(n3048), .ZN(n3015)
         );
  XNOR2_X1 U3807 ( .A(n3015), .B(n3198), .ZN(n3018) );
  OR2_X1 U3808 ( .A1(n3056), .A2(n3226), .ZN(n3017) );
  NAND2_X1 U3809 ( .A1(n4424), .A2(n2841), .ZN(n3016) );
  NAND2_X1 U3810 ( .A1(n3018), .A2(n3019), .ZN(n3042) );
  INV_X1 U3811 ( .A(n3018), .ZN(n3021) );
  INV_X1 U3812 ( .A(n3019), .ZN(n3020) );
  NAND2_X1 U3813 ( .A1(n3021), .A2(n3020), .ZN(n3044) );
  OAI22_X1 U3814 ( .A1(n4414), .A2(n3225), .B1(n3222), .B2(n3027), .ZN(n3022)
         );
  XNOR2_X1 U3815 ( .A(n3022), .B(n3223), .ZN(n3088) );
  OR2_X1 U3816 ( .A1(n4414), .A2(n3226), .ZN(n3025) );
  NAND2_X1 U3817 ( .A1(n3023), .A2(n2841), .ZN(n3024) );
  NAND2_X1 U3818 ( .A1(n3025), .A2(n3024), .ZN(n3087) );
  INV_X1 U3819 ( .A(n3087), .ZN(n3073) );
  XNOR2_X1 U3820 ( .A(n3088), .B(n3073), .ZN(n3026) );
  XNOR2_X1 U3821 ( .A(n3079), .B(n3026), .ZN(n3032) );
  OAI22_X1 U3822 ( .A1(n3902), .A2(n3388), .B1(n3387), .B2(n3056), .ZN(n3029)
         );
  NAND2_X1 U3823 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4337) );
  OAI21_X1 U3824 ( .B1(n3401), .B2(n3027), .A(n4337), .ZN(n3028) );
  AOI211_X1 U3825 ( .C1(n3030), .C2(n3403), .A(n3029), .B(n3028), .ZN(n3031)
         );
  OAI21_X1 U3826 ( .B1(n3032), .B2(n3406), .A(n3031), .ZN(U3221) );
  INV_X1 U3827 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3035) );
  AOI21_X1 U3828 ( .B1(n3034), .B2(n4554), .A(n3033), .ZN(n3037) );
  MUX2_X1 U3829 ( .A(n3035), .B(n3037), .S(n4572), .Z(n3036) );
  OAI21_X1 U3830 ( .B1(n3039), .B2(n4231), .A(n3036), .ZN(U3491) );
  INV_X1 U3831 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4037) );
  MUX2_X1 U3832 ( .A(n4037), .B(n3037), .S(n4590), .Z(n3038) );
  OAI21_X1 U3833 ( .B1(n3039), .B2(n4176), .A(n3038), .ZN(U3530) );
  INV_X1 U3834 ( .A(n3040), .ZN(n3045) );
  AOI21_X1 U3835 ( .B1(n3044), .B2(n3042), .A(n3041), .ZN(n3043) );
  AOI211_X1 U3836 ( .C1(n3045), .C2(n3044), .A(n3406), .B(n3043), .ZN(n3051)
         );
  OAI22_X1 U3837 ( .A1(n4414), .A2(n3388), .B1(n3387), .B2(n3046), .ZN(n3050)
         );
  NAND2_X1 U3838 ( .A1(REG3_REG_11__SCAN_IN), .A2(U3149), .ZN(n4326) );
  NAND2_X1 U3839 ( .A1(n3403), .A2(n4421), .ZN(n3047) );
  OAI211_X1 U3840 ( .C1(n3401), .C2(n3048), .A(n4326), .B(n3047), .ZN(n3049)
         );
  OR3_X1 U3841 ( .A1(n3051), .A2(n3050), .A3(n3049), .ZN(U3233) );
  OAI21_X1 U3842 ( .B1(n2099), .B2(n2098), .A(n4423), .ZN(n4429) );
  INV_X1 U3843 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3062) );
  INV_X1 U3844 ( .A(n4563), .ZN(n4543) );
  NAND2_X1 U3845 ( .A1(n3423), .A2(n3424), .ZN(n3485) );
  XNOR2_X1 U3846 ( .A(n3052), .B(n3485), .ZN(n3057) );
  INV_X1 U3847 ( .A(n3057), .ZN(n4431) );
  XOR2_X1 U3848 ( .A(n3485), .B(n3053), .Z(n3060) );
  AOI22_X1 U3849 ( .A1(n3570), .A2(n4411), .B1(n3054), .B2(n4446), .ZN(n3055)
         );
  OAI21_X1 U3850 ( .B1(n3056), .B2(n4472), .A(n3055), .ZN(n3059) );
  NOR2_X1 U3851 ( .A1(n3057), .A2(n4417), .ZN(n3058) );
  AOI211_X1 U3852 ( .C1(n3060), .C2(n4469), .A(n3059), .B(n3058), .ZN(n4434)
         );
  INV_X1 U3853 ( .A(n4434), .ZN(n3061) );
  AOI21_X1 U3854 ( .B1(n4543), .B2(n4431), .A(n3061), .ZN(n3064) );
  MUX2_X1 U3855 ( .A(n3062), .B(n3064), .S(n4590), .Z(n3063) );
  OAI21_X1 U3856 ( .B1(n4429), .B2(n4176), .A(n3063), .ZN(U3528) );
  INV_X1 U3857 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3065) );
  MUX2_X1 U3858 ( .A(n3065), .B(n3064), .S(n4572), .Z(n3066) );
  OAI21_X1 U3859 ( .B1(n4429), .B2(n4231), .A(n3066), .ZN(U3487) );
  INV_X1 U3860 ( .A(n3088), .ZN(n3090) );
  NAND2_X1 U3861 ( .A1(n3567), .A2(n2841), .ZN(n3068) );
  NAND2_X1 U3862 ( .A1(n3070), .A2(n2709), .ZN(n3067) );
  NAND2_X1 U3863 ( .A1(n3068), .A2(n3067), .ZN(n3069) );
  XNOR2_X1 U3864 ( .A(n3069), .B(n3198), .ZN(n3075) );
  INV_X1 U3865 ( .A(n3075), .ZN(n3072) );
  AOI22_X1 U3866 ( .A1(n3567), .A2(n3210), .B1(n2841), .B2(n3070), .ZN(n3074)
         );
  INV_X1 U3867 ( .A(n3074), .ZN(n3071) );
  NAND2_X1 U3868 ( .A1(n3072), .A2(n3071), .ZN(n3092) );
  OAI21_X1 U3869 ( .B1(n3090), .B2(n3073), .A(n3092), .ZN(n3078) );
  NOR2_X1 U3870 ( .A1(n3088), .A2(n3087), .ZN(n3076) );
  AND2_X1 U3871 ( .A1(n3075), .A2(n3074), .ZN(n3093) );
  AOI21_X1 U3872 ( .B1(n3076), .B2(n3092), .A(n3093), .ZN(n3077) );
  OAI22_X1 U3873 ( .A1(n3880), .A2(n3226), .B1(n3225), .B2(n3082), .ZN(n3122)
         );
  OAI22_X1 U3874 ( .A1(n3880), .A2(n3225), .B1(n3222), .B2(n3082), .ZN(n3080)
         );
  XOR2_X1 U3875 ( .A(n3223), .B(n3080), .Z(n3125) );
  XOR2_X1 U3876 ( .A(n3122), .B(n3125), .Z(n3081) );
  XNOR2_X1 U3877 ( .A(n3124), .B(n3081), .ZN(n3086) );
  OAI22_X1 U3878 ( .A1(n3902), .A2(n3387), .B1(n3388), .B2(n3309), .ZN(n3084)
         );
  NAND2_X1 U3879 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4360) );
  OAI21_X1 U3880 ( .B1(n3401), .B2(n3082), .A(n4360), .ZN(n3083) );
  AOI211_X1 U3881 ( .C1(n3908), .C2(n3403), .A(n3084), .B(n3083), .ZN(n3085)
         );
  OAI21_X1 U3882 ( .B1(n3086), .B2(n3406), .A(n3085), .ZN(U3212) );
  INV_X1 U3883 ( .A(n3079), .ZN(n3091) );
  OAI21_X1 U3884 ( .B1(n3079), .B2(n3088), .A(n3087), .ZN(n3089) );
  OAI21_X1 U3885 ( .B1(n3091), .B2(n3090), .A(n3089), .ZN(n3096) );
  INV_X1 U3886 ( .A(n3092), .ZN(n3094) );
  NOR2_X1 U3887 ( .A1(n3094), .A2(n3093), .ZN(n3095) );
  XNOR2_X1 U3888 ( .A(n3096), .B(n3095), .ZN(n3103) );
  AOI22_X1 U3889 ( .A1(n3399), .A2(n3568), .B1(n3398), .B2(n3566), .ZN(n3102)
         );
  NOR2_X1 U3890 ( .A1(STATE_REG_SCAN_IN), .A2(n3097), .ZN(n4350) );
  NOR2_X1 U3891 ( .A1(n3401), .A2(n3098), .ZN(n3099) );
  AOI211_X1 U3892 ( .C1(n3403), .C2(n3100), .A(n4350), .B(n3099), .ZN(n3101)
         );
  OAI211_X1 U3893 ( .C1(n3103), .C2(n3406), .A(n3102), .B(n3101), .ZN(U3231)
         );
  INV_X1 U3894 ( .A(D_REG_0__SCAN_IN), .ZN(n3106) );
  NOR2_X1 U3895 ( .A1(n2646), .A2(n4490), .ZN(n3105) );
  AOI22_X1 U3896 ( .A1(n4489), .A2(n3106), .B1(n3105), .B2(n3104), .ZN(U3458)
         );
  NAND2_X1 U3897 ( .A1(n2052), .A2(DATAI_29_), .ZN(n3410) );
  XNOR2_X1 U3898 ( .A(n3411), .B(n3410), .ZN(n3496) );
  XNOR2_X1 U3899 ( .A(n3109), .B(n3496), .ZN(n3947) );
  INV_X1 U3900 ( .A(n3410), .ZN(n3115) );
  AOI22_X1 U3901 ( .A1(n3945), .A2(n4463), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4466), .ZN(n3121) );
  NAND2_X1 U3902 ( .A1(n3112), .A2(n3111), .ZN(n3542) );
  OAI21_X1 U3903 ( .B1(n3668), .B2(n3542), .A(n3408), .ZN(n3113) );
  XNOR2_X1 U3904 ( .A(n3113), .B(n3496), .ZN(n3114) );
  NAND2_X1 U3905 ( .A1(n3114), .A2(n4469), .ZN(n3117) );
  AOI21_X1 U3906 ( .B1(n4237), .B2(B_REG_SCAN_IN), .A(n4472), .ZN(n3932) );
  AOI22_X1 U3907 ( .A1(n3478), .A2(n3932), .B1(n4446), .B2(n3115), .ZN(n3116)
         );
  OAI211_X1 U3908 ( .C1(n3671), .C2(n4449), .A(n3117), .B(n3116), .ZN(n3944)
         );
  NOR2_X1 U3909 ( .A1(n3118), .A2(n4482), .ZN(n3119) );
  OAI21_X1 U3910 ( .B1(n3944), .B2(n3119), .A(n4477), .ZN(n3120) );
  OAI211_X1 U3911 ( .C1(n3947), .C2(n3896), .A(n3121), .B(n3120), .ZN(U3354)
         );
  NAND2_X1 U3912 ( .A1(n3123), .A2(n3122), .ZN(n3129) );
  INV_X1 U3913 ( .A(n3124), .ZN(n3127) );
  INV_X1 U3914 ( .A(n3125), .ZN(n3126) );
  NAND2_X1 U3915 ( .A1(n3127), .A2(n3126), .ZN(n3128) );
  NAND2_X1 U3916 ( .A1(n3129), .A2(n3128), .ZN(n3132) );
  OAI22_X1 U3917 ( .A1(n3309), .A2(n3225), .B1(n3222), .B2(n3889), .ZN(n3130)
         );
  XNOR2_X1 U3918 ( .A(n3130), .B(n3223), .ZN(n3133) );
  OAI22_X1 U3919 ( .A1(n3882), .A2(n3226), .B1(n3225), .B2(n3870), .ZN(n3141)
         );
  OAI22_X1 U3920 ( .A1(n3882), .A2(n3225), .B1(n3222), .B2(n3870), .ZN(n3131)
         );
  XNOR2_X1 U3921 ( .A(n3131), .B(n3223), .ZN(n3142) );
  XOR2_X1 U3922 ( .A(n3141), .B(n3142), .Z(n3308) );
  INV_X1 U3923 ( .A(n3132), .ZN(n3135) );
  NAND2_X1 U3924 ( .A1(n3135), .A2(n3134), .ZN(n3305) );
  NAND2_X1 U3925 ( .A1(n3900), .A2(n3210), .ZN(n3138) );
  NAND2_X1 U3926 ( .A1(n3136), .A2(n2841), .ZN(n3137) );
  NAND2_X1 U3927 ( .A1(n3138), .A2(n3137), .ZN(n3397) );
  NAND2_X1 U3928 ( .A1(n3305), .A2(n3397), .ZN(n3139) );
  NAND2_X1 U3929 ( .A1(n3140), .A2(n3139), .ZN(n3144) );
  OAI22_X1 U3930 ( .A1(n3865), .A2(n3225), .B1(n3222), .B2(n3857), .ZN(n3145)
         );
  XNOR2_X1 U3931 ( .A(n3145), .B(n3223), .ZN(n3316) );
  OR2_X1 U3932 ( .A1(n3865), .A2(n3226), .ZN(n3148) );
  NAND2_X1 U3933 ( .A1(n3146), .A2(n2841), .ZN(n3147) );
  NAND2_X1 U3934 ( .A1(n3148), .A2(n3147), .ZN(n3315) );
  NOR2_X1 U3935 ( .A1(n3316), .A2(n3315), .ZN(n3150) );
  NAND2_X1 U3936 ( .A1(n3316), .A2(n3315), .ZN(n3149) );
  OAI22_X1 U3937 ( .A1(n3851), .A2(n3225), .B1(n3222), .B2(n3841), .ZN(n3151)
         );
  XNOR2_X1 U3938 ( .A(n3151), .B(n3198), .ZN(n3155) );
  OR2_X1 U3939 ( .A1(n3851), .A2(n3226), .ZN(n3153) );
  NAND2_X1 U3940 ( .A1(n3834), .A2(n2841), .ZN(n3152) );
  NOR2_X1 U3941 ( .A1(n3155), .A2(n3154), .ZN(n3375) );
  NAND2_X1 U3942 ( .A1(n3155), .A2(n3154), .ZN(n3373) );
  OAI22_X1 U3943 ( .A1(n3833), .A2(n3226), .B1(n3225), .B2(n3823), .ZN(n3157)
         );
  OAI22_X1 U3944 ( .A1(n3833), .A2(n3225), .B1(n3222), .B2(n3823), .ZN(n3156)
         );
  XNOR2_X1 U3945 ( .A(n3156), .B(n3223), .ZN(n3158) );
  XOR2_X1 U3946 ( .A(n3157), .B(n3158), .Z(n3279) );
  NAND2_X1 U3947 ( .A1(n3818), .A2(n2841), .ZN(n3161) );
  NAND2_X1 U3948 ( .A1(n3163), .A2(n2709), .ZN(n3160) );
  NAND2_X1 U3949 ( .A1(n3161), .A2(n3160), .ZN(n3162) );
  XNOR2_X1 U3950 ( .A(n3162), .B(n3223), .ZN(n3166) );
  NAND2_X1 U3951 ( .A1(n3818), .A2(n3210), .ZN(n3165) );
  NAND2_X1 U3952 ( .A1(n3163), .A2(n2841), .ZN(n3164) );
  NAND2_X1 U3953 ( .A1(n3165), .A2(n3164), .ZN(n3167) );
  NAND2_X1 U3954 ( .A1(n3166), .A2(n3167), .ZN(n3355) );
  INV_X1 U3955 ( .A(n3166), .ZN(n3169) );
  INV_X1 U3956 ( .A(n3167), .ZN(n3168) );
  NAND2_X1 U3957 ( .A1(n3169), .A2(n3168), .ZN(n3357) );
  OAI22_X1 U3958 ( .A1(n3793), .A2(n3225), .B1(n3222), .B2(n3780), .ZN(n3170)
         );
  XNOR2_X1 U3959 ( .A(n3170), .B(n3223), .ZN(n3285) );
  OR2_X1 U3960 ( .A1(n3793), .A2(n3226), .ZN(n3173) );
  NAND2_X1 U3961 ( .A1(n3171), .A2(n2841), .ZN(n3172) );
  NAND2_X1 U3962 ( .A1(n3173), .A2(n3172), .ZN(n3284) );
  NOR2_X1 U3963 ( .A1(n3285), .A2(n3284), .ZN(n3174) );
  OAI22_X1 U3964 ( .A1(n3775), .A2(n3225), .B1(n3222), .B2(n3368), .ZN(n3175)
         );
  XNOR2_X1 U3965 ( .A(n3175), .B(n3223), .ZN(n3177) );
  OAI22_X1 U3966 ( .A1(n3775), .A2(n3226), .B1(n3225), .B2(n3368), .ZN(n3176)
         );
  XNOR2_X1 U3967 ( .A(n3177), .B(n3176), .ZN(n3366) );
  NOR2_X1 U3968 ( .A1(n3177), .A2(n3176), .ZN(n3269) );
  NAND2_X1 U3969 ( .A1(n3761), .A2(n2841), .ZN(n3179) );
  NAND2_X1 U3970 ( .A1(n3272), .A2(n2709), .ZN(n3178) );
  NAND2_X1 U3971 ( .A1(n3179), .A2(n3178), .ZN(n3180) );
  XNOR2_X1 U3972 ( .A(n3180), .B(n3198), .ZN(n3183) );
  AND2_X1 U3973 ( .A1(n2841), .A2(n3272), .ZN(n3181) );
  AOI21_X1 U3974 ( .B1(n3761), .B2(n3210), .A(n3181), .ZN(n3184) );
  XNOR2_X1 U3975 ( .A(n3183), .B(n3184), .ZN(n3268) );
  NOR2_X1 U3976 ( .A1(n3269), .A2(n3268), .ZN(n3182) );
  INV_X1 U3977 ( .A(n3183), .ZN(n3186) );
  INV_X1 U3978 ( .A(n3184), .ZN(n3185) );
  NAND2_X1 U3979 ( .A1(n3186), .A2(n3185), .ZN(n3191) );
  AND2_X1 U3980 ( .A1(n2841), .A2(n3187), .ZN(n3188) );
  AOI21_X1 U3981 ( .B1(n3745), .B2(n3210), .A(n3188), .ZN(n3192) );
  OAI22_X1 U3982 ( .A1(n3707), .A2(n3225), .B1(n3222), .B2(n3728), .ZN(n3190)
         );
  XNOR2_X1 U3983 ( .A(n3190), .B(n3223), .ZN(n3325) );
  NAND2_X1 U3984 ( .A1(n3323), .A2(n3325), .ZN(n3195) );
  INV_X1 U3985 ( .A(n3192), .ZN(n3193) );
  NAND2_X1 U3986 ( .A1(n3194), .A2(n3193), .ZN(n3322) );
  NAND2_X1 U3987 ( .A1(n3195), .A2(n3322), .ZN(n3295) );
  NAND2_X1 U3988 ( .A1(n3724), .A2(n2841), .ZN(n3197) );
  NAND2_X1 U3989 ( .A1(n3200), .A2(n2709), .ZN(n3196) );
  NAND2_X1 U3990 ( .A1(n3197), .A2(n3196), .ZN(n3199) );
  XNOR2_X1 U3991 ( .A(n3199), .B(n3198), .ZN(n3202) );
  AND2_X1 U3992 ( .A1(n2841), .A2(n3200), .ZN(n3201) );
  AOI21_X1 U3993 ( .B1(n3724), .B2(n3210), .A(n3201), .ZN(n3203) );
  NAND2_X1 U3994 ( .A1(n3202), .A2(n3203), .ZN(n3293) );
  NAND2_X1 U3995 ( .A1(n3295), .A2(n3293), .ZN(n3206) );
  INV_X1 U3996 ( .A(n3202), .ZN(n3205) );
  INV_X1 U3997 ( .A(n3203), .ZN(n3204) );
  NAND2_X1 U3998 ( .A1(n3205), .A2(n3204), .ZN(n3294) );
  NAND2_X1 U3999 ( .A1(n3206), .A2(n3294), .ZN(n3386) );
  NAND2_X1 U4000 ( .A1(n3709), .A2(n2841), .ZN(n3208) );
  NAND2_X1 U4001 ( .A1(n3685), .A2(n2709), .ZN(n3207) );
  NAND2_X1 U4002 ( .A1(n3208), .A2(n3207), .ZN(n3209) );
  XNOR2_X1 U4003 ( .A(n3209), .B(n3223), .ZN(n3213) );
  NAND2_X1 U4004 ( .A1(n3709), .A2(n3210), .ZN(n3212) );
  NAND2_X1 U4005 ( .A1(n3685), .A2(n2841), .ZN(n3211) );
  NAND2_X1 U4006 ( .A1(n3212), .A2(n3211), .ZN(n3214) );
  AND2_X1 U4007 ( .A1(n3213), .A2(n3214), .ZN(n3384) );
  INV_X1 U4008 ( .A(n3213), .ZN(n3216) );
  INV_X1 U4009 ( .A(n3214), .ZN(n3215) );
  NAND2_X1 U4010 ( .A1(n3216), .A2(n3215), .ZN(n3383) );
  OAI22_X1 U4011 ( .A1(n3389), .A2(n3225), .B1(n3676), .B2(n3222), .ZN(n3217)
         );
  XNOR2_X1 U4012 ( .A(n3217), .B(n3223), .ZN(n3219) );
  OAI22_X1 U4013 ( .A1(n3389), .A2(n3226), .B1(n3676), .B2(n3225), .ZN(n3218)
         );
  XNOR2_X1 U4014 ( .A(n3219), .B(n3218), .ZN(n3260) );
  INV_X1 U4015 ( .A(n3218), .ZN(n3221) );
  INV_X1 U4016 ( .A(n3219), .ZN(n3220) );
  OAI22_X1 U4017 ( .A1(n3671), .A2(n3225), .B1(n3222), .B2(n3231), .ZN(n3224)
         );
  XNOR2_X1 U4018 ( .A(n3224), .B(n3223), .ZN(n3228) );
  OAI22_X1 U4019 ( .A1(n3671), .A2(n3226), .B1(n3225), .B2(n3231), .ZN(n3227)
         );
  XNOR2_X1 U4020 ( .A(n3228), .B(n3227), .ZN(n3229) );
  OAI22_X1 U4021 ( .A1(n3401), .A2(n3231), .B1(STATE_REG_SCAN_IN), .B2(n3230), 
        .ZN(n3234) );
  INV_X1 U4022 ( .A(n3411), .ZN(n3232) );
  OAI22_X1 U4023 ( .A1(n3232), .A2(n3388), .B1(n3389), .B2(n3387), .ZN(n3233)
         );
  AOI211_X1 U4024 ( .C1(n3238), .C2(n3403), .A(n3234), .B(n3233), .ZN(n3235)
         );
  NAND2_X1 U4025 ( .A1(n3236), .A2(n3235), .ZN(U3217) );
  INV_X1 U4026 ( .A(n3237), .ZN(n3242) );
  AOI22_X1 U4027 ( .A1(n3238), .A2(n4458), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4466), .ZN(n3239) );
  OAI21_X1 U4028 ( .B1(n3240), .B2(n3892), .A(n3239), .ZN(n3241) );
  AOI21_X1 U4029 ( .B1(n3242), .B2(n4477), .A(n3241), .ZN(n3243) );
  OAI21_X1 U4030 ( .B1(n3244), .B2(n3896), .A(n3243), .ZN(U3262) );
  NAND2_X1 U4031 ( .A1(n3245), .A2(n3344), .ZN(n3248) );
  AOI22_X1 U4032 ( .A1(n3273), .A2(n4460), .B1(REG3_REG_0__SCAN_IN), .B2(n3246), .ZN(n3247) );
  OAI211_X1 U4033 ( .C1(n2708), .C2(n3388), .A(n3248), .B(n3247), .ZN(U3229)
         );
  AOI21_X1 U4034 ( .B1(n3250), .B2(n3249), .A(n3406), .ZN(n3252) );
  NAND2_X1 U4035 ( .A1(n3252), .A2(n3251), .ZN(n3258) );
  AOI22_X1 U4036 ( .A1(n3399), .A2(n3573), .B1(n3398), .B2(n3571), .ZN(n3257)
         );
  NOR2_X1 U4037 ( .A1(STATE_REG_SCAN_IN), .A2(n4098), .ZN(n4284) );
  NOR2_X1 U4038 ( .A1(n3401), .A2(n3253), .ZN(n3254) );
  AOI211_X1 U4039 ( .C1(n3403), .C2(n3255), .A(n4284), .B(n3254), .ZN(n3256)
         );
  NAND3_X1 U4040 ( .A1(n3258), .A2(n3257), .A3(n3256), .ZN(U3210) );
  XNOR2_X1 U4041 ( .A(n3259), .B(n3260), .ZN(n3266) );
  INV_X1 U4042 ( .A(n3261), .ZN(n3677) );
  OAI22_X1 U40430 ( .A1(n3401), .A2(n3676), .B1(STATE_REG_SCAN_IN), .B2(n3262), 
        .ZN(n3264) );
  OAI22_X1 U4044 ( .A1(n3671), .A2(n3388), .B1(n3298), .B2(n3387), .ZN(n3263)
         );
  AOI211_X1 U4045 ( .C1(n3677), .C2(n3403), .A(n3264), .B(n3263), .ZN(n3265)
         );
  OAI21_X1 U4046 ( .B1(n3266), .B2(n3406), .A(n3265), .ZN(U3211) );
  INV_X1 U4047 ( .A(n3267), .ZN(n3364) );
  OAI21_X1 U4048 ( .B1(n3364), .B2(n3269), .A(n3268), .ZN(n3271) );
  NAND3_X1 U4049 ( .A1(n3271), .A2(n3344), .A3(n3270), .ZN(n3277) );
  AOI22_X1 U4050 ( .A1(n3398), .A2(n3745), .B1(n3399), .B2(n3564), .ZN(n3276)
         );
  AOI22_X1 U4051 ( .A1(n3273), .A2(n3272), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3275) );
  NAND2_X1 U4052 ( .A1(n3403), .A2(n3751), .ZN(n3274) );
  NAND4_X1 U4053 ( .A1(n3277), .A2(n3276), .A3(n3275), .A4(n3274), .ZN(U3213)
         );
  XOR2_X1 U4054 ( .A(n3279), .B(n3278), .Z(n3283) );
  AOI22_X1 U4055 ( .A1(n3399), .A2(n3565), .B1(n3398), .B2(n3818), .ZN(n3282)
         );
  NAND2_X1 U4056 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3658) );
  OAI21_X1 U4057 ( .B1(n3401), .B2(n3823), .A(n3658), .ZN(n3280) );
  AOI21_X1 U4058 ( .B1(n3824), .B2(n3403), .A(n3280), .ZN(n3281) );
  OAI211_X1 U4059 ( .C1(n3283), .C2(n3406), .A(n3282), .B(n3281), .ZN(U3216)
         );
  XNOR2_X1 U4060 ( .A(n3285), .B(n3284), .ZN(n3286) );
  XNOR2_X1 U4061 ( .A(n3287), .B(n3286), .ZN(n3292) );
  AOI22_X1 U4062 ( .A1(n3399), .A2(n3818), .B1(n3398), .B2(n3564), .ZN(n3291)
         );
  OAI22_X1 U4063 ( .A1(n3401), .A2(n3780), .B1(STATE_REG_SCAN_IN), .B2(n3288), 
        .ZN(n3289) );
  AOI21_X1 U4064 ( .B1(n3782), .B2(n3403), .A(n3289), .ZN(n3290) );
  OAI211_X1 U4065 ( .C1(n3292), .C2(n3406), .A(n3291), .B(n3290), .ZN(U3220)
         );
  NAND2_X1 U4066 ( .A1(n3294), .A2(n3293), .ZN(n3296) );
  XOR2_X1 U4067 ( .A(n3296), .B(n3295), .Z(n3303) );
  INV_X1 U4068 ( .A(n3297), .ZN(n3713) );
  OAI22_X1 U4069 ( .A1(n3298), .A2(n3388), .B1(n3387), .B2(n3707), .ZN(n3301)
         );
  OAI22_X1 U4070 ( .A1(n3401), .A2(n3712), .B1(STATE_REG_SCAN_IN), .B2(n3299), 
        .ZN(n3300) );
  AOI211_X1 U4071 ( .C1(n3713), .C2(n3403), .A(n3301), .B(n3300), .ZN(n3302)
         );
  OAI21_X1 U4072 ( .B1(n3303), .B2(n3406), .A(n3302), .ZN(U3222) );
  INV_X1 U4073 ( .A(n3304), .ZN(n3306) );
  OAI21_X1 U4074 ( .B1(n3306), .B2(n3397), .A(n3305), .ZN(n3307) );
  XOR2_X1 U4075 ( .A(n3308), .B(n3307), .Z(n3313) );
  OAI22_X1 U4076 ( .A1(n3309), .A2(n3387), .B1(n3388), .B2(n3865), .ZN(n3311)
         );
  NAND2_X1 U4077 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4378) );
  OAI21_X1 U4078 ( .B1(n3401), .B2(n3870), .A(n4378), .ZN(n3310) );
  AOI211_X1 U4079 ( .C1(n3871), .C2(n3403), .A(n3311), .B(n3310), .ZN(n3312)
         );
  OAI21_X1 U4080 ( .B1(n3313), .B2(n3406), .A(n3312), .ZN(U3223) );
  XNOR2_X1 U4081 ( .A(n3316), .B(n3315), .ZN(n3317) );
  XNOR2_X1 U4082 ( .A(n3314), .B(n3317), .ZN(n3321) );
  AOI22_X1 U4083 ( .A1(n3399), .A2(n3853), .B1(n3398), .B2(n3565), .ZN(n3320)
         );
  NOR2_X1 U4084 ( .A1(STATE_REG_SCAN_IN), .A2(n2481), .ZN(n4392) );
  NOR2_X1 U4085 ( .A1(n3401), .A2(n3857), .ZN(n3318) );
  AOI211_X1 U4086 ( .C1(n3403), .C2(n3858), .A(n4392), .B(n3318), .ZN(n3319)
         );
  OAI211_X1 U4087 ( .C1(n3321), .C2(n3406), .A(n3320), .B(n3319), .ZN(U3225)
         );
  NAND2_X1 U4088 ( .A1(n3322), .A2(n3323), .ZN(n3324) );
  XOR2_X1 U4089 ( .A(n3325), .B(n3324), .Z(n3331) );
  INV_X1 U4090 ( .A(n3326), .ZN(n3729) );
  OAI22_X1 U4091 ( .A1(n3722), .A2(n3387), .B1(n3388), .B2(n3694), .ZN(n3329)
         );
  OAI22_X1 U4092 ( .A1(n3401), .A2(n3728), .B1(STATE_REG_SCAN_IN), .B2(n3327), 
        .ZN(n3328) );
  AOI211_X1 U4093 ( .C1(n3729), .C2(n3403), .A(n3329), .B(n3328), .ZN(n3330)
         );
  OAI21_X1 U4094 ( .B1(n3331), .B2(n3406), .A(n3330), .ZN(U3226) );
  OAI21_X1 U4095 ( .B1(n3334), .B2(n3333), .A(n3332), .ZN(n3335) );
  NAND3_X1 U4096 ( .A1(n2090), .A2(n3344), .A3(n3335), .ZN(n3342) );
  AOI22_X1 U4097 ( .A1(n3398), .A2(n3574), .B1(n3399), .B2(n3919), .ZN(n3341)
         );
  NOR2_X1 U4098 ( .A1(n3401), .A2(n3336), .ZN(n3337) );
  AOI211_X1 U4099 ( .C1(n3403), .C2(n3339), .A(n3338), .B(n3337), .ZN(n3340)
         );
  NAND3_X1 U4100 ( .A1(n3342), .A2(n3341), .A3(n3340), .ZN(U3227) );
  OAI21_X1 U4101 ( .B1(n3343), .B2(n2279), .A(n2978), .ZN(n3345) );
  NAND2_X1 U4102 ( .A1(n3345), .A2(n3344), .ZN(n3352) );
  AOI22_X1 U4103 ( .A1(n3399), .A2(n3571), .B1(n3398), .B2(n4412), .ZN(n3351)
         );
  NOR2_X1 U4104 ( .A1(STATE_REG_SCAN_IN), .A2(n3346), .ZN(n4311) );
  NOR2_X1 U4105 ( .A1(n3401), .A2(n3347), .ZN(n3348) );
  AOI211_X1 U4106 ( .C1(n3403), .C2(n3349), .A(n4311), .B(n3348), .ZN(n3350)
         );
  NAND3_X1 U4107 ( .A1(n3352), .A2(n3351), .A3(n3350), .ZN(U3228) );
  INV_X1 U4108 ( .A(n3353), .ZN(n3358) );
  AOI21_X1 U4109 ( .B1(n3357), .B2(n3355), .A(n3354), .ZN(n3356) );
  AOI21_X1 U4110 ( .B1(n3358), .B2(n3357), .A(n3356), .ZN(n3363) );
  OAI22_X1 U4111 ( .A1(n3833), .A2(n3387), .B1(n3388), .B2(n3793), .ZN(n3361)
         );
  OAI22_X1 U4112 ( .A1(n3401), .A2(n3799), .B1(STATE_REG_SCAN_IN), .B2(n3359), 
        .ZN(n3360) );
  AOI211_X1 U4113 ( .C1(n3800), .C2(n3403), .A(n3361), .B(n3360), .ZN(n3362)
         );
  OAI21_X1 U4114 ( .B1(n3363), .B2(n3406), .A(n3362), .ZN(U3230) );
  AOI21_X1 U4115 ( .B1(n3366), .B2(n3365), .A(n3364), .ZN(n3372) );
  OAI22_X1 U4116 ( .A1(n3722), .A2(n3388), .B1(n3387), .B2(n3793), .ZN(n3370)
         );
  OAI22_X1 U4117 ( .A1(n3401), .A2(n3368), .B1(STATE_REG_SCAN_IN), .B2(n3367), 
        .ZN(n3369) );
  AOI211_X1 U4118 ( .C1(n3766), .C2(n3403), .A(n3370), .B(n3369), .ZN(n3371)
         );
  OAI21_X1 U4119 ( .B1(n3372), .B2(n3406), .A(n3371), .ZN(U3232) );
  INV_X1 U4120 ( .A(n3373), .ZN(n3374) );
  NOR2_X1 U4121 ( .A1(n3375), .A2(n3374), .ZN(n3376) );
  XNOR2_X1 U4122 ( .A(n3377), .B(n3376), .ZN(n3382) );
  AOI22_X1 U4123 ( .A1(n3398), .A2(n3795), .B1(n3399), .B2(n2493), .ZN(n3381)
         );
  NOR2_X1 U4124 ( .A1(STATE_REG_SCAN_IN), .A2(n3378), .ZN(n4401) );
  NOR2_X1 U4125 ( .A1(n3401), .A2(n3841), .ZN(n3379) );
  AOI211_X1 U4126 ( .C1(n3403), .C2(n3842), .A(n4401), .B(n3379), .ZN(n3380)
         );
  OAI211_X1 U4127 ( .C1(n3382), .C2(n3406), .A(n3381), .B(n3380), .ZN(U3235)
         );
  NOR2_X1 U4128 ( .A1(n2255), .A2(n3384), .ZN(n3385) );
  XNOR2_X1 U4129 ( .A(n3386), .B(n3385), .ZN(n3395) );
  INV_X1 U4130 ( .A(n3686), .ZN(n3393) );
  OAI22_X1 U4131 ( .A1(n3389), .A2(n3388), .B1(n3694), .B2(n3387), .ZN(n3392)
         );
  OAI22_X1 U4132 ( .A1(n3401), .A2(n3693), .B1(STATE_REG_SCAN_IN), .B2(n3390), 
        .ZN(n3391) );
  AOI211_X1 U4133 ( .C1(n3393), .C2(n3403), .A(n3392), .B(n3391), .ZN(n3394)
         );
  OAI21_X1 U4134 ( .B1(n3395), .B2(n3406), .A(n3394), .ZN(U3237) );
  NAND2_X1 U4135 ( .A1(n3305), .A2(n3304), .ZN(n3396) );
  XOR2_X1 U4136 ( .A(n3397), .B(n3396), .Z(n3407) );
  AOI22_X1 U4137 ( .A1(n3399), .A2(n3566), .B1(n3398), .B2(n3853), .ZN(n3405)
         );
  NOR2_X1 U4138 ( .A1(STATE_REG_SCAN_IN), .A2(n3400), .ZN(n4372) );
  NOR2_X1 U4139 ( .A1(n3401), .A2(n3889), .ZN(n3402) );
  AOI211_X1 U4140 ( .C1(n3403), .C2(n3890), .A(n4372), .B(n3402), .ZN(n3404)
         );
  OAI211_X1 U4141 ( .C1(n3407), .C2(n3406), .A(n3405), .B(n3404), .ZN(U3238)
         );
  INV_X1 U4142 ( .A(n3408), .ZN(n3409) );
  AOI21_X1 U4143 ( .B1(n3411), .B2(n3410), .A(n3409), .ZN(n3522) );
  OR2_X1 U4144 ( .A1(n3411), .A2(n3410), .ZN(n3417) );
  NAND2_X1 U4145 ( .A1(n2052), .A2(DATAI_30_), .ZN(n3938) );
  OR2_X1 U4146 ( .A1(n3478), .A2(n3938), .ZN(n3416) );
  NAND2_X1 U4147 ( .A1(n2559), .A2(REG1_REG_31__SCAN_IN), .ZN(n3415) );
  NAND2_X1 U4148 ( .A1(n2336), .A2(REG2_REG_31__SCAN_IN), .ZN(n3414) );
  NAND2_X1 U4149 ( .A1(n3412), .A2(REG0_REG_31__SCAN_IN), .ZN(n3413) );
  NAND3_X1 U4150 ( .A1(n3415), .A2(n3414), .A3(n3413), .ZN(n3933) );
  NAND2_X1 U4151 ( .A1(n2053), .A2(DATAI_31_), .ZN(n3931) );
  NAND2_X1 U4152 ( .A1(n3933), .A2(n3931), .ZN(n3481) );
  AND2_X1 U4153 ( .A1(n3416), .A2(n3481), .ZN(n3512) );
  NAND2_X1 U4154 ( .A1(n3417), .A2(n3512), .ZN(n3540) );
  AOI21_X1 U4155 ( .B1(n3522), .B2(n3542), .A(n3540), .ZN(n3546) );
  NOR2_X1 U4156 ( .A1(n3420), .A2(n2207), .ZN(n3530) );
  NAND2_X1 U4157 ( .A1(n3422), .A2(n3421), .ZN(n3460) );
  AND2_X1 U4158 ( .A1(n3460), .A2(n3523), .ZN(n3527) );
  INV_X1 U4159 ( .A(n3423), .ZN(n3434) );
  AND2_X1 U4160 ( .A1(n3425), .A2(n3424), .ZN(n3426) );
  AND2_X1 U4161 ( .A1(n3428), .A2(n3426), .ZN(n3465) );
  INV_X1 U4162 ( .A(n3427), .ZN(n3430) );
  OAI21_X1 U4163 ( .B1(n3430), .B2(n3429), .A(n3428), .ZN(n3431) );
  NAND4_X1 U4164 ( .A1(n3877), .A2(n3432), .A3(n3523), .A4(n3431), .ZN(n3433)
         );
  AOI21_X1 U4165 ( .B1(n3434), .B2(n3465), .A(n3433), .ZN(n3467) );
  INV_X1 U4166 ( .A(n3435), .ZN(n3436) );
  NAND4_X1 U4167 ( .A1(n3436), .A2(n3456), .A3(n3455), .A4(n3448), .ZN(n3462)
         );
  INV_X1 U4168 ( .A(n3491), .ZN(n3453) );
  NAND2_X1 U4169 ( .A1(n3577), .A2(n4474), .ZN(n3499) );
  OAI211_X1 U4170 ( .C1(n4240), .C2(n2199), .A(n3499), .B(n3437), .ZN(n3438)
         );
  NAND3_X1 U4171 ( .A1(n3439), .A2(n2597), .A3(n3438), .ZN(n3441) );
  OAI211_X1 U4172 ( .C1(n3443), .C2(n3442), .A(n3441), .B(n3440), .ZN(n3444)
         );
  NAND3_X1 U4173 ( .A1(n3446), .A2(n3445), .A3(n3444), .ZN(n3447) );
  NAND4_X1 U4174 ( .A1(n3450), .A2(n3449), .A3(n3448), .A4(n3447), .ZN(n3451)
         );
  NAND3_X1 U4175 ( .A1(n3453), .A2(n3452), .A3(n3451), .ZN(n3454) );
  NAND3_X1 U4176 ( .A1(n3456), .A2(n3455), .A3(n3454), .ZN(n3457) );
  AND3_X1 U4177 ( .A1(n3459), .A2(n3458), .A3(n3457), .ZN(n3461) );
  OAI22_X1 U4178 ( .A1(n3527), .A2(n3462), .B1(n3461), .B2(n3460), .ZN(n3463)
         );
  NAND3_X1 U4179 ( .A1(n3465), .A2(n3464), .A3(n3463), .ZN(n3466) );
  OAI211_X1 U4180 ( .C1(n3527), .C2(n3467), .A(n3526), .B(n3466), .ZN(n3468)
         );
  NAND3_X1 U4181 ( .A1(n3530), .A2(n2209), .A3(n3468), .ZN(n3469) );
  AND2_X1 U4182 ( .A1(n3470), .A2(n3469), .ZN(n3471) );
  OAI21_X1 U4183 ( .B1(n3737), .B2(n3471), .A(n3532), .ZN(n3472) );
  INV_X1 U4184 ( .A(n3472), .ZN(n3474) );
  OAI211_X1 U4185 ( .C1(n3475), .C2(n3474), .A(n3473), .B(n3538), .ZN(n3476)
         );
  NAND4_X1 U4186 ( .A1(n3522), .A2(n2188), .A3(n3477), .A4(n3476), .ZN(n3482)
         );
  NOR2_X1 U4187 ( .A1(n3933), .A2(n3931), .ZN(n3550) );
  INV_X1 U4188 ( .A(n3550), .ZN(n3480) );
  AND2_X1 U4189 ( .A1(n3478), .A2(n3938), .ZN(n3551) );
  INV_X1 U4190 ( .A(n3551), .ZN(n3479) );
  NAND2_X1 U4191 ( .A1(n3480), .A2(n3479), .ZN(n3514) );
  AOI22_X1 U4192 ( .A1(n3546), .A2(n3482), .B1(n3481), .B2(n3514), .ZN(n3555)
         );
  INV_X1 U4193 ( .A(n3665), .ZN(n3484) );
  NAND2_X1 U4194 ( .A1(n3809), .A2(n3807), .ZN(n3850) );
  NOR3_X1 U4195 ( .A1(n3484), .A2(n3850), .A3(n3483), .ZN(n3495) );
  NOR4_X1 U4196 ( .A1(n3830), .A2(n3486), .A3(n4416), .A4(n3485), .ZN(n3494)
         );
  NOR4_X1 U4197 ( .A1(n2134), .A2(n3489), .A3(n3488), .A4(n3487), .ZN(n3493)
         );
  INV_X1 U4198 ( .A(n3899), .ZN(n3903) );
  NOR4_X1 U4199 ( .A1(n3903), .A2(n2598), .A3(n3491), .A4(n4452), .ZN(n3492)
         );
  AND4_X1 U4200 ( .A1(n3495), .A2(n3494), .A3(n3493), .A4(n3492), .ZN(n3503)
         );
  INV_X1 U4201 ( .A(n3496), .ZN(n3502) );
  NAND2_X1 U4202 ( .A1(n3497), .A2(n3521), .ZN(n3691) );
  INV_X1 U4203 ( .A(n3739), .ZN(n3498) );
  OR2_X1 U4204 ( .A1(n3737), .A2(n3498), .ZN(n3773) );
  NAND2_X1 U4205 ( .A1(n4451), .A2(n3499), .ZN(n4520) );
  NOR4_X1 U4206 ( .A1(n3691), .A2(n3773), .A3(n3879), .A4(n4520), .ZN(n3500)
         );
  NAND4_X1 U4207 ( .A1(n3503), .A2(n3502), .A3(n3501), .A4(n3500), .ZN(n3520)
         );
  XNOR2_X1 U4208 ( .A(n3833), .B(n3823), .ZN(n3806) );
  INV_X1 U4209 ( .A(n3806), .ZN(n3814) );
  NAND2_X1 U4210 ( .A1(n3504), .A2(n3702), .ZN(n3720) );
  NAND2_X1 U4211 ( .A1(n3718), .A2(n3505), .ZN(n3742) );
  NOR4_X1 U4212 ( .A1(n3507), .A2(n3506), .A3(n3720), .A4(n3742), .ZN(n3517)
         );
  INV_X1 U4213 ( .A(n3508), .ZN(n3509) );
  NOR2_X1 U4214 ( .A1(n3510), .A2(n3509), .ZN(n3791) );
  NAND2_X1 U4215 ( .A1(n3689), .A2(n3511), .ZN(n3705) );
  INV_X1 U4216 ( .A(n3512), .ZN(n3513) );
  NOR4_X1 U4217 ( .A1(n3791), .A2(n3705), .A3(n3514), .A4(n3513), .ZN(n3516)
         );
  NAND3_X1 U4218 ( .A1(n3517), .A2(n3516), .A3(n3515), .ZN(n3518) );
  NOR4_X1 U4219 ( .A1(n3520), .A2(n3814), .A3(n3519), .A4(n3518), .ZN(n3553)
         );
  INV_X1 U4220 ( .A(n3931), .ZN(n3934) );
  INV_X1 U4221 ( .A(n3938), .ZN(n3941) );
  INV_X1 U4222 ( .A(n3933), .ZN(n3548) );
  NAND3_X1 U4223 ( .A1(n3522), .A2(n3665), .A3(n3521), .ZN(n3545) );
  INV_X1 U4224 ( .A(n3523), .ZN(n3524) );
  NOR3_X1 U4225 ( .A1(n3898), .A2(n3525), .A3(n3524), .ZN(n3528) );
  OAI21_X1 U4226 ( .B1(n3528), .B2(n3527), .A(n3526), .ZN(n3531) );
  AOI21_X1 U4227 ( .B1(n3531), .B2(n3530), .A(n3529), .ZN(n3534) );
  OAI21_X1 U4228 ( .B1(n3534), .B2(n3533), .A(n3532), .ZN(n3536) );
  NAND2_X1 U4229 ( .A1(n3536), .A2(n3535), .ZN(n3539) );
  INV_X1 U4230 ( .A(n3537), .ZN(n3690) );
  AOI21_X1 U4231 ( .B1(n3539), .B2(n3538), .A(n3690), .ZN(n3543) );
  NOR4_X1 U4232 ( .A1(n3543), .A2(n3542), .A3(n3541), .A4(n3540), .ZN(n3544)
         );
  AOI21_X1 U4233 ( .B1(n3546), .B2(n3545), .A(n3544), .ZN(n3547) );
  AOI21_X1 U4234 ( .B1(n3941), .B2(n3548), .A(n3547), .ZN(n3549) );
  AOI211_X1 U4235 ( .C1(n3934), .C2(n3551), .A(n3550), .B(n3549), .ZN(n3552)
         );
  MUX2_X1 U4236 ( .A(n3553), .B(n3552), .S(n4240), .Z(n3554) );
  MUX2_X1 U4237 ( .A(n3555), .B(n3554), .S(n4241), .Z(n3556) );
  XNOR2_X1 U4238 ( .A(n3556), .B(n4242), .ZN(n3562) );
  NOR2_X1 U4239 ( .A1(n3558), .A2(n3557), .ZN(n3560) );
  OAI21_X1 U4240 ( .B1(n3561), .B2(n4239), .A(B_REG_SCAN_IN), .ZN(n3559) );
  OAI22_X1 U4241 ( .A1(n3562), .A2(n3561), .B1(n3560), .B2(n3559), .ZN(U3239)
         );
  MUX2_X1 U4242 ( .A(n3933), .B(DATAO_REG_31__SCAN_IN), .S(n3576), .Z(U3581)
         );
  MUX2_X1 U4243 ( .A(DATAO_REG_28__SCAN_IN), .B(n3563), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4244 ( .A(DATAO_REG_27__SCAN_IN), .B(n3696), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4245 ( .A(DATAO_REG_26__SCAN_IN), .B(n3709), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4246 ( .A(DATAO_REG_25__SCAN_IN), .B(n3724), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4247 ( .A(DATAO_REG_24__SCAN_IN), .B(n3745), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4248 ( .A(DATAO_REG_22__SCAN_IN), .B(n3564), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4249 ( .A(DATAO_REG_19__SCAN_IN), .B(n3795), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4250 ( .A(DATAO_REG_18__SCAN_IN), .B(n3565), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4251 ( .A(DATAO_REG_17__SCAN_IN), .B(n2493), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4252 ( .A(DATAO_REG_16__SCAN_IN), .B(n3853), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4253 ( .A(n3900), .B(DATAO_REG_15__SCAN_IN), .S(n3576), .Z(U3565)
         );
  MUX2_X1 U4254 ( .A(DATAO_REG_14__SCAN_IN), .B(n3566), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4255 ( .A(n3567), .B(DATAO_REG_13__SCAN_IN), .S(n3576), .Z(U3563)
         );
  MUX2_X1 U4256 ( .A(DATAO_REG_12__SCAN_IN), .B(n3568), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4257 ( .A(DATAO_REG_11__SCAN_IN), .B(n3569), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4258 ( .A(n4412), .B(DATAO_REG_10__SCAN_IN), .S(n3576), .Z(U3560)
         );
  MUX2_X1 U4259 ( .A(n3570), .B(DATAO_REG_9__SCAN_IN), .S(n3576), .Z(U3559) );
  MUX2_X1 U4260 ( .A(n3571), .B(DATAO_REG_8__SCAN_IN), .S(n3576), .Z(U3558) );
  MUX2_X1 U4261 ( .A(DATAO_REG_7__SCAN_IN), .B(n3572), .S(U4043), .Z(U3557) );
  MUX2_X1 U4262 ( .A(n3573), .B(DATAO_REG_6__SCAN_IN), .S(n3576), .Z(U3556) );
  MUX2_X1 U4263 ( .A(n3574), .B(DATAO_REG_5__SCAN_IN), .S(n3576), .Z(U3555) );
  MUX2_X1 U4264 ( .A(DATAO_REG_4__SCAN_IN), .B(n3575), .S(U4043), .Z(U3554) );
  MUX2_X1 U4265 ( .A(n3919), .B(DATAO_REG_3__SCAN_IN), .S(n3576), .Z(U3553) );
  MUX2_X1 U4266 ( .A(DATAO_REG_2__SCAN_IN), .B(n2331), .S(U4043), .Z(U3552) );
  MUX2_X1 U4267 ( .A(DATAO_REG_1__SCAN_IN), .B(n2323), .S(U4043), .Z(U3551) );
  MUX2_X1 U4268 ( .A(DATAO_REG_0__SCAN_IN), .B(n3577), .S(U4043), .Z(U3550) );
  INV_X1 U4269 ( .A(n3578), .ZN(n3580) );
  OAI211_X1 U4270 ( .C1(n3580), .C2(n3579), .A(n4345), .B(n3593), .ZN(n3588)
         );
  OAI211_X1 U4271 ( .C1(n3583), .C2(n3582), .A(n4404), .B(n3581), .ZN(n3587)
         );
  AOI22_X1 U4272 ( .A1(n4402), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3586) );
  INV_X1 U4273 ( .A(n4409), .ZN(n3584) );
  NAND4_X1 U4274 ( .A1(n3588), .A2(n3587), .A3(n3586), .A4(n3585), .ZN(U3241)
         );
  AOI22_X1 U4275 ( .A1(n4402), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3589) );
  OAI21_X1 U4276 ( .B1(n3590), .B2(n4409), .A(n3589), .ZN(n3591) );
  INV_X1 U4277 ( .A(n3591), .ZN(n3602) );
  MUX2_X1 U4278 ( .A(n3925), .B(REG2_REG_2__SCAN_IN), .S(n4245), .Z(n3594) );
  NAND3_X1 U4279 ( .A1(n3594), .A2(n3593), .A3(n3592), .ZN(n3595) );
  NAND3_X1 U4280 ( .A1(n4345), .A2(n3596), .A3(n3595), .ZN(n3601) );
  OAI211_X1 U4281 ( .C1(n3599), .C2(n3598), .A(n4404), .B(n3597), .ZN(n3600)
         );
  NAND4_X1 U4282 ( .A1(n3603), .A2(n3602), .A3(n3601), .A4(n3600), .ZN(U3242)
         );
  INV_X1 U4283 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3621) );
  INV_X1 U4284 ( .A(n3654), .ZN(n4493) );
  AOI22_X1 U4285 ( .A1(n3654), .A2(REG1_REG_18__SCAN_IN), .B1(n3621), .B2(
        n4493), .ZN(n4406) );
  INV_X1 U4286 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4167) );
  INV_X1 U4287 ( .A(n3649), .ZN(n4498) );
  INV_X1 U4288 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U4289 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3649), .B1(n4498), .B2(
        n4174), .ZN(n4375) );
  INV_X1 U4290 ( .A(n4501), .ZN(n4356) );
  INV_X1 U4291 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U4292 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4501), .B1(n4356), .B2(
        n4042), .ZN(n4353) );
  NAND2_X1 U4293 ( .A1(n4300), .A2(REG1_REG_9__SCAN_IN), .ZN(n3612) );
  INV_X1 U4294 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3604) );
  MUX2_X1 U4295 ( .A(REG1_REG_9__SCAN_IN), .B(n3604), .S(n4300), .Z(n4302) );
  INV_X1 U4296 ( .A(n3605), .ZN(n3607) );
  INV_X1 U4297 ( .A(n4515), .ZN(n4269) );
  INV_X1 U4298 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4582) );
  AOI22_X1 U4299 ( .A1(REG1_REG_5__SCAN_IN), .A2(n4269), .B1(n4515), .B2(n4582), .ZN(n4260) );
  INV_X1 U4300 ( .A(n3634), .ZN(n4514) );
  NOR2_X1 U4301 ( .A1(n3608), .A2(n4514), .ZN(n3609) );
  INV_X1 U4302 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4273) );
  XNOR2_X1 U4303 ( .A(n4514), .B(n3608), .ZN(n4272) );
  INV_X1 U4304 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4584) );
  NAND2_X1 U4305 ( .A1(n3636), .A2(n3610), .ZN(n3611) );
  INV_X1 U4306 ( .A(n3636), .ZN(n4510) );
  NAND2_X1 U4307 ( .A1(n3611), .A2(n4296), .ZN(n4303) );
  NAND2_X1 U4308 ( .A1(n4302), .A2(n4303), .ZN(n4301) );
  NAND2_X1 U4309 ( .A1(n4507), .A2(n3613), .ZN(n3614) );
  INV_X1 U4310 ( .A(n4507), .ZN(n4319) );
  XNOR2_X1 U4311 ( .A(n3613), .B(n4319), .ZN(n4314) );
  NAND2_X1 U4312 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4314), .ZN(n4313) );
  INV_X1 U4313 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4588) );
  AOI22_X1 U4314 ( .A1(n4505), .A2(REG1_REG_11__SCAN_IN), .B1(n4588), .B2(
        n4334), .ZN(n4331) );
  NAND2_X1 U4315 ( .A1(n3644), .A2(n3615), .ZN(n3616) );
  NAND2_X1 U4316 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4341), .ZN(n4340) );
  NAND2_X1 U4317 ( .A1(n4499), .A2(n3617), .ZN(n3618) );
  NAND2_X1 U4318 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4364), .ZN(n4363) );
  NAND2_X1 U4319 ( .A1(n3618), .A2(n4363), .ZN(n4374) );
  NAND2_X1 U4320 ( .A1(n4375), .A2(n4374), .ZN(n4373) );
  NOR2_X1 U4321 ( .A1(n3650), .A2(n3619), .ZN(n3620) );
  AOI22_X1 U4322 ( .A1(REG1_REG_17__SCAN_IN), .A2(n4494), .B1(n3653), .B2(
        n4167), .ZN(n4393) );
  NAND2_X1 U4323 ( .A1(n4406), .A2(n4405), .ZN(n4403) );
  OAI21_X1 U4324 ( .B1(n3621), .B2(n4493), .A(n4403), .ZN(n3623) );
  XNOR2_X1 U4325 ( .A(n3659), .B(REG1_REG_19__SCAN_IN), .ZN(n3622) );
  XNOR2_X1 U4326 ( .A(n3623), .B(n3622), .ZN(n3663) );
  INV_X1 U4327 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4328 ( .A1(n3654), .A2(n3624), .B1(REG2_REG_18__SCAN_IN), .B2(
        n4493), .ZN(n4399) );
  INV_X1 U4329 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4330 ( .A1(REG2_REG_17__SCAN_IN), .A2(n3653), .B1(n4494), .B2(
        n3625), .ZN(n4390) );
  INV_X1 U4331 ( .A(n4499), .ZN(n4367) );
  INV_X1 U4332 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4333 ( .A1(n4505), .A2(REG2_REG_11__SCAN_IN), .B1(n3642), .B2(
        n4334), .ZN(n4325) );
  NAND2_X1 U4334 ( .A1(n4300), .A2(REG2_REG_9__SCAN_IN), .ZN(n3639) );
  MUX2_X1 U4335 ( .A(n2943), .B(REG2_REG_9__SCAN_IN), .S(n4300), .Z(n3626) );
  INV_X1 U4336 ( .A(n3626), .ZN(n4305) );
  AOI22_X1 U4337 ( .A1(n4280), .A2(REG2_REG_7__SCAN_IN), .B1(n3998), .B2(n4512), .ZN(n4288) );
  INV_X1 U4338 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4339 ( .A1(REG2_REG_5__SCAN_IN), .A2(n4515), .B1(n4269), .B2(n3632), .ZN(n4266) );
  INV_X1 U4340 ( .A(n3627), .ZN(n3629) );
  OAI22_X1 U4341 ( .A1(n3631), .A2(n3630), .B1(n3629), .B2(n3628), .ZN(n4265)
         );
  NAND2_X1 U4342 ( .A1(n4266), .A2(n4265), .ZN(n4264) );
  OAI21_X1 U4343 ( .B1(n4269), .B2(n3632), .A(n4264), .ZN(n3633) );
  NAND2_X1 U4344 ( .A1(n3634), .A2(n3633), .ZN(n3635) );
  XOR2_X1 U4345 ( .A(n3634), .B(n3633), .Z(n4277) );
  NAND2_X1 U4346 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4277), .ZN(n4276) );
  NAND2_X1 U4347 ( .A1(n3635), .A2(n4276), .ZN(n4287) );
  NAND2_X1 U4348 ( .A1(n4288), .A2(n4287), .ZN(n4286) );
  NAND2_X1 U4349 ( .A1(n3636), .A2(n3637), .ZN(n3638) );
  XNOR2_X1 U4350 ( .A(n3637), .B(n4510), .ZN(n4292) );
  NAND2_X1 U4351 ( .A1(n4507), .A2(n3640), .ZN(n3641) );
  XNOR2_X1 U4352 ( .A(n3640), .B(n4319), .ZN(n4316) );
  NAND2_X1 U4353 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4316), .ZN(n4315) );
  NAND2_X1 U4354 ( .A1(n3644), .A2(n3643), .ZN(n3645) );
  NOR2_X1 U4355 ( .A1(n4367), .A2(n3646), .ZN(n3647) );
  INV_X1 U4356 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4359) );
  NOR2_X1 U4357 ( .A1(n4359), .A2(n4358), .ZN(n4357) );
  NAND2_X1 U4358 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3649), .ZN(n3648) );
  OAI21_X1 U4359 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3649), .A(n3648), .ZN(n4369) );
  INV_X1 U4360 ( .A(n3650), .ZN(n4496) );
  NAND2_X1 U4361 ( .A1(n3651), .A2(n4496), .ZN(n3652) );
  INV_X1 U4362 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4379) );
  NAND2_X1 U4363 ( .A1(n4381), .A2(n4379), .ZN(n4380) );
  XNOR2_X1 U4364 ( .A(n3659), .B(REG2_REG_19__SCAN_IN), .ZN(n3655) );
  XNOR2_X1 U4365 ( .A(n3656), .B(n3655), .ZN(n3661) );
  NAND2_X1 U4366 ( .A1(n4402), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3657) );
  OAI211_X1 U4367 ( .C1(n4409), .C2(n3659), .A(n3658), .B(n3657), .ZN(n3660)
         );
  AOI21_X1 U4368 ( .B1(n3661), .B2(n4345), .A(n3660), .ZN(n3662) );
  OAI21_X1 U4369 ( .B1(n3663), .B2(n4270), .A(n3662), .ZN(U3259) );
  XNOR2_X1 U4370 ( .A(n3664), .B(n3665), .ZN(n3948) );
  INV_X1 U4371 ( .A(n3948), .ZN(n3682) );
  NOR2_X1 U4372 ( .A1(n3666), .A2(n3665), .ZN(n3667) );
  OR2_X1 U4373 ( .A1(n3668), .A2(n3667), .ZN(n3673) );
  AOI22_X1 U4374 ( .A1(n3709), .A2(n4411), .B1(n3669), .B2(n4446), .ZN(n3670)
         );
  OAI21_X1 U4375 ( .B1(n3671), .B2(n4472), .A(n3670), .ZN(n3672) );
  AOI21_X1 U4376 ( .B1(n3673), .B2(n4469), .A(n3672), .ZN(n3949) );
  INV_X1 U4377 ( .A(n3949), .ZN(n3680) );
  INV_X1 U4378 ( .A(n3674), .ZN(n3675) );
  OAI21_X1 U4379 ( .B1(n3684), .B2(n3676), .A(n3675), .ZN(n3951) );
  AOI22_X1 U4380 ( .A1(n3677), .A2(n4458), .B1(n4466), .B2(
        REG2_REG_27__SCAN_IN), .ZN(n3678) );
  OAI21_X1 U4381 ( .B1(n3951), .B2(n3892), .A(n3678), .ZN(n3679) );
  AOI21_X1 U4382 ( .B1(n3680), .B2(n4477), .A(n3679), .ZN(n3681) );
  OAI21_X1 U4383 ( .B1(n3682), .B2(n3896), .A(n3681), .ZN(U3263) );
  XNOR2_X1 U4384 ( .A(n3683), .B(n3691), .ZN(n4130) );
  AOI21_X1 U4385 ( .B1(n3685), .B2(n2055), .A(n3684), .ZN(n4128) );
  OAI22_X1 U4386 ( .A1(n4477), .A2(n3687), .B1(n3686), .B2(n4482), .ZN(n3688)
         );
  AOI21_X1 U4387 ( .B1(n4128), .B2(n4463), .A(n3688), .ZN(n3700) );
  OAI21_X1 U4388 ( .B1(n3704), .B2(n3690), .A(n3689), .ZN(n3692) );
  XNOR2_X1 U4389 ( .A(n3692), .B(n3691), .ZN(n3698) );
  OAI22_X1 U4390 ( .A1(n3694), .A2(n4449), .B1(n3693), .B2(n3881), .ZN(n3695)
         );
  AOI21_X1 U4391 ( .B1(n3696), .B2(n4447), .A(n3695), .ZN(n3697) );
  OAI21_X1 U4392 ( .B1(n3698), .B2(n4453), .A(n3697), .ZN(n4127) );
  NAND2_X1 U4393 ( .A1(n4127), .A2(n4477), .ZN(n3699) );
  OAI211_X1 U4394 ( .C1(n4130), .C2(n3896), .A(n3700), .B(n3699), .ZN(U3264)
         );
  XOR2_X1 U4395 ( .A(n3705), .B(n3701), .Z(n4134) );
  INV_X1 U4396 ( .A(n4134), .ZN(n3717) );
  INV_X1 U4397 ( .A(n3702), .ZN(n3703) );
  NOR2_X1 U4398 ( .A1(n3704), .A2(n3703), .ZN(n3706) );
  XNOR2_X1 U4399 ( .A(n3706), .B(n3705), .ZN(n3711) );
  OAI22_X1 U4400 ( .A1(n3707), .A2(n4449), .B1(n3712), .B2(n3881), .ZN(n3708)
         );
  AOI21_X1 U4401 ( .B1(n4447), .B2(n3709), .A(n3708), .ZN(n3710) );
  OAI21_X1 U4402 ( .B1(n3711), .B2(n4453), .A(n3710), .ZN(n4133) );
  OAI21_X1 U4403 ( .B1(n2118), .B2(n3712), .A(n2055), .ZN(n4197) );
  AOI22_X1 U4404 ( .A1(n4466), .A2(REG2_REG_25__SCAN_IN), .B1(n3713), .B2(
        n4458), .ZN(n3714) );
  OAI21_X1 U4405 ( .B1(n4197), .B2(n3892), .A(n3714), .ZN(n3715) );
  AOI21_X1 U4406 ( .B1(n4133), .B2(n4477), .A(n3715), .ZN(n3716) );
  OAI21_X1 U4407 ( .B1(n3717), .B2(n3896), .A(n3716), .ZN(U3265) );
  XNOR2_X1 U4408 ( .A(n2069), .B(n3720), .ZN(n4138) );
  INV_X1 U4409 ( .A(n4138), .ZN(n3733) );
  NAND2_X1 U4410 ( .A1(n3719), .A2(n3718), .ZN(n3721) );
  XNOR2_X1 U4411 ( .A(n3721), .B(n3720), .ZN(n3726) );
  OAI22_X1 U4412 ( .A1(n3722), .A2(n4449), .B1(n3881), .B2(n3728), .ZN(n3723)
         );
  AOI21_X1 U4413 ( .B1(n4447), .B2(n3724), .A(n3723), .ZN(n3725) );
  OAI21_X1 U4414 ( .B1(n3726), .B2(n4453), .A(n3725), .ZN(n4137) );
  OAI21_X1 U4415 ( .B1(n3748), .B2(n3728), .A(n3727), .ZN(n4201) );
  AOI22_X1 U4416 ( .A1(n4466), .A2(REG2_REG_24__SCAN_IN), .B1(n3729), .B2(
        n4458), .ZN(n3730) );
  OAI21_X1 U4417 ( .B1(n4201), .B2(n3892), .A(n3730), .ZN(n3731) );
  AOI21_X1 U4418 ( .B1(n4137), .B2(n4477), .A(n3731), .ZN(n3732) );
  OAI21_X1 U4419 ( .B1(n3733), .B2(n3896), .A(n3732), .ZN(U3266) );
  OR2_X1 U4420 ( .A1(n3734), .A2(n3760), .ZN(n3756) );
  NAND2_X1 U4421 ( .A1(n3756), .A2(n3735), .ZN(n3736) );
  XOR2_X1 U4422 ( .A(n3742), .B(n3736), .Z(n4142) );
  INV_X1 U4423 ( .A(n4142), .ZN(n3755) );
  INV_X1 U4424 ( .A(n3737), .ZN(n3738) );
  NAND2_X1 U4425 ( .A1(n3774), .A2(n3738), .ZN(n3740) );
  NAND2_X1 U4426 ( .A1(n3740), .A2(n3739), .ZN(n3759) );
  NAND2_X1 U4427 ( .A1(n3759), .A2(n3760), .ZN(n3758) );
  NAND2_X1 U4428 ( .A1(n3758), .A2(n3741), .ZN(n3743) );
  XNOR2_X1 U4429 ( .A(n3743), .B(n3742), .ZN(n3747) );
  OAI22_X1 U4430 ( .A1(n3775), .A2(n4449), .B1(n3881), .B2(n3750), .ZN(n3744)
         );
  AOI21_X1 U4431 ( .B1(n4447), .B2(n3745), .A(n3744), .ZN(n3746) );
  OAI21_X1 U4432 ( .B1(n3747), .B2(n4453), .A(n3746), .ZN(n4141) );
  INV_X1 U4433 ( .A(n3748), .ZN(n3749) );
  OAI21_X1 U4434 ( .B1(n2122), .B2(n3750), .A(n3749), .ZN(n4205) );
  AOI22_X1 U4435 ( .A1(n4466), .A2(REG2_REG_23__SCAN_IN), .B1(n3751), .B2(
        n4458), .ZN(n3752) );
  OAI21_X1 U4436 ( .B1(n4205), .B2(n3892), .A(n3752), .ZN(n3753) );
  AOI21_X1 U4437 ( .B1(n4141), .B2(n4477), .A(n3753), .ZN(n3754) );
  OAI21_X1 U4438 ( .B1(n3755), .B2(n3896), .A(n3754), .ZN(U3267) );
  INV_X1 U4439 ( .A(n3734), .ZN(n3757) );
  OAI21_X1 U4440 ( .B1(n3757), .B2(n2134), .A(n3756), .ZN(n4149) );
  OAI21_X1 U4441 ( .B1(n3760), .B2(n3759), .A(n3758), .ZN(n3765) );
  NAND2_X1 U4442 ( .A1(n3767), .A2(n4446), .ZN(n3763) );
  NAND2_X1 U4443 ( .A1(n3761), .A2(n4447), .ZN(n3762) );
  OAI211_X1 U4444 ( .C1(n3793), .C2(n4449), .A(n3763), .B(n3762), .ZN(n3764)
         );
  AOI21_X1 U4445 ( .B1(n3765), .B2(n4469), .A(n3764), .ZN(n4148) );
  AOI22_X1 U4446 ( .A1(n4466), .A2(REG2_REG_22__SCAN_IN), .B1(n3766), .B2(
        n4458), .ZN(n3769) );
  NAND2_X1 U4447 ( .A1(n3779), .A2(n3767), .ZN(n4145) );
  NAND3_X1 U4448 ( .A1(n4146), .A2(n4463), .A3(n4145), .ZN(n3768) );
  OAI211_X1 U4449 ( .C1(n4148), .C2(n4466), .A(n3769), .B(n3768), .ZN(n3770)
         );
  INV_X1 U4450 ( .A(n3770), .ZN(n3771) );
  OAI21_X1 U4451 ( .B1(n4149), .B2(n3896), .A(n3771), .ZN(U3268) );
  XOR2_X1 U4452 ( .A(n3773), .B(n3772), .Z(n4151) );
  INV_X1 U4453 ( .A(n4151), .ZN(n3786) );
  XNOR2_X1 U4454 ( .A(n3774), .B(n3773), .ZN(n3778) );
  OAI22_X1 U4455 ( .A1(n3775), .A2(n4472), .B1(n3881), .B2(n3780), .ZN(n3776)
         );
  AOI21_X1 U4456 ( .B1(n4411), .B2(n3818), .A(n3776), .ZN(n3777) );
  OAI21_X1 U4457 ( .B1(n3778), .B2(n4453), .A(n3777), .ZN(n4150) );
  INV_X1 U4458 ( .A(n3798), .ZN(n3781) );
  OAI21_X1 U4459 ( .B1(n3781), .B2(n3780), .A(n3779), .ZN(n4210) );
  AOI22_X1 U4460 ( .A1(n4466), .A2(REG2_REG_21__SCAN_IN), .B1(n3782), .B2(
        n4458), .ZN(n3783) );
  OAI21_X1 U4461 ( .B1(n4210), .B2(n3892), .A(n3783), .ZN(n3784) );
  AOI21_X1 U4462 ( .B1(n4150), .B2(n4477), .A(n3784), .ZN(n3785) );
  OAI21_X1 U4463 ( .B1(n3786), .B2(n3896), .A(n3785), .ZN(U3269) );
  XNOR2_X1 U4464 ( .A(n3787), .B(n3791), .ZN(n4155) );
  INV_X1 U4465 ( .A(n4155), .ZN(n3804) );
  INV_X1 U4466 ( .A(n3788), .ZN(n3789) );
  NAND2_X1 U4467 ( .A1(n3790), .A2(n3789), .ZN(n3792) );
  XNOR2_X1 U4468 ( .A(n3792), .B(n3791), .ZN(n3797) );
  OAI22_X1 U4469 ( .A1(n3793), .A2(n4472), .B1(n3881), .B2(n3799), .ZN(n3794)
         );
  AOI21_X1 U4470 ( .B1(n4411), .B2(n3795), .A(n3794), .ZN(n3796) );
  OAI21_X1 U4471 ( .B1(n3797), .B2(n4453), .A(n3796), .ZN(n4154) );
  OAI21_X1 U4472 ( .B1(n3821), .B2(n3799), .A(n3798), .ZN(n4214) );
  AOI22_X1 U4473 ( .A1(n4466), .A2(REG2_REG_20__SCAN_IN), .B1(n3800), .B2(
        n4458), .ZN(n3801) );
  OAI21_X1 U4474 ( .B1(n4214), .B2(n3892), .A(n3801), .ZN(n3802) );
  AOI21_X1 U4475 ( .B1(n4154), .B2(n4477), .A(n3802), .ZN(n3803) );
  OAI21_X1 U4476 ( .B1(n3804), .B2(n3896), .A(n3803), .ZN(U3270) );
  XNOR2_X1 U4477 ( .A(n3805), .B(n3806), .ZN(n4159) );
  INV_X1 U4478 ( .A(n4159), .ZN(n3828) );
  INV_X1 U4479 ( .A(n3807), .ZN(n3808) );
  OR2_X1 U4480 ( .A1(n3849), .A2(n3808), .ZN(n3810) );
  NAND2_X1 U4481 ( .A1(n3810), .A2(n3809), .ZN(n3832) );
  INV_X1 U4482 ( .A(n3811), .ZN(n3813) );
  OAI21_X1 U4483 ( .B1(n3832), .B2(n3813), .A(n3812), .ZN(n3815) );
  XNOR2_X1 U4484 ( .A(n3815), .B(n3814), .ZN(n3816) );
  NAND2_X1 U4485 ( .A1(n3816), .A2(n4469), .ZN(n3820) );
  AOI22_X1 U4486 ( .A1(n3818), .A2(n4447), .B1(n3817), .B2(n4446), .ZN(n3819)
         );
  OAI211_X1 U4487 ( .C1(n3851), .C2(n4449), .A(n3820), .B(n3819), .ZN(n4158)
         );
  INV_X1 U4488 ( .A(n3821), .ZN(n3822) );
  OAI21_X1 U4489 ( .B1(n3839), .B2(n3823), .A(n3822), .ZN(n4218) );
  AOI22_X1 U4490 ( .A1(n4466), .A2(REG2_REG_19__SCAN_IN), .B1(n3824), .B2(
        n4458), .ZN(n3825) );
  OAI21_X1 U4491 ( .B1(n4218), .B2(n3892), .A(n3825), .ZN(n3826) );
  AOI21_X1 U4492 ( .B1(n4158), .B2(n4477), .A(n3826), .ZN(n3827) );
  OAI21_X1 U4493 ( .B1(n3828), .B2(n3896), .A(n3827), .ZN(U3271) );
  XOR2_X1 U4494 ( .A(n3830), .B(n3829), .Z(n4164) );
  INV_X1 U4495 ( .A(n3830), .ZN(n3831) );
  XNOR2_X1 U4496 ( .A(n3832), .B(n3831), .ZN(n3838) );
  OR2_X1 U4497 ( .A1(n3833), .A2(n4472), .ZN(n3836) );
  NAND2_X1 U4498 ( .A1(n3834), .A2(n4446), .ZN(n3835) );
  OAI211_X1 U4499 ( .C1(n3865), .C2(n4449), .A(n3836), .B(n3835), .ZN(n3837)
         );
  AOI21_X1 U4500 ( .B1(n3838), .B2(n4469), .A(n3837), .ZN(n4163) );
  INV_X1 U4501 ( .A(n4163), .ZN(n3846) );
  INV_X1 U4502 ( .A(n3839), .ZN(n3840) );
  OAI211_X1 U4503 ( .C1(n2113), .C2(n3841), .A(n3840), .B(n4569), .ZN(n4162)
         );
  AOI22_X1 U4504 ( .A1(n4466), .A2(REG2_REG_18__SCAN_IN), .B1(n3842), .B2(
        n4458), .ZN(n3843) );
  OAI21_X1 U4505 ( .B1(n4162), .B2(n3844), .A(n3843), .ZN(n3845) );
  AOI21_X1 U4506 ( .B1(n3846), .B2(n4477), .A(n3845), .ZN(n3847) );
  OAI21_X1 U4507 ( .B1(n4164), .B2(n3896), .A(n3847), .ZN(U3272) );
  XNOR2_X1 U4508 ( .A(n3848), .B(n3850), .ZN(n4166) );
  INV_X1 U4509 ( .A(n4166), .ZN(n3862) );
  XOR2_X1 U4510 ( .A(n3850), .B(n3849), .Z(n3855) );
  OAI22_X1 U4511 ( .A1(n3851), .A2(n4472), .B1(n3881), .B2(n3857), .ZN(n3852)
         );
  AOI21_X1 U4512 ( .B1(n4411), .B2(n3853), .A(n3852), .ZN(n3854) );
  OAI21_X1 U4513 ( .B1(n3855), .B2(n4453), .A(n3854), .ZN(n4165) );
  OAI21_X1 U4514 ( .B1(n2114), .B2(n3857), .A(n3856), .ZN(n4223) );
  AOI22_X1 U4515 ( .A1(n4466), .A2(REG2_REG_17__SCAN_IN), .B1(n3858), .B2(
        n4458), .ZN(n3859) );
  OAI21_X1 U4516 ( .B1(n4223), .B2(n3892), .A(n3859), .ZN(n3860) );
  AOI21_X1 U4517 ( .B1(n4165), .B2(n4477), .A(n3860), .ZN(n3861) );
  OAI21_X1 U4518 ( .B1(n3862), .B2(n3896), .A(n3861), .ZN(U3273) );
  XNOR2_X1 U4519 ( .A(n3863), .B(n2137), .ZN(n4170) );
  INV_X1 U4520 ( .A(n4170), .ZN(n3875) );
  XNOR2_X1 U4521 ( .A(n3864), .B(n2137), .ZN(n3868) );
  OAI22_X1 U4522 ( .A1(n3865), .A2(n4472), .B1(n3881), .B2(n3870), .ZN(n3866)
         );
  AOI21_X1 U4523 ( .B1(n4411), .B2(n3900), .A(n3866), .ZN(n3867) );
  OAI21_X1 U4524 ( .B1(n3868), .B2(n4453), .A(n3867), .ZN(n4169) );
  OAI21_X1 U4525 ( .B1(n3887), .B2(n3870), .A(n3869), .ZN(n4227) );
  AOI22_X1 U4526 ( .A1(n4466), .A2(REG2_REG_16__SCAN_IN), .B1(n3871), .B2(
        n4458), .ZN(n3872) );
  OAI21_X1 U4527 ( .B1(n4227), .B2(n3892), .A(n3872), .ZN(n3873) );
  AOI21_X1 U4528 ( .B1(n4169), .B2(n4477), .A(n3873), .ZN(n3874) );
  OAI21_X1 U4529 ( .B1(n3875), .B2(n3896), .A(n3874), .ZN(U3274) );
  XNOR2_X1 U4530 ( .A(n3876), .B(n3879), .ZN(n4173) );
  INV_X1 U4531 ( .A(n4173), .ZN(n3895) );
  NAND2_X1 U4532 ( .A1(n3897), .A2(n3877), .ZN(n3878) );
  XOR2_X1 U4533 ( .A(n3879), .B(n3878), .Z(n3885) );
  NOR2_X1 U4534 ( .A1(n3880), .A2(n4449), .ZN(n3884) );
  OAI22_X1 U4535 ( .A1(n3882), .A2(n4472), .B1(n3881), .B2(n3889), .ZN(n3883)
         );
  AOI211_X1 U4536 ( .C1(n3885), .C2(n4469), .A(n3884), .B(n3883), .ZN(n3886)
         );
  INV_X1 U4537 ( .A(n3886), .ZN(n4172) );
  INV_X1 U4538 ( .A(n3887), .ZN(n3888) );
  OAI21_X1 U4539 ( .B1(n3909), .B2(n3889), .A(n3888), .ZN(n4232) );
  AOI22_X1 U4540 ( .A1(n4466), .A2(REG2_REG_15__SCAN_IN), .B1(n3890), .B2(
        n4458), .ZN(n3891) );
  OAI21_X1 U4541 ( .B1(n4232), .B2(n3892), .A(n3891), .ZN(n3893) );
  AOI21_X1 U4542 ( .B1(n4172), .B2(n4477), .A(n3893), .ZN(n3894) );
  OAI21_X1 U4543 ( .B1(n3896), .B2(n3895), .A(n3894), .ZN(U3275) );
  OAI21_X1 U4544 ( .B1(n3899), .B2(n3898), .A(n3897), .ZN(n3907) );
  AOI22_X1 U4545 ( .A1(n3900), .A2(n4447), .B1(n4446), .B2(n3910), .ZN(n3901)
         );
  OAI21_X1 U4546 ( .B1(n3902), .B2(n4449), .A(n3901), .ZN(n3906) );
  XNOR2_X1 U4547 ( .A(n3904), .B(n3903), .ZN(n4181) );
  NOR2_X1 U4548 ( .A1(n4181), .A2(n4417), .ZN(n3905) );
  AOI211_X1 U4549 ( .C1(n4469), .C2(n3907), .A(n3906), .B(n3905), .ZN(n4180)
         );
  AOI22_X1 U4550 ( .A1(n4466), .A2(REG2_REG_14__SCAN_IN), .B1(n3908), .B2(
        n4458), .ZN(n3913) );
  INV_X1 U4551 ( .A(n3909), .ZN(n4178) );
  NAND2_X1 U4552 ( .A1(n3911), .A2(n3910), .ZN(n4177) );
  NAND3_X1 U4553 ( .A1(n4178), .A2(n4463), .A3(n4177), .ZN(n3912) );
  OAI211_X1 U4554 ( .C1(n4181), .C2(n3914), .A(n3913), .B(n3912), .ZN(n3915)
         );
  INV_X1 U4555 ( .A(n3915), .ZN(n3916) );
  OAI21_X1 U4556 ( .B1(n4180), .B2(n4466), .A(n3916), .ZN(U3276) );
  OAI21_X1 U4557 ( .B1(n3918), .B2(n2598), .A(n3917), .ZN(n4533) );
  AOI22_X1 U4558 ( .A1(n3919), .A2(n4447), .B1(n3927), .B2(n4446), .ZN(n3920)
         );
  OAI21_X1 U4559 ( .B1(n2708), .B2(n4449), .A(n3920), .ZN(n3924) );
  NAND3_X1 U4560 ( .A1(n2598), .A2(n2597), .A3(n4455), .ZN(n3921) );
  AOI21_X1 U4561 ( .B1(n3922), .B2(n3921), .A(n4453), .ZN(n3923) );
  AOI211_X1 U4562 ( .C1(n4470), .C2(n4533), .A(n3924), .B(n3923), .ZN(n4530)
         );
  MUX2_X1 U4563 ( .A(n3925), .B(n4530), .S(n4477), .Z(n3930) );
  AOI22_X1 U4564 ( .A1(n4533), .A2(n4468), .B1(REG3_REG_2__SCAN_IN), .B2(n4458), .ZN(n3929) );
  NAND2_X1 U4565 ( .A1(n2109), .A2(n3927), .ZN(n4529) );
  NAND3_X1 U4566 ( .A1(n4463), .A2(n4528), .A3(n4529), .ZN(n3928) );
  NAND3_X1 U4567 ( .A1(n3930), .A2(n3929), .A3(n3928), .ZN(U3288) );
  NAND2_X1 U4568 ( .A1(n3939), .A2(n3938), .ZN(n3937) );
  XNOR2_X1 U4569 ( .A(n3937), .B(n3931), .ZN(n4246) );
  INV_X1 U4570 ( .A(n4246), .ZN(n4188) );
  AND2_X1 U4571 ( .A1(n3933), .A2(n3932), .ZN(n3940) );
  AOI21_X1 U4572 ( .B1(n3934), .B2(n4446), .A(n3940), .ZN(n4248) );
  INV_X1 U4573 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3935) );
  MUX2_X1 U4574 ( .A(n4248), .B(n3935), .S(n4587), .Z(n3936) );
  OAI21_X1 U4575 ( .B1(n4188), .B2(n4176), .A(n3936), .ZN(U3549) );
  OAI21_X1 U4576 ( .B1(n3939), .B2(n3938), .A(n3937), .ZN(n4249) );
  AOI21_X1 U4577 ( .B1(n3941), .B2(n4446), .A(n3940), .ZN(n4252) );
  INV_X1 U4578 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3942) );
  MUX2_X1 U4579 ( .A(n4252), .B(n3942), .S(n4587), .Z(n3943) );
  OAI21_X1 U4580 ( .B1(n4249), .B2(n4176), .A(n3943), .ZN(U3548) );
  OAI21_X1 U4581 ( .B1(n3947), .B2(n4557), .A(n3946), .ZN(n4191) );
  MUX2_X1 U4582 ( .A(REG1_REG_29__SCAN_IN), .B(n4191), .S(n4590), .Z(U3547) );
  NAND2_X1 U4583 ( .A1(n3948), .A2(n4554), .ZN(n3950) );
  OAI211_X1 U4584 ( .C1(n4548), .C2(n3951), .A(n3950), .B(n3949), .ZN(n4192)
         );
  MUX2_X1 U4585 ( .A(REG1_REG_27__SCAN_IN), .B(n4192), .S(n4590), .Z(U3545) );
  OAI22_X1 U4586 ( .A1(REG2_REG_11__SCAN_IN), .A2(keyinput122), .B1(
        REG1_REG_13__SCAN_IN), .B2(keyinput127), .ZN(n3952) );
  AOI221_X1 U4587 ( .B1(REG2_REG_11__SCAN_IN), .B2(keyinput122), .C1(
        keyinput127), .C2(REG1_REG_13__SCAN_IN), .A(n3952), .ZN(n3959) );
  OAI22_X1 U4588 ( .A1(REG2_REG_6__SCAN_IN), .A2(keyinput92), .B1(
        REG2_REG_13__SCAN_IN), .B2(keyinput120), .ZN(n3953) );
  AOI221_X1 U4589 ( .B1(REG2_REG_6__SCAN_IN), .B2(keyinput92), .C1(keyinput120), .C2(REG2_REG_13__SCAN_IN), .A(n3953), .ZN(n3958) );
  OAI22_X1 U4590 ( .A1(REG1_REG_22__SCAN_IN), .A2(keyinput90), .B1(
        DATAO_REG_22__SCAN_IN), .B2(keyinput103), .ZN(n3954) );
  AOI221_X1 U4591 ( .B1(REG1_REG_22__SCAN_IN), .B2(keyinput90), .C1(
        keyinput103), .C2(DATAO_REG_22__SCAN_IN), .A(n3954), .ZN(n3957) );
  OAI22_X1 U4592 ( .A1(REG1_REG_20__SCAN_IN), .A2(keyinput102), .B1(
        REG1_REG_6__SCAN_IN), .B2(keyinput97), .ZN(n3955) );
  AOI221_X1 U4593 ( .B1(REG1_REG_20__SCAN_IN), .B2(keyinput102), .C1(
        keyinput97), .C2(REG1_REG_6__SCAN_IN), .A(n3955), .ZN(n3956) );
  NAND4_X1 U4594 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n3956), .ZN(n3987)
         );
  OAI22_X1 U4595 ( .A1(DATAO_REG_30__SCAN_IN), .A2(keyinput70), .B1(
        DATAO_REG_29__SCAN_IN), .B2(keyinput68), .ZN(n3960) );
  AOI221_X1 U4596 ( .B1(DATAO_REG_30__SCAN_IN), .B2(keyinput70), .C1(
        keyinput68), .C2(DATAO_REG_29__SCAN_IN), .A(n3960), .ZN(n3967) );
  OAI22_X1 U4597 ( .A1(DATAO_REG_14__SCAN_IN), .A2(keyinput110), .B1(
        DATAO_REG_17__SCAN_IN), .B2(keyinput112), .ZN(n3961) );
  AOI221_X1 U4598 ( .B1(DATAO_REG_14__SCAN_IN), .B2(keyinput110), .C1(
        keyinput112), .C2(DATAO_REG_17__SCAN_IN), .A(n3961), .ZN(n3966) );
  OAI22_X1 U4599 ( .A1(ADDR_REG_9__SCAN_IN), .A2(keyinput81), .B1(
        ADDR_REG_13__SCAN_IN), .B2(keyinput125), .ZN(n3962) );
  AOI221_X1 U4600 ( .B1(ADDR_REG_9__SCAN_IN), .B2(keyinput81), .C1(keyinput125), .C2(ADDR_REG_13__SCAN_IN), .A(n3962), .ZN(n3965) );
  OAI22_X1 U4601 ( .A1(REG2_REG_24__SCAN_IN), .A2(keyinput119), .B1(
        ADDR_REG_1__SCAN_IN), .B2(keyinput100), .ZN(n3963) );
  AOI221_X1 U4602 ( .B1(REG2_REG_24__SCAN_IN), .B2(keyinput119), .C1(
        keyinput100), .C2(ADDR_REG_1__SCAN_IN), .A(n3963), .ZN(n3964) );
  NAND4_X1 U4603 ( .A1(n3967), .A2(n3966), .A3(n3965), .A4(n3964), .ZN(n3986)
         );
  OAI22_X1 U4604 ( .A1(REG0_REG_18__SCAN_IN), .A2(keyinput104), .B1(
        REG0_REG_17__SCAN_IN), .B2(keyinput82), .ZN(n3968) );
  AOI221_X1 U4605 ( .B1(REG0_REG_18__SCAN_IN), .B2(keyinput104), .C1(
        keyinput82), .C2(REG0_REG_17__SCAN_IN), .A(n3968), .ZN(n3975) );
  OAI22_X1 U4606 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput95), .B1(DATAI_8_), 
        .B2(keyinput118), .ZN(n3969) );
  AOI221_X1 U4607 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput95), .C1(keyinput118), .C2(DATAI_8_), .A(n3969), .ZN(n3974) );
  OAI22_X1 U4608 ( .A1(D_REG_18__SCAN_IN), .A2(keyinput121), .B1(
        D_REG_3__SCAN_IN), .B2(keyinput106), .ZN(n3970) );
  AOI221_X1 U4609 ( .B1(D_REG_18__SCAN_IN), .B2(keyinput121), .C1(keyinput106), 
        .C2(D_REG_3__SCAN_IN), .A(n3970), .ZN(n3973) );
  OAI22_X1 U4610 ( .A1(REG0_REG_23__SCAN_IN), .A2(keyinput88), .B1(keyinput111), .B2(REG0_REG_22__SCAN_IN), .ZN(n3971) );
  AOI221_X1 U4611 ( .B1(REG0_REG_23__SCAN_IN), .B2(keyinput88), .C1(
        REG0_REG_22__SCAN_IN), .C2(keyinput111), .A(n3971), .ZN(n3972) );
  NAND4_X1 U4612 ( .A1(n3975), .A2(n3974), .A3(n3973), .A4(n3972), .ZN(n3985)
         );
  OAI22_X1 U4613 ( .A1(IR_REG_1__SCAN_IN), .A2(keyinput93), .B1(
        REG3_REG_5__SCAN_IN), .B2(keyinput83), .ZN(n3976) );
  AOI221_X1 U4614 ( .B1(IR_REG_1__SCAN_IN), .B2(keyinput93), .C1(keyinput83), 
        .C2(REG3_REG_5__SCAN_IN), .A(n3976), .ZN(n3983) );
  OAI22_X1 U4615 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput101), .B1(keyinput69), 
        .B2(ADDR_REG_18__SCAN_IN), .ZN(n3977) );
  AOI221_X1 U4616 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput101), .C1(
        ADDR_REG_18__SCAN_IN), .C2(keyinput69), .A(n3977), .ZN(n3982) );
  OAI22_X1 U4617 ( .A1(REG3_REG_21__SCAN_IN), .A2(keyinput72), .B1(keyinput105), .B2(DATAI_19_), .ZN(n3978) );
  AOI221_X1 U4618 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput72), .C1(DATAI_19_), 
        .C2(keyinput105), .A(n3978), .ZN(n3981) );
  OAI22_X1 U4619 ( .A1(D_REG_1__SCAN_IN), .A2(keyinput109), .B1(DATAI_17_), 
        .B2(keyinput64), .ZN(n3979) );
  AOI221_X1 U4620 ( .B1(D_REG_1__SCAN_IN), .B2(keyinput109), .C1(keyinput64), 
        .C2(DATAI_17_), .A(n3979), .ZN(n3980) );
  NAND4_X1 U4621 ( .A1(n3983), .A2(n3982), .A3(n3981), .A4(n3980), .ZN(n3984)
         );
  NOR4_X1 U4622 ( .A1(n3987), .A2(n3986), .A3(n3985), .A4(n3984), .ZN(n4035)
         );
  INV_X1 U4623 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4229) );
  INV_X1 U4624 ( .A(REG0_REG_26__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4625 ( .A1(n4229), .A2(keyinput126), .B1(n3989), .B2(keyinput79), 
        .ZN(n3988) );
  OAI221_X1 U4626 ( .B1(n4229), .B2(keyinput126), .C1(n3989), .C2(keyinput79), 
        .A(n3988), .ZN(n3996) );
  INV_X1 U4627 ( .A(DATAI_15_), .ZN(n4497) );
  INV_X1 U4628 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4556) );
  AOI22_X1 U4629 ( .A1(n4497), .A2(keyinput65), .B1(keyinput73), .B2(n4556), 
        .ZN(n3990) );
  OAI221_X1 U4630 ( .B1(n4497), .B2(keyinput65), .C1(n4556), .C2(keyinput73), 
        .A(n3990), .ZN(n3995) );
  INV_X1 U4631 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4521) );
  AOI22_X1 U4632 ( .A1(n4484), .A2(keyinput123), .B1(keyinput76), .B2(n4521), 
        .ZN(n3991) );
  OAI221_X1 U4633 ( .B1(n4484), .B2(keyinput123), .C1(n4521), .C2(keyinput76), 
        .A(n3991), .ZN(n3994) );
  AOI22_X1 U4634 ( .A1(n4575), .A2(keyinput74), .B1(n4485), .B2(keyinput115), 
        .ZN(n3992) );
  OAI221_X1 U4635 ( .B1(n4575), .B2(keyinput74), .C1(n4485), .C2(keyinput115), 
        .A(n3992), .ZN(n3993) );
  NOR4_X1 U4636 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n4034)
         );
  AOI22_X1 U4637 ( .A1(D_REG_29__SCAN_IN), .A2(keyinput117), .B1(n3998), .B2(
        keyinput91), .ZN(n3997) );
  OAI221_X1 U4638 ( .B1(D_REG_29__SCAN_IN), .B2(keyinput117), .C1(n3998), .C2(
        keyinput91), .A(n3997), .ZN(n4007) );
  AOI22_X1 U4639 ( .A1(REG0_REG_3__SCAN_IN), .A2(keyinput86), .B1(
        REG0_REG_4__SCAN_IN), .B2(keyinput99), .ZN(n3999) );
  OAI221_X1 U4640 ( .B1(REG0_REG_3__SCAN_IN), .B2(keyinput86), .C1(
        REG0_REG_4__SCAN_IN), .C2(keyinput99), .A(n3999), .ZN(n4006) );
  INV_X1 U4641 ( .A(REG2_REG_10__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4642 ( .A1(n4359), .A2(keyinput94), .B1(keyinput66), .B2(n4001), 
        .ZN(n4000) );
  OAI221_X1 U4643 ( .B1(n4359), .B2(keyinput94), .C1(n4001), .C2(keyinput66), 
        .A(n4000), .ZN(n4005) );
  AOI22_X1 U4644 ( .A1(n2691), .A2(keyinput89), .B1(n4003), .B2(keyinput98), 
        .ZN(n4002) );
  OAI221_X1 U4645 ( .B1(n2691), .B2(keyinput89), .C1(n4003), .C2(keyinput98), 
        .A(n4002), .ZN(n4004) );
  NOR4_X1 U4646 ( .A1(n4007), .A2(n4006), .A3(n4005), .A4(n4004), .ZN(n4033)
         );
  INV_X1 U4647 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4010) );
  INV_X1 U4648 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4649 ( .A1(n4010), .A2(keyinput124), .B1(n4009), .B2(keyinput78), 
        .ZN(n4008) );
  OAI221_X1 U4650 ( .B1(n4010), .B2(keyinput124), .C1(n4009), .C2(keyinput78), 
        .A(n4008), .ZN(n4014) );
  INV_X1 U4651 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4652 ( .A1(n4039), .A2(keyinput116), .B1(n4012), .B2(keyinput77), 
        .ZN(n4011) );
  OAI221_X1 U4653 ( .B1(n4039), .B2(keyinput116), .C1(n4012), .C2(keyinput77), 
        .A(n4011), .ZN(n4013) );
  NOR2_X1 U4654 ( .A1(n4014), .A2(n4013), .ZN(n4031) );
  AOI22_X1 U4655 ( .A1(n4037), .A2(keyinput96), .B1(n4115), .B2(keyinput108), 
        .ZN(n4015) );
  OAI221_X1 U4656 ( .B1(n4037), .B2(keyinput96), .C1(n4115), .C2(keyinput108), 
        .A(n4015), .ZN(n4018) );
  INV_X1 U4657 ( .A(DATAI_18_), .ZN(n4492) );
  INV_X1 U4658 ( .A(DATAI_27_), .ZN(n4094) );
  AOI22_X1 U4659 ( .A1(n4492), .A2(keyinput75), .B1(keyinput114), .B2(n4094), 
        .ZN(n4016) );
  OAI221_X1 U4660 ( .B1(n4492), .B2(keyinput75), .C1(n4094), .C2(keyinput114), 
        .A(n4016), .ZN(n4017) );
  NOR2_X1 U4661 ( .A1(n4018), .A2(n4017), .ZN(n4030) );
  AOI22_X1 U4662 ( .A1(n2481), .A2(keyinput84), .B1(n3106), .B2(keyinput71), 
        .ZN(n4019) );
  OAI221_X1 U4663 ( .B1(n2481), .B2(keyinput84), .C1(n3106), .C2(keyinput71), 
        .A(n4019), .ZN(n4021) );
  XNOR2_X1 U4664 ( .A(n4062), .B(keyinput113), .ZN(n4020) );
  NOR2_X1 U4665 ( .A1(n4021), .A2(n4020), .ZN(n4029) );
  INV_X1 U4666 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U4667 ( .A1(n4061), .A2(keyinput67), .B1(keyinput80), .B2(n4135), 
        .ZN(n4022) );
  OAI221_X1 U4668 ( .B1(n4061), .B2(keyinput67), .C1(n4135), .C2(keyinput80), 
        .A(n4022), .ZN(n4027) );
  XNOR2_X1 U4669 ( .A(IR_REG_27__SCAN_IN), .B(keyinput87), .ZN(n4025) );
  XNOR2_X1 U4670 ( .A(IR_REG_9__SCAN_IN), .B(keyinput107), .ZN(n4024) );
  XNOR2_X1 U4671 ( .A(IR_REG_2__SCAN_IN), .B(keyinput85), .ZN(n4023) );
  NAND3_X1 U4672 ( .A1(n4025), .A2(n4024), .A3(n4023), .ZN(n4026) );
  NOR2_X1 U4673 ( .A1(n4027), .A2(n4026), .ZN(n4028) );
  AND4_X1 U4674 ( .A1(n4031), .A2(n4030), .A3(n4029), .A4(n4028), .ZN(n4032)
         );
  AND4_X1 U4675 ( .A1(n4035), .A2(n4034), .A3(n4033), .A4(n4032), .ZN(n4126)
         );
  AOI22_X1 U4676 ( .A1(n4037), .A2(keyinput32), .B1(n4229), .B2(keyinput62), 
        .ZN(n4036) );
  OAI221_X1 U4677 ( .B1(n4037), .B2(keyinput32), .C1(n4229), .C2(keyinput62), 
        .A(n4036), .ZN(n4046) );
  INV_X1 U4678 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4344) );
  AOI22_X1 U4679 ( .A1(n4039), .A2(keyinput52), .B1(n4344), .B2(keyinput56), 
        .ZN(n4038) );
  OAI221_X1 U4680 ( .B1(n4039), .B2(keyinput52), .C1(n4344), .C2(keyinput56), 
        .A(n4038), .ZN(n4045) );
  INV_X1 U4681 ( .A(DATAI_8_), .ZN(n4509) );
  AOI22_X1 U4682 ( .A1(n4484), .A2(keyinput59), .B1(keyinput54), .B2(n4509), 
        .ZN(n4040) );
  OAI221_X1 U4683 ( .B1(n4484), .B2(keyinput59), .C1(n4509), .C2(keyinput54), 
        .A(n4040), .ZN(n4044) );
  AOI22_X1 U4684 ( .A1(n2492), .A2(keyinput0), .B1(keyinput63), .B2(n4042), 
        .ZN(n4041) );
  OAI221_X1 U4685 ( .B1(n2492), .B2(keyinput0), .C1(n4042), .C2(keyinput63), 
        .A(n4041), .ZN(n4043) );
  NOR4_X1 U4686 ( .A1(n4046), .A2(n4045), .A3(n4044), .A4(n4043), .ZN(n4082)
         );
  AOI22_X1 U4687 ( .A1(ADDR_REG_18__SCAN_IN), .A2(keyinput5), .B1(
        ADDR_REG_13__SCAN_IN), .B2(keyinput61), .ZN(n4047) );
  OAI221_X1 U4688 ( .B1(ADDR_REG_18__SCAN_IN), .B2(keyinput5), .C1(
        ADDR_REG_13__SCAN_IN), .C2(keyinput61), .A(n4047), .ZN(n4054) );
  AOI22_X1 U4689 ( .A1(ADDR_REG_9__SCAN_IN), .A2(keyinput17), .B1(
        REG3_REG_0__SCAN_IN), .B2(keyinput37), .ZN(n4048) );
  OAI221_X1 U4690 ( .B1(ADDR_REG_9__SCAN_IN), .B2(keyinput17), .C1(
        REG3_REG_0__SCAN_IN), .C2(keyinput37), .A(n4048), .ZN(n4053) );
  AOI22_X1 U4691 ( .A1(D_REG_18__SCAN_IN), .A2(keyinput57), .B1(
        D_REG_1__SCAN_IN), .B2(keyinput45), .ZN(n4049) );
  OAI221_X1 U4692 ( .B1(D_REG_18__SCAN_IN), .B2(keyinput57), .C1(
        D_REG_1__SCAN_IN), .C2(keyinput45), .A(n4049), .ZN(n4052) );
  AOI22_X1 U4693 ( .A1(REG0_REG_7__SCAN_IN), .A2(keyinput9), .B1(
        IR_REG_1__SCAN_IN), .B2(keyinput29), .ZN(n4050) );
  OAI221_X1 U4694 ( .B1(REG0_REG_7__SCAN_IN), .B2(keyinput9), .C1(
        IR_REG_1__SCAN_IN), .C2(keyinput29), .A(n4050), .ZN(n4051) );
  NOR4_X1 U4695 ( .A1(n4054), .A2(n4053), .A3(n4052), .A4(n4051), .ZN(n4081)
         );
  AOI22_X1 U4696 ( .A1(n4575), .A2(keyinput10), .B1(n4492), .B2(keyinput11), 
        .ZN(n4055) );
  OAI221_X1 U4697 ( .B1(n4575), .B2(keyinput10), .C1(n4492), .C2(keyinput11), 
        .A(n4055), .ZN(n4059) );
  AOI22_X1 U4698 ( .A1(n4057), .A2(keyinput6), .B1(n3106), .B2(keyinput7), 
        .ZN(n4056) );
  OAI221_X1 U4699 ( .B1(n4057), .B2(keyinput6), .C1(n3106), .C2(keyinput7), 
        .A(n4056), .ZN(n4058) );
  NOR2_X1 U4700 ( .A1(n4059), .A2(n4058), .ZN(n4079) );
  AOI22_X1 U4701 ( .A1(n4061), .A2(keyinput3), .B1(keyinput33), .B2(n4273), 
        .ZN(n4060) );
  OAI221_X1 U4702 ( .B1(n4061), .B2(keyinput3), .C1(n4273), .C2(keyinput33), 
        .A(n4060), .ZN(n4064) );
  XNOR2_X1 U4703 ( .A(n4062), .B(keyinput49), .ZN(n4063) );
  NOR2_X1 U4704 ( .A1(n4064), .A2(n4063), .ZN(n4078) );
  INV_X1 U4705 ( .A(D_REG_29__SCAN_IN), .ZN(n4483) );
  AOI22_X1 U4706 ( .A1(n4135), .A2(keyinput16), .B1(n4483), .B2(keyinput53), 
        .ZN(n4065) );
  OAI221_X1 U4707 ( .B1(n4135), .B2(keyinput16), .C1(n4483), .C2(keyinput53), 
        .A(n4065), .ZN(n4069) );
  AOI22_X1 U4708 ( .A1(n2691), .A2(keyinput25), .B1(n4067), .B2(keyinput41), 
        .ZN(n4066) );
  OAI221_X1 U4709 ( .B1(n2691), .B2(keyinput25), .C1(n4067), .C2(keyinput41), 
        .A(n4066), .ZN(n4068) );
  NOR2_X1 U4710 ( .A1(n4069), .A2(n4068), .ZN(n4077) );
  INV_X1 U4711 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U4712 ( .A1(n4497), .A2(keyinput1), .B1(keyinput24), .B2(n4203), 
        .ZN(n4070) );
  OAI221_X1 U4713 ( .B1(n4497), .B2(keyinput1), .C1(n4203), .C2(keyinput24), 
        .A(n4070), .ZN(n4075) );
  XNOR2_X1 U4714 ( .A(IR_REG_27__SCAN_IN), .B(keyinput23), .ZN(n4073) );
  XNOR2_X1 U4715 ( .A(IR_REG_2__SCAN_IN), .B(keyinput21), .ZN(n4072) );
  XNOR2_X1 U4716 ( .A(keyinput19), .B(REG3_REG_5__SCAN_IN), .ZN(n4071) );
  NAND3_X1 U4717 ( .A1(n4073), .A2(n4072), .A3(n4071), .ZN(n4074) );
  NOR2_X1 U4718 ( .A1(n4075), .A2(n4074), .ZN(n4076) );
  AND4_X1 U4719 ( .A1(n4079), .A2(n4078), .A3(n4077), .A4(n4076), .ZN(n4080)
         );
  NAND3_X1 U4720 ( .A1(n4082), .A2(n4081), .A3(n4080), .ZN(n4125) );
  AOI22_X1 U4721 ( .A1(DATAO_REG_14__SCAN_IN), .A2(keyinput46), .B1(
        REG2_REG_11__SCAN_IN), .B2(keyinput58), .ZN(n4083) );
  OAI221_X1 U4722 ( .B1(DATAO_REG_14__SCAN_IN), .B2(keyinput46), .C1(
        REG2_REG_11__SCAN_IN), .C2(keyinput58), .A(n4083), .ZN(n4090) );
  AOI22_X1 U4723 ( .A1(D_REG_3__SCAN_IN), .A2(keyinput42), .B1(
        REG1_REG_29__SCAN_IN), .B2(keyinput34), .ZN(n4084) );
  OAI221_X1 U4724 ( .B1(D_REG_3__SCAN_IN), .B2(keyinput42), .C1(
        REG1_REG_29__SCAN_IN), .C2(keyinput34), .A(n4084), .ZN(n4089) );
  AOI22_X1 U4725 ( .A1(REG1_REG_22__SCAN_IN), .A2(keyinput26), .B1(
        REG2_REG_14__SCAN_IN), .B2(keyinput30), .ZN(n4085) );
  OAI221_X1 U4726 ( .B1(REG1_REG_22__SCAN_IN), .B2(keyinput26), .C1(
        REG2_REG_14__SCAN_IN), .C2(keyinput30), .A(n4085), .ZN(n4088) );
  AOI22_X1 U4727 ( .A1(REG2_REG_10__SCAN_IN), .A2(keyinput2), .B1(
        REG2_REG_20__SCAN_IN), .B2(keyinput14), .ZN(n4086) );
  OAI221_X1 U4728 ( .B1(REG2_REG_10__SCAN_IN), .B2(keyinput2), .C1(
        REG2_REG_20__SCAN_IN), .C2(keyinput14), .A(n4086), .ZN(n4087) );
  NOR4_X1 U4729 ( .A1(n4090), .A2(n4089), .A3(n4088), .A4(n4087), .ZN(n4123)
         );
  INV_X1 U4730 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U4731 ( .A1(n4485), .A2(keyinput51), .B1(keyinput47), .B2(n4092), 
        .ZN(n4091) );
  OAI221_X1 U4732 ( .B1(n4485), .B2(keyinput51), .C1(n4092), .C2(keyinput47), 
        .A(n4091), .ZN(n4102) );
  AOI22_X1 U4733 ( .A1(n4095), .A2(keyinput55), .B1(keyinput50), .B2(n4094), 
        .ZN(n4093) );
  OAI221_X1 U4734 ( .B1(n4095), .B2(keyinput55), .C1(n4094), .C2(keyinput50), 
        .A(n4093), .ZN(n4101) );
  INV_X1 U4735 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4539) );
  INV_X1 U4736 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4221) );
  AOI22_X1 U4737 ( .A1(n4539), .A2(keyinput22), .B1(n4221), .B2(keyinput18), 
        .ZN(n4096) );
  OAI221_X1 U4738 ( .B1(n4539), .B2(keyinput22), .C1(n4221), .C2(keyinput18), 
        .A(n4096), .ZN(n4100) );
  INV_X1 U4739 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4156) );
  AOI22_X1 U4740 ( .A1(n4156), .A2(keyinput38), .B1(n4098), .B2(keyinput31), 
        .ZN(n4097) );
  OAI221_X1 U4741 ( .B1(n4156), .B2(keyinput38), .C1(n4098), .C2(keyinput31), 
        .A(n4097), .ZN(n4099) );
  NOR4_X1 U4742 ( .A1(n4102), .A2(n4101), .A3(n4100), .A4(n4099), .ZN(n4122)
         );
  AOI22_X1 U4743 ( .A1(REG2_REG_25__SCAN_IN), .A2(keyinput13), .B1(
        REG3_REG_21__SCAN_IN), .B2(keyinput8), .ZN(n4103) );
  OAI221_X1 U4744 ( .B1(REG2_REG_25__SCAN_IN), .B2(keyinput13), .C1(
        REG3_REG_21__SCAN_IN), .C2(keyinput8), .A(n4103), .ZN(n4110) );
  AOI22_X1 U4745 ( .A1(ADDR_REG_1__SCAN_IN), .A2(keyinput36), .B1(
        REG0_REG_18__SCAN_IN), .B2(keyinput40), .ZN(n4104) );
  OAI221_X1 U4746 ( .B1(ADDR_REG_1__SCAN_IN), .B2(keyinput36), .C1(
        REG0_REG_18__SCAN_IN), .C2(keyinput40), .A(n4104), .ZN(n4109) );
  AOI22_X1 U4747 ( .A1(DATAO_REG_29__SCAN_IN), .A2(keyinput4), .B1(
        REG2_REG_6__SCAN_IN), .B2(keyinput28), .ZN(n4105) );
  OAI221_X1 U4748 ( .B1(DATAO_REG_29__SCAN_IN), .B2(keyinput4), .C1(
        REG2_REG_6__SCAN_IN), .C2(keyinput28), .A(n4105), .ZN(n4108) );
  AOI22_X1 U4749 ( .A1(REG0_REG_0__SCAN_IN), .A2(keyinput12), .B1(
        REG3_REG_17__SCAN_IN), .B2(keyinput20), .ZN(n4106) );
  OAI221_X1 U4750 ( .B1(REG0_REG_0__SCAN_IN), .B2(keyinput12), .C1(
        REG3_REG_17__SCAN_IN), .C2(keyinput20), .A(n4106), .ZN(n4107) );
  NOR4_X1 U4751 ( .A1(n4110), .A2(n4109), .A3(n4108), .A4(n4107), .ZN(n4121)
         );
  AOI22_X1 U4752 ( .A1(REG2_REG_19__SCAN_IN), .A2(keyinput60), .B1(
        REG0_REG_26__SCAN_IN), .B2(keyinput15), .ZN(n4111) );
  OAI221_X1 U4753 ( .B1(REG2_REG_19__SCAN_IN), .B2(keyinput60), .C1(
        REG0_REG_26__SCAN_IN), .C2(keyinput15), .A(n4111), .ZN(n4119) );
  AOI22_X1 U4754 ( .A1(REG0_REG_4__SCAN_IN), .A2(keyinput35), .B1(
        REG2_REG_7__SCAN_IN), .B2(keyinput27), .ZN(n4112) );
  OAI221_X1 U4755 ( .B1(REG0_REG_4__SCAN_IN), .B2(keyinput35), .C1(
        REG2_REG_7__SCAN_IN), .C2(keyinput27), .A(n4112), .ZN(n4118) );
  AOI22_X1 U4756 ( .A1(DATAO_REG_17__SCAN_IN), .A2(keyinput48), .B1(
        DATAO_REG_22__SCAN_IN), .B2(keyinput39), .ZN(n4113) );
  OAI221_X1 U4757 ( .B1(DATAO_REG_17__SCAN_IN), .B2(keyinput48), .C1(
        DATAO_REG_22__SCAN_IN), .C2(keyinput39), .A(n4113), .ZN(n4117) );
  AOI22_X1 U4758 ( .A1(IR_REG_9__SCAN_IN), .A2(keyinput43), .B1(n4115), .B2(
        keyinput44), .ZN(n4114) );
  OAI221_X1 U4759 ( .B1(IR_REG_9__SCAN_IN), .B2(keyinput43), .C1(n4115), .C2(
        keyinput44), .A(n4114), .ZN(n4116) );
  NOR4_X1 U4760 ( .A1(n4119), .A2(n4118), .A3(n4117), .A4(n4116), .ZN(n4120)
         );
  NAND4_X1 U4761 ( .A1(n4123), .A2(n4122), .A3(n4121), .A4(n4120), .ZN(n4124)
         );
  NOR3_X1 U4762 ( .A1(n4126), .A2(n4125), .A3(n4124), .ZN(n4132) );
  AOI21_X1 U4763 ( .B1(n4569), .B2(n4128), .A(n4127), .ZN(n4129) );
  OAI21_X1 U4764 ( .B1(n4130), .B2(n4557), .A(n4129), .ZN(n4193) );
  MUX2_X1 U4765 ( .A(REG1_REG_26__SCAN_IN), .B(n4193), .S(n4590), .Z(n4131) );
  XOR2_X1 U4766 ( .A(n4132), .B(n4131), .Z(U3544) );
  AOI21_X1 U4767 ( .B1(n4134), .B2(n4554), .A(n4133), .ZN(n4194) );
  MUX2_X1 U4768 ( .A(n4135), .B(n4194), .S(n4590), .Z(n4136) );
  OAI21_X1 U4769 ( .B1(n4176), .B2(n4197), .A(n4136), .ZN(U3543) );
  INV_X1 U4770 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4139) );
  AOI21_X1 U4771 ( .B1(n4138), .B2(n4554), .A(n4137), .ZN(n4198) );
  MUX2_X1 U4772 ( .A(n4139), .B(n4198), .S(n4590), .Z(n4140) );
  OAI21_X1 U4773 ( .B1(n4176), .B2(n4201), .A(n4140), .ZN(U3542) );
  INV_X1 U4774 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4143) );
  AOI21_X1 U4775 ( .B1(n4142), .B2(n4554), .A(n4141), .ZN(n4202) );
  MUX2_X1 U4776 ( .A(n4143), .B(n4202), .S(n4590), .Z(n4144) );
  OAI21_X1 U4777 ( .B1(n4176), .B2(n4205), .A(n4144), .ZN(U3541) );
  NAND3_X1 U4778 ( .A1(n4146), .A2(n4569), .A3(n4145), .ZN(n4147) );
  OAI211_X1 U4779 ( .C1(n4149), .C2(n4557), .A(n4148), .B(n4147), .ZN(n4206)
         );
  MUX2_X1 U4780 ( .A(REG1_REG_22__SCAN_IN), .B(n4206), .S(n4590), .Z(U3540) );
  INV_X1 U4781 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4152) );
  AOI21_X1 U4782 ( .B1(n4151), .B2(n4554), .A(n4150), .ZN(n4207) );
  MUX2_X1 U4783 ( .A(n4152), .B(n4207), .S(n4590), .Z(n4153) );
  OAI21_X1 U4784 ( .B1(n4176), .B2(n4210), .A(n4153), .ZN(U3539) );
  AOI21_X1 U4785 ( .B1(n4155), .B2(n4554), .A(n4154), .ZN(n4211) );
  MUX2_X1 U4786 ( .A(n4156), .B(n4211), .S(n4590), .Z(n4157) );
  OAI21_X1 U4787 ( .B1(n4176), .B2(n4214), .A(n4157), .ZN(U3538) );
  INV_X1 U4788 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4160) );
  AOI21_X1 U4789 ( .B1(n4159), .B2(n4554), .A(n4158), .ZN(n4215) );
  MUX2_X1 U4790 ( .A(n4160), .B(n4215), .S(n4590), .Z(n4161) );
  OAI21_X1 U4791 ( .B1(n4176), .B2(n4218), .A(n4161), .ZN(U3537) );
  OAI211_X1 U4792 ( .C1(n4164), .C2(n4557), .A(n4163), .B(n4162), .ZN(n4219)
         );
  MUX2_X1 U4793 ( .A(REG1_REG_18__SCAN_IN), .B(n4219), .S(n4590), .Z(U3536) );
  AOI21_X1 U4794 ( .B1(n4166), .B2(n4554), .A(n4165), .ZN(n4220) );
  MUX2_X1 U4795 ( .A(n4167), .B(n4220), .S(n4590), .Z(n4168) );
  OAI21_X1 U4796 ( .B1(n4176), .B2(n4223), .A(n4168), .ZN(U3535) );
  AOI21_X1 U4797 ( .B1(n4170), .B2(n4554), .A(n4169), .ZN(n4224) );
  MUX2_X1 U4798 ( .A(n2173), .B(n4224), .S(n4590), .Z(n4171) );
  OAI21_X1 U4799 ( .B1(n4176), .B2(n4227), .A(n4171), .ZN(U3534) );
  AOI21_X1 U4800 ( .B1(n4554), .B2(n4173), .A(n4172), .ZN(n4228) );
  MUX2_X1 U4801 ( .A(n4174), .B(n4228), .S(n4590), .Z(n4175) );
  OAI21_X1 U4802 ( .B1(n4176), .B2(n4232), .A(n4175), .ZN(U3533) );
  NAND3_X1 U4803 ( .A1(n4178), .A2(n4177), .A3(n4569), .ZN(n4179) );
  OAI211_X1 U4804 ( .C1(n4181), .C2(n4563), .A(n4180), .B(n4179), .ZN(n4233)
         );
  MUX2_X1 U4805 ( .A(REG1_REG_14__SCAN_IN), .B(n4233), .S(n4590), .Z(U3532) );
  NAND2_X1 U4806 ( .A1(n4182), .A2(n4554), .ZN(n4184) );
  OAI211_X1 U4807 ( .C1(n4548), .C2(n4185), .A(n4184), .B(n4183), .ZN(n4234)
         );
  MUX2_X1 U4808 ( .A(REG1_REG_13__SCAN_IN), .B(n4234), .S(n4590), .Z(U3531) );
  INV_X1 U4809 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4186) );
  MUX2_X1 U4810 ( .A(n4248), .B(n4186), .S(n4570), .Z(n4187) );
  OAI21_X1 U4811 ( .B1(n4188), .B2(n4231), .A(n4187), .ZN(U3517) );
  INV_X1 U4812 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4189) );
  MUX2_X1 U4813 ( .A(n4252), .B(n4189), .S(n4570), .Z(n4190) );
  OAI21_X1 U4814 ( .B1(n4249), .B2(n4231), .A(n4190), .ZN(U3516) );
  MUX2_X1 U4815 ( .A(REG0_REG_29__SCAN_IN), .B(n4191), .S(n4572), .Z(U3515) );
  MUX2_X1 U4816 ( .A(REG0_REG_27__SCAN_IN), .B(n4192), .S(n4572), .Z(U3513) );
  MUX2_X1 U4817 ( .A(REG0_REG_26__SCAN_IN), .B(n4193), .S(n4572), .Z(U3512) );
  INV_X1 U4818 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4195) );
  MUX2_X1 U4819 ( .A(n4195), .B(n4194), .S(n4572), .Z(n4196) );
  OAI21_X1 U4820 ( .B1(n4197), .B2(n4231), .A(n4196), .ZN(U3511) );
  INV_X1 U4821 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4199) );
  MUX2_X1 U4822 ( .A(n4199), .B(n4198), .S(n4572), .Z(n4200) );
  OAI21_X1 U4823 ( .B1(n4201), .B2(n4231), .A(n4200), .ZN(U3510) );
  MUX2_X1 U4824 ( .A(n4203), .B(n4202), .S(n4572), .Z(n4204) );
  OAI21_X1 U4825 ( .B1(n4205), .B2(n4231), .A(n4204), .ZN(U3509) );
  MUX2_X1 U4826 ( .A(REG0_REG_22__SCAN_IN), .B(n4206), .S(n4572), .Z(U3508) );
  INV_X1 U4827 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4208) );
  MUX2_X1 U4828 ( .A(n4208), .B(n4207), .S(n4572), .Z(n4209) );
  OAI21_X1 U4829 ( .B1(n4210), .B2(n4231), .A(n4209), .ZN(U3507) );
  INV_X1 U4830 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4212) );
  MUX2_X1 U4831 ( .A(n4212), .B(n4211), .S(n4572), .Z(n4213) );
  OAI21_X1 U4832 ( .B1(n4214), .B2(n4231), .A(n4213), .ZN(U3506) );
  INV_X1 U4833 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4216) );
  MUX2_X1 U4834 ( .A(n4216), .B(n4215), .S(n4572), .Z(n4217) );
  OAI21_X1 U4835 ( .B1(n4218), .B2(n4231), .A(n4217), .ZN(U3505) );
  MUX2_X1 U4836 ( .A(REG0_REG_18__SCAN_IN), .B(n4219), .S(n4572), .Z(U3503) );
  MUX2_X1 U4837 ( .A(n4221), .B(n4220), .S(n4572), .Z(n4222) );
  OAI21_X1 U4838 ( .B1(n4223), .B2(n4231), .A(n4222), .ZN(U3501) );
  INV_X1 U4839 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4225) );
  MUX2_X1 U4840 ( .A(n4225), .B(n4224), .S(n4572), .Z(n4226) );
  OAI21_X1 U4841 ( .B1(n4227), .B2(n4231), .A(n4226), .ZN(U3499) );
  MUX2_X1 U4842 ( .A(n4229), .B(n4228), .S(n4572), .Z(n4230) );
  OAI21_X1 U4843 ( .B1(n4232), .B2(n4231), .A(n4230), .ZN(U3497) );
  MUX2_X1 U4844 ( .A(REG0_REG_14__SCAN_IN), .B(n4233), .S(n4572), .Z(U3495) );
  MUX2_X1 U4845 ( .A(REG0_REG_13__SCAN_IN), .B(n4234), .S(n4572), .Z(U3493) );
  MUX2_X1 U4846 ( .A(DATAI_30_), .B(n4235), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4847 ( .A(DATAI_28_), .B(n4236), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U4848 ( .A(n4237), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4849 ( .A(n2646), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4850 ( .A(n4238), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U4851 ( .A(n4239), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U4852 ( .A(n4240), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4853 ( .A(DATAI_20_), .B(n4241), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4854 ( .A(n4242), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4855 ( .A(n4300), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U4856 ( .A(DATAI_4_), .B(n4243), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4857 ( .A(n4244), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4858 ( .A(n4245), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  AOI22_X1 U4859 ( .A1(n4246), .A2(n4463), .B1(n4466), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4247) );
  OAI21_X1 U4860 ( .B1(n4466), .B2(n4248), .A(n4247), .ZN(U3260) );
  INV_X1 U4861 ( .A(n4249), .ZN(n4250) );
  AOI22_X1 U4862 ( .A1(n4250), .A2(n4463), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4466), .ZN(n4251) );
  OAI21_X1 U4863 ( .B1(n4466), .B2(n4252), .A(n4251), .ZN(U3261) );
  INV_X1 U4864 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4573) );
  AOI21_X1 U4865 ( .B1(n4573), .B2(n4254), .A(n4253), .ZN(n4255) );
  XOR2_X1 U4866 ( .A(n4255), .B(n2228), .Z(n4257) );
  AOI22_X1 U4867 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4402), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4256) );
  OAI21_X1 U4868 ( .B1(n4258), .B2(n4257), .A(n4256), .ZN(U3240) );
  AOI211_X1 U4869 ( .C1(n4261), .C2(n4260), .A(n4259), .B(n4270), .ZN(n4263)
         );
  AOI211_X1 U4870 ( .C1(n4402), .C2(ADDR_REG_5__SCAN_IN), .A(n4263), .B(n4262), 
        .ZN(n4268) );
  OAI211_X1 U4871 ( .C1(n4266), .C2(n4265), .A(n4345), .B(n4264), .ZN(n4267)
         );
  OAI211_X1 U4872 ( .C1(n4409), .C2(n4269), .A(n4268), .B(n4267), .ZN(U3245)
         );
  AOI211_X1 U4873 ( .C1(n4273), .C2(n4272), .A(n4271), .B(n4270), .ZN(n4275)
         );
  AOI211_X1 U4874 ( .C1(n4402), .C2(ADDR_REG_6__SCAN_IN), .A(n4275), .B(n4274), 
        .ZN(n4279) );
  OAI211_X1 U4875 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4277), .A(n4345), .B(n4276), 
        .ZN(n4278) );
  OAI211_X1 U4876 ( .C1(n4409), .C2(n4514), .A(n4279), .B(n4278), .ZN(U3246)
         );
  AOI22_X1 U4877 ( .A1(n4280), .A2(n4584), .B1(REG1_REG_7__SCAN_IN), .B2(n4512), .ZN(n4282) );
  OAI21_X1 U4878 ( .B1(n4283), .B2(n4282), .A(n4404), .ZN(n4281) );
  AOI21_X1 U4879 ( .B1(n4283), .B2(n4282), .A(n4281), .ZN(n4285) );
  AOI211_X1 U4880 ( .C1(n4402), .C2(ADDR_REG_7__SCAN_IN), .A(n4285), .B(n4284), 
        .ZN(n4290) );
  OAI211_X1 U4881 ( .C1(n4288), .C2(n4287), .A(n4345), .B(n4286), .ZN(n4289)
         );
  OAI211_X1 U4882 ( .C1(n4409), .C2(n4512), .A(n4290), .B(n4289), .ZN(U3247)
         );
  OAI211_X1 U4883 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4292), .A(n4345), .B(n4291), 
        .ZN(n4294) );
  NAND2_X1 U4884 ( .A1(n4294), .A2(n4293), .ZN(n4295) );
  AOI21_X1 U4885 ( .B1(n4402), .B2(ADDR_REG_8__SCAN_IN), .A(n4295), .ZN(n4299)
         );
  OAI211_X1 U4886 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4297), .A(n4404), .B(n4296), 
        .ZN(n4298) );
  OAI211_X1 U4887 ( .C1(n4409), .C2(n4510), .A(n4299), .B(n4298), .ZN(U3248)
         );
  INV_X1 U4888 ( .A(n4300), .ZN(n4309) );
  OAI211_X1 U4889 ( .C1(n4303), .C2(n4302), .A(n4404), .B(n4301), .ZN(n4308)
         );
  OAI211_X1 U4890 ( .C1(n4306), .C2(n4305), .A(n4345), .B(n4304), .ZN(n4307)
         );
  OAI211_X1 U4891 ( .C1(n4409), .C2(n4309), .A(n4308), .B(n4307), .ZN(n4310)
         );
  AOI211_X1 U4892 ( .C1(n4402), .C2(ADDR_REG_9__SCAN_IN), .A(n4311), .B(n4310), 
        .ZN(n4312) );
  INV_X1 U4893 ( .A(n4312), .ZN(U3249) );
  OAI211_X1 U4894 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4314), .A(n4404), .B(n4313), .ZN(n4318) );
  OAI211_X1 U4895 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4316), .A(n4345), .B(n4315), .ZN(n4317) );
  OAI211_X1 U4896 ( .C1(n4409), .C2(n4319), .A(n4318), .B(n4317), .ZN(n4320)
         );
  AOI211_X1 U4897 ( .C1(n4402), .C2(ADDR_REG_10__SCAN_IN), .A(n4321), .B(n4320), .ZN(n4322) );
  INV_X1 U4898 ( .A(n4322), .ZN(U3250) );
  OAI211_X1 U4899 ( .C1(n4325), .C2(n4324), .A(n4345), .B(n4323), .ZN(n4327)
         );
  NAND2_X1 U4900 ( .A1(n4327), .A2(n4326), .ZN(n4328) );
  AOI21_X1 U4901 ( .B1(n4402), .B2(ADDR_REG_11__SCAN_IN), .A(n4328), .ZN(n4333) );
  OAI211_X1 U4902 ( .C1(n4331), .C2(n4330), .A(n4404), .B(n4329), .ZN(n4332)
         );
  OAI211_X1 U4903 ( .C1(n4409), .C2(n4334), .A(n4333), .B(n4332), .ZN(U3251)
         );
  OAI211_X1 U4904 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4336), .A(n4345), .B(n4335), .ZN(n4338) );
  NAND2_X1 U4905 ( .A1(n4338), .A2(n4337), .ZN(n4339) );
  AOI21_X1 U4906 ( .B1(n4402), .B2(ADDR_REG_12__SCAN_IN), .A(n4339), .ZN(n4343) );
  OAI211_X1 U4907 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4341), .A(n4404), .B(n4340), .ZN(n4342) );
  OAI211_X1 U4908 ( .C1(n4409), .C2(n4504), .A(n4343), .B(n4342), .ZN(U3252)
         );
  AOI22_X1 U4909 ( .A1(REG2_REG_13__SCAN_IN), .A2(n4501), .B1(n4356), .B2(
        n4344), .ZN(n4348) );
  OAI21_X1 U4910 ( .B1(n4348), .B2(n4347), .A(n4345), .ZN(n4346) );
  AOI21_X1 U4911 ( .B1(n4348), .B2(n4347), .A(n4346), .ZN(n4349) );
  AOI211_X1 U4912 ( .C1(n4402), .C2(ADDR_REG_13__SCAN_IN), .A(n4350), .B(n4349), .ZN(n4355) );
  OAI211_X1 U4913 ( .C1(n4353), .C2(n4352), .A(n4404), .B(n4351), .ZN(n4354)
         );
  OAI211_X1 U4914 ( .C1(n4409), .C2(n4356), .A(n4355), .B(n4354), .ZN(U3253)
         );
  AOI211_X1 U4915 ( .C1(n4359), .C2(n4358), .A(n4357), .B(n4397), .ZN(n4362)
         );
  INV_X1 U4916 ( .A(n4360), .ZN(n4361) );
  AOI211_X1 U4917 ( .C1(n4402), .C2(ADDR_REG_14__SCAN_IN), .A(n4362), .B(n4361), .ZN(n4366) );
  OAI211_X1 U4918 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4364), .A(n4404), .B(n4363), .ZN(n4365) );
  OAI211_X1 U4919 ( .C1(n4409), .C2(n4367), .A(n4366), .B(n4365), .ZN(U3254)
         );
  AOI211_X1 U4920 ( .C1(n4370), .C2(n4369), .A(n4368), .B(n4397), .ZN(n4371)
         );
  AOI211_X1 U4921 ( .C1(n4402), .C2(ADDR_REG_15__SCAN_IN), .A(n4372), .B(n4371), .ZN(n4377) );
  OAI211_X1 U4922 ( .C1(n4375), .C2(n4374), .A(n4404), .B(n4373), .ZN(n4376)
         );
  OAI211_X1 U4923 ( .C1(n4409), .C2(n4498), .A(n4377), .B(n4376), .ZN(U3255)
         );
  INV_X1 U4924 ( .A(n4378), .ZN(n4383) );
  AOI221_X1 U4925 ( .B1(n4381), .B2(n4380), .C1(n4379), .C2(n4380), .A(n4397), 
        .ZN(n4382) );
  AOI211_X1 U4926 ( .C1(n4402), .C2(ADDR_REG_16__SCAN_IN), .A(n4383), .B(n4382), .ZN(n4387) );
  OAI221_X1 U4927 ( .B1(n4385), .B2(REG1_REG_16__SCAN_IN), .C1(n4385), .C2(
        n4384), .A(n4404), .ZN(n4386) );
  OAI211_X1 U4928 ( .C1(n4409), .C2(n4496), .A(n4387), .B(n4386), .ZN(U3256)
         );
  AOI221_X1 U4929 ( .B1(n4390), .B2(n4389), .C1(n4388), .C2(n4389), .A(n4397), 
        .ZN(n4391) );
  AOI211_X1 U4930 ( .C1(n4402), .C2(ADDR_REG_17__SCAN_IN), .A(n4392), .B(n4391), .ZN(n4396) );
  OAI221_X1 U4931 ( .B1(n4394), .B2(n2073), .C1(n4394), .C2(n4393), .A(n4404), 
        .ZN(n4395) );
  OAI211_X1 U4932 ( .C1(n4409), .C2(n4494), .A(n4396), .B(n4395), .ZN(U3257)
         );
  AOI211_X1 U4933 ( .C1(n4399), .C2(n4398), .A(n2063), .B(n4397), .ZN(n4400)
         );
  AOI211_X1 U4934 ( .C1(ADDR_REG_18__SCAN_IN), .C2(n4402), .A(n4401), .B(n4400), .ZN(n4408) );
  OAI211_X1 U4935 ( .C1(n4406), .C2(n4405), .A(n4404), .B(n4403), .ZN(n4407)
         );
  OAI211_X1 U4936 ( .C1(n4409), .C2(n4493), .A(n4408), .B(n4407), .ZN(U3258)
         );
  XOR2_X1 U4937 ( .A(n4416), .B(n4410), .Z(n4420) );
  AOI22_X1 U4938 ( .A1(n4412), .A2(n4411), .B1(n4424), .B2(n4446), .ZN(n4413)
         );
  OAI21_X1 U4939 ( .B1(n4414), .B2(n4472), .A(n4413), .ZN(n4419) );
  XOR2_X1 U4940 ( .A(n4416), .B(n4415), .Z(n4564) );
  NOR2_X1 U4941 ( .A1(n4564), .A2(n4417), .ZN(n4418) );
  AOI211_X1 U4942 ( .C1(n4420), .C2(n4469), .A(n4419), .B(n4418), .ZN(n4565)
         );
  AOI22_X1 U4943 ( .A1(n4421), .A2(n4458), .B1(REG2_REG_11__SCAN_IN), .B2(
        n4466), .ZN(n4427) );
  INV_X1 U4944 ( .A(n4564), .ZN(n4425) );
  AOI21_X1 U4945 ( .B1(n4424), .B2(n4423), .A(n4422), .ZN(n4568) );
  AOI22_X1 U4946 ( .A1(n4425), .A2(n4468), .B1(n4463), .B2(n4568), .ZN(n4426)
         );
  OAI211_X1 U4947 ( .C1(n4466), .C2(n4565), .A(n4427), .B(n4426), .ZN(U3279)
         );
  AOI22_X1 U4948 ( .A1(n4428), .A2(n4458), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4466), .ZN(n4433) );
  INV_X1 U4949 ( .A(n4429), .ZN(n4430) );
  AOI22_X1 U4950 ( .A1(n4431), .A2(n4468), .B1(n4463), .B2(n4430), .ZN(n4432)
         );
  OAI211_X1 U4951 ( .C1(n4466), .C2(n4434), .A(n4433), .B(n4432), .ZN(U3280)
         );
  AOI22_X1 U4952 ( .A1(n4435), .A2(n4458), .B1(REG2_REG_8__SCAN_IN), .B2(n4466), .ZN(n4441) );
  INV_X1 U4953 ( .A(n4436), .ZN(n4439) );
  INV_X1 U4954 ( .A(n4437), .ZN(n4438) );
  AOI22_X1 U4955 ( .A1(n4439), .A2(n4468), .B1(n4463), .B2(n4438), .ZN(n4440)
         );
  OAI211_X1 U4956 ( .C1(n4466), .C2(n4442), .A(n4441), .B(n4440), .ZN(U3282)
         );
  OR2_X1 U4957 ( .A1(n4452), .A2(n4443), .ZN(n4444) );
  AND2_X1 U4958 ( .A1(n4445), .A2(n4444), .ZN(n4526) );
  AOI22_X1 U4959 ( .A1(n2331), .A2(n4447), .B1(n4446), .B2(n4459), .ZN(n4448)
         );
  OAI21_X1 U4960 ( .B1(n4450), .B2(n4449), .A(n4448), .ZN(n4457) );
  NAND2_X1 U4961 ( .A1(n4452), .A2(n4451), .ZN(n4454) );
  AOI21_X1 U4962 ( .B1(n4455), .B2(n4454), .A(n4453), .ZN(n4456) );
  AOI211_X1 U4963 ( .C1(n4526), .C2(n4470), .A(n4457), .B(n4456), .ZN(n4523)
         );
  AOI22_X1 U4964 ( .A1(REG3_REG_1__SCAN_IN), .A2(n4458), .B1(
        REG2_REG_1__SCAN_IN), .B2(n4466), .ZN(n4465) );
  NAND2_X1 U4965 ( .A1(n4460), .A2(n4459), .ZN(n4461) );
  NAND2_X1 U4966 ( .A1(n2109), .A2(n4461), .ZN(n4522) );
  INV_X1 U4967 ( .A(n4522), .ZN(n4462) );
  AOI22_X1 U4968 ( .A1(n4463), .A2(n4462), .B1(n4526), .B2(n4468), .ZN(n4464)
         );
  OAI211_X1 U4969 ( .C1(n4466), .C2(n4523), .A(n4465), .B(n4464), .ZN(U3289)
         );
  INV_X1 U4970 ( .A(REG3_REG_0__SCAN_IN), .ZN(n4481) );
  AOI22_X1 U4971 ( .A1(n4468), .A2(n4520), .B1(REG2_REG_0__SCAN_IN), .B2(n4466), .ZN(n4480) );
  OAI21_X1 U4972 ( .B1(n4470), .B2(n4469), .A(n4520), .ZN(n4471) );
  OAI21_X1 U4973 ( .B1(n2708), .B2(n4472), .A(n4471), .ZN(n4518) );
  NOR2_X1 U4974 ( .A1(n4474), .A2(n4473), .ZN(n4519) );
  INV_X1 U4975 ( .A(n4519), .ZN(n4476) );
  NOR2_X1 U4976 ( .A1(n4476), .A2(n4475), .ZN(n4478) );
  OAI21_X1 U4977 ( .B1(n4518), .B2(n4478), .A(n4477), .ZN(n4479) );
  OAI211_X1 U4978 ( .C1(n4482), .C2(n4481), .A(n4480), .B(n4479), .ZN(U3290)
         );
  AND2_X1 U4979 ( .A1(D_REG_31__SCAN_IN), .A2(n4489), .ZN(U3291) );
  AND2_X1 U4980 ( .A1(D_REG_30__SCAN_IN), .A2(n4489), .ZN(U3292) );
  INV_X1 U4981 ( .A(n4489), .ZN(n4488) );
  NOR2_X1 U4982 ( .A1(n4488), .A2(n4483), .ZN(U3293) );
  AND2_X1 U4983 ( .A1(D_REG_28__SCAN_IN), .A2(n4489), .ZN(U3294) );
  AND2_X1 U4984 ( .A1(D_REG_27__SCAN_IN), .A2(n4489), .ZN(U3295) );
  AND2_X1 U4985 ( .A1(D_REG_26__SCAN_IN), .A2(n4489), .ZN(U3296) );
  AND2_X1 U4986 ( .A1(D_REG_25__SCAN_IN), .A2(n4489), .ZN(U3297) );
  AND2_X1 U4987 ( .A1(D_REG_24__SCAN_IN), .A2(n4489), .ZN(U3298) );
  AND2_X1 U4988 ( .A1(D_REG_23__SCAN_IN), .A2(n4489), .ZN(U3299) );
  NOR2_X1 U4989 ( .A1(n4488), .A2(n4484), .ZN(U3300) );
  NOR2_X1 U4990 ( .A1(n4488), .A2(n4485), .ZN(U3301) );
  AND2_X1 U4991 ( .A1(D_REG_20__SCAN_IN), .A2(n4489), .ZN(U3302) );
  AND2_X1 U4992 ( .A1(D_REG_19__SCAN_IN), .A2(n4489), .ZN(U3303) );
  NOR2_X1 U4993 ( .A1(n4488), .A2(n4486), .ZN(U3304) );
  AND2_X1 U4994 ( .A1(D_REG_17__SCAN_IN), .A2(n4489), .ZN(U3305) );
  AND2_X1 U4995 ( .A1(D_REG_16__SCAN_IN), .A2(n4489), .ZN(U3306) );
  AND2_X1 U4996 ( .A1(D_REG_15__SCAN_IN), .A2(n4489), .ZN(U3307) );
  AND2_X1 U4997 ( .A1(D_REG_14__SCAN_IN), .A2(n4489), .ZN(U3308) );
  AND2_X1 U4998 ( .A1(D_REG_13__SCAN_IN), .A2(n4489), .ZN(U3309) );
  AND2_X1 U4999 ( .A1(D_REG_12__SCAN_IN), .A2(n4489), .ZN(U3310) );
  AND2_X1 U5000 ( .A1(D_REG_11__SCAN_IN), .A2(n4489), .ZN(U3311) );
  AND2_X1 U5001 ( .A1(D_REG_10__SCAN_IN), .A2(n4489), .ZN(U3312) );
  AND2_X1 U5002 ( .A1(D_REG_9__SCAN_IN), .A2(n4489), .ZN(U3313) );
  AND2_X1 U5003 ( .A1(D_REG_8__SCAN_IN), .A2(n4489), .ZN(U3314) );
  AND2_X1 U5004 ( .A1(D_REG_7__SCAN_IN), .A2(n4489), .ZN(U3315) );
  AND2_X1 U5005 ( .A1(D_REG_6__SCAN_IN), .A2(n4489), .ZN(U3316) );
  AND2_X1 U5006 ( .A1(D_REG_5__SCAN_IN), .A2(n4489), .ZN(U3317) );
  AND2_X1 U5007 ( .A1(D_REG_4__SCAN_IN), .A2(n4489), .ZN(U3318) );
  NOR2_X1 U5008 ( .A1(n4488), .A2(n4487), .ZN(U3319) );
  AND2_X1 U5009 ( .A1(D_REG_2__SCAN_IN), .A2(n4489), .ZN(U3320) );
  OAI21_X1 U5010 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4490), .ZN(
        n4491) );
  INV_X1 U5011 ( .A(n4491), .ZN(U3329) );
  AOI22_X1 U5012 ( .A1(STATE_REG_SCAN_IN), .A2(n4493), .B1(n4492), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5013 ( .A1(STATE_REG_SCAN_IN), .A2(n4494), .B1(n2492), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5014 ( .A(DATAI_16_), .ZN(n4495) );
  AOI22_X1 U5015 ( .A1(STATE_REG_SCAN_IN), .A2(n4496), .B1(n4495), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5016 ( .A1(STATE_REG_SCAN_IN), .A2(n4498), .B1(n4497), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5017 ( .A1(U3149), .A2(n4499), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4500) );
  INV_X1 U5018 ( .A(n4500), .ZN(U3338) );
  OAI22_X1 U5019 ( .A1(U3149), .A2(n4501), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4502) );
  INV_X1 U5020 ( .A(n4502), .ZN(U3339) );
  AOI22_X1 U5021 ( .A1(STATE_REG_SCAN_IN), .A2(n4504), .B1(n4503), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5022 ( .A1(U3149), .A2(n4505), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4506) );
  INV_X1 U5023 ( .A(n4506), .ZN(U3341) );
  OAI22_X1 U5024 ( .A1(U3149), .A2(n4507), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4508) );
  INV_X1 U5025 ( .A(n4508), .ZN(U3342) );
  AOI22_X1 U5026 ( .A1(STATE_REG_SCAN_IN), .A2(n4510), .B1(n4509), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5027 ( .A(DATAI_7_), .ZN(n4511) );
  AOI22_X1 U5028 ( .A1(STATE_REG_SCAN_IN), .A2(n4512), .B1(n4511), .B2(U3149), 
        .ZN(U3345) );
  INV_X1 U5029 ( .A(DATAI_6_), .ZN(n4513) );
  AOI22_X1 U5030 ( .A1(STATE_REG_SCAN_IN), .A2(n4514), .B1(n4513), .B2(U3149), 
        .ZN(U3346) );
  OAI22_X1 U5031 ( .A1(U3149), .A2(n4515), .B1(DATAI_5_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4516) );
  INV_X1 U5032 ( .A(n4516), .ZN(U3347) );
  OAI22_X1 U5033 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4517) );
  INV_X1 U5034 ( .A(n4517), .ZN(U3352) );
  AOI211_X1 U5035 ( .C1(n4543), .C2(n4520), .A(n4519), .B(n4518), .ZN(n4574)
         );
  AOI22_X1 U5036 ( .A1(n4572), .A2(n4574), .B1(n4521), .B2(n4570), .ZN(U3467)
         );
  NOR2_X1 U5037 ( .A1(n4522), .A2(n4548), .ZN(n4525) );
  INV_X1 U5038 ( .A(n4523), .ZN(n4524) );
  AOI211_X1 U5039 ( .C1(n4526), .C2(n4543), .A(n4525), .B(n4524), .ZN(n4576)
         );
  INV_X1 U5040 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4527) );
  AOI22_X1 U5041 ( .A1(n4572), .A2(n4576), .B1(n4527), .B2(n4570), .ZN(U3469)
         );
  AND3_X1 U5042 ( .A1(n4529), .A2(n4569), .A3(n4528), .ZN(n4532) );
  INV_X1 U5043 ( .A(n4530), .ZN(n4531) );
  AOI211_X1 U5044 ( .C1(n4543), .C2(n4533), .A(n4532), .B(n4531), .ZN(n4577)
         );
  INV_X1 U5045 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4534) );
  AOI22_X1 U5046 ( .A1(n4572), .A2(n4577), .B1(n4534), .B2(n4570), .ZN(U3471)
         );
  AOI22_X1 U5047 ( .A1(n4536), .A2(n4543), .B1(n4569), .B2(n4535), .ZN(n4537)
         );
  AND2_X1 U5048 ( .A1(n4538), .A2(n4537), .ZN(n4579) );
  AOI22_X1 U5049 ( .A1(n4572), .A2(n4579), .B1(n4539), .B2(n4570), .ZN(U3473)
         );
  INV_X1 U5050 ( .A(n4540), .ZN(n4542) );
  AOI211_X1 U5051 ( .C1(n4544), .C2(n4543), .A(n4542), .B(n4541), .ZN(n4581)
         );
  INV_X1 U5052 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4545) );
  AOI22_X1 U5053 ( .A1(n4572), .A2(n4581), .B1(n4545), .B2(n4570), .ZN(U3475)
         );
  OAI21_X1 U5054 ( .B1(n4548), .B2(n4547), .A(n4546), .ZN(n4549) );
  AOI21_X1 U5055 ( .B1(n4550), .B2(n4554), .A(n4549), .ZN(n4583) );
  INV_X1 U5056 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4551) );
  AOI22_X1 U5057 ( .A1(n4572), .A2(n4583), .B1(n4551), .B2(n4570), .ZN(U3477)
         );
  AOI211_X1 U5058 ( .C1(n4555), .C2(n4554), .A(n4553), .B(n4552), .ZN(n4585)
         );
  AOI22_X1 U5059 ( .A1(n4572), .A2(n4585), .B1(n4556), .B2(n4570), .ZN(U3481)
         );
  NOR2_X1 U5060 ( .A1(n4558), .A2(n4557), .ZN(n4559) );
  AOI211_X1 U5061 ( .C1(n4569), .C2(n4561), .A(n4560), .B(n4559), .ZN(n4586)
         );
  INV_X1 U5062 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4562) );
  AOI22_X1 U5063 ( .A1(n4572), .A2(n4586), .B1(n4562), .B2(n4570), .ZN(U3485)
         );
  NOR2_X1 U5064 ( .A1(n4564), .A2(n4563), .ZN(n4567) );
  INV_X1 U5065 ( .A(n4565), .ZN(n4566) );
  AOI211_X1 U5066 ( .C1(n4569), .C2(n4568), .A(n4567), .B(n4566), .ZN(n4589)
         );
  INV_X1 U5067 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4571) );
  AOI22_X1 U5068 ( .A1(n4572), .A2(n4589), .B1(n4571), .B2(n4570), .ZN(U3489)
         );
  AOI22_X1 U5069 ( .A1(n4590), .A2(n4574), .B1(n4573), .B2(n4587), .ZN(U3518)
         );
  AOI22_X1 U5070 ( .A1(n4590), .A2(n4576), .B1(n4575), .B2(n4587), .ZN(U3519)
         );
  AOI22_X1 U5071 ( .A1(n4590), .A2(n4577), .B1(n2699), .B2(n4587), .ZN(U3520)
         );
  AOI22_X1 U5072 ( .A1(n4590), .A2(n4579), .B1(n4578), .B2(n4587), .ZN(U3521)
         );
  AOI22_X1 U5073 ( .A1(n4590), .A2(n4581), .B1(n4580), .B2(n4587), .ZN(U3522)
         );
  AOI22_X1 U5074 ( .A1(n4590), .A2(n4583), .B1(n4582), .B2(n4587), .ZN(U3523)
         );
  AOI22_X1 U5075 ( .A1(n4590), .A2(n4585), .B1(n4584), .B2(n4587), .ZN(U3525)
         );
  AOI22_X1 U5076 ( .A1(n4590), .A2(n4586), .B1(n3604), .B2(n4587), .ZN(U3527)
         );
  AOI22_X1 U5077 ( .A1(n4590), .A2(n4589), .B1(n4588), .B2(n4587), .ZN(U3529)
         );
  CLKBUF_X1 U2409 ( .A(n2337), .Z(n3412) );
  INV_X2 U2885 ( .A(n4477), .ZN(n4466) );
endmodule

