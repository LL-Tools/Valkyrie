

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361;

  NOR2_X2 U4877 ( .A1(n9755), .A2(n9635), .ZN(n9626) );
  NAND2_X1 U4878 ( .A1(n8736), .A2(n8719), .ZN(n8713) );
  NAND2_X1 U4879 ( .A1(n8305), .A2(n5725), .ZN(n9600) );
  XNOR2_X1 U4880 ( .A(n5548), .B(n5547), .ZN(n7683) );
  INV_X1 U4881 ( .A(n10006), .ZN(n10090) );
  CLKBUF_X2 U4883 ( .A(n6754), .Z(n6929) );
  INV_X1 U4884 ( .A(n7647), .ZN(n10076) );
  OR2_X1 U4885 ( .A1(n6570), .A2(n10194), .ZN(n8146) );
  NAND2_X1 U4886 ( .A1(n6023), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6047) );
  XNOR2_X1 U4887 ( .A(n5053), .B(n5052), .ZN(n6716) );
  NAND2_X1 U4888 ( .A1(n5244), .A2(n5243), .ZN(n8330) );
  NAND2_X1 U4889 ( .A1(n5242), .A2(n5241), .ZN(n5244) );
  NAND2_X1 U4890 ( .A1(n5884), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5886) );
  NOR2_X1 U4892 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5041) );
  INV_X1 U4893 ( .A(n4400), .ZN(n4382) );
  NAND2_X1 U4894 ( .A1(n9490), .A2(n7019), .ZN(n5823) );
  NAND2_X1 U4895 ( .A1(n5786), .A2(n7653), .ZN(n5815) );
  CLKBUF_X3 U4896 ( .A(n7033), .Z(n5192) );
  NAND2_X1 U4897 ( .A1(n8533), .A2(n10226), .ZN(n6445) );
  NOR2_X1 U4898 ( .A1(n5915), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U4899 ( .A1(n9419), .A2(n9421), .ZN(n9336) );
  NAND2_X1 U4900 ( .A1(n10016), .A2(n5365), .ZN(n5789) );
  NAND2_X1 U4901 ( .A1(n9989), .A2(n10006), .ZN(n5788) );
  INV_X1 U4902 ( .A(n8657), .ZN(n8367) );
  AND2_X1 U4903 ( .A1(n8408), .A2(n6667), .ZN(n4509) );
  INV_X1 U4904 ( .A(n8726), .ZN(n8496) );
  INV_X1 U4905 ( .A(n4373), .ZN(n4374) );
  INV_X1 U4906 ( .A(n8644), .ZN(n8633) );
  OR2_X1 U4907 ( .A1(n6373), .A2(n4760), .ZN(n6568) );
  NAND2_X1 U4908 ( .A1(n6511), .A2(n6496), .ZN(n8707) );
  OAI21_X1 U4909 ( .B1(n9443), .B2(n9327), .A(n9326), .ZN(n9328) );
  CLKBUF_X2 U4910 ( .A(n5397), .Z(n4388) );
  CLKBUF_X3 U4911 ( .A(n5674), .Z(n5690) );
  INV_X1 U4912 ( .A(n9474), .ZN(n9612) );
  CLKBUF_X2 U4913 ( .A(n6733), .Z(n4387) );
  INV_X1 U4914 ( .A(n5364), .ZN(n10016) );
  INV_X1 U4915 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5050) );
  NAND2_X1 U4916 ( .A1(n6288), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6317) );
  NAND2_X1 U4917 ( .A1(n9430), .A2(n9429), .ZN(n9434) );
  AND2_X1 U4918 ( .A1(n4628), .A2(n4627), .ZN(n8165) );
  AOI211_X1 U4919 ( .C1(n10106), .C2(n9750), .A(n9749), .B(n9748), .ZN(n9751)
         );
  AND2_X1 U4920 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9872), .ZN(n10345) );
  NAND2_X1 U4921 ( .A1(n6252), .A2(n6251), .ZN(n8666) );
  NAND2_X1 U4922 ( .A1(n8393), .A2(n6378), .ZN(n8893) );
  INV_X2 U4923 ( .A(n10033), .ZN(n10047) );
  INV_X1 U4924 ( .A(n6396), .ZN(n4373) );
  BUF_X1 U4925 ( .A(n5957), .Z(n6396) );
  AND2_X1 U4926 ( .A1(n5003), .A2(n4419), .ZN(n4372) );
  INV_X1 U4927 ( .A(n5397), .ZN(n5604) );
  OAI211_X4 U4928 ( .C1(n6257), .C2(P2_REG3_REG_3__SCAN_IN), .A(n5948), .B(
        n4502), .ZN(n8535) );
  AND2_X2 U4929 ( .A1(n4850), .A2(n4468), .ZN(n9951) );
  OAI21_X2 U4930 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10322), .ZN(n10320) );
  NAND2_X2 U4931 ( .A1(n7634), .A2(n5823), .ZN(n7552) );
  XNOR2_X2 U4932 ( .A(n5668), .B(n5667), .ZN(n9042) );
  INV_X2 U4933 ( .A(n4373), .ZN(n4375) );
  NAND2_X2 U4934 ( .A1(n9875), .A2(n9876), .ZN(n9877) );
  NAND2_X1 U4935 ( .A1(n5783), .A2(n8043), .ZN(n8044) );
  AOI21_X2 U4936 ( .B1(n4571), .B2(n4569), .A(n7982), .ZN(n8045) );
  CLKBUF_X1 U4937 ( .A(n6570), .Z(n4376) );
  NAND4_X1 U4939 ( .A1(n5925), .A2(n5924), .A3(n5923), .A4(n5922), .ZN(n6570)
         );
  NAND2_X2 U4940 ( .A1(n5929), .A2(n5928), .ZN(n8538) );
  INV_X1 U4941 ( .A(n5333), .ZN(n4378) );
  INV_X2 U4942 ( .A(n5333), .ZN(n4379) );
  INV_X1 U4943 ( .A(n5333), .ZN(n5347) );
  NAND2_X2 U4944 ( .A1(n4846), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5348) );
  NAND2_X2 U4945 ( .A1(n8191), .A2(n8190), .ZN(n8193) );
  NAND2_X2 U4946 ( .A1(n4946), .A2(n4945), .ZN(n8273) );
  INV_X1 U4947 ( .A(n6328), .ZN(n6374) );
  INV_X1 U4948 ( .A(n8532), .ZN(n7528) );
  NAND4_X2 U4949 ( .A1(n5999), .A2(n5998), .A3(n5997), .A4(n5996), .ZN(n8532)
         );
  OR2_X2 U4950 ( .A1(n8974), .A2(n8419), .ZN(n6544) );
  NOR2_X2 U4951 ( .A1(n6717), .A2(n6908), .ZN(n6754) );
  XNOR2_X2 U4952 ( .A(n6317), .B(n6316), .ZN(n6373) );
  NOR2_X2 U4953 ( .A1(n9599), .A2(n8306), .ZN(n9581) );
  NAND2_X2 U4954 ( .A1(n5566), .A2(n5565), .ZN(n9778) );
  OAI22_X2 U4955 ( .A1(n8258), .A2(n8257), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n8256), .ZN(n8259) );
  XNOR2_X2 U4956 ( .A(n5440), .B(n5439), .ZN(n9322) );
  XNOR2_X2 U4957 ( .A(n8379), .B(n4452), .ZN(n8918) );
  XOR2_X2 U4958 ( .A(n9874), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10344) );
  NOR2_X4 U4959 ( .A1(n10346), .A2(n9873), .ZN(n9874) );
  NAND2_X2 U4960 ( .A1(n6122), .A2(n6121), .ZN(n8980) );
  XNOR2_X2 U4961 ( .A(n5640), .B(n5639), .ZN(n8054) );
  OAI21_X2 U4962 ( .B1(n5610), .B2(n5609), .A(n5170), .ZN(n5640) );
  XNOR2_X2 U4963 ( .A(n5443), .B(n4407), .ZN(n7058) );
  INV_X2 U4964 ( .A(n8620), .ZN(n4760) );
  OAI21_X2 U4965 ( .B1(n5275), .B2(n4897), .A(n5148), .ZN(n5548) );
  OAI21_X2 U4966 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10319), .ZN(n10350) );
  NAND2_X1 U4967 ( .A1(n8310), .A2(n8309), .ZN(n9551) );
  AOI21_X1 U4968 ( .B1(n4740), .B2(n4741), .A(n4739), .ZN(n4738) );
  NAND2_X1 U4969 ( .A1(n8279), .A2(n8278), .ZN(n9594) );
  NAND2_X1 U4970 ( .A1(n9458), .A2(n6858), .ZN(n9382) );
  NAND2_X1 U4971 ( .A1(n6523), .A2(n6522), .ZN(n8644) );
  NAND2_X1 U4972 ( .A1(n6243), .A2(n6242), .ZN(n8930) );
  INV_X1 U4973 ( .A(n8666), .ZN(n8439) );
  NAND2_X1 U4974 ( .A1(n5579), .A2(n5578), .ZN(n9773) );
  NOR2_X2 U4975 ( .A1(n8080), .A2(n8997), .ZN(n8842) );
  AND2_X1 U4976 ( .A1(n5508), .A2(n5507), .ZN(n9809) );
  INV_X1 U4977 ( .A(n7887), .ZN(n4381) );
  NAND2_X1 U4978 ( .A1(n6444), .A2(n7884), .ZN(n7937) );
  NAND2_X1 U4979 ( .A1(n7933), .A2(n8532), .ZN(n6000) );
  NAND2_X2 U4980 ( .A1(n6428), .A2(n6445), .ZN(n7851) );
  NAND2_X1 U4981 ( .A1(n9994), .A2(n10017), .ZN(n7699) );
  NAND2_X1 U4982 ( .A1(n4568), .A2(n5789), .ZN(n10035) );
  INV_X4 U4983 ( .A(n6917), .ZN(n6947) );
  INV_X1 U4984 ( .A(n9487), .ZN(n9967) );
  INV_X1 U4985 ( .A(n8533), .ZN(n7958) );
  NAND2_X1 U4986 ( .A1(n5094), .A2(n5093), .ZN(n5393) );
  INV_X1 U4987 ( .A(n5313), .ZN(n5818) );
  NAND2_X1 U4988 ( .A1(n7801), .A2(n6434), .ZN(n6546) );
  NOR2_X1 U4989 ( .A1(n7217), .A2(n4966), .ZN(n7653) );
  INV_X2 U4990 ( .A(n10041), .ZN(n7554) );
  INV_X2 U4991 ( .A(n8535), .ZN(n7957) );
  INV_X2 U4992 ( .A(n9493), .ZN(n5553) );
  NAND2_X2 U4993 ( .A1(n6373), .A2(n6374), .ZN(n6567) );
  INV_X1 U4994 ( .A(n5262), .ZN(n8327) );
  NAND2_X1 U4995 ( .A1(n5226), .A2(n5222), .ZN(n5880) );
  CLKBUF_X2 U4996 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n10173) );
  INV_X2 U4997 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  AOI21_X1 U4998 ( .B1(n6669), .B2(n6670), .A(n6668), .ZN(n6672) );
  NAND2_X1 U4999 ( .A1(n8380), .A2(n4452), .ZN(n8381) );
  OR2_X1 U5000 ( .A1(n6665), .A2(n6666), .ZN(n4511) );
  NAND2_X1 U5001 ( .A1(n4737), .A2(n4738), .ZN(n6387) );
  NAND2_X1 U5002 ( .A1(n8652), .A2(n8651), .ZN(n8650) );
  NAND2_X1 U5003 ( .A1(n4918), .A2(n4916), .ZN(n9430) );
  NAND2_X1 U5004 ( .A1(n9382), .A2(n4919), .ZN(n4918) );
  AND2_X1 U5005 ( .A1(n8656), .A2(n4420), .ZN(n4742) );
  NAND2_X1 U5006 ( .A1(n8731), .A2(n6351), .ZN(n8720) );
  NOR2_X1 U5007 ( .A1(n9600), .A2(n4595), .ZN(n4594) );
  CLKBUF_X1 U5008 ( .A(n8747), .Z(n8766) );
  OAI21_X1 U5009 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10325), .ZN(n10323) );
  OAI21_X2 U5010 ( .B1(n8786), .B2(n6162), .A(n6161), .ZN(n8764) );
  NAND2_X1 U5011 ( .A1(n4983), .A2(n4982), .ZN(n9635) );
  CLKBUF_X1 U5012 ( .A(n8461), .Z(n4513) );
  NAND2_X1 U5013 ( .A1(n5670), .A2(n5669), .ZN(n9743) );
  AOI21_X1 U5014 ( .B1(n4412), .B2(n4919), .A(n4917), .ZN(n4916) );
  NAND2_X1 U5015 ( .A1(n6222), .A2(n6221), .ZN(n8940) );
  INV_X1 U5016 ( .A(n6877), .ZN(n4917) );
  NAND2_X1 U5017 ( .A1(n6211), .A2(n6210), .ZN(n8945) );
  NAND2_X1 U5018 ( .A1(n6168), .A2(n6167), .ZN(n8970) );
  NAND2_X2 U5019 ( .A1(n6156), .A2(n6155), .ZN(n8974) );
  XNOR2_X1 U5020 ( .A(n5573), .B(n5572), .ZN(n7753) );
  AND2_X2 U5021 ( .A1(n8842), .A2(n8846), .ZN(n8843) );
  MUX2_X1 U5022 ( .A(n5476), .B(n5475), .S(n6972), .Z(n5522) );
  NAND2_X1 U5023 ( .A1(n5555), .A2(n5554), .ZN(n9783) );
  NAND2_X1 U5024 ( .A1(n5281), .A2(n5280), .ZN(n9790) );
  NAND2_X1 U5025 ( .A1(n5152), .A2(n5151), .ZN(n5573) );
  NAND2_X1 U5026 ( .A1(n5144), .A2(n5143), .ZN(n5275) );
  NAND2_X1 U5027 ( .A1(n6065), .A2(n6064), .ZN(n9002) );
  OR2_X1 U5028 ( .A1(n7815), .A2(n7814), .ZN(n7813) );
  NAND2_X1 U5029 ( .A1(n6074), .A2(n6073), .ZN(n8134) );
  NAND2_X1 U5030 ( .A1(n5464), .A2(n5463), .ZN(n9816) );
  NAND2_X1 U5031 ( .A1(n4617), .A2(n6034), .ZN(n10263) );
  NAND2_X1 U5032 ( .A1(n5451), .A2(n5450), .ZN(n7815) );
  NAND2_X1 U5033 ( .A1(n5485), .A2(n5484), .ZN(n9819) );
  NAND2_X1 U5034 ( .A1(n4676), .A2(n5118), .ZN(n5461) );
  OAI21_X1 U5035 ( .B1(n9947), .B2(n8266), .A(n9348), .ZN(n4871) );
  NAND2_X1 U5036 ( .A1(n5418), .A2(n5417), .ZN(n9976) );
  NAND2_X1 U5037 ( .A1(n5115), .A2(n4677), .ZN(n4676) );
  NAND2_X1 U5038 ( .A1(n7147), .A2(n7146), .ZN(n7171) );
  NAND2_X1 U5039 ( .A1(n5391), .A2(n5390), .ZN(n9994) );
  AND2_X1 U5040 ( .A1(n4625), .A2(n4624), .ZN(n7147) );
  AND2_X2 U5041 ( .A1(n7066), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NAND2_X1 U5042 ( .A1(n4721), .A2(n5984), .ZN(n7854) );
  NAND2_X1 U5043 ( .A1(n5393), .A2(n5097), .ZN(n4899) );
  NAND2_X1 U5044 ( .A1(n5376), .A2(n5375), .ZN(n10006) );
  XNOR2_X1 U5045 ( .A(n5393), .B(n5392), .ZN(n7038) );
  CLKBUF_X1 U5046 ( .A(n7019), .Z(n10069) );
  NAND2_X1 U5047 ( .A1(n5869), .A2(n7754), .ZN(n7006) );
  NAND4_X1 U5048 ( .A1(n5317), .A2(n5316), .A3(n5315), .A4(n5314), .ZN(n7217)
         );
  AND2_X1 U5049 ( .A1(n5362), .A2(n4499), .ZN(n4498) );
  OAI211_X1 U5050 ( .C1(n5333), .C2(n7046), .A(n5332), .B(n5331), .ZN(n7553)
         );
  CLKBUF_X1 U5051 ( .A(n7852), .Z(n10282) );
  XNOR2_X1 U5052 ( .A(n5888), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6951) );
  CLKBUF_X1 U5053 ( .A(n6177), .Z(n6406) );
  NAND2_X1 U5054 ( .A1(n5887), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U5055 ( .A1(n5056), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U5056 ( .A1(n7110), .A2(n7111), .ZN(n9938) );
  NAND2_X1 U5057 ( .A1(n4385), .A2(n5192), .ZN(n6177) );
  NAND2_X1 U5058 ( .A1(n5322), .A2(n5192), .ZN(n5333) );
  NAND2_X1 U5059 ( .A1(n6362), .A2(n9040), .ZN(n7284) );
  XNOR2_X1 U5060 ( .A(n6324), .B(n6323), .ZN(n7917) );
  NAND2_X1 U5061 ( .A1(n5051), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U5062 ( .A1(n5875), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U5063 ( .A1(n5907), .A2(n5906), .ZN(n5975) );
  XNOR2_X1 U5064 ( .A(n5374), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7101) );
  NAND2_X1 U5065 ( .A1(n4551), .A2(n5049), .ZN(n5875) );
  NAND2_X1 U5066 ( .A1(n5921), .A2(n5920), .ZN(n9040) );
  XNOR2_X1 U5067 ( .A(n6319), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6328) );
  NAND2_X2 U5068 ( .A1(n7033), .A2(P1_U3084), .ZN(n7914) );
  INV_X1 U5069 ( .A(n5880), .ZN(n4551) );
  MUX2_X1 U5070 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5918), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5921) );
  MUX2_X1 U5071 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5229), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5233) );
  NAND2_X1 U5072 ( .A1(n9031), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4561) );
  NAND2_X1 U5073 ( .A1(n5243), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5238) );
  NAND2_X2 U5074 ( .A1(n4518), .A2(P1_U3084), .ZN(n8332) );
  NAND2_X1 U5075 ( .A1(n6318), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6319) );
  XNOR2_X1 U5076 ( .A(n5359), .B(n5358), .ZN(n9935) );
  NOR2_X1 U5077 ( .A1(n5372), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5388) );
  NAND2_X1 U5078 ( .A1(n5366), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U5079 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5240), .ZN(n5241) );
  MUX2_X1 U5080 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5309), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5311) );
  NOR2_X1 U5081 ( .A1(n9899), .A2(n9864), .ZN(n10316) );
  NOR2_X1 U5082 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5895) );
  INV_X1 U5083 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5052) );
  INV_X1 U5084 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5223) );
  INV_X1 U5085 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6116) );
  INV_X1 U5086 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5885) );
  INV_X1 U5087 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5898) );
  NOR2_X1 U5088 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5047) );
  NOR2_X1 U5089 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5046) );
  NOR2_X1 U5090 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5045) );
  INV_X4 U5091 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X2 U5092 ( .A1(n5035), .A2(n9731), .ZN(n9560) );
  XNOR2_X2 U5093 ( .A(n4997), .B(n5313), .ZN(n7650) );
  OR2_X2 U5094 ( .A1(n10146), .A2(n6574), .ZN(n7801) );
  NAND2_X1 U5095 ( .A1(n6376), .A2(n4760), .ZN(n4383) );
  NAND2_X1 U5096 ( .A1(n6376), .A2(n4760), .ZN(n4384) );
  NAND2_X2 U5097 ( .A1(n6376), .A2(n4760), .ZN(n8351) );
  AND4_X2 U5098 ( .A1(n5405), .A2(n5404), .A3(n5403), .A4(n5402), .ZN(n9988)
         );
  NAND2_X2 U5099 ( .A1(n6362), .A2(n9040), .ZN(n4385) );
  OR2_X2 U5100 ( .A1(n8698), .A2(n8697), .ZN(n8700) );
  XNOR2_X2 U5101 ( .A(n6321), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8620) );
  BUF_X1 U5102 ( .A(n8948), .Z(n4386) );
  INV_X4 U5103 ( .A(n6758), .ZN(n6917) );
  AOI21_X2 U5104 ( .B1(n6387), .B2(n6557), .A(n6386), .ZN(n8380) );
  NAND2_X1 U5105 ( .A1(n4537), .A2(n7006), .ZN(n6733) );
  OAI21_X2 U5106 ( .B1(n8058), .B2(n8063), .A(n6031), .ZN(n8101) );
  OAI211_X2 U5107 ( .C1(n4805), .C2(n4381), .A(n4803), .B(n6014), .ZN(n8058)
         );
  AOI22_X2 U5108 ( .A1(n8038), .A2(n8037), .B1(n8036), .B2(n9482), .ZN(n8191)
         );
  OAI22_X2 U5109 ( .A1(n7979), .A2(n7978), .B1(n8005), .B2(n9483), .ZN(n8038)
         );
  NOR2_X1 U5110 ( .A1(n4591), .A2(n5007), .ZN(n4589) );
  INV_X1 U5111 ( .A(n4592), .ZN(n4591) );
  INV_X1 U5112 ( .A(n5575), .ZN(n5161) );
  NAND2_X1 U5113 ( .A1(n6279), .A2(n6278), .ZN(n6288) );
  INV_X1 U5114 ( .A(n6318), .ZN(n6279) );
  AOI21_X1 U5115 ( .B1(n4910), .B2(n4901), .A(n4909), .ZN(n4900) );
  INV_X1 U5116 ( .A(n6896), .ZN(n4901) );
  OAI211_X1 U5117 ( .C1(n5215), .C2(n5214), .A(n5213), .B(n5212), .ZN(n5249)
         );
  NAND2_X1 U5118 ( .A1(n5215), .A2(n5211), .ZN(n5258) );
  NAND2_X1 U5119 ( .A1(n5460), .A2(n5124), .ZN(n4879) );
  NOR2_X2 U5120 ( .A1(n8386), .A2(n8914), .ZN(n8628) );
  MUX2_X1 U5121 ( .A(n6427), .B(n6426), .S(n4382), .Z(n6447) );
  AOI21_X1 U5122 ( .B1(n5622), .B2(n5621), .A(n5011), .ZN(n5628) );
  OAI21_X1 U5123 ( .B1(n5763), .B2(n5779), .A(n5778), .ZN(n5755) );
  INV_X1 U5124 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4795) );
  AOI21_X1 U5125 ( .B1(n4594), .B2(n8304), .A(n5012), .ZN(n4592) );
  NAND2_X1 U5126 ( .A1(n5777), .A2(n8305), .ZN(n5012) );
  INV_X1 U5127 ( .A(n4594), .ZN(n4593) );
  AND2_X1 U5128 ( .A1(n5785), .A2(n7736), .ZN(n7706) );
  NAND2_X1 U5129 ( .A1(n5696), .A2(n5196), .ZN(n5215) );
  AND2_X1 U5130 ( .A1(n5697), .A2(n5695), .ZN(n5196) );
  NOR2_X1 U5131 ( .A1(n4688), .A2(n4683), .ZN(n4682) );
  INV_X1 U5132 ( .A(n5143), .ZN(n4683) );
  INV_X1 U5133 ( .A(n4689), .ZN(n4688) );
  NAND2_X1 U5134 ( .A1(n6650), .A2(n6651), .ZN(n4781) );
  NOR2_X1 U5135 ( .A1(n4517), .A2(n4414), .ZN(n4516) );
  NOR2_X1 U5136 ( .A1(n4659), .A2(n4658), .ZN(n4657) );
  NOR2_X1 U5137 ( .A1(n4660), .A2(n7410), .ZN(n4658) );
  INV_X1 U5138 ( .A(n7414), .ZN(n4659) );
  OR2_X1 U5139 ( .A1(n8919), .A2(n6710), .ZN(n6526) );
  NAND2_X1 U5140 ( .A1(n4755), .A2(n4753), .ZN(n8685) );
  AND2_X1 U5141 ( .A1(n6352), .A2(n4754), .ZN(n4753) );
  INV_X1 U5142 ( .A(n4821), .ZN(n4819) );
  OAI21_X1 U5143 ( .B1(n8791), .B2(n4747), .A(n4745), .ZN(n8747) );
  INV_X1 U5144 ( .A(n4748), .ZN(n4747) );
  AND2_X1 U5145 ( .A1(n6346), .A2(n4746), .ZN(n4745) );
  NAND2_X1 U5146 ( .A1(n4748), .A2(n6420), .ZN(n4746) );
  NAND2_X1 U5147 ( .A1(n8639), .A2(n6380), .ZN(n8386) );
  INV_X1 U5148 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U5149 ( .A1(n9370), .A2(n9337), .ZN(n4520) );
  XNOR2_X1 U5150 ( .A(n6759), .B(n6945), .ZN(n7583) );
  INV_X1 U5151 ( .A(n4905), .ZN(n4904) );
  OAI21_X1 U5152 ( .B1(n9362), .B2(n4909), .A(n6914), .ZN(n4905) );
  INV_X1 U5153 ( .A(n4910), .ZN(n4902) );
  NOR2_X1 U5154 ( .A1(n5273), .A2(n5272), .ZN(n5769) );
  AND2_X1 U5155 ( .A1(n8323), .A2(n8322), .ZN(n5806) );
  NOR2_X1 U5156 ( .A1(n4951), .A2(n4403), .ZN(n4949) );
  NAND2_X1 U5157 ( .A1(n9783), .A2(n9696), .ZN(n4954) );
  OR2_X1 U5158 ( .A1(n9783), .A2(n8240), .ZN(n5781) );
  OR2_X1 U5159 ( .A1(n9804), .A2(n9481), .ZN(n8192) );
  AND2_X1 U5160 ( .A1(n4372), .A2(n7983), .ZN(n4569) );
  NAND2_X1 U5161 ( .A1(n7735), .A2(n7706), .ZN(n7812) );
  AND2_X1 U5162 ( .A1(n5364), .A2(n10082), .ZN(n5001) );
  NAND2_X1 U5163 ( .A1(n7561), .A2(n7560), .ZN(n9982) );
  AND2_X1 U5164 ( .A1(n7910), .A2(n7754), .ZN(n6971) );
  NAND2_X1 U5165 ( .A1(n4691), .A2(n4695), .ZN(n5682) );
  AOI21_X1 U5166 ( .B1(n4699), .B2(n4697), .A(n4696), .ZN(n4695) );
  INV_X1 U5167 ( .A(n5667), .ZN(n4696) );
  AOI21_X1 U5168 ( .B1(n4877), .B2(n4876), .A(n4875), .ZN(n4874) );
  INV_X1 U5169 ( .A(n5129), .ZN(n4875) );
  INV_X1 U5170 ( .A(n5124), .ZN(n4876) );
  NAND2_X1 U5171 ( .A1(n4507), .A2(n5020), .ZN(n5115) );
  NAND2_X1 U5172 ( .A1(n5426), .A2(n4508), .ZN(n4507) );
  AND2_X1 U5173 ( .A1(n5441), .A2(n5425), .ZN(n4508) );
  AND2_X1 U5174 ( .A1(n8448), .A2(n6641), .ZN(n4533) );
  INV_X1 U5175 ( .A(n6373), .ZN(n6354) );
  INV_X1 U5176 ( .A(n10175), .ZN(n8904) );
  INV_X1 U5177 ( .A(n6523), .ZN(n4739) );
  AOI21_X1 U5178 ( .B1(n8644), .B2(n4799), .A(n4442), .ZN(n4798) );
  INV_X1 U5179 ( .A(n6253), .ZN(n4799) );
  NAND2_X1 U5180 ( .A1(n6526), .A2(n6525), .ZN(n6385) );
  OR2_X1 U5181 ( .A1(n8950), .A2(n8427), .ZN(n8696) );
  OR2_X1 U5182 ( .A1(n8963), .A2(n8428), .ZN(n6497) );
  AND2_X2 U5183 ( .A1(n6502), .A2(n6497), .ZN(n8759) );
  OR2_X1 U5184 ( .A1(n10269), .A2(n6328), .ZN(n8903) );
  NAND2_X1 U5185 ( .A1(n6389), .A2(n6388), .ZN(n8914) );
  NAND2_X1 U5186 ( .A1(n6312), .A2(n10186), .ZN(n10175) );
  INV_X1 U5187 ( .A(n7281), .ZN(n6312) );
  XNOR2_X1 U5188 ( .A(n5914), .B(n5913), .ZN(n6362) );
  OR2_X1 U5189 ( .A1(n5919), .A2(n6283), .ZN(n5914) );
  NOR2_X1 U5190 ( .A1(n6288), .A2(n6281), .ZN(n6285) );
  AND2_X1 U5191 ( .A1(n6895), .A2(n9361), .ZN(n6896) );
  AND2_X1 U5192 ( .A1(n9358), .A2(n6890), .ZN(n4477) );
  CLKBUF_X1 U5193 ( .A(n5339), .Z(n4480) );
  BUF_X1 U5194 ( .A(n6715), .Z(n7001) );
  AND2_X1 U5195 ( .A1(n9931), .A2(n9930), .ZN(n9934) );
  NAND2_X1 U5196 ( .A1(n4863), .A2(n4866), .ZN(n4858) );
  NOR2_X1 U5197 ( .A1(n4861), .A2(n4860), .ZN(n4859) );
  NAND2_X1 U5198 ( .A1(n9528), .A2(n4852), .ZN(n4851) );
  INV_X1 U5199 ( .A(n8251), .ZN(n4852) );
  AOI21_X1 U5200 ( .B1(n4397), .B2(n4942), .A(n4439), .ZN(n4939) );
  NAND2_X1 U5201 ( .A1(n4941), .A2(n4942), .ZN(n4940) );
  INV_X1 U5202 ( .A(n8276), .ZN(n4941) );
  OR2_X1 U5203 ( .A1(n4439), .A2(n8276), .ZN(n9623) );
  NOR2_X1 U5204 ( .A1(n4985), .A2(n9758), .ZN(n4982) );
  INV_X1 U5205 ( .A(n8267), .ZN(n8270) );
  INV_X1 U5206 ( .A(n5361), .ZN(n5528) );
  INV_X1 U5207 ( .A(n10119), .ZN(n10106) );
  XNOR2_X1 U5208 ( .A(n5220), .B(n5219), .ZN(n9030) );
  NAND2_X1 U5209 ( .A1(n5217), .A2(n5216), .ZN(n5220) );
  NAND2_X1 U5210 ( .A1(n5863), .A2(n5862), .ZN(n6999) );
  OR2_X1 U5211 ( .A1(n5861), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n5862) );
  XNOR2_X1 U5212 ( .A(n5597), .B(n5596), .ZN(n7912) );
  INV_X1 U5213 ( .A(n8519), .ZN(n10153) );
  NAND2_X1 U5214 ( .A1(n4606), .A2(n7917), .ZN(n6563) );
  NAND2_X1 U5215 ( .A1(n4609), .A2(n4418), .ZN(n4608) );
  INV_X1 U5216 ( .A(n9462), .ZN(n9437) );
  NAND2_X1 U5217 ( .A1(n4843), .A2(n4847), .ZN(n9909) );
  NAND2_X1 U5218 ( .A1(n9906), .A2(n9905), .ZN(n4847) );
  NOR2_X1 U5219 ( .A1(n7263), .A2(n4629), .ZN(n7673) );
  NOR2_X1 U5220 ( .A1(n7267), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4629) );
  MUX2_X1 U5221 ( .A(n6437), .B(n6436), .S(n4400), .Z(n6439) );
  INV_X1 U5222 ( .A(n6444), .ZN(n4711) );
  NOR2_X1 U5223 ( .A1(n7884), .A2(n4382), .ZN(n4709) );
  INV_X1 U5224 ( .A(n4614), .ZN(n4613) );
  OAI21_X1 U5225 ( .B1(n6509), .B2(n8719), .A(n6507), .ZN(n4614) );
  INV_X1 U5226 ( .A(n6516), .ZN(n4616) );
  INV_X1 U5227 ( .A(n4602), .ZN(n4601) );
  OAI21_X1 U5228 ( .B1(n8651), .B2(n4603), .A(n4382), .ZN(n4602) );
  NAND2_X1 U5229 ( .A1(n4393), .A2(n8669), .ZN(n4603) );
  NAND2_X1 U5230 ( .A1(n8102), .A2(n6552), .ZN(n4558) );
  INV_X1 U5231 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n9075) );
  AOI21_X1 U5232 ( .B1(n5627), .B2(n6972), .A(n4885), .ZN(n4884) );
  NAND2_X1 U5233 ( .A1(n8300), .A2(n4886), .ZN(n4885) );
  INV_X1 U5234 ( .A(n5666), .ZN(n4887) );
  NOR2_X1 U5235 ( .A1(n9641), .A2(n5011), .ZN(n5010) );
  INV_X1 U5236 ( .A(n5148), .ZN(n4687) );
  NOR2_X1 U5237 ( .A1(n4427), .A2(n4896), .ZN(n4895) );
  INV_X1 U5238 ( .A(n5151), .ZN(n4896) );
  AND2_X1 U5239 ( .A1(n4690), .A2(n5149), .ZN(n4689) );
  NAND2_X1 U5240 ( .A1(n4897), .A2(n5148), .ZN(n4690) );
  NAND2_X1 U5241 ( .A1(n5287), .A2(n5286), .ZN(n5144) );
  INV_X1 U5242 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5138) );
  INV_X1 U5243 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4824) );
  INV_X1 U5244 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4827) );
  INV_X1 U5245 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4826) );
  INV_X1 U5246 ( .A(n6628), .ZN(n4786) );
  NAND2_X1 U5247 ( .A1(n4536), .A2(n4535), .ZN(n4534) );
  NAND2_X1 U5248 ( .A1(n6652), .A2(n6653), .ZN(n4535) );
  NAND2_X2 U5249 ( .A1(n4759), .A2(n6569), .ZN(n6589) );
  INV_X1 U5250 ( .A(n8352), .ZN(n6673) );
  NAND2_X1 U5251 ( .A1(n8633), .A2(n4394), .ZN(n4720) );
  INV_X1 U5252 ( .A(n5958), .ZN(n5995) );
  INV_X1 U5253 ( .A(n8565), .ZN(n4660) );
  INV_X1 U5254 ( .A(n7489), .ZN(n4663) );
  NOR2_X1 U5255 ( .A1(n7468), .A2(n4665), .ZN(n4664) );
  INV_X1 U5256 ( .A(n7464), .ZN(n4665) );
  NAND2_X1 U5257 ( .A1(n4674), .A2(n8657), .ZN(n6523) );
  NOR2_X2 U5258 ( .A1(n8671), .A2(n8930), .ZN(n4494) );
  NOR2_X1 U5259 ( .A1(n8940), .A2(n8945), .ZN(n4831) );
  AND2_X1 U5260 ( .A1(n6512), .A2(n6516), .ZN(n6542) );
  NAND2_X1 U5261 ( .A1(n6497), .A2(n8732), .ZN(n4756) );
  NAND2_X1 U5262 ( .A1(n4836), .A2(n4835), .ZN(n4834) );
  NOR2_X1 U5263 ( .A1(n8980), .A2(n8984), .ZN(n4836) );
  AND2_X1 U5264 ( .A1(n7964), .A2(n4815), .ZN(n4809) );
  NOR2_X1 U5265 ( .A1(n8114), .A2(n4840), .ZN(n4839) );
  AND2_X1 U5266 ( .A1(n6335), .A2(n6445), .ZN(n4734) );
  INV_X1 U5267 ( .A(n7851), .ZN(n6548) );
  NAND2_X1 U5268 ( .A1(n7917), .A2(n6328), .ZN(n6569) );
  INV_X1 U5269 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U5270 ( .A1(n6289), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6309) );
  INV_X1 U5271 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U5272 ( .A1(n6277), .A2(n6276), .ZN(n6318) );
  INV_X1 U5273 ( .A(n7240), .ZN(n4915) );
  NAND2_X1 U5274 ( .A1(n6896), .A2(n4405), .ZN(n4906) );
  INV_X1 U5275 ( .A(n9429), .ZN(n4541) );
  AND2_X1 U5276 ( .A1(n6907), .A2(n6906), .ZN(n6914) );
  NAND2_X1 U5277 ( .A1(n4547), .A2(n6844), .ZN(n4546) );
  INV_X1 U5278 ( .A(n6841), .ZN(n4547) );
  NAND2_X1 U5279 ( .A1(n4413), .A2(n4548), .ZN(n4543) );
  INV_X1 U5280 ( .A(n6844), .ZN(n4548) );
  AOI211_X1 U5281 ( .C1(n5772), .C2(n5771), .A(n7913), .B(n5806), .ZN(n5813)
         );
  INV_X1 U5282 ( .A(n5806), .ZN(n5852) );
  OR2_X1 U5283 ( .A1(n7180), .A2(n4864), .ZN(n4863) );
  INV_X1 U5284 ( .A(n4867), .ZN(n4864) );
  OR2_X1 U5285 ( .A1(n9731), .A2(n8313), .ZN(n5774) );
  AND2_X1 U5286 ( .A1(n5775), .A2(n9550), .ZN(n8309) );
  NOR2_X1 U5287 ( .A1(n9739), .A2(n4974), .ZN(n4973) );
  INV_X1 U5288 ( .A(n4975), .ZN(n4974) );
  INV_X1 U5289 ( .A(n8303), .ZN(n4595) );
  NAND2_X1 U5290 ( .A1(n8298), .A2(n5010), .ZN(n5009) );
  NOR2_X1 U5291 ( .A1(n8295), .A2(n4583), .ZN(n4582) );
  AND2_X1 U5292 ( .A1(n9773), .A2(n9666), .ZN(n8295) );
  OR2_X1 U5293 ( .A1(n4971), .A2(n9795), .ZN(n4968) );
  OR2_X1 U5294 ( .A1(n9790), .A2(n9798), .ZN(n4971) );
  OR2_X1 U5295 ( .A1(n9816), .A2(n9483), .ZN(n7983) );
  NAND2_X1 U5296 ( .A1(n10120), .A2(n4981), .ZN(n4980) );
  OR2_X1 U5297 ( .A1(n7747), .A2(n9967), .ZN(n5785) );
  OR2_X1 U5298 ( .A1(n9976), .A2(n7739), .ZN(n7736) );
  NAND2_X1 U5299 ( .A1(n10105), .A2(n9988), .ZN(n9969) );
  AND2_X1 U5300 ( .A1(n5789), .A2(n5825), .ZN(n4999) );
  NAND2_X1 U5301 ( .A1(n10041), .A2(n7647), .ZN(n5825) );
  NAND2_X1 U5302 ( .A1(n4997), .A2(n5313), .ZN(n5816) );
  NAND2_X1 U5303 ( .A1(n6716), .A2(n6971), .ZN(n7007) );
  AND2_X1 U5304 ( .A1(n5777), .A2(n5776), .ZN(n8307) );
  OR2_X1 U5305 ( .A1(n7016), .A2(n6973), .ZN(n7191) );
  OAI21_X1 U5306 ( .B1(n5875), .B2(n5874), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5876) );
  NAND2_X1 U5307 ( .A1(n5177), .A2(n5176), .ZN(n5630) );
  AOI21_X1 U5308 ( .B1(n4446), .B2(n4874), .A(n4399), .ZN(n4873) );
  INV_X1 U5309 ( .A(SI_12_), .ZN(n5120) );
  XNOR2_X1 U5310 ( .A(n5116), .B(SI_11_), .ZN(n5477) );
  NAND2_X1 U5311 ( .A1(n4899), .A2(n4898), .ZN(n5426) );
  AND2_X1 U5312 ( .A1(n5104), .A2(n5099), .ZN(n4898) );
  NAND2_X1 U5313 ( .A1(n5092), .A2(n4404), .ZN(n5093) );
  NAND2_X1 U5314 ( .A1(n4775), .A2(n4781), .ZN(n4774) );
  NAND2_X1 U5315 ( .A1(n6123), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6139) );
  AND2_X1 U5316 ( .A1(n8533), .A2(n8351), .ZN(n6591) );
  NOR2_X1 U5317 ( .A1(n4534), .A2(n4778), .ZN(n4770) );
  INV_X1 U5318 ( .A(n4534), .ZN(n8415) );
  OR2_X1 U5319 ( .A1(n6645), .A2(n6644), .ZN(n6646) );
  NAND2_X1 U5320 ( .A1(n8425), .A2(n8424), .ZN(n8490) );
  AND2_X1 U5321 ( .A1(n7518), .A2(n6597), .ZN(n4792) );
  INV_X1 U5322 ( .A(n7917), .ZN(n6561) );
  NAND2_X1 U5323 ( .A1(n8077), .A2(n4553), .ZN(n6554) );
  NOR2_X1 U5324 ( .A1(n4554), .A2(n8809), .ZN(n4553) );
  NAND2_X1 U5325 ( .A1(n4555), .A2(n8857), .ZN(n4554) );
  NOR2_X1 U5326 ( .A1(n8835), .A2(n4556), .ZN(n4555) );
  NOR2_X1 U5327 ( .A1(n6558), .A2(n4563), .ZN(n4562) );
  NOR2_X1 U5328 ( .A1(n4565), .A2(n8707), .ZN(n4564) );
  INV_X1 U5329 ( .A(n6559), .ZN(n4567) );
  INV_X1 U5330 ( .A(n4657), .ZN(n4655) );
  OR2_X1 U5331 ( .A1(n7453), .A2(n7452), .ZN(n7450) );
  OR2_X1 U5332 ( .A1(n7778), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7780) );
  NOR2_X1 U5333 ( .A1(n8595), .A2(n8610), .ZN(n8608) );
  NAND2_X1 U5334 ( .A1(n6394), .A2(n6393), .ZN(n8627) );
  NAND2_X1 U5335 ( .A1(n4634), .A2(n4433), .ZN(n8378) );
  NAND2_X1 U5336 ( .A1(n8650), .A2(n4798), .ZN(n4634) );
  NAND2_X1 U5337 ( .A1(n4798), .A2(n8633), .ZN(n4797) );
  OR2_X1 U5338 ( .A1(n8930), .A2(n8666), .ZN(n6253) );
  NAND2_X1 U5339 ( .A1(n4743), .A2(n4742), .ZN(n8654) );
  NAND2_X1 U5340 ( .A1(n8668), .A2(n6241), .ZN(n8652) );
  OR2_X1 U5341 ( .A1(n8673), .A2(n8689), .ZN(n6241) );
  NOR2_X1 U5342 ( .A1(n8713), .A2(n4829), .ZN(n8680) );
  INV_X1 U5343 ( .A(n4831), .ZN(n4829) );
  NOR2_X1 U5344 ( .A1(n8713), .A2(n8945), .ZN(n6370) );
  AOI21_X2 U5345 ( .B1(n4406), .B2(n8764), .A(n4479), .ZN(n8712) );
  NAND2_X1 U5346 ( .A1(n4636), .A2(n4637), .ZN(n4479) );
  AOI21_X1 U5347 ( .B1(n4817), .B2(n6197), .A(n6196), .ZN(n4637) );
  INV_X1 U5348 ( .A(n4638), .ZN(n4635) );
  OR2_X1 U5349 ( .A1(n8970), .A2(n8779), .ZN(n4821) );
  NOR2_X1 U5350 ( .A1(n8759), .A2(n4819), .ZN(n4818) );
  OR2_X1 U5351 ( .A1(n8764), .A2(n6176), .ZN(n4820) );
  AND2_X1 U5352 ( .A1(n8747), .A2(n6348), .ZN(n8750) );
  NAND2_X1 U5353 ( .A1(n4749), .A2(n6544), .ZN(n4748) );
  INV_X1 U5354 ( .A(n4751), .ZN(n4749) );
  AOI21_X1 U5355 ( .B1(n8803), .B2(n6418), .A(n4752), .ZN(n4751) );
  INV_X1 U5356 ( .A(n6543), .ZN(n4752) );
  OR2_X1 U5357 ( .A1(n8980), .A2(n8505), .ZN(n6418) );
  AOI21_X1 U5358 ( .B1(n8077), .B2(n6099), .A(n4802), .ZN(n4801) );
  OAI21_X1 U5359 ( .B1(n8836), .B2(n6344), .A(n6481), .ZN(n8810) );
  NAND2_X1 U5360 ( .A1(n6085), .A2(n6084), .ZN(n8076) );
  OR2_X1 U5361 ( .A1(n8076), .A2(n8077), .ZN(n8074) );
  NOR2_X1 U5362 ( .A1(n8879), .A2(n6340), .ZN(n6341) );
  OR2_X1 U5363 ( .A1(n10263), .A2(n7967), .ZN(n6458) );
  AND2_X1 U5364 ( .A1(n8879), .A2(n8873), .ZN(n4815) );
  NAND2_X1 U5365 ( .A1(n8068), .A2(n4839), .ZN(n8890) );
  AND2_X2 U5366 ( .A1(n7927), .A2(n10239), .ZN(n8068) );
  NAND2_X1 U5367 ( .A1(n6008), .A2(n6007), .ZN(n6025) );
  AND2_X1 U5368 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n6007) );
  NAND2_X1 U5369 ( .A1(n6404), .A2(n7036), .ZN(n4721) );
  OR2_X1 U5370 ( .A1(n5968), .A2(n7954), .ZN(n5969) );
  NAND2_X1 U5371 ( .A1(n7957), .A2(n10150), .ZN(n7952) );
  OR2_X1 U5372 ( .A1(n7279), .A2(n6363), .ZN(n8882) );
  OR2_X1 U5373 ( .A1(n7279), .A2(n6364), .ZN(n8880) );
  AND2_X1 U5374 ( .A1(n6442), .A2(n7952), .ZN(n7797) );
  INV_X1 U5375 ( .A(n8882), .ZN(n8815) );
  NAND2_X1 U5376 ( .A1(n8537), .A2(n8124), .ZN(n6571) );
  INV_X1 U5377 ( .A(n8880), .ZN(n8816) );
  NAND2_X1 U5378 ( .A1(n8381), .A2(n8384), .ZN(n4730) );
  INV_X1 U5379 ( .A(n8382), .ZN(n4728) );
  NAND2_X1 U5380 ( .A1(n6265), .A2(n6264), .ZN(n8919) );
  INV_X1 U5381 ( .A(n8673), .ZN(n8935) );
  NAND2_X1 U5382 ( .A1(n6089), .A2(n6088), .ZN(n8997) );
  INV_X1 U5383 ( .A(n8225), .ZN(n6305) );
  INV_X1 U5384 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6284) );
  INV_X1 U5385 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U5386 ( .A1(n6166), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6321) );
  AND2_X1 U5387 ( .A1(n6781), .A2(n7720), .ZN(n4501) );
  NAND2_X1 U5388 ( .A1(n6737), .A2(n6738), .ZN(n6739) );
  NAND2_X1 U5389 ( .A1(n6896), .A2(n6897), .ZN(n4903) );
  OR2_X1 U5390 ( .A1(n9372), .A2(n9337), .ZN(n4932) );
  NAND2_X1 U5391 ( .A1(n5339), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4995) );
  AND2_X1 U5392 ( .A1(n7996), .A2(n4410), .ZN(n4925) );
  INV_X1 U5393 ( .A(n7553), .ZN(n7019) );
  INV_X1 U5394 ( .A(n5714), .ZN(n4894) );
  OAI21_X1 U5395 ( .B1(n9934), .B2(n7083), .A(n7084), .ZN(n7100) );
  NAND2_X1 U5396 ( .A1(n5448), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5415) );
  OR2_X1 U5397 ( .A1(n7097), .A2(n7096), .ZN(n4625) );
  OR2_X1 U5398 ( .A1(n7176), .A2(n9210), .ZN(n5032) );
  INV_X1 U5399 ( .A(n4863), .ZN(n4862) );
  NAND2_X1 U5400 ( .A1(n8168), .A2(n8172), .ZN(n4841) );
  AND2_X1 U5401 ( .A1(n9522), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4855) );
  NOR2_X1 U5402 ( .A1(n9518), .A2(n4622), .ZN(n9536) );
  AND2_X1 U5403 ( .A1(n9522), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n4622) );
  OR2_X1 U5404 ( .A1(n9536), .A2(n9535), .ZN(n4621) );
  INV_X1 U5405 ( .A(n9952), .ZN(n4849) );
  AND2_X1 U5406 ( .A1(n4596), .A2(n4594), .ZN(n9599) );
  AOI21_X1 U5407 ( .B1(n4390), .B2(n8275), .A(n4431), .ZN(n4942) );
  NAND2_X1 U5408 ( .A1(n9656), .A2(n9655), .ZN(n8298) );
  INV_X1 U5409 ( .A(n5009), .ZN(n9640) );
  NAND2_X1 U5410 ( .A1(n9654), .A2(n9667), .ZN(n4944) );
  NAND2_X1 U5411 ( .A1(n4572), .A2(n4573), .ZN(n9656) );
  AOI21_X1 U5412 ( .B1(n4575), .B2(n4581), .A(n4574), .ZN(n4573) );
  NAND2_X1 U5413 ( .A1(n4575), .A2(n9694), .ZN(n4572) );
  INV_X1 U5414 ( .A(n8296), .ZN(n4574) );
  INV_X1 U5415 ( .A(n4582), .ZN(n4581) );
  AOI21_X1 U5416 ( .B1(n4580), .B2(n4582), .A(n4579), .ZN(n4578) );
  INV_X1 U5417 ( .A(n9695), .ZN(n4580) );
  NOR2_X1 U5418 ( .A1(n9773), .A2(n9697), .ZN(n8272) );
  NOR2_X1 U5419 ( .A1(n9688), .A2(n9773), .ZN(n9677) );
  OR2_X1 U5420 ( .A1(n4579), .A2(n8295), .ZN(n9681) );
  NAND2_X1 U5421 ( .A1(n9694), .A2(n9695), .ZN(n9693) );
  NAND2_X1 U5422 ( .A1(n4447), .A2(n4954), .ZN(n4951) );
  NAND2_X1 U5423 ( .A1(n4401), .A2(n8269), .ZN(n4953) );
  AND2_X1 U5424 ( .A1(n5780), .A2(n8293), .ZN(n9695) );
  NAND2_X1 U5425 ( .A1(n4401), .A2(n4954), .ZN(n4950) );
  NAND2_X1 U5426 ( .A1(n5781), .A2(n8292), .ZN(n9702) );
  INV_X1 U5427 ( .A(n4956), .ZN(n4955) );
  OAI22_X1 U5428 ( .A1(n8229), .A2(n4962), .B1(n8228), .B2(n9468), .ZN(n4956)
         );
  AND2_X1 U5429 ( .A1(n4457), .A2(n8192), .ZN(n4961) );
  AND2_X1 U5430 ( .A1(n5743), .A2(n5729), .ZN(n8229) );
  AND4_X1 U5431 ( .A1(n5516), .A2(n5515), .A3(n5514), .A4(n5513), .ZN(n8048)
         );
  NAND2_X1 U5432 ( .A1(n7901), .A2(n5733), .ZN(n5003) );
  AND2_X1 U5433 ( .A1(n7811), .A2(n7901), .ZN(n5005) );
  AND2_X1 U5434 ( .A1(n7983), .A2(n7981), .ZN(n7978) );
  INV_X1 U5435 ( .A(n7708), .ZN(n7696) );
  NAND2_X1 U5436 ( .A1(n7565), .A2(n7564), .ZN(n7689) );
  AND2_X1 U5437 ( .A1(n10025), .A2(n10090), .ZN(n10003) );
  CLKBUF_X1 U5438 ( .A(n9982), .Z(n9983) );
  NOR2_X1 U5439 ( .A1(n10024), .A2(n5365), .ZN(n10025) );
  INV_X1 U5440 ( .A(n9715), .ZN(n10040) );
  OR2_X1 U5441 ( .A1(n7010), .A2(n9492), .ZN(n10018) );
  INV_X1 U5442 ( .A(n10018), .ZN(n10037) );
  NAND2_X1 U5443 ( .A1(n5251), .A2(n5250), .ZN(n9726) );
  OAI211_X1 U5444 ( .C1(n8163), .C2(P1_B_REG_SCAN_IN), .A(n6951), .B(n6950), 
        .ZN(n7188) );
  INV_X1 U5445 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5237) );
  INV_X1 U5446 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5221) );
  XNOR2_X1 U5447 ( .A(n5258), .B(n5257), .ZN(n8329) );
  XNOR2_X1 U5448 ( .A(n5685), .B(n5684), .ZN(n9039) );
  NAND2_X1 U5449 ( .A1(n5682), .A2(n5681), .ZN(n5685) );
  XNOR2_X1 U5450 ( .A(n5652), .B(n5651), .ZN(n8222) );
  OAI21_X1 U5451 ( .B1(n5630), .B2(n5181), .A(n5180), .ZN(n5652) );
  XNOR2_X1 U5452 ( .A(n4653), .B(n5577), .ZN(n7909) );
  OAI21_X1 U5453 ( .B1(n5573), .B2(n5572), .A(n5574), .ZN(n4653) );
  OR2_X1 U5454 ( .A1(n5494), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5525) );
  XNOR2_X1 U5455 ( .A(n5430), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7232) );
  NAND2_X1 U5456 ( .A1(n5429), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U5457 ( .A1(n5305), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4872) );
  NOR2_X1 U5458 ( .A1(n9871), .A2(n9870), .ZN(n9872) );
  NAND2_X1 U5459 ( .A1(n7532), .A2(n6608), .ZN(n7547) );
  AND2_X1 U5460 ( .A1(n6209), .A2(n6208), .ZN(n8427) );
  INV_X1 U5461 ( .A(n8769), .ZN(n8428) );
  NAND2_X1 U5462 ( .A1(n6189), .A2(n6188), .ZN(n8741) );
  INV_X1 U5463 ( .A(n8526), .ZN(n8854) );
  NAND3_X1 U5464 ( .A1(n6684), .A2(n8908), .A3(n6676), .ZN(n8519) );
  AND2_X1 U5465 ( .A1(n7257), .A2(n6679), .ZN(n10151) );
  NAND2_X1 U5466 ( .A1(n6273), .A2(n6272), .ZN(n8635) );
  NAND2_X1 U5467 ( .A1(n7389), .A2(n7390), .ZN(n7388) );
  NOR2_X1 U5468 ( .A1(n8596), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8607) );
  OAI21_X1 U5469 ( .B1(n8619), .B2(n8618), .A(n4670), .ZN(n4669) );
  AND2_X1 U5470 ( .A1(n8617), .A2(n10166), .ZN(n4670) );
  INV_X1 U5471 ( .A(n4668), .ZN(n4667) );
  AOI21_X1 U5472 ( .B1(n10164), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n8621), .ZN(
        n4668) );
  NAND2_X1 U5473 ( .A1(n6408), .A2(n6407), .ZN(n8899) );
  OAI21_X1 U5474 ( .B1(n4728), .B2(n4730), .A(n4729), .ZN(n8917) );
  AOI21_X1 U5475 ( .B1(n8915), .B2(n8895), .A(n8390), .ZN(n8391) );
  NAND2_X1 U5476 ( .A1(n8378), .A2(n8377), .ZN(n8379) );
  OR2_X1 U5477 ( .A1(n8919), .A2(n8635), .ZN(n8377) );
  OR2_X1 U5478 ( .A1(n5954), .A2(n7056), .ZN(n5931) );
  AND2_X1 U5479 ( .A1(n6377), .A2(n7538), .ZN(n8895) );
  NAND2_X1 U5480 ( .A1(n4728), .A2(n4729), .ZN(n4727) );
  NAND2_X1 U5481 ( .A1(n4730), .A2(n4729), .ZN(n4726) );
  NAND2_X1 U5482 ( .A1(n7753), .A2(n5347), .ZN(n5566) );
  NOR2_X1 U5483 ( .A1(n5036), .A2(n6991), .ZN(n6992) );
  INV_X1 U5484 ( .A(n9770), .ZN(n9369) );
  AND2_X1 U5485 ( .A1(n5607), .A2(n5606), .ZN(n9478) );
  NAND2_X1 U5486 ( .A1(n6980), .A2(n6979), .ZN(n9462) );
  INV_X1 U5487 ( .A(n8216), .ZN(n9798) );
  AND2_X1 U5488 ( .A1(n7731), .A2(n10106), .ZN(n9470) );
  OR2_X1 U5489 ( .A1(n5604), .A2(n5353), .ZN(n5033) );
  CLKBUF_X1 U5490 ( .A(n5322), .Z(n9493) );
  NAND2_X1 U5491 ( .A1(n7081), .A2(n7080), .ZN(n7119) );
  NOR2_X1 U5492 ( .A1(n7123), .A2(n4626), .ZN(n7097) );
  NOR2_X1 U5493 ( .A1(n7130), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4626) );
  OAI21_X1 U5494 ( .B1(n7673), .B2(n7672), .A(n4465), .ZN(n7863) );
  NOR2_X1 U5495 ( .A1(n9520), .A2(n9519), .ZN(n9518) );
  NAND2_X1 U5496 ( .A1(n10033), .A2(n10007), .ZN(n9710) );
  INV_X1 U5497 ( .A(n7754), .ZN(n10011) );
  INV_X1 U5498 ( .A(n9710), .ZN(n10050) );
  INV_X1 U5499 ( .A(n9573), .ZN(n10028) );
  OR2_X1 U5500 ( .A1(n9757), .A2(n10110), .ZN(n4490) );
  NOR2_X1 U5501 ( .A1(n9884), .A2(n10353), .ZN(n10342) );
  NOR2_X1 U5502 ( .A1(n7887), .A2(n4709), .ZN(n4708) );
  NAND2_X1 U5503 ( .A1(n4706), .A2(n4408), .ZN(n4705) );
  AND2_X1 U5504 ( .A1(n4802), .A2(n6479), .ZN(n4600) );
  AOI21_X1 U5505 ( .B1(n4382), .B2(n8686), .A(n4616), .ZN(n4615) );
  NOR2_X1 U5506 ( .A1(n8301), .A2(n9641), .ZN(n4886) );
  AND2_X1 U5507 ( .A1(n5741), .A2(n4568), .ZN(n5742) );
  NAND2_X1 U5508 ( .A1(n5624), .A2(n8297), .ZN(n5763) );
  INV_X1 U5509 ( .A(n6661), .ZN(n4517) );
  OAI21_X1 U5510 ( .B1(n6517), .B2(n4604), .A(n4601), .ZN(n4605) );
  NAND2_X1 U5511 ( .A1(n8656), .A2(n4393), .ZN(n4604) );
  NAND2_X1 U5512 ( .A1(n6351), .A2(n4756), .ZN(n4754) );
  NOR2_X1 U5513 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6152) );
  NOR2_X1 U5514 ( .A1(n4698), .A2(n4693), .ZN(n4692) );
  INV_X1 U5515 ( .A(n5176), .ZN(n4693) );
  INV_X1 U5516 ( .A(n4699), .ZN(n4698) );
  INV_X1 U5517 ( .A(n4701), .ZN(n4697) );
  INV_X1 U5518 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5145) );
  INV_X1 U5519 ( .A(SI_16_), .ZN(n5139) );
  INV_X1 U5520 ( .A(SI_15_), .ZN(n5133) );
  NAND2_X1 U5521 ( .A1(n5126), .A2(n5125), .ZN(n5129) );
  INV_X1 U5522 ( .A(SI_13_), .ZN(n5125) );
  NOR2_X1 U5523 ( .A1(n5119), .A2(n4678), .ZN(n4677) );
  INV_X1 U5524 ( .A(n5114), .ZN(n4678) );
  INV_X1 U5525 ( .A(n5477), .ZN(n5119) );
  OAI21_X1 U5526 ( .B1(n7033), .B2(n5096), .A(n5095), .ZN(n5098) );
  OAI21_X1 U5527 ( .B1(n5305), .B2(n5087), .A(n5086), .ZN(n5088) );
  AND2_X1 U5528 ( .A1(n6105), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6123) );
  NOR2_X1 U5529 ( .A1(n6551), .A2(n4558), .ZN(n4557) );
  NOR2_X1 U5530 ( .A1(n8879), .A2(n4560), .ZN(n4559) );
  NOR2_X1 U5531 ( .A1(n8651), .A2(n4643), .ZN(n4566) );
  NAND2_X1 U5532 ( .A1(n4657), .A2(n4660), .ZN(n4656) );
  AND3_X1 U5533 ( .A1(n4680), .A2(n8632), .A3(n8633), .ZN(n4740) );
  INV_X1 U5534 ( .A(n4742), .ZN(n4741) );
  OR2_X1 U5535 ( .A1(n8930), .A2(n8439), .ZN(n6519) );
  AND2_X1 U5536 ( .A1(n6212), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6223) );
  INV_X1 U5537 ( .A(n6213), .ZN(n6212) );
  OR2_X1 U5538 ( .A1(n8940), .A2(n8699), .ZN(n4640) );
  OR2_X1 U5539 ( .A1(n8940), .A2(n8440), .ZN(n6512) );
  NAND2_X1 U5540 ( .A1(n6169), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6180) );
  INV_X1 U5541 ( .A(n6171), .ZN(n6169) );
  OR2_X1 U5542 ( .A1(n6157), .A2(n9173), .ZN(n6171) );
  NAND2_X1 U5543 ( .A1(n6124), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6157) );
  INV_X1 U5544 ( .A(n6139), .ZN(n6124) );
  AND2_X1 U5545 ( .A1(n6343), .A2(n8855), .ZN(n6081) );
  INV_X1 U5546 ( .A(n7797), .ZN(n7802) );
  NAND2_X1 U5547 ( .A1(n10144), .A2(n7959), .ZN(n6425) );
  NAND2_X1 U5548 ( .A1(n8534), .A2(n10218), .ZN(n6443) );
  AND2_X1 U5549 ( .A1(n4795), .A2(n9075), .ZN(n4793) );
  INV_X1 U5550 ( .A(SI_22_), .ZN(n9253) );
  INV_X1 U5551 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6278) );
  INV_X1 U5552 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9131) );
  INV_X1 U5553 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9173) );
  INV_X1 U5554 ( .A(n9391), .ZN(n4922) );
  AND2_X1 U5555 ( .A1(n4920), .A2(n6871), .ZN(n4919) );
  NAND2_X1 U5556 ( .A1(n9391), .A2(n4921), .ZN(n4920) );
  AND2_X1 U5557 ( .A1(n5846), .A2(n5255), .ZN(n5709) );
  INV_X1 U5558 ( .A(n5665), .ZN(n4880) );
  OR2_X1 U5559 ( .A1(n9570), .A2(n9582), .ZN(n5775) );
  NAND2_X1 U5560 ( .A1(n7232), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4866) );
  INV_X1 U5561 ( .A(n5032), .ZN(n4861) );
  INV_X1 U5562 ( .A(n4866), .ZN(n4860) );
  AOI21_X1 U5563 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n8167), .A(n8166), .ZN(
        n8168) );
  NAND2_X1 U5564 ( .A1(n4588), .A2(n4590), .ZN(n8310) );
  AOI21_X1 U5565 ( .B1(n4592), .B2(n4593), .A(n4445), .ZN(n4590) );
  NOR2_X1 U5566 ( .A1(n9743), .A2(n9750), .ZN(n4975) );
  INV_X1 U5567 ( .A(n9610), .ZN(n4937) );
  NAND3_X1 U5568 ( .A1(n8298), .A2(n5010), .A3(n5663), .ZN(n5008) );
  AND2_X1 U5569 ( .A1(n4578), .A2(n4576), .ZN(n4575) );
  INV_X1 U5570 ( .A(n9664), .ZN(n4576) );
  NAND2_X1 U5571 ( .A1(n9369), .A2(n4987), .ZN(n4986) );
  OR2_X1 U5572 ( .A1(n9763), .A2(n4986), .ZN(n4985) );
  NOR2_X1 U5573 ( .A1(n8229), .A2(n4959), .ZN(n4958) );
  INV_X1 U5574 ( .A(n4961), .ZN(n4959) );
  NAND2_X1 U5575 ( .A1(n10076), .A2(n7554), .ZN(n5829) );
  NAND2_X1 U5576 ( .A1(n9626), .A2(n4424), .ZN(n5035) );
  NAND2_X1 U5577 ( .A1(n7659), .A2(n10069), .ZN(n7643) );
  NAND2_X1 U5578 ( .A1(n5682), .A2(n5191), .ZN(n5696) );
  NOR2_X1 U5579 ( .A1(n5651), .A2(n4702), .ZN(n4701) );
  INV_X1 U5580 ( .A(n5180), .ZN(n4702) );
  AND2_X1 U5581 ( .A1(n5681), .A2(n5189), .ZN(n5667) );
  AOI21_X1 U5582 ( .B1(n4701), .B2(n5181), .A(n4700), .ZN(n4699) );
  INV_X1 U5583 ( .A(n5186), .ZN(n4700) );
  NAND2_X1 U5584 ( .A1(n4550), .A2(n4549), .ZN(n5051) );
  AOI21_X1 U5585 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_20__SCAN_IN), .ZN(n4549) );
  OR2_X1 U5586 ( .A1(n5161), .A2(n5160), .ZN(n5594) );
  AND2_X1 U5587 ( .A1(n4895), .A2(n4686), .ZN(n4685) );
  NAND2_X1 U5588 ( .A1(n4689), .A2(n4687), .ZN(n4686) );
  INV_X1 U5589 ( .A(n5274), .ZN(n4897) );
  XNOR2_X1 U5590 ( .A(n5150), .B(SI_18_), .ZN(n5547) );
  XNOR2_X1 U5591 ( .A(n5146), .B(SI_17_), .ZN(n5274) );
  NAND2_X1 U5592 ( .A1(n5124), .A2(n5123), .ZN(n5460) );
  INV_X1 U5593 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4828) );
  INV_X1 U5594 ( .A(n8635), .ZN(n6710) );
  NOR2_X1 U5595 ( .A1(n8095), .A2(n4786), .ZN(n4785) );
  NAND2_X1 U5596 ( .A1(n8397), .A2(n8398), .ZN(n8396) );
  INV_X1 U5597 ( .A(n7664), .ZN(n4764) );
  XNOR2_X1 U5598 ( .A(n6589), .B(n10194), .ZN(n7250) );
  CLKBUF_X1 U5599 ( .A(n8007), .Z(n4506) );
  AND2_X1 U5600 ( .A1(n8470), .A2(n8471), .ZN(n4495) );
  INV_X1 U5601 ( .A(n6663), .ZN(n4510) );
  INV_X1 U5602 ( .A(n8699), .ZN(n8440) );
  AOI21_X1 U5603 ( .B1(n7546), .B2(n4767), .A(n4425), .ZN(n4766) );
  INV_X1 U5604 ( .A(n6608), .ZN(n4767) );
  INV_X1 U5605 ( .A(n7546), .ZN(n4768) );
  NAND2_X1 U5606 ( .A1(n4506), .A2(n6627), .ZN(n8008) );
  XNOR2_X1 U5607 ( .A(n6574), .B(n6589), .ZN(n6577) );
  NAND2_X1 U5608 ( .A1(n6647), .A2(n4783), .ZN(n4782) );
  INV_X1 U5609 ( .A(n6648), .ZN(n4783) );
  AND2_X1 U5610 ( .A1(n6677), .A2(n8904), .ZN(n6684) );
  AND2_X1 U5611 ( .A1(n6532), .A2(n6531), .ZN(n4717) );
  OAI21_X1 U5612 ( .B1(n7411), .B2(n4660), .A(n4657), .ZN(n8579) );
  AOI21_X1 U5613 ( .B1(n4664), .B2(n7420), .A(n4663), .ZN(n4662) );
  NAND2_X1 U5614 ( .A1(n7465), .A2(n4664), .ZN(n7491) );
  INV_X1 U5615 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6117) );
  OAI21_X1 U5616 ( .B1(n8021), .B2(n8020), .A(n8022), .ZN(n8025) );
  AOI21_X1 U5617 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8598), .A(n8597), .ZN(
        n8612) );
  AND2_X1 U5618 ( .A1(n6355), .A2(n6267), .ZN(n8364) );
  AND2_X1 U5619 ( .A1(n4743), .A2(n4420), .ZN(n8655) );
  NAND2_X1 U5620 ( .A1(n8657), .A2(n8816), .ZN(n4531) );
  OR2_X1 U5621 ( .A1(n6234), .A2(n8437), .ZN(n6246) );
  NAND2_X1 U5622 ( .A1(n8935), .A2(n4831), .ZN(n4830) );
  NOR2_X1 U5623 ( .A1(n8970), .A2(n4834), .ZN(n4832) );
  INV_X1 U5624 ( .A(n4834), .ZN(n4833) );
  NAND2_X1 U5625 ( .A1(n8843), .A2(n4836), .ZN(n8795) );
  NAND2_X1 U5626 ( .A1(n8843), .A2(n8826), .ZN(n8828) );
  INV_X1 U5627 ( .A(n8809), .ZN(n8811) );
  OR2_X1 U5628 ( .A1(n6076), .A2(n6066), .ZN(n6091) );
  NAND2_X1 U5629 ( .A1(n6090), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6107) );
  INV_X1 U5630 ( .A(n6091), .ZN(n6090) );
  INV_X1 U5631 ( .A(n6343), .ZN(n8857) );
  INV_X1 U5632 ( .A(n6458), .ZN(n4725) );
  AND3_X1 U5633 ( .A1(n4422), .A2(n10274), .A3(n8068), .ZN(n8130) );
  NAND2_X1 U5634 ( .A1(n4810), .A2(n4811), .ZN(n8127) );
  INV_X1 U5635 ( .A(n4812), .ZN(n4811) );
  OAI21_X1 U5636 ( .B1(n5015), .B2(n4813), .A(n6062), .ZN(n4812) );
  AND2_X1 U5637 ( .A1(n4422), .A2(n8068), .ZN(n8889) );
  INV_X1 U5638 ( .A(n6025), .ZN(n6023) );
  AND2_X1 U5639 ( .A1(n6000), .A2(n4423), .ZN(n4807) );
  AND2_X1 U5640 ( .A1(n5985), .A2(n6000), .ZN(n4808) );
  NAND2_X1 U5641 ( .A1(n5971), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6006) );
  AND2_X1 U5642 ( .A1(n4822), .A2(n10212), .ZN(n7947) );
  AND3_X1 U5643 ( .A1(n6574), .A2(n10188), .A3(n10194), .ZN(n4822) );
  NAND2_X1 U5644 ( .A1(n4823), .A2(n6574), .ZN(n7838) );
  INV_X1 U5645 ( .A(n8144), .ZN(n4823) );
  NAND2_X1 U5646 ( .A1(n5946), .A2(n5945), .ZN(n7796) );
  CLKBUF_X1 U5647 ( .A(n7800), .Z(n7841) );
  NAND2_X1 U5648 ( .A1(n10194), .A2(n10188), .ZN(n8144) );
  INV_X1 U5649 ( .A(n8070), .ZN(n4840) );
  INV_X1 U5650 ( .A(n10282), .ZN(n10265) );
  INV_X1 U5651 ( .A(n8908), .ZN(n9007) );
  NOR2_X1 U5652 ( .A1(n8907), .A2(n8906), .ZN(n9008) );
  OR2_X1 U5653 ( .A1(n6309), .A2(n6308), .ZN(n6310) );
  XNOR2_X1 U5654 ( .A(n4758), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U5655 ( .A1(n4757), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4758) );
  INV_X1 U5656 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6316) );
  AND2_X1 U5657 ( .A1(n6001), .A2(n5991), .ZN(n7360) );
  NAND2_X1 U5658 ( .A1(n4914), .A2(n7239), .ZN(n4913) );
  INV_X1 U5659 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9249) );
  AND2_X1 U5660 ( .A1(n6726), .A2(n6725), .ZN(n9372) );
  AOI22_X1 U5661 ( .A1(n6758), .A2(n7626), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6727), .ZN(n6728) );
  NAND2_X1 U5662 ( .A1(n6736), .A2(n7626), .ZN(n6732) );
  NOR2_X1 U5663 ( .A1(n4389), .A2(n4541), .ZN(n4540) );
  NAND2_X1 U5664 ( .A1(n4906), .A2(n4904), .ZN(n4907) );
  INV_X1 U5665 ( .A(n6914), .ZN(n6915) );
  OR2_X1 U5666 ( .A1(n5454), .A2(n5264), .ZN(n5486) );
  NAND2_X1 U5667 ( .A1(n7040), .A2(n6977), .ZN(n7016) );
  NOR2_X1 U5668 ( .A1(n9444), .A2(n9445), .ZN(n4929) );
  NAND2_X1 U5669 ( .A1(n4544), .A2(n4434), .ZN(n9457) );
  INV_X1 U5670 ( .A(n4892), .ZN(n4891) );
  OAI211_X1 U5671 ( .C1(n5805), .C2(n5722), .A(n4409), .B(n4893), .ZN(n4892)
         );
  NAND2_X1 U5672 ( .A1(n5769), .A2(n5715), .ZN(n4893) );
  NAND2_X1 U5673 ( .A1(n5227), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5228) );
  NOR2_X1 U5674 ( .A1(n9940), .A2(n4623), .ZN(n7073) );
  AND2_X1 U5675 ( .A1(n9935), .A2(n7070), .ZN(n4623) );
  OR2_X1 U5676 ( .A1(n7101), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4869) );
  NAND2_X1 U5677 ( .A1(n7073), .A2(n7072), .ZN(n7091) );
  NOR2_X1 U5678 ( .A1(n7126), .A2(n4868), .ZN(n7105) );
  AND2_X1 U5679 ( .A1(n7130), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4868) );
  INV_X1 U5680 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9268) );
  AND2_X1 U5681 ( .A1(n7267), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4856) );
  AOI21_X1 U5682 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7866), .A(n7865), .ZN(
        n7869) );
  NOR2_X1 U5683 ( .A1(n8169), .A2(n8170), .ZN(n8245) );
  AND2_X1 U5684 ( .A1(n5774), .A2(n5847), .ZN(n9549) );
  AND2_X1 U5685 ( .A1(n8285), .A2(n8283), .ZN(n8284) );
  AND2_X1 U5686 ( .A1(n9561), .A2(n5703), .ZN(n9569) );
  INV_X1 U5687 ( .A(n8307), .ZN(n9589) );
  XNOR2_X1 U5688 ( .A(n4402), .B(n9623), .ZN(n4486) );
  NOR2_X1 U5689 ( .A1(n9688), .A2(n4986), .ZN(n9668) );
  NOR2_X1 U5690 ( .A1(n4949), .A2(n4437), .ZN(n4945) );
  INV_X1 U5691 ( .A(n9702), .ZN(n9714) );
  OAI21_X1 U5692 ( .B1(n8291), .B2(n8290), .A(n8289), .ZN(n9713) );
  INV_X1 U5693 ( .A(n4968), .ZN(n4967) );
  NOR2_X1 U5694 ( .A1(n4968), .A2(n8214), .ZN(n8287) );
  OR2_X1 U5695 ( .A1(n5285), .A2(n8290), .ZN(n8238) );
  NAND2_X1 U5696 ( .A1(n4969), .A2(n4970), .ZN(n8231) );
  NOR2_X1 U5697 ( .A1(n9795), .A2(n9798), .ZN(n4970) );
  AND2_X1 U5698 ( .A1(n8202), .A2(n8201), .ZN(n8209) );
  OAI21_X1 U5699 ( .B1(n8045), .B2(n8044), .A(n8043), .ZN(n8046) );
  NAND2_X1 U5700 ( .A1(n4992), .A2(n8039), .ZN(n8200) );
  INV_X1 U5701 ( .A(n8046), .ZN(n4992) );
  INV_X1 U5702 ( .A(n9809), .ZN(n8036) );
  AND2_X1 U5703 ( .A1(n7988), .A2(n9809), .ZN(n8040) );
  AND4_X1 U5704 ( .A1(n5503), .A2(n5502), .A3(n5501), .A4(n5500), .ZN(n8189)
         );
  NOR2_X1 U5705 ( .A1(n7904), .A2(n9816), .ZN(n7988) );
  NAND3_X1 U5706 ( .A1(n4979), .A2(n7876), .A3(n4978), .ZN(n7904) );
  NOR2_X1 U5707 ( .A1(n4980), .A2(n9819), .ZN(n4978) );
  NAND2_X1 U5708 ( .A1(n7812), .A2(n7811), .ZN(n5004) );
  INV_X1 U5709 ( .A(n4980), .ZN(n4977) );
  AND2_X1 U5710 ( .A1(n7813), .A2(n5784), .ZN(n7708) );
  NAND2_X1 U5711 ( .A1(n5432), .A2(n5431), .ZN(n7747) );
  NOR2_X1 U5712 ( .A1(n7713), .A2(n4980), .ZN(n7745) );
  AND4_X1 U5713 ( .A1(n5459), .A2(n5458), .A3(n5457), .A4(n5456), .ZN(n7814)
         );
  NAND2_X1 U5714 ( .A1(n7705), .A2(n7704), .ZN(n7735) );
  AND2_X1 U5715 ( .A1(n9968), .A2(n7703), .ZN(n7704) );
  AOI21_X1 U5716 ( .B1(n7702), .B2(n7701), .A(n7700), .ZN(n7703) );
  NOR2_X1 U5717 ( .A1(n7713), .A2(n9976), .ZN(n9977) );
  NAND2_X1 U5718 ( .A1(n5419), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U5719 ( .A1(n7690), .A2(n7691), .ZN(n9966) );
  AND2_X2 U5720 ( .A1(n5791), .A2(n7736), .ZN(n9968) );
  NOR2_X2 U5721 ( .A1(n7698), .A2(n7563), .ZN(n9990) );
  NAND3_X1 U5722 ( .A1(n10069), .A2(n5819), .A3(n4426), .ZN(n10024) );
  NAND2_X1 U5723 ( .A1(n7009), .A2(n7008), .ZN(n10034) );
  OR3_X1 U5724 ( .A1(n7016), .A2(n7199), .A3(n7015), .ZN(n7575) );
  NAND2_X1 U5725 ( .A1(n5642), .A2(n5641), .ZN(n9758) );
  INV_X1 U5726 ( .A(n10121), .ZN(n10004) );
  OR2_X1 U5727 ( .A1(n10034), .A2(n10126), .ZN(n10093) );
  OR2_X1 U5728 ( .A1(n7574), .A2(n7573), .ZN(n10121) );
  OR2_X1 U5729 ( .A1(n7574), .A2(n6971), .ZN(n10119) );
  NAND2_X1 U5730 ( .A1(n6716), .A2(n7913), .ZN(n7574) );
  AND2_X1 U5731 ( .A1(n7001), .A2(n6999), .ZN(n6976) );
  XNOR2_X1 U5732 ( .A(n5249), .B(n5248), .ZN(n8326) );
  CLKBUF_X1 U5733 ( .A(n5870), .Z(n9926) );
  XNOR2_X1 U5734 ( .A(n5698), .B(n5697), .ZN(n8341) );
  AND2_X1 U5735 ( .A1(n5696), .A2(n5695), .ZN(n5698) );
  NAND2_X1 U5736 ( .A1(n5883), .A2(n5884), .ZN(n8163) );
  NAND2_X1 U5737 ( .A1(n5879), .A2(n5878), .ZN(n5883) );
  NAND2_X1 U5738 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5877), .ZN(n5878) );
  AND2_X1 U5739 ( .A1(n5176), .A2(n5175), .ZN(n5639) );
  XNOR2_X1 U5740 ( .A(n5275), .B(n5274), .ZN(n7436) );
  AND2_X1 U5741 ( .A1(n5496), .A2(n5525), .ZN(n8256) );
  OAI21_X1 U5742 ( .B1(n5461), .B2(n4878), .A(n4874), .ZN(n5493) );
  NAND2_X1 U5743 ( .A1(n5115), .A2(n5114), .ZN(n5478) );
  OR2_X1 U5744 ( .A1(n5394), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5448) );
  INV_X1 U5745 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5446) );
  XNOR2_X1 U5746 ( .A(n5413), .B(n5414), .ZN(n7044) );
  NAND2_X1 U5747 ( .A1(n4899), .A2(n5099), .ZN(n5414) );
  BUF_X1 U5748 ( .A(n7032), .Z(n4518) );
  NAND2_X1 U5749 ( .A1(n9878), .A2(n9879), .ZN(n9880) );
  NAND2_X1 U5750 ( .A1(n4790), .A2(n4788), .ZN(n7534) );
  OR2_X1 U5751 ( .A1(n4792), .A2(n4791), .ZN(n4790) );
  INV_X1 U5752 ( .A(n6601), .ZN(n4791) );
  NAND2_X1 U5753 ( .A1(n9039), .A2(n6404), .ZN(n4675) );
  AND2_X1 U5754 ( .A1(n5956), .A2(n4416), .ZN(n4492) );
  NAND2_X1 U5755 ( .A1(n8416), .A2(n8415), .ZN(n8414) );
  NAND2_X1 U5756 ( .A1(n4776), .A2(n4774), .ZN(n8416) );
  NAND2_X1 U5757 ( .A1(n4513), .A2(n4777), .ZN(n4776) );
  NOR2_X1 U5758 ( .A1(n8362), .A2(n8361), .ZN(n8363) );
  AND2_X1 U5759 ( .A1(n6696), .A2(n6695), .ZN(n8371) );
  AND2_X1 U5760 ( .A1(n8355), .A2(n8359), .ZN(n8372) );
  INV_X1 U5761 ( .A(n8527), .ZN(n8881) );
  INV_X1 U5762 ( .A(n8525), .ZN(n8401) );
  NAND2_X1 U5763 ( .A1(n6233), .A2(n6232), .ZN(n8673) );
  INV_X1 U5764 ( .A(n8534), .ZN(n10144) );
  OR2_X1 U5765 ( .A1(n6591), .A2(n6590), .ZN(n6592) );
  CLKBUF_X1 U5766 ( .A(n7438), .Z(n7500) );
  NAND2_X1 U5767 ( .A1(n4766), .A2(n4765), .ZN(n7666) );
  OR2_X1 U5768 ( .A1(n7532), .A2(n4768), .ZN(n4765) );
  NAND2_X1 U5769 ( .A1(n6572), .A2(n4384), .ZN(n7541) );
  AOI21_X1 U5770 ( .B1(n4773), .B2(n8415), .A(n4772), .ZN(n4771) );
  INV_X1 U5771 ( .A(n4536), .ZN(n4772) );
  NAND2_X1 U5772 ( .A1(n8008), .A2(n6628), .ZN(n8096) );
  NAND2_X1 U5773 ( .A1(n6199), .A2(n6198), .ZN(n8950) );
  NAND2_X1 U5774 ( .A1(n4779), .A2(n4782), .ZN(n8503) );
  OR2_X1 U5775 ( .A1(n4513), .A2(n8460), .ZN(n4779) );
  OR2_X1 U5776 ( .A1(n8516), .A2(n8882), .ZN(n10148) );
  OR2_X1 U5777 ( .A1(n8516), .A2(n8880), .ZN(n10145) );
  NAND2_X1 U5778 ( .A1(n6104), .A2(n6103), .ZN(n8992) );
  INV_X1 U5779 ( .A(n6566), .ZN(n4704) );
  AOI22_X1 U5780 ( .A1(n8381), .A2(n6403), .B1(n6528), .B2(n6402), .ZN(n6411)
         );
  AND3_X1 U5781 ( .A1(n4567), .A2(n6555), .A3(n4562), .ZN(n6560) );
  OR2_X1 U5782 ( .A1(n6143), .A2(n6142), .ZN(n8523) );
  AND2_X1 U5783 ( .A1(n5947), .A2(n5949), .ZN(n4502) );
  INV_X2 U5784 ( .A(P2_U3966), .ZN(n8536) );
  NAND2_X1 U5785 ( .A1(n5976), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U5786 ( .A1(n7388), .A2(n7373), .ZN(n7289) );
  NAND2_X1 U5787 ( .A1(n7411), .A2(n7410), .ZN(n8566) );
  OR2_X1 U5788 ( .A1(n7407), .A2(n7408), .ZN(n7475) );
  OR2_X1 U5789 ( .A1(n7421), .A2(n7420), .ZN(n7465) );
  NAND2_X1 U5790 ( .A1(n7465), .A2(n7464), .ZN(n7469) );
  NAND2_X1 U5791 ( .A1(n7484), .A2(n7483), .ZN(n7765) );
  AND2_X1 U5792 ( .A1(n7775), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7785) );
  NAND2_X1 U5793 ( .A1(n7137), .A2(n7136), .ZN(n10164) );
  OR2_X1 U5794 ( .A1(n4428), .A2(n8608), .ZN(n8596) );
  XNOR2_X1 U5795 ( .A(n8622), .B(n8899), .ZN(n8901) );
  INV_X1 U5796 ( .A(n8627), .ZN(n8912) );
  AOI21_X1 U5797 ( .B1(n6368), .B2(n8886), .A(n6367), .ZN(n8922) );
  OAI21_X1 U5798 ( .B1(n8650), .B2(n8633), .A(n4798), .ZN(n6274) );
  NAND2_X1 U5799 ( .A1(n8645), .A2(n8644), .ZN(n8643) );
  INV_X1 U5800 ( .A(n8636), .ZN(n8637) );
  XNOR2_X1 U5801 ( .A(n8634), .B(n8633), .ZN(n8638) );
  AOI22_X1 U5802 ( .A1(n8635), .A2(n8816), .B1(n8815), .B2(n8666), .ZN(n8636)
         );
  AOI21_X1 U5803 ( .B1(n4532), .B2(n8886), .A(n4529), .ZN(n8932) );
  NAND2_X1 U5804 ( .A1(n4531), .A2(n4530), .ZN(n4529) );
  OAI21_X1 U5805 ( .B1(n8655), .B2(n8656), .A(n8654), .ZN(n4532) );
  NAND2_X1 U5806 ( .A1(n8689), .A2(n8815), .ZN(n4530) );
  AND2_X1 U5807 ( .A1(n8691), .A2(n8690), .ZN(n8943) );
  INV_X1 U5808 ( .A(n6370), .ZN(n8701) );
  OAI21_X1 U5809 ( .B1(n8712), .B2(n4647), .A(n4644), .ZN(n8679) );
  NAND2_X1 U5810 ( .A1(n4648), .A2(n4646), .ZN(n8706) );
  AND2_X1 U5811 ( .A1(n4648), .A2(n4411), .ZN(n8708) );
  NAND2_X1 U5812 ( .A1(n8712), .A2(n6350), .ZN(n4648) );
  INV_X1 U5813 ( .A(n8950), .ZN(n8719) );
  NOR2_X1 U5814 ( .A1(n8750), .A2(n6349), .ZN(n8733) );
  NAND2_X1 U5815 ( .A1(n4816), .A2(n4392), .ZN(n8730) );
  NAND2_X1 U5816 ( .A1(n8764), .A2(n4818), .ZN(n4816) );
  NAND2_X1 U5817 ( .A1(n4820), .A2(n4821), .ZN(n8760) );
  NAND2_X1 U5818 ( .A1(n4820), .A2(n4818), .ZN(n8962) );
  AND2_X1 U5819 ( .A1(n8753), .A2(n8752), .ZN(n8968) );
  OR3_X1 U5820 ( .A1(n8750), .A2(n8821), .A3(n8749), .ZN(n8753) );
  NAND2_X1 U5821 ( .A1(n4744), .A2(n4748), .ZN(n8767) );
  NAND2_X1 U5822 ( .A1(n8791), .A2(n4750), .ZN(n4744) );
  NAND2_X1 U5823 ( .A1(n8074), .A2(n6099), .ZN(n8833) );
  NAND2_X1 U5824 ( .A1(n4724), .A2(n6458), .ZN(n7965) );
  NAND2_X1 U5825 ( .A1(n8877), .A2(n6341), .ZN(n4724) );
  NAND2_X1 U5826 ( .A1(n7963), .A2(n7964), .ZN(n7962) );
  NAND2_X1 U5827 ( .A1(n4814), .A2(n5015), .ZN(n7963) );
  NAND2_X1 U5828 ( .A1(n8101), .A2(n4815), .ZN(n4814) );
  NAND2_X1 U5829 ( .A1(n8068), .A2(n8070), .ZN(n8113) );
  NAND2_X1 U5830 ( .A1(n4735), .A2(n6445), .ZN(n7936) );
  INV_X1 U5831 ( .A(n7854), .ZN(n10226) );
  OR2_X1 U5832 ( .A1(n10175), .A2(n8903), .ZN(n8891) );
  INV_X1 U5833 ( .A(n8393), .ZN(n8866) );
  INV_X1 U5834 ( .A(n8893), .ZN(n8825) );
  AND2_X2 U5835 ( .A1(n9008), .A2(n8908), .ZN(n10314) );
  AND2_X1 U5836 ( .A1(n9045), .A2(n8160), .ZN(n10182) );
  AND2_X1 U5837 ( .A1(n6680), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10186) );
  NOR2_X1 U5838 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n4796) );
  CLKBUF_X1 U5839 ( .A(n6362), .Z(n6363) );
  INV_X1 U5840 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9044) );
  INV_X1 U5841 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8227) );
  OR2_X1 U5842 ( .A1(n6287), .A2(n6286), .ZN(n8225) );
  XNOR2_X1 U5843 ( .A(n6291), .B(n6290), .ZN(n8160) );
  INV_X1 U5844 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U5845 ( .A1(n6311), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6291) );
  INV_X1 U5846 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8057) );
  INV_X1 U5847 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7943) );
  INV_X1 U5848 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7918) );
  INV_X1 U5849 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6323) );
  INV_X1 U5850 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n9077) );
  INV_X1 U5851 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7516) );
  INV_X1 U5852 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7387) );
  INV_X1 U5853 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7224) );
  INV_X1 U5854 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7153) );
  INV_X1 U5855 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9060) );
  INV_X1 U5856 ( .A(n4552), .ZN(n6032) );
  INV_X1 U5857 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9052) );
  NOR2_X1 U5858 ( .A1(n7001), .A2(n7000), .ZN(n7066) );
  NAND2_X1 U5859 ( .A1(n7038), .A2(n4379), .ZN(n5396) );
  AND4_X1 U5860 ( .A1(n5538), .A2(n5537), .A3(n5536), .A4(n5535), .ZN(n9384)
         );
  CLKBUF_X1 U5861 ( .A(n7612), .Z(n7616) );
  CLKBUF_X1 U5862 ( .A(n7205), .Z(n7206) );
  CLKBUF_X1 U5863 ( .A(n7428), .Z(n7600) );
  NAND2_X1 U5864 ( .A1(n9356), .A2(n6896), .ZN(n4908) );
  INV_X1 U5865 ( .A(n4930), .ZN(n9446) );
  NAND2_X1 U5866 ( .A1(n4923), .A2(n9379), .ZN(n9392) );
  OR2_X1 U5867 ( .A1(n9382), .A2(n9380), .ZN(n4923) );
  AND4_X1 U5868 ( .A1(n5424), .A2(n5423), .A3(n5422), .A4(n5421), .ZN(n7739)
         );
  AND4_X2 U5869 ( .A1(n4996), .A2(n4995), .A3(n4994), .A4(n4993), .ZN(n5313)
         );
  NAND2_X1 U5870 ( .A1(n5340), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4994) );
  NAND2_X1 U5871 ( .A1(n5674), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4996) );
  NAND2_X1 U5872 ( .A1(n7909), .A2(n4379), .ZN(n5579) );
  INV_X1 U5873 ( .A(n9467), .ZN(n9440) );
  INV_X1 U5874 ( .A(n9470), .ZN(n9456) );
  AND2_X1 U5875 ( .A1(n6982), .A2(n6965), .ZN(n9448) );
  INV_X1 U5876 ( .A(n9479), .ZN(n9468) );
  NAND2_X1 U5877 ( .A1(n5028), .A2(n5856), .ZN(n5867) );
  NOR2_X1 U5878 ( .A1(n5855), .A2(n5854), .ZN(n5856) );
  CLKBUF_X1 U5879 ( .A(n5890), .Z(n9920) );
  AND4_X1 U5880 ( .A1(n5271), .A2(n5270), .A3(n5269), .A4(n5268), .ZN(n8313)
         );
  AND4_X1 U5881 ( .A1(n5468), .A2(n5467), .A3(n5466), .A4(n5465), .ZN(n9483)
         );
  INV_X1 U5882 ( .A(n4625), .ZN(n7143) );
  NAND2_X1 U5883 ( .A1(n7144), .A2(n7145), .ZN(n4624) );
  NAND2_X1 U5884 ( .A1(n4865), .A2(n4867), .ZN(n7179) );
  NAND2_X1 U5885 ( .A1(n7177), .A2(n5032), .ZN(n4865) );
  NAND2_X1 U5886 ( .A1(n7861), .A2(n7860), .ZN(n4627) );
  NAND2_X1 U5887 ( .A1(n7863), .A2(n7862), .ZN(n4628) );
  OR2_X1 U5888 ( .A1(n9515), .A2(n4855), .ZN(n4854) );
  INV_X1 U5889 ( .A(n4621), .ZN(n9534) );
  NAND2_X1 U5890 ( .A1(n9532), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n4620) );
  NAND2_X1 U5891 ( .A1(n4850), .A2(n4851), .ZN(n9953) );
  INV_X1 U5892 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8266) );
  AND2_X1 U5893 ( .A1(n5235), .A2(n5234), .ZN(n8323) );
  XNOR2_X1 U5894 ( .A(n9723), .B(n9541), .ZN(n9725) );
  INV_X1 U5895 ( .A(n9726), .ZN(n9542) );
  NAND2_X1 U5896 ( .A1(n5260), .A2(n5259), .ZN(n9731) );
  NAND2_X1 U5897 ( .A1(n4596), .A2(n8303), .ZN(n9601) );
  OR2_X1 U5898 ( .A1(n9649), .A2(n4940), .ZN(n4935) );
  NAND2_X1 U5899 ( .A1(n4938), .A2(n4942), .ZN(n9622) );
  NAND2_X1 U5900 ( .A1(n9649), .A2(n4390), .ZN(n4938) );
  NAND2_X1 U5901 ( .A1(n5632), .A2(n5631), .ZN(n9755) );
  NAND2_X1 U5902 ( .A1(n4485), .A2(n4483), .ZN(n9753) );
  INV_X1 U5903 ( .A(n4484), .ZN(n4483) );
  NAND2_X1 U5904 ( .A1(n4486), .A2(n10043), .ZN(n4485) );
  OAI22_X1 U5905 ( .A1(n9625), .A2(n10018), .B1(n10040), .B2(n9624), .ZN(n4484) );
  NAND2_X1 U5906 ( .A1(n8298), .A2(n8297), .ZN(n9642) );
  OR2_X1 U5907 ( .A1(n9649), .A2(n8275), .ZN(n4943) );
  NAND2_X1 U5908 ( .A1(n5599), .A2(n5598), .ZN(n9770) );
  NAND2_X1 U5909 ( .A1(n4577), .A2(n4578), .ZN(n9663) );
  OR2_X1 U5910 ( .A1(n9694), .A2(n4581), .ZN(n4577) );
  NAND2_X1 U5911 ( .A1(n8293), .A2(n9693), .ZN(n9680) );
  NAND2_X1 U5912 ( .A1(n4947), .A2(n4951), .ZN(n9687) );
  NAND2_X1 U5913 ( .A1(n8270), .A2(n4948), .ZN(n4947) );
  INV_X1 U5914 ( .A(n4950), .ZN(n4948) );
  NAND2_X1 U5915 ( .A1(n4952), .A2(n4401), .ZN(n9703) );
  OR2_X1 U5916 ( .A1(n8270), .A2(n8269), .ZN(n4952) );
  AOI21_X1 U5917 ( .B1(n8193), .B2(n4961), .A(n4960), .ZN(n8230) );
  AND2_X1 U5918 ( .A1(n5531), .A2(n5530), .ZN(n8216) );
  NAND2_X1 U5919 ( .A1(n4571), .A2(n4372), .ZN(n4570) );
  NAND2_X1 U5920 ( .A1(n9983), .A2(n7562), .ZN(n7686) );
  AND2_X1 U5921 ( .A1(n7568), .A2(n4387), .ZN(n10020) );
  NAND2_X1 U5922 ( .A1(n5002), .A2(n5789), .ZN(n10012) );
  NAND2_X1 U5923 ( .A1(n5740), .A2(n4568), .ZN(n5002) );
  NAND2_X1 U5924 ( .A1(n5564), .A2(n4500), .ZN(n4499) );
  AND2_X2 U5925 ( .A1(n7200), .A2(n7192), .ZN(n10129) );
  AND2_X1 U5926 ( .A1(n6976), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7040) );
  NAND2_X1 U5927 ( .A1(n7040), .A2(n7188), .ZN(n10062) );
  NOR2_X1 U5928 ( .A1(n4396), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4587) );
  INV_X1 U5929 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8224) );
  INV_X1 U5930 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7977) );
  INV_X1 U5931 ( .A(n5868), .ZN(n7913) );
  INV_X1 U5932 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7911) );
  INV_X1 U5933 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9250) );
  XNOR2_X1 U5934 ( .A(n5059), .B(n5049), .ZN(n7754) );
  INV_X1 U5935 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9137) );
  INV_X1 U5936 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9300) );
  INV_X1 U5937 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7155) );
  INV_X1 U5938 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9107) );
  INV_X1 U5939 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9046) );
  INV_X1 U5940 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9049) );
  INV_X1 U5941 ( .A(n7178), .ZN(n7176) );
  INV_X1 U5942 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5061) );
  XNOR2_X1 U5943 ( .A(n5327), .B(n5326), .ZN(n7046) );
  NAND2_X1 U5944 ( .A1(n5050), .A2(n5043), .ZN(n4844) );
  NAND2_X1 U5945 ( .A1(n5329), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n4845) );
  XNOR2_X1 U5946 ( .A(n5308), .B(n5303), .ZN(n4528) );
  NOR2_X1 U5947 ( .A1(n10315), .A2(n9865), .ZN(n10357) );
  XNOR2_X1 U5948 ( .A(n9877), .B(n4527), .ZN(n10343) );
  XNOR2_X1 U5949 ( .A(n9880), .B(n4526), .ZN(n10348) );
  NOR2_X1 U5950 ( .A1(n10340), .A2(n4472), .ZN(n10339) );
  NOR2_X1 U5951 ( .A1(n10339), .A2(n10338), .ZN(n10337) );
  AND2_X1 U5952 ( .A1(n4525), .A2(n4524), .ZN(n10336) );
  NAND2_X1 U5953 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n4524) );
  INV_X1 U5954 ( .A(n10337), .ZN(n4525) );
  NAND2_X1 U5955 ( .A1(n10336), .A2(n10335), .ZN(n10334) );
  OAI21_X1 U5956 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10334), .ZN(n10332) );
  NAND2_X1 U5957 ( .A1(n10332), .A2(n10333), .ZN(n10331) );
  NAND2_X1 U5958 ( .A1(n10331), .A2(n4522), .ZN(n10329) );
  NAND2_X1 U5959 ( .A1(n7471), .A2(n4523), .ZN(n4522) );
  INV_X1 U5960 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n4523) );
  OAI21_X1 U5961 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10328), .ZN(n10326) );
  NAND2_X1 U5962 ( .A1(n7547), .A2(n7546), .ZN(n7545) );
  OAI21_X1 U5963 ( .B1(n6691), .B2(n8459), .A(n6690), .ZN(n6692) );
  NAND2_X1 U5964 ( .A1(n4672), .A2(n4760), .ZN(n4671) );
  AOI21_X1 U5965 ( .B1(n4669), .B2(n8620), .A(n4667), .ZN(n4666) );
  OAI22_X1 U5966 ( .A1(n8615), .A2(n10165), .B1(n8616), .B2(n10167), .ZN(n4672) );
  INV_X1 U5967 ( .A(n8391), .ZN(n8392) );
  INV_X1 U5968 ( .A(n4733), .ZN(n4732) );
  NAND2_X1 U5969 ( .A1(n10288), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4731) );
  NOR2_X1 U5970 ( .A1(n4733), .A2(n4729), .ZN(n4649) );
  AOI211_X1 U5971 ( .C1(n9778), .C2(n9470), .A(n9351), .B(n9350), .ZN(n9352)
         );
  AOI222_X1 U5972 ( .A1(n9994), .A2(n10050), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n10047), .C1(n10009), .C2(n9993), .ZN(n9999) );
  NAND2_X1 U5973 ( .A1(n4489), .A2(n4487), .ZN(P1_U3547) );
  OR2_X1 U5974 ( .A1(n10143), .A2(n4488), .ZN(n4487) );
  INV_X1 U5975 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n4488) );
  OAI21_X1 U5976 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9888), .A(n10349), .ZN(
        n9890) );
  OR2_X1 U5977 ( .A1(n8757), .A2(n8428), .ZN(n5019) );
  NAND2_X1 U5978 ( .A1(n6896), .A2(n6905), .ZN(n4389) );
  AND2_X1 U5979 ( .A1(n4436), .A2(n4944), .ZN(n4390) );
  INV_X1 U5980 ( .A(n4997), .ZN(n5819) );
  AND2_X1 U5981 ( .A1(n9626), .A2(n4973), .ZN(n4391) );
  AND2_X1 U5982 ( .A1(n4635), .A2(n5019), .ZN(n4392) );
  OR2_X1 U5983 ( .A1(n8935), .A2(n8689), .ZN(n4393) );
  INV_X1 U5984 ( .A(n5019), .ZN(n4817) );
  OR2_X1 U5985 ( .A1(n8632), .A2(n4382), .ZN(n4394) );
  INV_X1 U5986 ( .A(n6350), .ZN(n4645) );
  AND4_X1 U5987 ( .A1(n4452), .A2(n4566), .A3(n6556), .A4(n4564), .ZN(n4395)
         );
  OR2_X1 U5988 ( .A1(n9750), .A2(n9625), .ZN(n8302) );
  NAND2_X1 U5989 ( .A1(n5237), .A2(n5240), .ZN(n4396) );
  NOR2_X1 U5990 ( .A1(n8276), .A2(n4390), .ZN(n4397) );
  AND4_X1 U5991 ( .A1(n5900), .A2(n5901), .A3(n6320), .A4(n6116), .ZN(n4398)
         );
  INV_X1 U5992 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5913) );
  AND2_X1 U5993 ( .A1(n5132), .A2(SI_14_), .ZN(n4399) );
  XNOR2_X1 U5994 ( .A(n5131), .B(SI_14_), .ZN(n5492) );
  NAND2_X1 U5995 ( .A1(n4963), .A2(n7694), .ZN(n7695) );
  INV_X1 U5996 ( .A(n7626), .ZN(n4966) );
  AND2_X1 U5997 ( .A1(n6373), .A2(n6419), .ZN(n4400) );
  OR2_X1 U5998 ( .A1(n8268), .A2(n9436), .ZN(n4401) );
  INV_X1 U5999 ( .A(n4537), .ZN(n7017) );
  NAND2_X1 U6000 ( .A1(n5868), .A2(n7910), .ZN(n4537) );
  AND2_X1 U6001 ( .A1(n5009), .A2(n8299), .ZN(n4402) );
  AND2_X1 U6002 ( .A1(n9778), .A2(n9717), .ZN(n4403) );
  NAND2_X1 U6003 ( .A1(n5383), .A2(n5091), .ZN(n4404) );
  AND2_X1 U6004 ( .A1(n6897), .A2(n6905), .ZN(n4405) );
  INV_X1 U6005 ( .A(n4878), .ZN(n4877) );
  INV_X1 U6006 ( .A(n4962), .ZN(n4960) );
  NAND2_X1 U6007 ( .A1(n9798), .A2(n9480), .ZN(n4962) );
  AND2_X1 U6008 ( .A1(n4818), .A2(n6197), .ZN(n4406) );
  INV_X1 U6009 ( .A(n9688), .ZN(n4983) );
  AND2_X1 U6010 ( .A1(n5114), .A2(n5111), .ZN(n4407) );
  AND4_X1 U6011 ( .A1(n6552), .A2(n4400), .A3(n6545), .A4(n6457), .ZN(n4408)
         );
  OR3_X1 U6012 ( .A1(n5713), .A2(n5847), .A3(n5716), .ZN(n4409) );
  NAND2_X1 U6013 ( .A1(n4935), .A2(n4939), .ZN(n9608) );
  NAND2_X1 U6014 ( .A1(n6829), .A2(n6828), .ZN(n4410) );
  NAND2_X1 U6015 ( .A1(n8719), .A2(n8427), .ZN(n4411) );
  INV_X1 U6016 ( .A(n8293), .ZN(n4583) );
  NAND2_X1 U6017 ( .A1(n4943), .A2(n4944), .ZN(n9633) );
  NAND2_X1 U6018 ( .A1(n8193), .A2(n8192), .ZN(n8207) );
  INV_X1 U6019 ( .A(n4647), .ZN(n4646) );
  NAND2_X1 U6020 ( .A1(n8707), .A2(n4411), .ZN(n4647) );
  OR2_X1 U6021 ( .A1(n4922), .A2(n9380), .ZN(n4412) );
  AND2_X1 U6022 ( .A1(n4546), .A2(n6854), .ZN(n4413) );
  AND3_X1 U6023 ( .A1(n6660), .A2(n6659), .A3(n8734), .ZN(n4414) );
  INV_X1 U6024 ( .A(n10263), .ZN(n4838) );
  AND2_X1 U6025 ( .A1(n5129), .A2(n5128), .ZN(n4415) );
  OR2_X1 U6026 ( .A1(n4385), .A2(n7385), .ZN(n4416) );
  INV_X1 U6027 ( .A(n8835), .ZN(n4802) );
  XOR2_X1 U6028 ( .A(n6925), .B(n6924), .Z(n4417) );
  NAND2_X1 U6029 ( .A1(n9763), .A2(n9667), .ZN(n8297) );
  INV_X1 U6030 ( .A(n8297), .ZN(n5011) );
  NAND2_X1 U6031 ( .A1(n5701), .A2(n5700), .ZN(n9570) );
  INV_X1 U6032 ( .A(n9570), .ZN(n4972) );
  AND2_X1 U6033 ( .A1(n6537), .A2(n4382), .ZN(n4418) );
  OR2_X1 U6034 ( .A1(n9819), .A2(n8000), .ZN(n4419) );
  NAND2_X1 U6035 ( .A1(n6664), .A2(n6663), .ZN(n8467) );
  OR2_X1 U6036 ( .A1(n8673), .A2(n8475), .ZN(n4420) );
  AND2_X1 U6037 ( .A1(n6534), .A2(n4400), .ZN(n4421) );
  AND2_X1 U6038 ( .A1(n4839), .A2(n4838), .ZN(n4422) );
  NOR2_X1 U6039 ( .A1(n8533), .A2(n7854), .ZN(n4423) );
  INV_X1 U6040 ( .A(n8228), .ZN(n9795) );
  AND2_X1 U6041 ( .A1(n5290), .A2(n5289), .ZN(n8228) );
  AND4_X1 U6042 ( .A1(n5659), .A2(n5658), .A3(n5657), .A4(n5656), .ZN(n9625)
         );
  AND2_X1 U6043 ( .A1(n4973), .A2(n4972), .ZN(n4424) );
  AND2_X1 U6044 ( .A1(n6611), .A2(n6610), .ZN(n4425) );
  INV_X1 U6045 ( .A(n9773), .ZN(n4987) );
  NAND2_X1 U6046 ( .A1(n6263), .A2(n6262), .ZN(n8657) );
  AND2_X1 U6047 ( .A1(n10076), .A2(n4966), .ZN(n4426) );
  OR2_X1 U6048 ( .A1(n5572), .A2(n5161), .ZN(n4427) );
  INV_X1 U6049 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5049) );
  INV_X1 U6050 ( .A(n9739), .ZN(n9587) );
  NAND2_X1 U6051 ( .A1(n5687), .A2(n5686), .ZN(n9739) );
  NAND2_X1 U6052 ( .A1(n6135), .A2(n6134), .ZN(n8984) );
  NAND2_X1 U6053 ( .A1(n9626), .A2(n4975), .ZN(n4976) );
  AND2_X1 U6054 ( .A1(n8595), .A2(n8610), .ZN(n4428) );
  INV_X1 U6055 ( .A(n4493), .ZN(n8639) );
  NAND2_X1 U6056 ( .A1(n4494), .A2(n4674), .ZN(n4493) );
  INV_X1 U6057 ( .A(n7964), .ZN(n4813) );
  AND2_X1 U6058 ( .A1(n5000), .A2(n5787), .ZN(n4429) );
  AND2_X1 U6059 ( .A1(n4641), .A2(n4640), .ZN(n4430) );
  INV_X1 U6060 ( .A(n9750), .ZN(n8277) );
  NAND2_X1 U6061 ( .A1(n5654), .A2(n5653), .ZN(n9750) );
  AND2_X1 U6062 ( .A1(n9758), .A2(n9657), .ZN(n4431) );
  AND2_X1 U6063 ( .A1(n6544), .A2(n6418), .ZN(n4750) );
  AND2_X1 U6064 ( .A1(n4726), .A2(n4727), .ZN(n4432) );
  OR2_X1 U6065 ( .A1(n9743), .A2(n9612), .ZN(n8305) );
  INV_X1 U6066 ( .A(n5007), .ZN(n5006) );
  AND2_X1 U6067 ( .A1(n4797), .A2(n6385), .ZN(n4433) );
  INV_X1 U6068 ( .A(n9804), .ZN(n8188) );
  NAND2_X1 U6069 ( .A1(n5498), .A2(n5497), .ZN(n9804) );
  AND2_X1 U6070 ( .A1(n4543), .A2(n6851), .ZN(n4434) );
  INV_X1 U6071 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5043) );
  NOR2_X1 U6072 ( .A1(n8532), .A2(n7933), .ZN(n4435) );
  OR2_X1 U6073 ( .A1(n9758), .A2(n9657), .ZN(n4436) );
  INV_X1 U6074 ( .A(n8384), .ZN(n8385) );
  INV_X1 U6075 ( .A(n4984), .ZN(n9650) );
  NOR2_X1 U6076 ( .A1(n9688), .A2(n4985), .ZN(n4984) );
  AND2_X1 U6077 ( .A1(n9692), .A2(n8271), .ZN(n4437) );
  AND2_X1 U6078 ( .A1(n5792), .A2(n9969), .ZN(n7688) );
  OR2_X1 U6079 ( .A1(n4639), .A2(n4819), .ZN(n4438) );
  NAND2_X1 U6080 ( .A1(n8384), .A2(n8821), .ZN(n4729) );
  NOR2_X1 U6081 ( .A1(n9755), .A2(n9476), .ZN(n4439) );
  OR2_X1 U6082 ( .A1(n9773), .A2(n9666), .ZN(n8294) );
  INV_X1 U6083 ( .A(n8294), .ZN(n4579) );
  NAND2_X1 U6084 ( .A1(n5221), .A2(n5885), .ZN(n4440) );
  NOR2_X1 U6085 ( .A1(n8705), .A2(n8496), .ZN(n4441) );
  NOR2_X1 U6086 ( .A1(n8924), .A2(n8657), .ZN(n4442) );
  INV_X1 U6087 ( .A(n5017), .ZN(n4787) );
  OR2_X1 U6088 ( .A1(n5038), .A2(n7596), .ZN(n4443) );
  INV_X1 U6089 ( .A(n4778), .ZN(n4777) );
  NAND2_X1 U6090 ( .A1(n4782), .A2(n4781), .ZN(n4778) );
  AND2_X1 U6091 ( .A1(n4908), .A2(n4910), .ZN(n4444) );
  AND2_X1 U6092 ( .A1(n9589), .A2(n5777), .ZN(n4445) );
  AND2_X1 U6093 ( .A1(n4878), .A2(n5492), .ZN(n4446) );
  INV_X1 U6094 ( .A(n5330), .ZN(n4846) );
  NAND2_X1 U6095 ( .A1(n9702), .A2(n4953), .ZN(n4447) );
  AND2_X1 U6096 ( .A1(n8741), .A2(n8751), .ZN(n6196) );
  OR2_X1 U6097 ( .A1(n6652), .A2(n6653), .ZN(n4536) );
  NAND2_X1 U6098 ( .A1(n5955), .A2(n4492), .ZN(n10150) );
  AND2_X1 U6099 ( .A1(n4874), .A2(n5492), .ZN(n4448) );
  AND3_X1 U6100 ( .A1(n6152), .A2(n5899), .A3(n6117), .ZN(n4449) );
  OR2_X1 U6101 ( .A1(n4838), .A2(n7967), .ZN(n4450) );
  AND2_X1 U6102 ( .A1(n4644), .A2(n4643), .ZN(n4451) );
  AND2_X1 U6103 ( .A1(n6529), .A2(n6530), .ZN(n4452) );
  AND2_X1 U6104 ( .A1(n5612), .A2(n5611), .ZN(n9654) );
  INV_X1 U6105 ( .A(n9654), .ZN(n9763) );
  AND2_X1 U6106 ( .A1(n6448), .A2(n4400), .ZN(n4453) );
  AND2_X1 U6107 ( .A1(n6557), .A2(n6524), .ZN(n4454) );
  AND2_X1 U6108 ( .A1(n7721), .A2(n4915), .ZN(n4455) );
  AND2_X1 U6109 ( .A1(n6627), .A2(n4787), .ZN(n4456) );
  INV_X1 U6110 ( .A(n6905), .ZN(n4909) );
  NAND2_X1 U6111 ( .A1(n8216), .A2(n9384), .ZN(n4457) );
  INV_X1 U6112 ( .A(n8199), .ZN(n4991) );
  OR2_X1 U6113 ( .A1(n9804), .A2(n8189), .ZN(n8199) );
  AND2_X1 U6114 ( .A1(n6533), .A2(n4421), .ZN(n4458) );
  AND2_X1 U6115 ( .A1(n4656), .A2(n8578), .ZN(n4459) );
  AND2_X1 U6116 ( .A1(n4903), .A2(n9362), .ZN(n4910) );
  OR2_X1 U6117 ( .A1(n4785), .A2(n5017), .ZN(n4460) );
  AND2_X1 U6118 ( .A1(n4854), .A2(n4853), .ZN(n4461) );
  INV_X1 U6119 ( .A(n9988), .ZN(n5406) );
  AND4_X1 U6120 ( .A1(n6471), .A2(n6470), .A3(n6469), .A4(n6468), .ZN(n4462)
         );
  AND2_X1 U6121 ( .A1(n6464), .A2(n6463), .ZN(n4463) );
  OR2_X1 U6122 ( .A1(n4403), .A2(n4950), .ZN(n4464) );
  NAND2_X1 U6123 ( .A1(n5352), .A2(n5825), .ZN(n5740) );
  OR2_X1 U6124 ( .A1(n9995), .A2(n10105), .ZN(n7713) );
  INV_X1 U6125 ( .A(n7713), .ZN(n4979) );
  NAND2_X1 U6126 ( .A1(n8200), .A2(n8199), .ZN(n8208) );
  NAND2_X1 U6127 ( .A1(n5004), .A2(n7813), .ZN(n7902) );
  INV_X1 U6128 ( .A(n6716), .ZN(n5869) );
  INV_X1 U6129 ( .A(n8974), .ZN(n4835) );
  INV_X1 U6130 ( .A(n9379), .ZN(n4921) );
  NAND2_X1 U6131 ( .A1(n4675), .A2(n6254), .ZN(n8924) );
  INV_X1 U6132 ( .A(n8924), .ZN(n4674) );
  NAND2_X1 U6133 ( .A1(n8843), .A2(n4833), .ZN(n4837) );
  OR2_X1 U6134 ( .A1(n7676), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4465) );
  INV_X1 U6135 ( .A(n9528), .ZN(n4853) );
  AND2_X1 U6136 ( .A1(n6459), .A2(n8876), .ZN(n8102) );
  OR2_X1 U6137 ( .A1(n9587), .A2(n9456), .ZN(n4466) );
  OR2_X1 U6138 ( .A1(n7676), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4467) );
  AND2_X1 U6139 ( .A1(n4851), .A2(n4849), .ZN(n4468) );
  AND2_X1 U6140 ( .A1(n4924), .A2(n4410), .ZN(n4469) );
  NAND2_X1 U6141 ( .A1(n6568), .A2(n6413), .ZN(n8886) );
  INV_X1 U6142 ( .A(n8886), .ZN(n8821) );
  INV_X1 U6143 ( .A(n9976), .ZN(n4981) );
  AND2_X2 U6144 ( .A1(n9008), .A2(n9007), .ZN(n10290) );
  NAND2_X1 U6145 ( .A1(n7140), .A2(n7139), .ZN(n7177) );
  AND2_X1 U6146 ( .A1(n7085), .A2(n9926), .ZN(n9957) );
  INV_X1 U6147 ( .A(n9957), .ZN(n4632) );
  AND2_X1 U6148 ( .A1(n5970), .A2(n5969), .ZN(n7850) );
  NAND2_X1 U6149 ( .A1(n6716), .A2(n10011), .ZN(n6972) );
  INV_X1 U6150 ( .A(n6972), .ZN(n4883) );
  NAND4_X1 U6151 ( .A1(n5357), .A2(n5033), .A3(n5356), .A4(n5355), .ZN(n5364)
         );
  AND2_X1 U6152 ( .A1(n6615), .A2(n6614), .ZN(n4470) );
  AND2_X1 U6153 ( .A1(n9496), .A2(n7071), .ZN(n9962) );
  AND2_X1 U6154 ( .A1(n4865), .A2(n4862), .ZN(n4471) );
  INV_X1 U6155 ( .A(n4933), .ZN(n7659) );
  NAND2_X1 U6156 ( .A1(n5819), .A2(n4966), .ZN(n4933) );
  AND2_X1 U6157 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n4472) );
  NOR2_X1 U6158 ( .A1(n8251), .A2(n4855), .ZN(n4473) );
  AND2_X1 U6159 ( .A1(n7440), .A2(n6597), .ZN(n4474) );
  INV_X1 U6160 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n4527) );
  INV_X1 U6161 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5877) );
  INV_X1 U6162 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4619) );
  INV_X1 U6163 ( .A(n9935), .ZN(n4500) );
  INV_X1 U6164 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n4526) );
  OR2_X1 U6165 ( .A1(n7010), .A2(n5808), .ZN(n4475) );
  OAI211_X1 U6166 ( .C1(n9338), .C2(n4932), .A(n4931), .B(n4417), .ZN(n4930)
         );
  OAI21_X2 U6167 ( .B1(n5718), .B2(n8308), .A(n5724), .ZN(n5719) );
  XNOR2_X1 U6168 ( .A(n5228), .B(n4911), .ZN(n5890) );
  NAND2_X1 U6169 ( .A1(n4890), .A2(n5723), .ZN(n4889) );
  NAND3_X1 U6170 ( .A1(n5721), .A2(n4894), .A3(n4891), .ZN(n4890) );
  NAND2_X2 U6171 ( .A1(n4476), .A2(n5788), .ZN(n7698) );
  NAND2_X1 U6172 ( .A1(n4584), .A2(n4429), .ZN(n4476) );
  NAND2_X1 U6173 ( .A1(n4884), .A2(n4882), .ZN(n4881) );
  AND2_X1 U6174 ( .A1(n5349), .A2(n4482), .ZN(n4481) );
  INV_X1 U6175 ( .A(n8436), .ZN(n6669) );
  NAND2_X1 U6176 ( .A1(n4684), .A2(n4689), .ZN(n5152) );
  NOR2_X1 U6177 ( .A1(n8467), .A2(n4495), .ZN(n6665) );
  NOR2_X1 U6178 ( .A1(n7234), .A2(n7233), .ZN(n7266) );
  NOR2_X1 U6179 ( .A1(n9506), .A2(n8248), .ZN(n9517) );
  AOI21_X1 U6180 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9956), .A(n9951), .ZN(
        n8253) );
  NAND2_X1 U6181 ( .A1(n4491), .A2(n4473), .ZN(n4850) );
  NAND2_X1 U6182 ( .A1(n9901), .A2(n9919), .ZN(n9906) );
  NAND2_X1 U6183 ( .A1(n7078), .A2(n4848), .ZN(n9901) );
  INV_X1 U6184 ( .A(n9515), .ZN(n4491) );
  NOR2_X1 U6185 ( .A1(n7677), .A2(n7678), .ZN(n7865) );
  NOR2_X1 U6186 ( .A1(n7869), .A2(n7868), .ZN(n8166) );
  NOR2_X1 U6187 ( .A1(n7128), .A2(n7127), .ZN(n7126) );
  NOR2_X1 U6188 ( .A1(n8168), .A2(n8172), .ZN(n8246) );
  NAND2_X1 U6189 ( .A1(n4742), .A2(n8669), .ZN(n4680) );
  NAND2_X1 U6190 ( .A1(n9360), .A2(n4477), .ZN(n6895) );
  NAND2_X1 U6191 ( .A1(n4519), .A2(n9420), .ZN(n6922) );
  NAND2_X1 U6192 ( .A1(n4780), .A2(n8502), .ZN(n4775) );
  NAND2_X1 U6193 ( .A1(n4478), .A2(n4714), .ZN(n4713) );
  NAND2_X1 U6194 ( .A1(n4598), .A2(n8811), .ZN(n4478) );
  NAND2_X1 U6195 ( .A1(n4718), .A2(n4717), .ZN(n4609) );
  NAND2_X1 U6196 ( .A1(n4707), .A2(n6461), .ZN(n4706) );
  AOI21_X1 U6197 ( .B1(n6441), .B2(n6440), .A(n4711), .ZN(n4710) );
  INV_X1 U6198 ( .A(n6176), .ZN(n4639) );
  NOR2_X1 U6199 ( .A1(n6563), .A2(n4716), .ZN(n4715) );
  NAND2_X1 U6200 ( .A1(n6508), .A2(n4613), .ZN(n4612) );
  NAND2_X1 U6201 ( .A1(n4638), .A2(n6197), .ZN(n4636) );
  OAI21_X1 U6202 ( .B1(n6521), .B2(n4720), .A(n4454), .ZN(n4719) );
  OAI211_X1 U6203 ( .C1(n6510), .C2(n8707), .A(n4615), .B(n4611), .ZN(n4610)
         );
  AOI21_X1 U6204 ( .B1(n4939), .B2(n4940), .A(n4937), .ZN(n4936) );
  OR2_X1 U6205 ( .A1(n8267), .A2(n4464), .ZN(n4946) );
  AOI21_X1 U6206 ( .B1(n7689), .B2(n7687), .A(n5021), .ZN(n7690) );
  NAND2_X1 U6207 ( .A1(n7734), .A2(n7693), .ZN(n4963) );
  OAI22_X2 U6208 ( .A1(n9594), .A2(n8280), .B1(n9598), .B2(n9612), .ZN(n9590)
         );
  NOR2_X2 U6209 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5224) );
  OR2_X1 U6211 ( .A1(n5351), .A2(n5061), .ZN(n4482) );
  NAND2_X1 U6212 ( .A1(n4957), .A2(n4955), .ZN(n8267) );
  OAI22_X1 U6213 ( .A1(n8273), .A2(n8272), .B1(n9666), .B2(n4987), .ZN(n9662)
         );
  NAND3_X1 U6214 ( .A1(n9741), .A2(n4515), .A3(n9740), .ZN(n9828) );
  NAND3_X1 U6215 ( .A1(n10002), .A2(n9985), .A3(n7563), .ZN(n7565) );
  AND2_X1 U6216 ( .A1(n5787), .A2(n5788), .ZN(n10002) );
  NAND2_X1 U6217 ( .A1(n4551), .A2(n5882), .ZN(n5884) );
  NAND2_X1 U6218 ( .A1(n9831), .A2(n10143), .ZN(n4489) );
  NAND2_X1 U6219 ( .A1(n9756), .A2(n4490), .ZN(n9831) );
  NAND2_X1 U6220 ( .A1(n5074), .A2(n5073), .ZN(n5346) );
  NAND2_X1 U6221 ( .A1(n8461), .A2(n4770), .ZN(n4769) );
  NAND2_X1 U6222 ( .A1(n7920), .A2(n7919), .ZN(n8007) );
  AND3_X2 U6223 ( .A1(n4846), .A2(n4845), .A3(n4844), .ZN(n9910) );
  NAND2_X1 U6224 ( .A1(n9909), .A2(n7117), .ZN(n7081) );
  INV_X1 U6225 ( .A(n8381), .ZN(n4652) );
  NAND2_X1 U6226 ( .A1(n7058), .A2(n6404), .ZN(n4617) );
  NAND2_X1 U6227 ( .A1(n5442), .A2(n5441), .ZN(n5443) );
  AOI21_X1 U6228 ( .B1(n4540), .B2(n9430), .A(n4907), .ZN(n4542) );
  OAI21_X1 U6229 ( .B1(n9431), .B2(n4389), .A(n4542), .ZN(n9419) );
  NOR2_X1 U6230 ( .A1(n4521), .A2(n4520), .ZN(n4519) );
  OAI21_X1 U6231 ( .B1(n4650), .B2(n4649), .A(n4731), .ZN(P2_U3517) );
  NAND2_X1 U6232 ( .A1(n4673), .A2(n5083), .ZN(n5382) );
  NOR2_X4 U6233 ( .A1(n5022), .A2(n8741), .ZN(n8736) );
  INV_X1 U6234 ( .A(n4494), .ZN(n8658) );
  MUX2_X2 U6235 ( .A(n5412), .B(n5411), .S(n6972), .Z(n5472) );
  MUX2_X2 U6236 ( .A(n5593), .B(n5592), .S(n6972), .Z(n5625) );
  NAND2_X1 U6237 ( .A1(n5352), .A2(n4999), .ZN(n4584) );
  AOI21_X2 U6238 ( .B1(n4496), .B2(n5563), .A(n5562), .ZN(n5591) );
  NAND3_X1 U6239 ( .A1(n5546), .A2(n5545), .A3(n8229), .ZN(n4496) );
  NAND2_X1 U6240 ( .A1(n4633), .A2(n5081), .ZN(n4673) );
  AOI21_X1 U6241 ( .B1(n4887), .B2(n4881), .A(n4880), .ZN(n5680) );
  OAI21_X1 U6242 ( .B1(n4890), .B2(n4475), .A(n4889), .ZN(n4888) );
  AND2_X4 U6243 ( .A1(n8327), .A2(n5261), .ZN(n5339) );
  NAND2_X1 U6244 ( .A1(n9546), .A2(n5026), .ZN(n9547) );
  NAND2_X1 U6245 ( .A1(n5275), .A2(n5148), .ZN(n4684) );
  INV_X1 U6246 ( .A(n9336), .ZN(n4521) );
  AND2_X2 U6247 ( .A1(n4930), .A2(n4929), .ZN(n9443) );
  AND2_X2 U6248 ( .A1(n9420), .A2(n9336), .ZN(n9338) );
  NAND2_X1 U6249 ( .A1(n4605), .A2(n4497), .ZN(n6520) );
  NAND3_X1 U6250 ( .A1(n6517), .A2(n6556), .A3(n6516), .ZN(n4497) );
  AOI21_X2 U6251 ( .B1(n5985), .B2(n4807), .A(n4435), .ZN(n4806) );
  NAND2_X1 U6252 ( .A1(n4612), .A2(n6511), .ZN(n4611) );
  NAND2_X1 U6253 ( .A1(n4610), .A2(n6512), .ZN(n6515) );
  NAND2_X1 U6254 ( .A1(n4609), .A2(n4458), .ZN(n4607) );
  NAND2_X1 U6255 ( .A1(n4713), .A2(n4712), .ZN(n6499) );
  NAND2_X1 U6256 ( .A1(n4642), .A2(n4430), .ZN(n8670) );
  NAND2_X1 U6257 ( .A1(n4671), .A2(n4666), .ZN(P2_U3264) );
  OAI21_X1 U6258 ( .B1(n4651), .B2(n4733), .A(n10290), .ZN(n4650) );
  NOR2_X1 U6259 ( .A1(n4715), .A2(n4704), .ZN(n4703) );
  OAI21_X1 U6260 ( .B1(n4710), .B2(n4453), .A(n4708), .ZN(n6451) );
  NOR3_X1 U6261 ( .A1(n9404), .A2(n9372), .A3(n4417), .ZN(n9373) );
  OR2_X1 U6262 ( .A1(n9742), .A2(n10110), .ZN(n4515) );
  NAND2_X2 U6263 ( .A1(n8274), .A2(n5030), .ZN(n9649) );
  NAND2_X1 U6264 ( .A1(n5233), .A2(n5232), .ZN(n5870) );
  NOR2_X1 U6265 ( .A1(n9584), .A2(n9583), .ZN(n9741) );
  NAND2_X2 U6266 ( .A1(n5363), .A2(n4498), .ZN(n5365) );
  NAND2_X1 U6267 ( .A1(n4597), .A2(n8302), .ZN(n4596) );
  NOR2_X1 U6268 ( .A1(n9581), .A2(n9589), .ZN(n9580) );
  NAND2_X1 U6269 ( .A1(n6787), .A2(n7721), .ZN(n7242) );
  NAND2_X1 U6270 ( .A1(n6782), .A2(n4501), .ZN(n6787) );
  NAND2_X1 U6271 ( .A1(n6821), .A2(n4927), .ZN(n4926) );
  NAND2_X1 U6272 ( .A1(n4538), .A2(n7213), .ZN(n8334) );
  NAND2_X1 U6273 ( .A1(n4539), .A2(n6740), .ZN(n7214) );
  NOR2_X1 U6274 ( .A1(n8163), .A2(n8223), .ZN(n5889) );
  NAND2_X1 U6275 ( .A1(n6754), .A2(n7217), .ZN(n6729) );
  NOR2_X2 U6276 ( .A1(n9340), .A2(n9339), .ZN(n9401) );
  NAND2_X1 U6277 ( .A1(n8851), .A2(n6473), .ZN(n8078) );
  NAND2_X1 U6278 ( .A1(n7883), .A2(n6337), .ZN(n8060) );
  NAND3_X1 U6279 ( .A1(n4503), .A2(n6565), .A3(n4703), .ZN(P2_U3244) );
  NAND3_X1 U6280 ( .A1(n6416), .A2(n7280), .A3(n6415), .ZN(n4503) );
  NAND2_X1 U6281 ( .A1(n4505), .A2(n5077), .ZN(n4633) );
  NAND2_X1 U6282 ( .A1(n5166), .A2(n5165), .ZN(n5610) );
  NAND2_X1 U6283 ( .A1(n4681), .A2(n4685), .ZN(n5595) );
  NAND2_X1 U6284 ( .A1(n5630), .A2(n4701), .ZN(n4694) );
  NAND2_X1 U6285 ( .A1(n4694), .A2(n4699), .ZN(n5668) );
  OAI21_X1 U6286 ( .B1(n8264), .B2(n8263), .A(n4632), .ZN(n4504) );
  INV_X1 U6287 ( .A(n4504), .ZN(n4631) );
  OAI21_X1 U6288 ( .B1(n8918), .B2(n10206), .A(n8916), .ZN(n4733) );
  NAND2_X1 U6289 ( .A1(n5075), .A2(n5346), .ZN(n4505) );
  NAND2_X1 U6290 ( .A1(n8450), .A2(n6646), .ZN(n8461) );
  NOR2_X2 U6291 ( .A1(n4511), .A2(n4509), .ZN(n8436) );
  XNOR2_X1 U6292 ( .A(n6664), .B(n4510), .ZN(n8408) );
  NOR2_X2 U6293 ( .A1(n6672), .A2(n6671), .ZN(n6707) );
  NAND2_X1 U6294 ( .A1(n4769), .A2(n4771), .ZN(n8481) );
  NAND2_X1 U6295 ( .A1(n8460), .A2(n4782), .ZN(n4780) );
  NAND2_X1 U6296 ( .A1(n6922), .A2(n6923), .ZN(n4931) );
  NAND3_X1 U6297 ( .A1(n9335), .A2(n9334), .A3(n4466), .ZN(P1_U3212) );
  NAND2_X1 U6298 ( .A1(n7168), .A2(n7167), .ZN(n7166) );
  NAND2_X1 U6299 ( .A1(n7214), .A2(n7215), .ZN(n4538) );
  NAND2_X1 U6300 ( .A1(n5876), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5879) );
  INV_X1 U6301 ( .A(n6742), .ZN(n4539) );
  OR2_X2 U6302 ( .A1(n6878), .A2(n6877), .ZN(n9431) );
  NOR3_X2 U6303 ( .A1(n9401), .A2(n9400), .A3(n9399), .ZN(n9404) );
  NOR2_X2 U6304 ( .A1(n9338), .A2(n9337), .ZN(n9400) );
  OAI21_X1 U6305 ( .B1(n9356), .B2(n4902), .A(n4900), .ZN(n6913) );
  INV_X1 U6307 ( .A(n9609), .ZN(n4597) );
  NAND2_X2 U6308 ( .A1(n5396), .A2(n5395), .ZN(n10105) );
  AND2_X2 U6309 ( .A1(n8151), .A2(n8145), .ZN(n7842) );
  NAND2_X2 U6310 ( .A1(n8146), .A2(n8147), .ZN(n8151) );
  AND3_X1 U6311 ( .A1(n5908), .A2(n5910), .A3(n5911), .ZN(n4736) );
  NAND2_X2 U6312 ( .A1(n6345), .A2(n6423), .ZN(n8791) );
  NAND2_X1 U6313 ( .A1(n6331), .A2(n7797), .ZN(n7799) );
  NAND2_X1 U6314 ( .A1(n4732), .A2(n4432), .ZN(n9011) );
  NAND2_X1 U6315 ( .A1(n5595), .A2(n5162), .ZN(n5166) );
  AND2_X2 U6316 ( .A1(n4825), .A2(n4512), .ZN(n7032) );
  NAND3_X1 U6317 ( .A1(n4824), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4512) );
  NAND2_X1 U6318 ( .A1(n7848), .A2(n6548), .ZN(n4735) );
  INV_X2 U6319 ( .A(n10150), .ZN(n10212) );
  NAND2_X1 U6320 ( .A1(n7675), .A2(n4467), .ZN(n7677) );
  NAND2_X1 U6321 ( .A1(n7100), .A2(n4869), .ZN(n7128) );
  NOR2_X1 U6322 ( .A1(n9517), .A2(n9516), .ZN(n9515) );
  NAND2_X2 U6323 ( .A1(n5311), .A2(n5310), .ZN(n7079) );
  AND3_X2 U6324 ( .A1(n4552), .A2(n6276), .A3(n5905), .ZN(n5919) );
  AND2_X1 U6325 ( .A1(n6596), .A2(n6601), .ZN(n4789) );
  OAI22_X2 U6326 ( .A1(n8481), .A2(n8480), .B1(n6656), .B2(n6655), .ZN(n8425)
         );
  INV_X4 U6327 ( .A(n5954), .ZN(n6404) );
  NAND2_X2 U6328 ( .A1(n4385), .A2(n4518), .ZN(n5954) );
  NAND3_X1 U6329 ( .A1(n4514), .A2(n5823), .A3(n7632), .ZN(n5352) );
  NAND2_X1 U6330 ( .A1(n5815), .A2(n5018), .ZN(n4514) );
  AND2_X2 U6331 ( .A1(n4912), .A2(n5222), .ZN(n5231) );
  OAI21_X2 U6332 ( .B1(n5524), .B2(n5523), .A(n5137), .ZN(n5287) );
  INV_X1 U6333 ( .A(n4774), .ZN(n4773) );
  OAI21_X2 U6334 ( .B1(n8490), .B2(n6662), .A(n4516), .ZN(n6664) );
  NAND2_X1 U6335 ( .A1(n4545), .A2(n6844), .ZN(n8177) );
  NAND2_X1 U6336 ( .A1(n6793), .A2(n4913), .ZN(n7428) );
  AND3_X2 U6337 ( .A1(n5231), .A2(n5230), .A3(n5237), .ZN(n5239) );
  INV_X2 U6338 ( .A(n8330), .ZN(n5261) );
  NAND2_X2 U6339 ( .A1(n6916), .A2(n6915), .ZN(n9420) );
  NAND2_X1 U6340 ( .A1(n7105), .A2(n7104), .ZN(n7140) );
  NAND2_X1 U6341 ( .A1(n4842), .A2(n4841), .ZN(n8169) );
  AOI21_X1 U6342 ( .B1(n4630), .B2(n10011), .A(n4871), .ZN(n4870) );
  NAND2_X1 U6343 ( .A1(n7272), .A2(n7271), .ZN(n7675) );
  NOR2_X1 U6344 ( .A1(n8245), .A2(n8246), .ZN(n8247) );
  XNOR2_X2 U6345 ( .A(n5348), .B(P1_IR_REG_3__SCAN_IN), .ZN(n7115) );
  OAI21_X1 U6346 ( .B1(n8262), .B2(n9533), .A(n4631), .ZN(n4630) );
  NAND2_X1 U6347 ( .A1(n5330), .A2(n4619), .ZN(n5372) );
  AND2_X4 U6348 ( .A1(n5328), .A2(n5043), .ZN(n5330) );
  NOR2_X1 U6349 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10345), .ZN(n9873) );
  INV_X1 U6350 ( .A(n8246), .ZN(n4842) );
  OAI21_X1 U6351 ( .B1(n8265), .B2(n10011), .A(n4870), .ZN(P1_U3260) );
  NOR2_X1 U6352 ( .A1(n7266), .A2(n4856), .ZN(n7272) );
  AND2_X2 U6353 ( .A1(n4794), .A2(n5950), .ZN(n4552) );
  OAI21_X1 U6354 ( .B1(n8877), .B2(n4725), .A(n4722), .ZN(n8136) );
  NAND2_X2 U6355 ( .A1(n8687), .A2(n6512), .ZN(n8665) );
  NAND2_X1 U6356 ( .A1(n5628), .A2(n4883), .ZN(n4882) );
  NAND2_X1 U6357 ( .A1(n5608), .A2(n8296), .ZN(n5622) );
  OAI22_X2 U6358 ( .A1(n8078), .A2(n6098), .B1(n8853), .B2(n8997), .ZN(n8836)
         );
  OAI21_X1 U6359 ( .B1(n5867), .B2(n4888), .A(n5866), .ZN(n5893) );
  INV_X4 U6360 ( .A(n5975), .ZN(n5994) );
  OAI21_X2 U6361 ( .B1(n5680), .B2(n9600), .A(n5679), .ZN(n5717) );
  XNOR2_X1 U6362 ( .A(n4528), .B(n5304), .ZN(n7056) );
  OAI21_X2 U6363 ( .B1(n8446), .B2(n6642), .A(n4533), .ZN(n8450) );
  NAND2_X1 U6364 ( .A1(n4762), .A2(n4761), .ZN(n7830) );
  NAND2_X1 U6365 ( .A1(n4679), .A2(n4873), .ZN(n5524) );
  NAND2_X2 U6366 ( .A1(n4537), .A2(n6715), .ZN(n6908) );
  INV_X1 U6367 ( .A(n7001), .ZN(n6727) );
  OAI21_X2 U6368 ( .B1(n7428), .B2(n4443), .A(n5016), .ZN(n7612) );
  INV_X2 U6369 ( .A(n5479), .ZN(n5226) );
  NAND2_X2 U6370 ( .A1(n5044), .A2(n5330), .ZN(n5479) );
  NAND2_X2 U6371 ( .A1(n9431), .A2(n9434), .ZN(n9356) );
  NAND2_X1 U6372 ( .A1(n8087), .A2(n4413), .ZN(n4544) );
  NAND2_X1 U6373 ( .A1(n8087), .A2(n6841), .ZN(n4545) );
  NAND2_X1 U6374 ( .A1(n5880), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4550) );
  NAND3_X1 U6375 ( .A1(n4552), .A2(n6276), .A3(n5916), .ZN(n5917) );
  NAND4_X1 U6376 ( .A1(n5905), .A2(n6276), .A3(n4552), .A4(n5913), .ZN(n4757)
         );
  NOR2_X2 U6377 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n6280) );
  NAND2_X1 U6378 ( .A1(n7958), .A2(n7854), .ZN(n6428) );
  NAND4_X1 U6379 ( .A1(n6553), .A2(n6550), .A3(n4559), .A4(n4557), .ZN(n4556)
         );
  NAND3_X1 U6380 ( .A1(n4381), .A2(n6335), .A3(n8063), .ZN(n4560) );
  XNOR2_X2 U6381 ( .A(n4561), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5907) );
  NAND3_X1 U6382 ( .A1(n6557), .A2(n8633), .A3(n4395), .ZN(n4563) );
  NAND3_X1 U6383 ( .A1(n8759), .A2(n8732), .A3(n4645), .ZN(n4565) );
  INV_X1 U6384 ( .A(n5001), .ZN(n4568) );
  NAND2_X1 U6385 ( .A1(n7812), .A2(n5005), .ZN(n4571) );
  XNOR2_X1 U6386 ( .A(n4570), .B(n7978), .ZN(n7903) );
  NAND2_X1 U6387 ( .A1(n7698), .A2(n7702), .ZN(n7705) );
  AND2_X2 U6388 ( .A1(n5044), .A2(n5222), .ZN(n4585) );
  AND2_X1 U6389 ( .A1(n5222), .A2(n4911), .ZN(n4586) );
  NAND4_X2 U6390 ( .A1(n4912), .A2(n4585), .A3(n4587), .A4(n5330), .ZN(n5243)
         );
  NAND4_X1 U6391 ( .A1(n4912), .A2(n4586), .A3(n5044), .A4(n5330), .ZN(n5236)
         );
  NAND2_X1 U6392 ( .A1(n5008), .A2(n5006), .ZN(n9609) );
  NAND2_X1 U6393 ( .A1(n5008), .A2(n4589), .ZN(n4588) );
  NAND2_X1 U6394 ( .A1(n4599), .A2(n6483), .ZN(n4598) );
  NAND2_X1 U6395 ( .A1(n6480), .A2(n4600), .ZN(n4599) );
  NAND3_X1 U6396 ( .A1(n4608), .A2(n4607), .A3(n6540), .ZN(n4606) );
  NAND2_X2 U6397 ( .A1(n6457), .A2(n6458), .ZN(n8879) );
  NAND3_X1 U6398 ( .A1(n4705), .A2(n4462), .A3(n4618), .ZN(n6472) );
  NAND3_X1 U6399 ( .A1(n4706), .A2(n6462), .A3(n4463), .ZN(n4618) );
  AND2_X2 U6400 ( .A1(n4621), .A2(n4620), .ZN(n9959) );
  AND3_X1 U6401 ( .A1(n9938), .A2(n9937), .A3(n9936), .ZN(n9940) );
  OAI22_X2 U6402 ( .A1(n8165), .A2(n8164), .B1(n8167), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n8255) );
  XNOR2_X1 U6403 ( .A(n4633), .B(n5360), .ZN(n7029) );
  NOR2_X1 U6404 ( .A1(n8759), .A2(n4438), .ZN(n4638) );
  NAND2_X1 U6405 ( .A1(n8712), .A2(n4451), .ZN(n4642) );
  NAND3_X1 U6406 ( .A1(n4644), .A2(n4647), .A3(n4643), .ZN(n4641) );
  INV_X2 U6407 ( .A(n6542), .ZN(n4643) );
  AOI21_X2 U6408 ( .B1(n4646), .B2(n4645), .A(n4441), .ZN(n4644) );
  OR3_X2 U6409 ( .A1(n4728), .A2(n8385), .A3(n4652), .ZN(n4651) );
  INV_X1 U6410 ( .A(n7411), .ZN(n4654) );
  OAI21_X1 U6411 ( .B1(n4654), .B2(n4655), .A(n4459), .ZN(n7416) );
  NAND2_X1 U6412 ( .A1(n4661), .A2(n4662), .ZN(n7487) );
  NAND2_X1 U6413 ( .A1(n7421), .A2(n4664), .ZN(n4661) );
  MUX2_X1 U6414 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n7845), .S(n7304), .Z(n7390)
         );
  NOR2_X2 U6415 ( .A1(n5941), .A2(n5950), .ZN(n7304) );
  NAND2_X1 U6416 ( .A1(n8025), .A2(n8024), .ZN(n8593) );
  NAND2_X1 U6417 ( .A1(n7780), .A2(n7761), .ZN(n8021) );
  NAND2_X1 U6418 ( .A1(n4448), .A2(n5461), .ZN(n4679) );
  NAND2_X1 U6419 ( .A1(n5144), .A2(n4682), .ZN(n4681) );
  NAND2_X1 U6420 ( .A1(n5177), .A2(n4692), .ZN(n4691) );
  NAND3_X1 U6421 ( .A1(n6454), .A2(n6453), .A3(n8876), .ZN(n4707) );
  AND2_X1 U6422 ( .A1(n6485), .A2(n6543), .ZN(n4712) );
  AND2_X1 U6423 ( .A1(n8790), .A2(n6484), .ZN(n4714) );
  NAND3_X1 U6424 ( .A1(n6568), .A2(n6567), .A3(n7280), .ZN(n4716) );
  AND2_X2 U6425 ( .A1(n4398), .A2(n4449), .ZN(n6276) );
  NAND3_X1 U6426 ( .A1(n4719), .A2(n6527), .A3(n4452), .ZN(n4718) );
  INV_X1 U6427 ( .A(n4723), .ZN(n4722) );
  OAI21_X1 U6428 ( .B1(n6341), .B2(n4725), .A(n6545), .ZN(n4723) );
  NAND2_X1 U6429 ( .A1(n8136), .A2(n6553), .ZN(n6342) );
  NAND2_X1 U6430 ( .A1(n4734), .A2(n4735), .ZN(n7883) );
  NAND2_X2 U6431 ( .A1(n4736), .A2(n5909), .ZN(n8537) );
  NAND2_X1 U6432 ( .A1(n8665), .A2(n4740), .ZN(n4737) );
  NAND2_X1 U6433 ( .A1(n8665), .A2(n6556), .ZN(n4743) );
  OAI21_X1 U6434 ( .B1(n8791), .B2(n8803), .A(n6418), .ZN(n8778) );
  NAND2_X1 U6435 ( .A1(n8750), .A2(n6351), .ZN(n4755) );
  OR2_X2 U6436 ( .A1(n8750), .A2(n4756), .ZN(n8731) );
  NAND3_X1 U6437 ( .A1(n6568), .A2(n6374), .A3(n6567), .ZN(n4759) );
  NAND2_X1 U6438 ( .A1(n7532), .A2(n4763), .ZN(n4762) );
  AOI21_X1 U6439 ( .B1(n4763), .B2(n4768), .A(n4470), .ZN(n4761) );
  AND2_X1 U6440 ( .A1(n4766), .A2(n4764), .ZN(n4763) );
  NAND2_X1 U6441 ( .A1(n8007), .A2(n4456), .ZN(n4784) );
  NAND2_X1 U6442 ( .A1(n4784), .A2(n4460), .ZN(n8397) );
  NAND2_X1 U6443 ( .A1(n4792), .A2(n7440), .ZN(n7517) );
  NAND2_X1 U6444 ( .A1(n7438), .A2(n6596), .ZN(n7440) );
  NAND2_X1 U6445 ( .A1(n7438), .A2(n4789), .ZN(n4788) );
  AND3_X1 U6446 ( .A1(n4794), .A2(n5950), .A3(n4795), .ZN(n6165) );
  AND3_X1 U6447 ( .A1(n4794), .A2(n5950), .A3(n4793), .ZN(n6277) );
  AND2_X4 U6448 ( .A1(n5927), .A2(n5898), .ZN(n5950) );
  AND4_X2 U6449 ( .A1(n5895), .A2(n5897), .A3(n5896), .A4(n5894), .ZN(n4794)
         );
  NAND2_X1 U6450 ( .A1(n5919), .A2(n4796), .ZN(n9031) );
  NAND2_X1 U6451 ( .A1(n8650), .A2(n6253), .ZN(n8645) );
  NAND2_X1 U6452 ( .A1(n4800), .A2(n4801), .ZN(n6114) );
  NAND2_X1 U6453 ( .A1(n8076), .A2(n6099), .ZN(n4800) );
  NAND2_X1 U6454 ( .A1(n4805), .A2(n4806), .ZN(n7888) );
  NAND2_X1 U6455 ( .A1(n4804), .A2(n7887), .ZN(n4803) );
  INV_X1 U6456 ( .A(n4806), .ZN(n4804) );
  NAND2_X1 U6457 ( .A1(n4808), .A2(n7850), .ZN(n4805) );
  OAI21_X1 U6458 ( .B1(n7850), .B2(n4423), .A(n5985), .ZN(n7926) );
  NAND2_X1 U6459 ( .A1(n8101), .A2(n4809), .ZN(n4810) );
  NAND2_X1 U6460 ( .A1(n7947), .A2(n10218), .ZN(n7949) );
  INV_X1 U6461 ( .A(n6574), .ZN(n10201) );
  NAND3_X1 U6462 ( .A1(n4828), .A2(n4827), .A3(n4826), .ZN(n4825) );
  OR2_X2 U6463 ( .A1(n8713), .A2(n4830), .ZN(n8671) );
  NAND2_X1 U6464 ( .A1(n8843), .A2(n4832), .ZN(n8771) );
  INV_X1 U6465 ( .A(n4837), .ZN(n8781) );
  MUX2_X1 U6466 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9904), .S(n9910), .Z(n4843)
         );
  OR2_X1 U6467 ( .A1(n7079), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4848) );
  INV_X1 U6468 ( .A(n4854), .ZN(n9529) );
  NAND2_X1 U6469 ( .A1(n7177), .A2(n4859), .ZN(n4857) );
  NAND2_X1 U6470 ( .A1(n4857), .A2(n4858), .ZN(n7234) );
  OR2_X1 U6471 ( .A1(n7178), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4867) );
  NOR2_X4 U6472 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5328) );
  OAI211_X1 U6473 ( .C1(n5305), .C2(n5325), .A(n4872), .B(n5323), .ZN(n5071)
         );
  OAI21_X1 U6474 ( .B1(n7033), .B2(n5325), .A(n4872), .ZN(n5326) );
  OAI21_X1 U6475 ( .B1(n5461), .B2(n5460), .A(n5124), .ZN(n5504) );
  NAND2_X1 U6476 ( .A1(n4879), .A2(n4415), .ZN(n4878) );
  NAND2_X1 U6477 ( .A1(n8334), .A2(n8335), .ZN(n8333) );
  NOR2_X1 U6478 ( .A1(n5479), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U6479 ( .A1(n5236), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5229) );
  INV_X1 U6480 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4911) );
  NOR2_X2 U6481 ( .A1(n5881), .A2(n4440), .ZN(n4912) );
  NAND4_X1 U6482 ( .A1(n5225), .A2(n5224), .A3(n5223), .A4(n5872), .ZN(n5881)
         );
  NAND2_X1 U6483 ( .A1(n6787), .A2(n4455), .ZN(n4914) );
  OAI21_X1 U6484 ( .B1(n9382), .B2(n4412), .A(n4919), .ZN(n6878) );
  NAND2_X1 U6485 ( .A1(n4926), .A2(n4925), .ZN(n7995) );
  CLKBUF_X1 U6486 ( .A(n4926), .Z(n4924) );
  NAND2_X1 U6487 ( .A1(n6821), .A2(n7613), .ZN(n7788) );
  NOR2_X1 U6488 ( .A1(n7787), .A2(n4928), .ZN(n4927) );
  INV_X1 U6489 ( .A(n7613), .ZN(n4928) );
  NAND2_X2 U6490 ( .A1(n5890), .A2(n5870), .ZN(n5322) );
  NAND2_X1 U6491 ( .A1(n4934), .A2(n4936), .ZN(n8279) );
  NAND2_X1 U6492 ( .A1(n9649), .A2(n4939), .ZN(n4934) );
  INV_X1 U6493 ( .A(n8273), .ZN(n9676) );
  NAND2_X1 U6494 ( .A1(n8193), .A2(n4958), .ZN(n4957) );
  NAND3_X1 U6495 ( .A1(n9982), .A2(n7687), .A3(n7562), .ZN(n7691) );
  NAND2_X2 U6496 ( .A1(n5829), .A2(n5825), .ZN(n7556) );
  AND4_X2 U6497 ( .A1(n5341), .A2(n5342), .A3(n5344), .A4(n5343), .ZN(n10041)
         );
  NAND3_X1 U6498 ( .A1(n4963), .A2(n7694), .A3(n7696), .ZN(n7817) );
  OAI21_X2 U6499 ( .B1(n9590), .B2(n8307), .A(n8284), .ZN(n9546) );
  NAND2_X2 U6500 ( .A1(n4964), .A2(n4998), .ZN(n4997) );
  INV_X1 U6501 ( .A(n4965), .ZN(n4964) );
  OAI21_X1 U6502 ( .B1(n5333), .B2(n7056), .A(n5312), .ZN(n4965) );
  INV_X1 U6503 ( .A(n8214), .ZN(n4969) );
  NAND3_X1 U6504 ( .A1(n4969), .A2(n4967), .A3(n9711), .ZN(n9704) );
  NOR2_X1 U6505 ( .A1(n8214), .A2(n9798), .ZN(n8194) );
  NAND2_X1 U6506 ( .A1(n9626), .A2(n8277), .ZN(n9613) );
  INV_X1 U6507 ( .A(n4976), .ZN(n9595) );
  NAND3_X1 U6508 ( .A1(n4979), .A2(n7876), .A3(n4977), .ZN(n7823) );
  NAND2_X1 U6509 ( .A1(n4990), .A2(n4988), .ZN(n8237) );
  INV_X1 U6510 ( .A(n4989), .ZN(n4988) );
  OAI21_X1 U6511 ( .B1(n8039), .B2(n4991), .A(n8201), .ZN(n4989) );
  NAND2_X1 U6512 ( .A1(n8046), .A2(n8199), .ZN(n4990) );
  NAND2_X1 U6513 ( .A1(n5397), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U6514 ( .A1(n5361), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4998) );
  NAND2_X1 U6515 ( .A1(n5001), .A2(n5789), .ZN(n5000) );
  OAI21_X1 U6516 ( .B1(n8301), .B2(n8299), .A(n8300), .ZN(n5007) );
  NAND2_X1 U6517 ( .A1(n8040), .A2(n8188), .ZN(n8214) );
  XNOR2_X1 U6518 ( .A(n5088), .B(SI_6_), .ZN(n5385) );
  NAND2_X1 U6519 ( .A1(n6369), .A2(n10226), .ZN(n7853) );
  NAND2_X1 U6520 ( .A1(n8376), .A2(n8363), .ZN(n8374) );
  INV_X1 U6521 ( .A(n6913), .ZN(n6916) );
  CLKBUF_X1 U6522 ( .A(n7883), .Z(n7934) );
  CLKBUF_X1 U6523 ( .A(n7799), .Z(n7953) );
  NAND4_X2 U6524 ( .A1(n5939), .A2(n5938), .A3(n5937), .A4(n5936), .ZN(n10146)
         );
  OR2_X1 U6525 ( .A1(n10017), .A2(n9994), .ZN(n7569) );
  AND2_X1 U6526 ( .A1(n5792), .A2(n7569), .ZN(n7702) );
  OR2_X1 U6527 ( .A1(n8127), .A2(n8138), .ZN(n8856) );
  OR2_X2 U6528 ( .A1(n8771), .A2(n8963), .ZN(n5022) );
  INV_X1 U6529 ( .A(n10105), .ZN(n5407) );
  INV_X1 U6530 ( .A(n7949), .ZN(n6369) );
  NAND2_X1 U6531 ( .A1(n5339), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5367) );
  XNOR2_X1 U6532 ( .A(n6387), .B(n6385), .ZN(n6368) );
  AOI21_X1 U6533 ( .B1(n8394), .B2(n8393), .A(n8392), .ZN(n8395) );
  INV_X1 U6534 ( .A(n8917), .ZN(n8394) );
  OAI21_X1 U6535 ( .B1(n8286), .B2(n8285), .A(n9546), .ZN(n9568) );
  INV_X1 U6536 ( .A(n5907), .ZN(n9034) );
  OAI211_X1 U6537 ( .C1(n9568), .C2(n10110), .A(n8318), .B(n8317), .ZN(n8319)
         );
  AND2_X4 U6538 ( .A1(n7017), .A2(n6715), .ZN(n6758) );
  NAND2_X1 U6539 ( .A1(n7553), .A2(n7655), .ZN(n7634) );
  NAND2_X1 U6540 ( .A1(n7033), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6541 ( .A1(n5305), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5086) );
  OR3_X1 U6542 ( .A1(n9551), .A2(n9548), .A3(n10014), .ZN(n9559) );
  OAI21_X2 U6543 ( .B1(n9966), .B2(n9968), .A(n7692), .ZN(n7734) );
  OR2_X1 U6544 ( .A1(n9704), .A2(n9778), .ZN(n9688) );
  AOI21_X2 U6545 ( .B1(n8060), .B2(n5014), .A(n5013), .ZN(n8877) );
  OR2_X1 U6546 ( .A1(n7032), .A2(n5078), .ZN(n5079) );
  OAI21_X1 U6547 ( .B1(n7032), .B2(n5061), .A(n5060), .ZN(n5076) );
  NAND2_X1 U6548 ( .A1(n7032), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5060) );
  AND2_X1 U6549 ( .A1(n8102), .A2(n6339), .ZN(n5013) );
  AND2_X1 U6550 ( .A1(n8102), .A2(n6338), .ZN(n5014) );
  AND2_X1 U6551 ( .A1(n6052), .A2(n4450), .ZN(n5015) );
  AND2_X1 U6552 ( .A1(n6811), .A2(n7597), .ZN(n5016) );
  INV_X1 U6553 ( .A(n5950), .ZN(n5951) );
  AND2_X1 U6554 ( .A1(n6632), .A2(n6631), .ZN(n5017) );
  AND2_X1 U6555 ( .A1(n5816), .A2(n7634), .ZN(n5018) );
  NAND2_X1 U6556 ( .A1(n7003), .A2(n7002), .ZN(n10043) );
  INV_X1 U6557 ( .A(n10043), .ZN(n10014) );
  AND2_X1 U6558 ( .A1(n4407), .A2(n5427), .ZN(n5020) );
  AND2_X1 U6559 ( .A1(n5407), .A2(n9988), .ZN(n5021) );
  AND2_X1 U6560 ( .A1(n9557), .A2(n9556), .ZN(n5023) );
  AND2_X1 U6561 ( .A1(n6970), .A2(n9448), .ZN(n5024) );
  OR2_X1 U6562 ( .A1(n8923), .A2(n8850), .ZN(n5025) );
  OR2_X1 U6563 ( .A1(n4972), .A2(n9582), .ZN(n5026) );
  NAND2_X1 U6564 ( .A1(n6993), .A2(n6992), .ZN(n5027) );
  AND2_X1 U6565 ( .A1(n5811), .A2(n5810), .ZN(n5028) );
  OR2_X1 U6566 ( .A1(n8313), .A2(n10018), .ZN(n5029) );
  OR2_X1 U6567 ( .A1(n9369), .A2(n9478), .ZN(n5030) );
  NOR2_X1 U6568 ( .A1(n6705), .A2(n6704), .ZN(n5031) );
  OR2_X1 U6569 ( .A1(n7001), .A2(n6730), .ZN(n5034) );
  AND2_X1 U6570 ( .A1(n9570), .A2(n9470), .ZN(n5036) );
  INV_X1 U6571 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5085) );
  AND2_X1 U6572 ( .A1(n5509), .A2(n5487), .ZN(n5037) );
  INV_X1 U6573 ( .A(n8194), .ZN(n8213) );
  INV_X1 U6574 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n5096) );
  INV_X1 U6575 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5080) );
  INV_X1 U6576 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5087) );
  INV_X1 U6577 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5307) );
  INV_X1 U6578 ( .A(n8765), .ZN(n6346) );
  INV_X1 U6579 ( .A(n8077), .ZN(n6098) );
  AND2_X1 U6580 ( .A1(n7598), .A2(n7599), .ZN(n5038) );
  NAND2_X2 U6581 ( .A1(n7575), .A2(n10031), .ZN(n10033) );
  INV_X1 U6582 ( .A(n7937), .ZN(n6335) );
  INV_X1 U6583 ( .A(n8872), .ZN(n8393) );
  NOR2_X1 U6584 ( .A1(n5620), .A2(n5619), .ZN(n5621) );
  NAND2_X1 U6585 ( .A1(n5775), .A2(n5777), .ZN(n5708) );
  INV_X1 U6586 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5901) );
  OR2_X1 U6587 ( .A1(n7596), .A2(n6806), .ZN(n6811) );
  AOI21_X1 U6588 ( .B1(n5717), .B2(n5776), .A(n5708), .ZN(n5712) );
  XNOR2_X1 U6589 ( .A(n6589), .B(n10150), .ZN(n6582) );
  INV_X1 U6590 ( .A(n6200), .ZN(n6202) );
  AND2_X1 U6591 ( .A1(n4645), .A2(n8721), .ZN(n6351) );
  AND2_X1 U6592 ( .A1(n6542), .A2(n6496), .ZN(n6353) );
  INV_X1 U6593 ( .A(n6990), .ZN(n6991) );
  OAI22_X1 U6594 ( .A1(n10016), .A2(n6917), .B1(n10082), .B2(n6908), .ZN(n6759) );
  OR2_X1 U6595 ( .A1(n7138), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7139) );
  OR2_X1 U6596 ( .A1(n7010), .A2(n6971), .ZN(n6977) );
  AND2_X1 U6597 ( .A1(n5681), .A2(n5683), .ZN(n5191) );
  INV_X1 U6598 ( .A(SI_23_), .ZN(n5172) );
  AND2_X1 U6599 ( .A1(n5594), .A2(n5596), .ZN(n5162) );
  INV_X1 U6600 ( .A(n5547), .ZN(n5149) );
  INV_X1 U6601 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U6602 ( .A1(n7033), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6603 ( .A1(n5305), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U6604 ( .A1(n6584), .A2(n6583), .ZN(n6585) );
  NOR2_X1 U6605 ( .A1(n7443), .A2(n6595), .ZN(n6596) );
  NAND2_X1 U6606 ( .A1(n6202), .A2(n6201), .ZN(n6213) );
  INV_X1 U6607 ( .A(n8433), .ZN(n6668) );
  OR2_X1 U6608 ( .A1(n6266), .A2(n8365), .ZN(n6355) );
  OR2_X1 U6609 ( .A1(n6255), .A2(n6709), .ZN(n6266) );
  NAND2_X1 U6610 ( .A1(n6223), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U6611 ( .A1(n6244), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6255) );
  AOI22_X1 U6612 ( .A1(n8635), .A2(n8815), .B1(n8624), .B2(n8521), .ZN(n8384)
         );
  OR2_X1 U6613 ( .A1(n8801), .A2(n8811), .ZN(n8813) );
  INV_X1 U6614 ( .A(n5671), .ZN(n5688) );
  AND2_X1 U6615 ( .A1(n6940), .A2(n6939), .ZN(n9327) );
  INV_X1 U6616 ( .A(n9451), .ZN(n9464) );
  INV_X1 U6617 ( .A(n5239), .ZN(n5232) );
  INV_X1 U6618 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9383) );
  INV_X1 U6619 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6620 ( .A1(n5640), .A2(n5639), .ZN(n5177) );
  NAND2_X1 U6621 ( .A1(n5140), .A2(n5139), .ZN(n5143) );
  NAND2_X1 U6622 ( .A1(n5134), .A2(n5133), .ZN(n5137) );
  NAND2_X1 U6623 ( .A1(n5121), .A2(n5120), .ZN(n5124) );
  NOR2_X1 U6624 ( .A1(n6703), .A2(n6699), .ZN(n6700) );
  OR2_X1 U6625 ( .A1(n7279), .A2(n6686), .ZN(n8902) );
  NAND2_X1 U6626 ( .A1(n6354), .A2(n6328), .ZN(n7279) );
  INV_X1 U6627 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9161) );
  INV_X1 U6628 ( .A(n8351), .ZN(n7538) );
  NAND2_X1 U6629 ( .A1(n6366), .A2(n6365), .ZN(n6367) );
  INV_X1 U6630 ( .A(n10280), .ZN(n10264) );
  INV_X1 U6631 ( .A(n8528), .ZN(n7967) );
  OR2_X1 U6632 ( .A1(n6329), .A2(n8620), .ZN(n8913) );
  NAND2_X1 U6633 ( .A1(n6309), .A2(n6308), .ZN(n6311) );
  OR2_X1 U6634 ( .A1(n9326), .A2(n9327), .ZN(n6941) );
  NAND2_X1 U6635 ( .A1(n5645), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5655) );
  OR2_X1 U6636 ( .A1(n6986), .A2(n6985), .ZN(n9451) );
  OR2_X1 U6637 ( .A1(n6984), .A2(n6983), .ZN(n9467) );
  NAND2_X1 U6638 ( .A1(n5567), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U6639 ( .A1(n7079), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7078) );
  INV_X1 U6640 ( .A(n7268), .ZN(n7676) );
  INV_X1 U6641 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9463) );
  NAND3_X1 U6642 ( .A1(n10126), .A2(n7040), .A3(n7913), .ZN(n10031) );
  INV_X1 U6643 ( .A(n8309), .ZN(n8285) );
  AND2_X1 U6644 ( .A1(n7011), .A2(n9492), .ZN(n9715) );
  INV_X1 U6645 ( .A(n7910), .ZN(n7573) );
  INV_X1 U6646 ( .A(n5881), .ZN(n5882) );
  AND2_X1 U6647 ( .A1(n5143), .A2(n5142), .ZN(n5286) );
  INV_X1 U6648 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5325) );
  INV_X1 U6649 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9899) );
  AND2_X1 U6650 ( .A1(n6305), .A2(n6313), .ZN(n6307) );
  AND2_X1 U6651 ( .A1(n7917), .A2(n4760), .ZN(n6686) );
  OR2_X1 U6652 ( .A1(n8640), .A2(n6257), .ZN(n6263) );
  INV_X1 U6653 ( .A(n5976), .ZN(n6359) );
  INV_X1 U6654 ( .A(n10165), .ZN(n10163) );
  INV_X1 U6655 ( .A(n10166), .ZN(n8588) );
  INV_X1 U6656 ( .A(n10167), .ZN(n10162) );
  AND2_X1 U6657 ( .A1(n6452), .A2(n8104), .ZN(n8063) );
  AND2_X1 U6658 ( .A1(n6315), .A2(n6314), .ZN(n8908) );
  OR2_X1 U6659 ( .A1(n6567), .A2(n6686), .ZN(n10280) );
  AND2_X1 U6660 ( .A1(n8913), .A2(n10269), .ZN(n10206) );
  INV_X1 U6661 ( .A(n10206), .ZN(n10287) );
  AND2_X1 U6662 ( .A1(n6295), .A2(n6313), .ZN(n10174) );
  XNOR2_X1 U6663 ( .A(n6294), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6313) );
  AND2_X1 U6664 ( .A1(n6980), .A2(n6975), .ZN(n7731) );
  AND4_X1 U6665 ( .A1(n5707), .A2(n5706), .A3(n5705), .A4(n5704), .ZN(n9582)
         );
  AND4_X1 U6666 ( .A1(n5618), .A2(n5617), .A3(n5616), .A4(n5615), .ZN(n9667)
         );
  INV_X1 U6667 ( .A(n5690), .ZN(n5571) );
  AND2_X1 U6668 ( .A1(n7085), .A2(n9492), .ZN(n9932) );
  INV_X1 U6669 ( .A(n9932), .ZN(n9950) );
  INV_X1 U6670 ( .A(n9947), .ZN(n9961) );
  INV_X1 U6671 ( .A(n8323), .ZN(n9723) );
  NAND2_X1 U6672 ( .A1(n8302), .A2(n8303), .ZN(n9610) );
  AND2_X1 U6673 ( .A1(n5778), .A2(n8297), .ZN(n9655) );
  AND3_X1 U6674 ( .A1(n8231), .A2(n10004), .A3(n8195), .ZN(n9794) );
  AND2_X1 U6675 ( .A1(n7217), .A2(n7626), .ZN(n7652) );
  AOI21_X1 U6676 ( .B1(n6953), .B2(n6952), .A(n7043), .ZN(n7199) );
  INV_X1 U6677 ( .A(n10093), .ZN(n10110) );
  OR2_X1 U6678 ( .A1(n6972), .A2(n7573), .ZN(n9824) );
  INV_X1 U6679 ( .A(n9824), .ZN(n10126) );
  NOR2_X1 U6680 ( .A1(n7191), .A2(n7190), .ZN(n7200) );
  AND2_X1 U6681 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9883), .ZN(n9884) );
  AND2_X1 U6682 ( .A1(n6307), .A2(n6306), .ZN(n7281) );
  NAND2_X1 U6683 ( .A1(n6683), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10161) );
  INV_X1 U6684 ( .A(n10151), .ZN(n8459) );
  INV_X1 U6685 ( .A(n6692), .ZN(n6693) );
  INV_X1 U6686 ( .A(n8427), .ZN(n8734) );
  NAND2_X1 U6687 ( .A1(n7286), .A2(n6363), .ZN(n10166) );
  OR2_X1 U6688 ( .A1(n7302), .A2(n8383), .ZN(n10167) );
  OR2_X1 U6689 ( .A1(n8618), .A2(n6363), .ZN(n10165) );
  AND2_X1 U6690 ( .A1(n6372), .A2(n8891), .ZN(n8872) );
  NAND2_X1 U6691 ( .A1(n8393), .A2(n6330), .ZN(n8850) );
  INV_X1 U6692 ( .A(n10314), .ZN(n10311) );
  INV_X1 U6693 ( .A(n10290), .ZN(n10288) );
  NOR2_X1 U6694 ( .A1(n10175), .A2(n10174), .ZN(n10180) );
  INV_X1 U6695 ( .A(n10180), .ZN(n10183) );
  INV_X1 U6696 ( .A(n5906), .ZN(n9038) );
  INV_X1 U6697 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8244) );
  INV_X1 U6698 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7158) );
  NAND2_X1 U6699 ( .A1(n9330), .A2(n5024), .ZN(n6996) );
  INV_X1 U6700 ( .A(n9448), .ZN(n9472) );
  INV_X1 U6701 ( .A(n9962), .ZN(n9533) );
  OR2_X1 U6702 ( .A1(P1_U3083), .A2(n7066), .ZN(n9947) );
  NAND2_X1 U6703 ( .A1(n10033), .A2(n10020), .ZN(n9722) );
  INV_X1 U6704 ( .A(n10143), .ZN(n10141) );
  AND2_X2 U6705 ( .A1(n7200), .A2(n7199), .ZN(n10143) );
  OR3_X1 U6706 ( .A1(n9813), .A2(n9812), .A3(n9811), .ZN(n9842) );
  INV_X1 U6707 ( .A(n10129), .ZN(n10127) );
  INV_X1 U6708 ( .A(n10062), .ZN(n10061) );
  AND2_X1 U6709 ( .A1(n9857), .A2(n8163), .ZN(n7043) );
  INV_X1 U6710 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7915) );
  INV_X1 U6711 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9159) );
  INV_X1 U6712 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7065) );
  NOR2_X1 U6713 ( .A1(n10355), .A2(n10354), .ZN(n10353) );
  NOR2_X1 U6714 ( .A1(n10342), .A2(n10341), .ZN(n10340) );
  AND2_X1 U6715 ( .A1(n7281), .A2(n10186), .ZN(P2_U3966) );
  NAND2_X1 U6716 ( .A1(n6694), .A2(n6693), .ZN(P2_U3242) );
  NAND2_X1 U6717 ( .A1(n5025), .A2(n6384), .ZN(P2_U3268) );
  NOR2_X1 U6718 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5042) );
  NOR2_X2 U6719 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5040) );
  NOR2_X2 U6720 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5039) );
  AND4_X2 U6721 ( .A1(n5042), .A2(n5041), .A3(n5040), .A4(n5039), .ZN(n5044)
         );
  NOR2_X1 U6722 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5048) );
  AND4_X2 U6723 ( .A1(n5048), .A2(n5047), .A3(n5046), .A4(n5045), .ZN(n5222)
         );
  INV_X2 U6724 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U6725 ( .A1(n5054), .A2(n5223), .ZN(n5056) );
  INV_X1 U6726 ( .A(n5054), .ZN(n5055) );
  NAND2_X1 U6727 ( .A1(n5055), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n5057) );
  AND2_X2 U6728 ( .A1(n5057), .A2(n5056), .ZN(n5868) );
  NAND2_X1 U6729 ( .A1(n5869), .A2(n5868), .ZN(n7010) );
  XNOR2_X2 U6730 ( .A(n5872), .B(n5058), .ZN(n7910) );
  NAND2_X1 U6731 ( .A1(n5880), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5059) );
  OR2_X1 U6732 ( .A1(n7910), .A2(n7754), .ZN(n5808) );
  XNOR2_X1 U6733 ( .A(n5076), .B(SI_3_), .ZN(n5345) );
  INV_X1 U6734 ( .A(n5345), .ZN(n5075) );
  INV_X4 U6735 ( .A(n7032), .ZN(n5305) );
  INV_X1 U6736 ( .A(SI_2_), .ZN(n5323) );
  NOR2_X1 U6737 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5064) );
  AND2_X1 U6738 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5301) );
  INV_X1 U6739 ( .A(n5301), .ZN(n5063) );
  NAND2_X1 U6740 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5062) );
  OAI21_X1 U6741 ( .B1(n5064), .B2(n5063), .A(n5062), .ZN(n5065) );
  NAND2_X1 U6742 ( .A1(n5305), .A2(n5065), .ZN(n5070) );
  NOR2_X1 U6743 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5067) );
  NAND2_X1 U6744 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5302) );
  NAND2_X1 U6745 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5066) );
  OAI21_X1 U6746 ( .B1(n5067), .B2(n5302), .A(n5066), .ZN(n5068) );
  NAND2_X1 U6747 ( .A1(n7032), .A2(n5068), .ZN(n5069) );
  NAND2_X1 U6748 ( .A1(n5070), .A2(n5069), .ZN(n5324) );
  NAND2_X1 U6749 ( .A1(n5071), .A2(n5324), .ZN(n5074) );
  INV_X1 U6750 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U6751 ( .A1(n5305), .A2(n9048), .ZN(n5072) );
  OAI211_X1 U6752 ( .C1(n5305), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5072), .B(
        SI_2_), .ZN(n5073) );
  NAND2_X1 U6753 ( .A1(n5076), .A2(SI_3_), .ZN(n5077) );
  INV_X1 U6754 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5078) );
  OAI21_X1 U6755 ( .B1(n5305), .B2(n5080), .A(n5079), .ZN(n5082) );
  XNOR2_X1 U6756 ( .A(n5082), .B(SI_4_), .ZN(n5360) );
  INV_X1 U6757 ( .A(n5360), .ZN(n5081) );
  NAND2_X1 U6758 ( .A1(n5082), .A2(SI_4_), .ZN(n5083) );
  OAI21_X1 U6759 ( .B1(n5305), .B2(n5085), .A(n5084), .ZN(n5090) );
  XNOR2_X1 U6760 ( .A(n5090), .B(SI_5_), .ZN(n5371) );
  INV_X1 U6761 ( .A(n5371), .ZN(n5381) );
  NAND2_X1 U6762 ( .A1(n5088), .A2(SI_6_), .ZN(n5091) );
  NAND2_X1 U6763 ( .A1(n5385), .A2(n5091), .ZN(n5092) );
  AND2_X1 U6764 ( .A1(n5092), .A2(n5381), .ZN(n5089) );
  NAND2_X1 U6765 ( .A1(n5382), .A2(n5089), .ZN(n5094) );
  NAND2_X1 U6766 ( .A1(n5090), .A2(SI_5_), .ZN(n5383) );
  BUF_X4 U6767 ( .A(n5305), .Z(n7033) );
  XNOR2_X1 U6768 ( .A(n5098), .B(SI_7_), .ZN(n5392) );
  INV_X1 U6769 ( .A(n5392), .ZN(n5097) );
  NAND2_X1 U6770 ( .A1(n5098), .A2(SI_7_), .ZN(n5099) );
  MUX2_X1 U6771 ( .A(n9052), .B(n9049), .S(n7033), .Z(n5101) );
  INV_X1 U6772 ( .A(SI_8_), .ZN(n5100) );
  NAND2_X1 U6773 ( .A1(n5101), .A2(n5100), .ZN(n5425) );
  INV_X1 U6774 ( .A(n5101), .ZN(n5102) );
  NAND2_X1 U6775 ( .A1(n5102), .A2(SI_8_), .ZN(n5103) );
  NAND2_X1 U6776 ( .A1(n5425), .A2(n5103), .ZN(n5413) );
  INV_X1 U6777 ( .A(n5413), .ZN(n5104) );
  INV_X1 U6778 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5105) );
  MUX2_X1 U6779 ( .A(n5105), .B(n9046), .S(n5192), .Z(n5112) );
  INV_X1 U6780 ( .A(SI_9_), .ZN(n5106) );
  NAND2_X1 U6781 ( .A1(n5112), .A2(n5106), .ZN(n5441) );
  INV_X1 U6782 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5107) );
  MUX2_X1 U6783 ( .A(n5107), .B(n7065), .S(n7033), .Z(n5109) );
  INV_X1 U6784 ( .A(SI_10_), .ZN(n5108) );
  NAND2_X1 U6785 ( .A1(n5109), .A2(n5108), .ZN(n5114) );
  INV_X1 U6786 ( .A(n5109), .ZN(n5110) );
  NAND2_X1 U6787 ( .A1(n5110), .A2(SI_10_), .ZN(n5111) );
  INV_X1 U6788 ( .A(n5112), .ZN(n5113) );
  NAND2_X1 U6789 ( .A1(n5113), .A2(SI_9_), .ZN(n5427) );
  MUX2_X1 U6790 ( .A(n9060), .B(n9107), .S(n5192), .Z(n5116) );
  INV_X1 U6791 ( .A(n5116), .ZN(n5117) );
  NAND2_X1 U6792 ( .A1(n5117), .A2(SI_11_), .ZN(n5118) );
  MUX2_X1 U6793 ( .A(n7153), .B(n7155), .S(n7033), .Z(n5121) );
  INV_X1 U6794 ( .A(n5121), .ZN(n5122) );
  NAND2_X1 U6795 ( .A1(n5122), .A2(SI_12_), .ZN(n5123) );
  MUX2_X1 U6796 ( .A(n7158), .B(n9300), .S(n7033), .Z(n5126) );
  INV_X1 U6797 ( .A(n5126), .ZN(n5127) );
  NAND2_X1 U6798 ( .A1(n5127), .A2(SI_13_), .ZN(n5128) );
  MUX2_X1 U6799 ( .A(n5130), .B(n9137), .S(n5192), .Z(n5131) );
  INV_X1 U6800 ( .A(n5131), .ZN(n5132) );
  MUX2_X1 U6801 ( .A(n7224), .B(n9159), .S(n5192), .Z(n5134) );
  INV_X1 U6802 ( .A(n5134), .ZN(n5135) );
  NAND2_X1 U6803 ( .A1(n5135), .A2(SI_15_), .ZN(n5136) );
  NAND2_X1 U6804 ( .A1(n5137), .A2(n5136), .ZN(n5523) );
  MUX2_X1 U6805 ( .A(n7387), .B(n5138), .S(n5192), .Z(n5140) );
  INV_X1 U6806 ( .A(n5140), .ZN(n5141) );
  NAND2_X1 U6807 ( .A1(n5141), .A2(SI_16_), .ZN(n5142) );
  MUX2_X1 U6808 ( .A(n7516), .B(n5145), .S(n5192), .Z(n5146) );
  INV_X1 U6809 ( .A(n5146), .ZN(n5147) );
  NAND2_X1 U6810 ( .A1(n5147), .A2(SI_17_), .ZN(n5148) );
  MUX2_X1 U6811 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5192), .Z(n5150) );
  NAND2_X1 U6812 ( .A1(n5150), .A2(SI_18_), .ZN(n5151) );
  MUX2_X1 U6813 ( .A(n9077), .B(n9250), .S(n5192), .Z(n5154) );
  INV_X1 U6814 ( .A(SI_19_), .ZN(n5153) );
  NAND2_X1 U6815 ( .A1(n5154), .A2(n5153), .ZN(n5574) );
  INV_X1 U6816 ( .A(n5154), .ZN(n5155) );
  NAND2_X1 U6817 ( .A1(n5155), .A2(SI_19_), .ZN(n5156) );
  NAND2_X1 U6818 ( .A1(n5574), .A2(n5156), .ZN(n5572) );
  MUX2_X1 U6819 ( .A(n7918), .B(n7911), .S(n5192), .Z(n5159) );
  INV_X1 U6820 ( .A(n5159), .ZN(n5157) );
  NAND2_X1 U6821 ( .A1(n5157), .A2(SI_20_), .ZN(n5575) );
  INV_X1 U6822 ( .A(SI_20_), .ZN(n5158) );
  NAND2_X1 U6823 ( .A1(n5159), .A2(n5158), .ZN(n5576) );
  AND2_X1 U6824 ( .A1(n5574), .A2(n5576), .ZN(n5160) );
  MUX2_X1 U6825 ( .A(n7943), .B(n7915), .S(n5192), .Z(n5163) );
  XNOR2_X1 U6826 ( .A(n5163), .B(SI_21_), .ZN(n5596) );
  INV_X1 U6827 ( .A(n5163), .ZN(n5164) );
  NAND2_X1 U6828 ( .A1(n5164), .A2(SI_21_), .ZN(n5165) );
  MUX2_X1 U6829 ( .A(n8244), .B(n7977), .S(n5192), .Z(n5167) );
  NAND2_X1 U6830 ( .A1(n5167), .A2(n9253), .ZN(n5170) );
  INV_X1 U6831 ( .A(n5167), .ZN(n5168) );
  NAND2_X1 U6832 ( .A1(n5168), .A2(SI_22_), .ZN(n5169) );
  NAND2_X1 U6833 ( .A1(n5170), .A2(n5169), .ZN(n5609) );
  INV_X1 U6834 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5171) );
  MUX2_X1 U6835 ( .A(n8057), .B(n5171), .S(n5192), .Z(n5173) );
  NAND2_X1 U6836 ( .A1(n5173), .A2(n5172), .ZN(n5176) );
  INV_X1 U6837 ( .A(n5173), .ZN(n5174) );
  NAND2_X1 U6838 ( .A1(n5174), .A2(SI_23_), .ZN(n5175) );
  MUX2_X1 U6839 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n5192), .Z(n5179) );
  INV_X1 U6840 ( .A(SI_24_), .ZN(n5178) );
  XNOR2_X1 U6841 ( .A(n5179), .B(n5178), .ZN(n5629) );
  INV_X1 U6842 ( .A(n5629), .ZN(n5181) );
  NAND2_X1 U6843 ( .A1(n5179), .A2(SI_24_), .ZN(n5180) );
  MUX2_X1 U6844 ( .A(n8227), .B(n8224), .S(n5192), .Z(n5183) );
  INV_X1 U6845 ( .A(SI_25_), .ZN(n5182) );
  NAND2_X1 U6846 ( .A1(n5183), .A2(n5182), .ZN(n5186) );
  INV_X1 U6847 ( .A(n5183), .ZN(n5184) );
  NAND2_X1 U6848 ( .A1(n5184), .A2(SI_25_), .ZN(n5185) );
  NAND2_X1 U6849 ( .A1(n5186), .A2(n5185), .ZN(n5651) );
  INV_X1 U6850 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9855) );
  MUX2_X1 U6851 ( .A(n9044), .B(n9855), .S(n5192), .Z(n5187) );
  INV_X1 U6852 ( .A(SI_26_), .ZN(n9105) );
  NAND2_X1 U6853 ( .A1(n5187), .A2(n9105), .ZN(n5681) );
  INV_X1 U6854 ( .A(n5187), .ZN(n5188) );
  NAND2_X1 U6855 ( .A1(n5188), .A2(SI_26_), .ZN(n5189) );
  INV_X1 U6856 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9041) );
  MUX2_X1 U6857 ( .A(n9041), .B(n9131), .S(n5192), .Z(n5194) );
  INV_X1 U6858 ( .A(SI_27_), .ZN(n5190) );
  NAND2_X1 U6859 ( .A1(n5194), .A2(n5190), .ZN(n5683) );
  INV_X1 U6860 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8342) );
  INV_X1 U6861 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5193) );
  MUX2_X1 U6862 ( .A(n8342), .B(n5193), .S(n5192), .Z(n5198) );
  XNOR2_X1 U6863 ( .A(n5198), .B(SI_28_), .ZN(n5697) );
  INV_X1 U6864 ( .A(n5194), .ZN(n5195) );
  NAND2_X1 U6865 ( .A1(n5195), .A2(SI_27_), .ZN(n5695) );
  INV_X1 U6866 ( .A(SI_28_), .ZN(n5197) );
  NAND2_X1 U6867 ( .A1(n5198), .A2(n5197), .ZN(n5211) );
  INV_X1 U6868 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8331) );
  INV_X1 U6869 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9292) );
  MUX2_X1 U6870 ( .A(n8331), .B(n9292), .S(n4518), .Z(n5256) );
  INV_X1 U6871 ( .A(SI_29_), .ZN(n5203) );
  NAND2_X1 U6872 ( .A1(n5256), .A2(n5203), .ZN(n5209) );
  INV_X1 U6873 ( .A(n5209), .ZN(n5199) );
  INV_X1 U6874 ( .A(n5256), .ZN(n5202) );
  NAND2_X1 U6875 ( .A1(n5202), .A2(SI_29_), .ZN(n5201) );
  OAI21_X1 U6876 ( .B1(n5258), .B2(n5199), .A(n5201), .ZN(n5200) );
  MUX2_X1 U6877 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n4518), .Z(n5204) );
  NAND2_X1 U6878 ( .A1(n5200), .A2(n5204), .ZN(n5217) );
  NAND2_X1 U6879 ( .A1(n5201), .A2(n5204), .ZN(n5214) );
  OAI21_X1 U6880 ( .B1(n5204), .B2(n5203), .A(n5202), .ZN(n5206) );
  INV_X1 U6881 ( .A(n5204), .ZN(n5210) );
  OAI21_X1 U6882 ( .B1(SI_29_), .B2(n5210), .A(n5256), .ZN(n5205) );
  NAND2_X1 U6883 ( .A1(n5206), .A2(n5205), .ZN(n5207) );
  OAI21_X1 U6884 ( .B1(n5214), .B2(n5211), .A(n5207), .ZN(n5208) );
  INV_X1 U6885 ( .A(n5208), .ZN(n5213) );
  NAND4_X1 U6886 ( .A1(n5215), .A2(n5211), .A3(n5210), .A4(n5209), .ZN(n5212)
         );
  NAND2_X1 U6887 ( .A1(n5249), .A2(SI_30_), .ZN(n5216) );
  MUX2_X1 U6888 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n4518), .Z(n5218) );
  XNOR2_X1 U6889 ( .A(n5218), .B(SI_31_), .ZN(n5219) );
  NOR2_X1 U6890 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5225) );
  NAND2_X1 U6891 ( .A1(n5231), .A2(n5226), .ZN(n5227) );
  NAND2_X1 U6892 ( .A1(n9030), .A2(n5347), .ZN(n5235) );
  NAND2_X1 U6893 ( .A1(n5322), .A2(n4518), .ZN(n5351) );
  INV_X1 U6894 ( .A(n5351), .ZN(n5361) );
  INV_X4 U6895 ( .A(n5528), .ZN(n5699) );
  NAND2_X1 U6896 ( .A1(n5699), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n5234) );
  XNOR2_X2 U6897 ( .A(n5238), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5262) );
  OAI21_X1 U6898 ( .B1(n5239), .B2(n5050), .A(P1_IR_REG_29__SCAN_IN), .ZN(
        n5242) );
  AND2_X2 U6899 ( .A1(n8327), .A2(n8330), .ZN(n5340) );
  BUF_X4 U6900 ( .A(n5340), .Z(n5646) );
  NAND2_X1 U6901 ( .A1(n5646), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U6902 ( .A1(n4480), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5246) );
  AND2_X2 U6903 ( .A1(n5262), .A2(n8330), .ZN(n5397) );
  NAND2_X1 U6904 ( .A1(n4388), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5245) );
  NAND3_X1 U6905 ( .A1(n5247), .A2(n5246), .A3(n5245), .ZN(n8322) );
  OR2_X1 U6906 ( .A1(n7913), .A2(n7910), .ZN(n7002) );
  NOR3_X1 U6907 ( .A1(n5806), .A2(n5869), .A3(n7002), .ZN(n5723) );
  INV_X1 U6908 ( .A(n8322), .ZN(n5254) );
  AND2_X1 U6909 ( .A1(n9723), .A2(n5254), .ZN(n5805) );
  INV_X1 U6910 ( .A(SI_30_), .ZN(n5248) );
  NAND2_X1 U6911 ( .A1(n8326), .A2(n5347), .ZN(n5251) );
  NAND2_X1 U6912 ( .A1(n5699), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5250) );
  INV_X1 U6913 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9200) );
  NAND2_X1 U6914 ( .A1(n4480), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U6915 ( .A1(n5646), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5252) );
  OAI211_X1 U6916 ( .C1(n5604), .C2(n9200), .A(n5253), .B(n5252), .ZN(n9554)
         );
  INV_X1 U6917 ( .A(n9554), .ZN(n5710) );
  NAND2_X1 U6918 ( .A1(n9726), .A2(n5710), .ZN(n5846) );
  NAND2_X1 U6919 ( .A1(n9726), .A2(n5254), .ZN(n5255) );
  INV_X1 U6920 ( .A(n5709), .ZN(n5273) );
  AOI21_X1 U6921 ( .B1(n6972), .B2(n5273), .A(n5806), .ZN(n5722) );
  XNOR2_X1 U6922 ( .A(n5256), .B(SI_29_), .ZN(n5257) );
  NAND2_X1 U6923 ( .A1(n8329), .A2(n4379), .ZN(n5260) );
  NAND2_X1 U6924 ( .A1(n5699), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U6925 ( .A1(n4388), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6926 ( .A1(n4480), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5270) );
  AND2_X4 U6927 ( .A1(n5262), .A2(n5261), .ZN(n5674) );
  INV_X1 U6928 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9374) );
  AND2_X2 U6929 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5366) );
  NAND2_X1 U6930 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n5263) );
  NOR2_X2 U6931 ( .A1(n5398), .A2(n5263), .ZN(n5419) );
  NAND2_X1 U6932 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n5264) );
  OR2_X2 U6933 ( .A1(n5486), .A2(n9268), .ZN(n5509) );
  NAND2_X1 U6934 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n5265) );
  NOR2_X2 U6935 ( .A1(n5509), .A2(n5265), .ZN(n5511) );
  NAND2_X1 U6936 ( .A1(n5511), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5532) );
  OR2_X2 U6937 ( .A1(n5532), .A2(n9463), .ZN(n5534) );
  NOR2_X2 U6938 ( .A1(n5534), .A2(n9383), .ZN(n5291) );
  AND2_X2 U6939 ( .A1(n5291), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5556) );
  AND2_X2 U6940 ( .A1(n5556), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5567) );
  INV_X1 U6941 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5580) );
  OR2_X2 U6942 ( .A1(n5581), .A2(n5580), .ZN(n5600) );
  NOR2_X2 U6943 ( .A1(n9249), .A2(n5600), .ZN(n5613) );
  AND2_X2 U6944 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n5613), .ZN(n5643) );
  AND2_X2 U6945 ( .A1(n5643), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5645) );
  NOR2_X2 U6946 ( .A1(n9374), .A2(n5655), .ZN(n5672) );
  NAND2_X1 U6947 ( .A1(n5672), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U6948 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n5688), .ZN(n5702) );
  INV_X1 U6949 ( .A(n5702), .ZN(n5266) );
  NAND2_X1 U6950 ( .A1(n5266), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9561) );
  INV_X1 U6951 ( .A(n9561), .ZN(n5267) );
  NAND2_X1 U6952 ( .A1(n5674), .A2(n5267), .ZN(n5269) );
  NAND2_X1 U6953 ( .A1(n5646), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6954 ( .A1(n9731), .A2(n8313), .ZN(n5847) );
  INV_X1 U6955 ( .A(n5847), .ZN(n5272) );
  NOR2_X1 U6956 ( .A1(n5774), .A2(n6972), .ZN(n5715) );
  NAND2_X1 U6957 ( .A1(n7436), .A2(n4379), .ZN(n5281) );
  NOR2_X1 U6958 ( .A1(n5479), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5481) );
  INV_X1 U6959 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5276) );
  AND2_X1 U6960 ( .A1(n5481), .A2(n5276), .ZN(n5505) );
  INV_X1 U6961 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U6962 ( .A1(n5505), .A2(n5277), .ZN(n5494) );
  OAI21_X1 U6963 ( .B1(n5525), .B2(P1_IR_REG_15__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5288) );
  INV_X1 U6964 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6965 ( .A1(n5288), .A2(n5278), .ZN(n5279) );
  NAND2_X1 U6966 ( .A1(n5279), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5550) );
  XNOR2_X1 U6967 ( .A(n5550), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9532) );
  AOI22_X1 U6968 ( .A1(n9532), .A2(n5553), .B1(n5699), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n5280) );
  NOR2_X1 U6969 ( .A1(n5291), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5282) );
  OR2_X1 U6970 ( .A1(n5556), .A2(n5282), .ZN(n9395) );
  AOI22_X1 U6971 ( .A1(n4388), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n4480), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U6972 ( .A1(n5646), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5283) );
  OAI211_X1 U6973 ( .C1(n9395), .C2(n5571), .A(n5284), .B(n5283), .ZN(n9716)
         );
  INV_X1 U6974 ( .A(n9716), .ZN(n9436) );
  NAND2_X1 U6975 ( .A1(n9790), .A2(n9436), .ZN(n8289) );
  INV_X1 U6976 ( .A(n8289), .ZN(n5285) );
  NOR2_X1 U6977 ( .A1(n9790), .A2(n9436), .ZN(n8290) );
  XNOR2_X1 U6978 ( .A(n5287), .B(n5286), .ZN(n7277) );
  NAND2_X1 U6979 ( .A1(n7277), .A2(n4379), .ZN(n5290) );
  XNOR2_X1 U6980 ( .A(n5288), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9522) );
  AOI22_X1 U6981 ( .A1(n9522), .A2(n5553), .B1(n5699), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n5289) );
  AND2_X1 U6982 ( .A1(n5534), .A2(n9383), .ZN(n5292) );
  OR2_X1 U6983 ( .A1(n5292), .A2(n5291), .ZN(n9387) );
  NAND2_X1 U6984 ( .A1(n4480), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5293) );
  OAI21_X1 U6985 ( .B1(n9387), .B2(n5571), .A(n5293), .ZN(n5294) );
  INV_X1 U6986 ( .A(n5294), .ZN(n5298) );
  NAND2_X1 U6987 ( .A1(n4388), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5296) );
  NAND2_X1 U6988 ( .A1(n5646), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5295) );
  AND2_X1 U6989 ( .A1(n5296), .A2(n5295), .ZN(n5297) );
  NAND2_X1 U6990 ( .A1(n5298), .A2(n5297), .ZN(n9479) );
  NAND2_X1 U6991 ( .A1(n8228), .A2(n9479), .ZN(n5743) );
  INV_X1 U6992 ( .A(n5743), .ZN(n5299) );
  NAND2_X1 U6993 ( .A1(n9795), .A2(n9468), .ZN(n5729) );
  INV_X1 U6994 ( .A(n5729), .ZN(n8235) );
  MUX2_X1 U6995 ( .A(n5299), .B(n8235), .S(n6972), .Z(n5300) );
  NOR2_X1 U6996 ( .A1(n8238), .A2(n5300), .ZN(n5563) );
  NAND2_X1 U6997 ( .A1(n7033), .A2(n5301), .ZN(n5320) );
  OAI21_X1 U6998 ( .B1(n7033), .B2(n5302), .A(n5320), .ZN(n5304) );
  INV_X1 U6999 ( .A(SI_1_), .ZN(n5303) );
  OAI21_X1 U7000 ( .B1(n7033), .B2(n5307), .A(n5306), .ZN(n5308) );
  INV_X2 U7001 ( .A(n5322), .ZN(n5564) );
  NAND2_X1 U7002 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5309) );
  INV_X1 U7003 ( .A(n5328), .ZN(n5310) );
  INV_X1 U7004 ( .A(n7079), .ZN(n9891) );
  NAND2_X1 U7005 ( .A1(n5564), .A2(n9891), .ZN(n5312) );
  INV_X1 U7006 ( .A(n7650), .ZN(n5786) );
  NAND2_X1 U7007 ( .A1(n5674), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U7008 ( .A1(n5397), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U7009 ( .A1(n5340), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U7010 ( .A1(n5339), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5314) );
  INV_X1 U7011 ( .A(SI_0_), .ZN(n5319) );
  INV_X1 U7012 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5318) );
  OAI21_X1 U7013 ( .B1(n4518), .B2(n5319), .A(n5318), .ZN(n5321) );
  AND2_X1 U7014 ( .A1(n5321), .A2(n5320), .ZN(n9858) );
  MUX2_X1 U7015 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9858), .S(n5322), .Z(n7626) );
  XNOR2_X1 U7016 ( .A(n5324), .B(n5323), .ZN(n5327) );
  NAND2_X1 U7017 ( .A1(n5361), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5332) );
  NOR2_X1 U7018 ( .A1(n5328), .A2(n5050), .ZN(n5329) );
  NAND2_X1 U7019 ( .A1(n5564), .A2(n9910), .ZN(n5331) );
  NAND2_X1 U7020 ( .A1(n5397), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5337) );
  NAND2_X1 U7021 ( .A1(n5674), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U7022 ( .A1(n5340), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U7023 ( .A1(n5339), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5334) );
  AND4_X2 U7024 ( .A1(n5337), .A2(n5336), .A3(n5335), .A4(n5334), .ZN(n7655)
         );
  NAND2_X1 U7025 ( .A1(n5397), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5344) );
  INV_X1 U7026 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U7027 ( .A1(n5674), .A2(n5338), .ZN(n5343) );
  NAND2_X1 U7028 ( .A1(n5339), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U7029 ( .A1(n5340), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5341) );
  XNOR2_X1 U7030 ( .A(n5346), .B(n5345), .ZN(n7030) );
  NAND2_X1 U7031 ( .A1(n4378), .A2(n7030), .ZN(n5350) );
  NAND2_X1 U7032 ( .A1(n5564), .A2(n7115), .ZN(n5349) );
  INV_X1 U7033 ( .A(n7556), .ZN(n7632) );
  INV_X2 U7034 ( .A(n7655), .ZN(n9490) );
  NAND2_X1 U7035 ( .A1(n5339), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5357) );
  INV_X1 U7036 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U7037 ( .A1(n5646), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5356) );
  NOR2_X1 U7038 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5354) );
  NOR2_X1 U7039 ( .A1(n5366), .A2(n5354), .ZN(n10030) );
  NAND2_X1 U7040 ( .A1(n5674), .A2(n10030), .ZN(n5355) );
  NAND2_X1 U7041 ( .A1(n5372), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5359) );
  INV_X1 U7042 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U7043 ( .A1(n7029), .A2(n5347), .ZN(n5363) );
  NAND2_X1 U7044 ( .A1(n5361), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5362) );
  INV_X1 U7045 ( .A(n5365), .ZN(n10082) );
  NAND2_X1 U7046 ( .A1(n5397), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U7047 ( .A1(n5646), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5369) );
  OAI21_X1 U7048 ( .B1(n5366), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5398), .ZN(
        n7591) );
  INV_X1 U7049 ( .A(n7591), .ZN(n10008) );
  NAND2_X1 U7050 ( .A1(n5690), .A2(n10008), .ZN(n5368) );
  NAND4_X4 U7051 ( .A1(n5370), .A2(n5369), .A3(n5368), .A4(n5367), .ZN(n10038)
         );
  XNOR2_X1 U7052 ( .A(n5382), .B(n5371), .ZN(n7036) );
  NAND2_X1 U7053 ( .A1(n7036), .A2(n4379), .ZN(n5376) );
  INV_X1 U7054 ( .A(n5388), .ZN(n5373) );
  NAND2_X1 U7055 ( .A1(n5373), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5374) );
  AOI22_X1 U7056 ( .A1(n5361), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5564), .B2(
        n7101), .ZN(n5375) );
  NAND2_X1 U7057 ( .A1(n10038), .A2(n10090), .ZN(n5787) );
  INV_X1 U7058 ( .A(n10038), .ZN(n9989) );
  NAND2_X1 U7059 ( .A1(n5339), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U7060 ( .A1(n5397), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5379) );
  XNOR2_X1 U7061 ( .A(n5398), .B(P1_REG3_REG_6__SCAN_IN), .ZN(n9993) );
  NAND2_X1 U7062 ( .A1(n5674), .A2(n9993), .ZN(n5378) );
  NAND2_X1 U7063 ( .A1(n5646), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5377) );
  AND4_X2 U7064 ( .A1(n5380), .A2(n5379), .A3(n5378), .A4(n5377), .ZN(n10017)
         );
  NAND2_X1 U7065 ( .A1(n5382), .A2(n5381), .ZN(n5384) );
  NAND2_X1 U7066 ( .A1(n5384), .A2(n5383), .ZN(n5386) );
  XNOR2_X1 U7067 ( .A(n5385), .B(n5386), .ZN(n7037) );
  NAND2_X1 U7068 ( .A1(n7037), .A2(n4379), .ZN(n5391) );
  INV_X1 U7069 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U7070 ( .A1(n5388), .A2(n5387), .ZN(n5394) );
  NAND2_X1 U7071 ( .A1(n5394), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5389) );
  XNOR2_X1 U7072 ( .A(n5389), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7130) );
  AOI22_X1 U7073 ( .A1(n5361), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5553), .B2(
        n7130), .ZN(n5390) );
  NAND2_X1 U7074 ( .A1(n7569), .A2(n7699), .ZN(n7563) );
  XNOR2_X1 U7075 ( .A(n5415), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7138) );
  AOI22_X1 U7076 ( .A1(n5361), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5564), .B2(
        n7138), .ZN(n5395) );
  NAND2_X1 U7077 ( .A1(n5397), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U7078 ( .A1(n5339), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5404) );
  INV_X1 U7079 ( .A(n5398), .ZN(n5399) );
  AOI21_X1 U7080 ( .B1(n5399), .B2(P1_REG3_REG_6__SCAN_IN), .A(
        P1_REG3_REG_7__SCAN_IN), .ZN(n5400) );
  OR2_X1 U7081 ( .A1(n5400), .A2(n5419), .ZN(n7576) );
  INV_X1 U7082 ( .A(n7576), .ZN(n5401) );
  NAND2_X1 U7083 ( .A1(n5674), .A2(n5401), .ZN(n5403) );
  NAND2_X1 U7084 ( .A1(n5646), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U7085 ( .A1(n5407), .A2(n5406), .ZN(n5792) );
  INV_X1 U7086 ( .A(n7702), .ZN(n5408) );
  OAI21_X1 U7087 ( .B1(n9990), .B2(n5408), .A(n9969), .ZN(n5412) );
  INV_X1 U7088 ( .A(n7698), .ZN(n5409) );
  OAI211_X1 U7089 ( .C1(n5409), .C2(n7563), .A(n9969), .B(n7699), .ZN(n5410)
         );
  NAND2_X1 U7090 ( .A1(n5410), .A2(n5792), .ZN(n5411) );
  INV_X1 U7091 ( .A(n5472), .ZN(n5438) );
  NAND2_X1 U7092 ( .A1(n7044), .A2(n4379), .ZN(n5418) );
  NAND2_X1 U7093 ( .A1(n5415), .A2(n5446), .ZN(n5416) );
  NAND2_X1 U7094 ( .A1(n5416), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5428) );
  XNOR2_X1 U7095 ( .A(n5428), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7178) );
  AOI22_X1 U7096 ( .A1(n5699), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7178), .B2(
        n5553), .ZN(n5417) );
  NAND2_X1 U7097 ( .A1(n4388), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U7098 ( .A1(n5646), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5423) );
  OR2_X1 U7099 ( .A1(n5419), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5420) );
  AND2_X1 U7100 ( .A1(n5454), .A2(n5420), .ZN(n9975) );
  NAND2_X1 U7101 ( .A1(n5690), .A2(n9975), .ZN(n5422) );
  NAND2_X1 U7102 ( .A1(n5339), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U7103 ( .A1(n9976), .A2(n7739), .ZN(n5791) );
  NAND2_X1 U7104 ( .A1(n5426), .A2(n5425), .ZN(n5440) );
  AND2_X1 U7105 ( .A1(n5441), .A2(n5427), .ZN(n5439) );
  NAND2_X1 U7106 ( .A1(n9322), .A2(n4379), .ZN(n5432) );
  INV_X1 U7107 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U7108 ( .A1(n5428), .A2(n5445), .ZN(n5429) );
  AOI22_X1 U7109 ( .A1(n7232), .A2(n5553), .B1(n5699), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U7110 ( .A1(n5339), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U7111 ( .A1(n4388), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5435) );
  XNOR2_X1 U7112 ( .A(n5454), .B(P1_REG3_REG_9__SCAN_IN), .ZN(n7746) );
  NAND2_X1 U7113 ( .A1(n5690), .A2(n7746), .ZN(n5434) );
  NAND2_X1 U7114 ( .A1(n5646), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5433) );
  NAND4_X1 U7115 ( .A1(n5436), .A2(n5435), .A3(n5434), .A4(n5433), .ZN(n9487)
         );
  INV_X1 U7116 ( .A(n7706), .ZN(n5437) );
  AOI21_X1 U7117 ( .B1(n5438), .B2(n5791), .A(n5437), .ZN(n5470) );
  NAND2_X1 U7118 ( .A1(n5440), .A2(n5439), .ZN(n5442) );
  NAND2_X1 U7119 ( .A1(n7058), .A2(n4379), .ZN(n5451) );
  INV_X1 U7120 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5444) );
  NAND3_X1 U7121 ( .A1(n5446), .A2(n5445), .A3(n5444), .ZN(n5447) );
  OAI21_X1 U7122 ( .B1(n5448), .B2(n5447), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5449) );
  XNOR2_X1 U7123 ( .A(n5449), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7267) );
  AOI22_X1 U7124 ( .A1(n5699), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5553), .B2(
        n7267), .ZN(n5450) );
  NAND2_X1 U7125 ( .A1(n5339), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7126 ( .A1(n4388), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5458) );
  INV_X1 U7127 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5453) );
  INV_X1 U7128 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5452) );
  OAI21_X1 U7129 ( .B1(n5454), .B2(n5453), .A(n5452), .ZN(n5455) );
  AND2_X1 U7130 ( .A1(n5455), .A2(n5486), .ZN(n7714) );
  NAND2_X1 U7131 ( .A1(n5690), .A2(n7714), .ZN(n5457) );
  NAND2_X1 U7132 ( .A1(n5646), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U7133 ( .A1(n7815), .A2(n7814), .ZN(n5784) );
  NAND2_X1 U7134 ( .A1(n7747), .A2(n9967), .ZN(n7707) );
  AND2_X1 U7135 ( .A1(n5784), .A2(n7707), .ZN(n7811) );
  INV_X1 U7136 ( .A(n7811), .ZN(n5469) );
  XNOR2_X1 U7137 ( .A(n5461), .B(n5460), .ZN(n7152) );
  NAND2_X1 U7138 ( .A1(n7152), .A2(n4379), .ZN(n5464) );
  OR2_X1 U7139 ( .A1(n5481), .A2(n5050), .ZN(n5462) );
  XNOR2_X1 U7140 ( .A(n5462), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7866) );
  AOI22_X1 U7141 ( .A1(n5699), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5553), .B2(
        n7866), .ZN(n5463) );
  NAND2_X1 U7142 ( .A1(n4388), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U7143 ( .A1(n5646), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5467) );
  XNOR2_X1 U7144 ( .A(n5509), .B(P1_REG3_REG_12__SCAN_IN), .ZN(n8002) );
  NAND2_X1 U7145 ( .A1(n5690), .A2(n8002), .ZN(n5466) );
  NAND2_X1 U7146 ( .A1(n5339), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5465) );
  OAI21_X1 U7147 ( .B1(n5470), .B2(n5469), .A(n7983), .ZN(n5476) );
  INV_X1 U7148 ( .A(n7736), .ZN(n5471) );
  OAI211_X1 U7149 ( .C1(n5472), .C2(n5471), .A(n7707), .B(n5791), .ZN(n5473)
         );
  NAND3_X1 U7150 ( .A1(n5473), .A2(n7813), .A3(n5785), .ZN(n5474) );
  NAND2_X1 U7151 ( .A1(n9816), .A2(n9483), .ZN(n7981) );
  NAND3_X1 U7152 ( .A1(n5474), .A2(n7981), .A3(n5784), .ZN(n5475) );
  XNOR2_X1 U7153 ( .A(n5478), .B(n5477), .ZN(n7062) );
  NAND2_X1 U7154 ( .A1(n7062), .A2(n4379), .ZN(n5485) );
  NAND2_X1 U7155 ( .A1(n5479), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5480) );
  MUX2_X1 U7156 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5480), .S(
        P1_IR_REG_11__SCAN_IN), .Z(n5483) );
  INV_X1 U7157 ( .A(n5481), .ZN(n5482) );
  NAND2_X1 U7158 ( .A1(n5483), .A2(n5482), .ZN(n7268) );
  AOI22_X1 U7159 ( .A1(n5699), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5553), .B2(
        n7676), .ZN(n5484) );
  NAND2_X1 U7160 ( .A1(n5339), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U7161 ( .A1(n4388), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U7162 ( .A1(n5486), .A2(n9268), .ZN(n5487) );
  NAND2_X1 U7163 ( .A1(n5690), .A2(n5037), .ZN(n5489) );
  NAND2_X1 U7164 ( .A1(n5646), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5488) );
  NAND4_X1 U7165 ( .A1(n5491), .A2(n5490), .A3(n5489), .A4(n5488), .ZN(n9485)
         );
  OR2_X1 U7166 ( .A1(n9819), .A2(n9485), .ZN(n7899) );
  NAND2_X1 U7167 ( .A1(n9819), .A2(n9485), .ZN(n7897) );
  NAND2_X1 U7168 ( .A1(n7899), .A2(n7897), .ZN(n7818) );
  OAI21_X1 U7169 ( .B1(n7813), .B2(n6972), .A(n7818), .ZN(n5521) );
  INV_X1 U7170 ( .A(n9485), .ZN(n8000) );
  NAND2_X1 U7171 ( .A1(n9819), .A2(n8000), .ZN(n7901) );
  NAND2_X1 U7172 ( .A1(n7981), .A2(n7901), .ZN(n5731) );
  XNOR2_X1 U7173 ( .A(n5493), .B(n5492), .ZN(n7164) );
  NAND2_X1 U7174 ( .A1(n7164), .A2(n5347), .ZN(n5498) );
  NAND2_X1 U7175 ( .A1(n5494), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5495) );
  MUX2_X1 U7176 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5495), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5496) );
  AOI22_X1 U7177 ( .A1(n5699), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5553), .B2(
        n8256), .ZN(n5497) );
  NAND2_X1 U7178 ( .A1(n5339), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U7179 ( .A1(n4388), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5502) );
  OR2_X1 U7180 ( .A1(n5511), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5499) );
  AND2_X1 U7181 ( .A1(n5499), .A2(n5532), .ZN(n8181) );
  NAND2_X1 U7182 ( .A1(n5674), .A2(n8181), .ZN(n5501) );
  NAND2_X1 U7183 ( .A1(n5646), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U7184 ( .A1(n9804), .A2(n8189), .ZN(n5782) );
  XNOR2_X1 U7185 ( .A(n5504), .B(n4415), .ZN(n7157) );
  NAND2_X1 U7186 ( .A1(n7157), .A2(n4379), .ZN(n5508) );
  OR2_X1 U7187 ( .A1(n5505), .A2(n5050), .ZN(n5506) );
  XNOR2_X1 U7188 ( .A(n5506), .B(P1_IR_REG_13__SCAN_IN), .ZN(n8167) );
  AOI22_X1 U7189 ( .A1(n5699), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5564), .B2(
        n8167), .ZN(n5507) );
  NAND2_X1 U7190 ( .A1(n4388), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7191 ( .A1(n4480), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5515) );
  INV_X1 U7192 ( .A(n5509), .ZN(n5510) );
  AOI21_X1 U7193 ( .B1(n5510), .B2(P1_REG3_REG_12__SCAN_IN), .A(
        P1_REG3_REG_13__SCAN_IN), .ZN(n5512) );
  NOR2_X1 U7194 ( .A1(n5512), .A2(n5511), .ZN(n8092) );
  NAND2_X1 U7195 ( .A1(n5690), .A2(n8092), .ZN(n5514) );
  NAND2_X1 U7196 ( .A1(n5646), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U7197 ( .A1(n8036), .A2(n8048), .ZN(n8043) );
  NAND2_X1 U7198 ( .A1(n5782), .A2(n8043), .ZN(n5540) );
  AOI21_X1 U7199 ( .B1(n7983), .B2(n5731), .A(n5540), .ZN(n5519) );
  OR2_X1 U7200 ( .A1(n8036), .A2(n8048), .ZN(n5783) );
  NAND2_X1 U7201 ( .A1(n8199), .A2(n5783), .ZN(n5539) );
  NAND2_X1 U7202 ( .A1(n7983), .A2(n4419), .ZN(n5517) );
  AND2_X1 U7203 ( .A1(n5517), .A2(n7981), .ZN(n5518) );
  NOR2_X1 U7204 ( .A1(n5539), .A2(n5518), .ZN(n5744) );
  MUX2_X1 U7205 ( .A(n5519), .B(n5744), .S(n6972), .Z(n5520) );
  OAI21_X1 U7206 ( .B1(n5522), .B2(n5521), .A(n5520), .ZN(n5544) );
  XNOR2_X1 U7207 ( .A(n5524), .B(n5523), .ZN(n7222) );
  NAND2_X1 U7208 ( .A1(n7222), .A2(n5347), .ZN(n5531) );
  NAND2_X1 U7209 ( .A1(n5525), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5527) );
  INV_X1 U7210 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5526) );
  XNOR2_X1 U7211 ( .A(n5527), .B(n5526), .ZN(n9505) );
  OAI22_X1 U7212 ( .A1(n9505), .A2(n9493), .B1(n5528), .B2(n9159), .ZN(n5529)
         );
  INV_X1 U7213 ( .A(n5529), .ZN(n5530) );
  NAND2_X1 U7214 ( .A1(n4388), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7215 ( .A1(n4480), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U7216 ( .A1(n5532), .A2(n9463), .ZN(n5533) );
  AND2_X1 U7217 ( .A1(n5534), .A2(n5533), .ZN(n9461) );
  NAND2_X1 U7218 ( .A1(n5690), .A2(n9461), .ZN(n5536) );
  NAND2_X1 U7219 ( .A1(n5646), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5535) );
  OR2_X1 U7220 ( .A1(n9798), .A2(n9384), .ZN(n8202) );
  NAND2_X1 U7221 ( .A1(n9798), .A2(n9384), .ZN(n8201) );
  NAND2_X1 U7222 ( .A1(n5539), .A2(n5782), .ZN(n5542) );
  NAND2_X1 U7223 ( .A1(n5540), .A2(n8199), .ZN(n5541) );
  MUX2_X1 U7224 ( .A(n5542), .B(n5541), .S(n6972), .Z(n5543) );
  NAND3_X1 U7225 ( .A1(n5544), .A2(n8209), .A3(n5543), .ZN(n5546) );
  MUX2_X1 U7226 ( .A(n8201), .B(n8202), .S(n6972), .Z(n5545) );
  NAND2_X1 U7227 ( .A1(n7683), .A2(n4379), .ZN(n5555) );
  INV_X1 U7228 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U7229 ( .A1(n5550), .A2(n5549), .ZN(n5551) );
  NAND2_X1 U7230 ( .A1(n5551), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5552) );
  XNOR2_X1 U7231 ( .A(n5552), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9956) );
  AOI22_X1 U7232 ( .A1(n9956), .A2(n5553), .B1(n5699), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n5554) );
  NOR2_X1 U7233 ( .A1(n5556), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5557) );
  OR2_X1 U7234 ( .A1(n5567), .A2(n5557), .ZN(n9707) );
  AOI22_X1 U7235 ( .A1(n4388), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n5646), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7236 ( .A1(n4480), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5558) );
  OAI211_X1 U7237 ( .C1(n9707), .C2(n5571), .A(n5559), .B(n5558), .ZN(n9696)
         );
  INV_X1 U7238 ( .A(n9696), .ZN(n8240) );
  NAND2_X1 U7239 ( .A1(n9783), .A2(n8240), .ZN(n8292) );
  NAND2_X1 U7240 ( .A1(n8292), .A2(n8289), .ZN(n5561) );
  INV_X1 U7241 ( .A(n8290), .ZN(n5560) );
  NAND2_X1 U7242 ( .A1(n5781), .A2(n5560), .ZN(n5757) );
  MUX2_X1 U7243 ( .A(n5561), .B(n5757), .S(n6972), .Z(n5562) );
  AOI22_X1 U7244 ( .A1(n5699), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5564), .B2(
        n10011), .ZN(n5565) );
  OR2_X1 U7245 ( .A1(n5567), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7246 ( .A1(n5581), .A2(n5568), .ZN(n9689) );
  AOI22_X1 U7247 ( .A1(n4388), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n5646), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7248 ( .A1(n4480), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5569) );
  OAI211_X1 U7249 ( .C1(n9689), .C2(n5571), .A(n5570), .B(n5569), .ZN(n9717)
         );
  INV_X1 U7250 ( .A(n9717), .ZN(n8271) );
  OR2_X1 U7251 ( .A1(n9778), .A2(n8271), .ZN(n5780) );
  NAND2_X1 U7252 ( .A1(n5780), .A2(n5781), .ZN(n5590) );
  AND2_X1 U7253 ( .A1(n5576), .A2(n5575), .ZN(n5577) );
  NAND2_X1 U7254 ( .A1(n5699), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7255 ( .A1(n5581), .A2(n5580), .ZN(n5582) );
  AND2_X1 U7256 ( .A1(n5600), .A2(n5582), .ZN(n9678) );
  NAND2_X1 U7257 ( .A1(n9678), .A2(n5690), .ZN(n5588) );
  INV_X1 U7258 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U7259 ( .A1(n4480), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U7260 ( .A1(n5646), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5583) );
  OAI211_X1 U7261 ( .C1(n5604), .C2(n5585), .A(n5584), .B(n5583), .ZN(n5586)
         );
  INV_X1 U7262 ( .A(n5586), .ZN(n5587) );
  NAND2_X1 U7263 ( .A1(n5588), .A2(n5587), .ZN(n9697) );
  INV_X1 U7264 ( .A(n9697), .ZN(n9666) );
  INV_X1 U7265 ( .A(n8295), .ZN(n5589) );
  NAND2_X1 U7266 ( .A1(n9778), .A2(n8271), .ZN(n8293) );
  OAI211_X1 U7267 ( .C1(n5591), .C2(n5590), .A(n5589), .B(n8293), .ZN(n5593)
         );
  NAND2_X1 U7268 ( .A1(n8293), .A2(n8292), .ZN(n5759) );
  AND2_X1 U7269 ( .A1(n8294), .A2(n5780), .ZN(n5756) );
  OAI21_X1 U7270 ( .B1(n5591), .B2(n5759), .A(n5756), .ZN(n5592) );
  NAND2_X1 U7271 ( .A1(n5625), .A2(n8294), .ZN(n5608) );
  NAND2_X1 U7272 ( .A1(n5595), .A2(n5594), .ZN(n5597) );
  NAND2_X1 U7273 ( .A1(n7912), .A2(n5347), .ZN(n5599) );
  NAND2_X1 U7274 ( .A1(n5699), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5598) );
  AOI21_X1 U7275 ( .B1(n5600), .B2(n9249), .A(n5613), .ZN(n9670) );
  NAND2_X1 U7276 ( .A1(n9670), .A2(n5674), .ZN(n5607) );
  INV_X1 U7277 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U7278 ( .A1(n4480), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U7279 ( .A1(n5646), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5601) );
  OAI211_X1 U7280 ( .C1(n5604), .C2(n5603), .A(n5602), .B(n5601), .ZN(n5605)
         );
  INV_X1 U7281 ( .A(n5605), .ZN(n5606) );
  NAND2_X1 U7282 ( .A1(n9770), .A2(n9478), .ZN(n8296) );
  XNOR2_X1 U7283 ( .A(n5610), .B(n5609), .ZN(n7976) );
  NAND2_X1 U7284 ( .A1(n7976), .A2(n5347), .ZN(n5612) );
  NAND2_X1 U7285 ( .A1(n5699), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7286 ( .A1(n4480), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U7287 ( .A1(n4388), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5617) );
  NOR2_X1 U7288 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n5613), .ZN(n5614) );
  NOR2_X1 U7289 ( .A1(n5643), .A2(n5614), .ZN(n9652) );
  NAND2_X1 U7290 ( .A1(n5674), .A2(n9652), .ZN(n5616) );
  NAND2_X1 U7291 ( .A1(n5646), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5615) );
  OR2_X1 U7292 ( .A1(n9763), .A2(n9667), .ZN(n5778) );
  INV_X1 U7293 ( .A(n5778), .ZN(n5620) );
  OR2_X1 U7294 ( .A1(n9770), .A2(n9478), .ZN(n5779) );
  INV_X1 U7295 ( .A(n5779), .ZN(n5619) );
  NAND2_X1 U7296 ( .A1(n5779), .A2(n8295), .ZN(n5623) );
  AND2_X1 U7297 ( .A1(n5623), .A2(n8296), .ZN(n5624) );
  INV_X1 U7298 ( .A(n5763), .ZN(n5626) );
  AOI21_X1 U7299 ( .B1(n5626), .B2(n5625), .A(n5755), .ZN(n5627) );
  XNOR2_X1 U7300 ( .A(n5630), .B(n5629), .ZN(n8159) );
  NAND2_X1 U7301 ( .A1(n8159), .A2(n5347), .ZN(n5632) );
  NAND2_X1 U7302 ( .A1(n5699), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U7303 ( .A1(n4388), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7304 ( .A1(n4480), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5637) );
  INV_X1 U7305 ( .A(n5645), .ZN(n5633) );
  INV_X1 U7306 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9405) );
  NAND2_X1 U7307 ( .A1(n5633), .A2(n9405), .ZN(n5634) );
  AND2_X1 U7308 ( .A1(n5634), .A2(n5655), .ZN(n9627) );
  NAND2_X1 U7309 ( .A1(n5690), .A2(n9627), .ZN(n5636) );
  NAND2_X1 U7310 ( .A1(n5646), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5635) );
  NAND4_X1 U7311 ( .A1(n5638), .A2(n5637), .A3(n5636), .A4(n5635), .ZN(n9476)
         );
  INV_X1 U7312 ( .A(n9476), .ZN(n9643) );
  OR2_X1 U7313 ( .A1(n9755), .A2(n9643), .ZN(n8300) );
  AND2_X1 U7314 ( .A1(n9755), .A2(n9643), .ZN(n8301) );
  NAND2_X1 U7315 ( .A1(n8054), .A2(n4378), .ZN(n5642) );
  NAND2_X1 U7316 ( .A1(n5699), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U7317 ( .A1(n4388), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7318 ( .A1(n4480), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5649) );
  NOR2_X1 U7319 ( .A1(n5643), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5644) );
  NOR2_X1 U7320 ( .A1(n5645), .A2(n5644), .ZN(n9637) );
  NAND2_X1 U7321 ( .A1(n5690), .A2(n9637), .ZN(n5648) );
  NAND2_X1 U7322 ( .A1(n5646), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5647) );
  NAND4_X1 U7323 ( .A1(n5650), .A2(n5649), .A3(n5648), .A4(n5647), .ZN(n9657)
         );
  INV_X1 U7324 ( .A(n9657), .ZN(n9624) );
  OR2_X1 U7325 ( .A1(n9758), .A2(n9624), .ZN(n8299) );
  NAND2_X1 U7326 ( .A1(n9758), .A2(n9624), .ZN(n5660) );
  NAND2_X1 U7327 ( .A1(n8299), .A2(n5660), .ZN(n9641) );
  NAND2_X1 U7328 ( .A1(n8222), .A2(n4379), .ZN(n5654) );
  NAND2_X1 U7329 ( .A1(n5699), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U7330 ( .A1(n4388), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U7331 ( .A1(n4480), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5658) );
  AOI21_X1 U7332 ( .B1(n5655), .B2(n9374), .A(n5672), .ZN(n9617) );
  NAND2_X1 U7333 ( .A1(n5674), .A2(n9617), .ZN(n5657) );
  NAND2_X1 U7334 ( .A1(n5646), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U7335 ( .A1(n9750), .A2(n9625), .ZN(n8303) );
  INV_X1 U7336 ( .A(n8301), .ZN(n5663) );
  INV_X1 U7337 ( .A(n5660), .ZN(n5661) );
  NAND2_X1 U7338 ( .A1(n8300), .A2(n5661), .ZN(n5662) );
  NAND3_X1 U7339 ( .A1(n8303), .A2(n5663), .A3(n5662), .ZN(n5839) );
  OAI211_X1 U7340 ( .C1(n8301), .C2(n8299), .A(n8302), .B(n8300), .ZN(n5664)
         );
  MUX2_X1 U7341 ( .A(n5839), .B(n5664), .S(n6972), .Z(n5666) );
  MUX2_X1 U7342 ( .A(n8302), .B(n8303), .S(n6972), .Z(n5665) );
  NAND2_X1 U7343 ( .A1(n9042), .A2(n5347), .ZN(n5670) );
  NAND2_X1 U7344 ( .A1(n5699), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U7345 ( .A1(n4388), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U7346 ( .A1(n4480), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5677) );
  OAI21_X1 U7347 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n5672), .A(n5671), .ZN(
        n5673) );
  INV_X1 U7348 ( .A(n5673), .ZN(n9596) );
  NAND2_X1 U7349 ( .A1(n5674), .A2(n9596), .ZN(n5676) );
  NAND2_X1 U7350 ( .A1(n5646), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5675) );
  NAND4_X1 U7351 ( .A1(n5678), .A2(n5677), .A3(n5676), .A4(n5675), .ZN(n9474)
         );
  NAND2_X1 U7352 ( .A1(n9743), .A2(n9612), .ZN(n5725) );
  MUX2_X1 U7353 ( .A(n8305), .B(n5725), .S(n6972), .Z(n5679) );
  AND2_X1 U7354 ( .A1(n5683), .A2(n5695), .ZN(n5684) );
  NAND2_X1 U7355 ( .A1(n9039), .A2(n5347), .ZN(n5687) );
  NAND2_X1 U7356 ( .A1(n5699), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U7357 ( .A1(n4388), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U7358 ( .A1(n5646), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5693) );
  OAI21_X1 U7359 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(n5688), .A(n5702), .ZN(
        n5689) );
  INV_X1 U7360 ( .A(n5689), .ZN(n9585) );
  NAND2_X1 U7361 ( .A1(n5690), .A2(n9585), .ZN(n5692) );
  NAND2_X1 U7362 ( .A1(n4480), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5691) );
  AND4_X2 U7363 ( .A1(n5694), .A2(n5693), .A3(n5692), .A4(n5691), .ZN(n9602)
         );
  NAND2_X1 U7364 ( .A1(n9739), .A2(n9602), .ZN(n5776) );
  NAND2_X1 U7365 ( .A1(n8341), .A2(n4379), .ZN(n5701) );
  NAND2_X1 U7366 ( .A1(n5699), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7367 ( .A1(n4388), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U7368 ( .A1(n4480), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5706) );
  INV_X1 U7369 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6987) );
  NAND2_X1 U7370 ( .A1(n5702), .A2(n6987), .ZN(n5703) );
  NAND2_X1 U7371 ( .A1(n5674), .A2(n9569), .ZN(n5705) );
  NAND2_X1 U7372 ( .A1(n5646), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5704) );
  OR2_X2 U7373 ( .A1(n9739), .A2(n9602), .ZN(n5777) );
  INV_X1 U7374 ( .A(n5777), .ZN(n8308) );
  NAND2_X1 U7375 ( .A1(n9570), .A2(n9582), .ZN(n9550) );
  NAND4_X1 U7376 ( .A1(n5709), .A2(n4883), .A3(n9550), .A4(n5847), .ZN(n5711)
         );
  OR2_X1 U7377 ( .A1(n9726), .A2(n5710), .ZN(n5850) );
  AOI21_X1 U7378 ( .B1(n8322), .B2(n5850), .A(n8323), .ZN(n5713) );
  INV_X1 U7379 ( .A(n5713), .ZN(n5771) );
  OAI22_X1 U7380 ( .A1(n5712), .A2(n5711), .B1(n5771), .B2(n6972), .ZN(n5714)
         );
  NAND2_X1 U7381 ( .A1(n5774), .A2(n6972), .ZN(n5716) );
  INV_X1 U7382 ( .A(n5716), .ZN(n5720) );
  INV_X1 U7383 ( .A(n5717), .ZN(n5718) );
  AND2_X1 U7384 ( .A1(n9550), .A2(n5776), .ZN(n5724) );
  NAND4_X1 U7385 ( .A1(n5771), .A2(n5720), .A3(n5775), .A4(n5719), .ZN(n5721)
         );
  INV_X1 U7386 ( .A(n5724), .ZN(n5728) );
  INV_X1 U7387 ( .A(n5725), .ZN(n5726) );
  AND2_X1 U7388 ( .A1(n5777), .A2(n5726), .ZN(n5727) );
  NOR2_X1 U7389 ( .A1(n5728), .A2(n5727), .ZN(n5842) );
  NOR2_X1 U7390 ( .A1(n5763), .A2(n4583), .ZN(n5814) );
  AND2_X1 U7391 ( .A1(n8289), .A2(n5729), .ZN(n5730) );
  NAND2_X1 U7392 ( .A1(n8292), .A2(n5730), .ZN(n5753) );
  AND2_X1 U7393 ( .A1(n8201), .A2(n5782), .ZN(n5749) );
  INV_X1 U7394 ( .A(n5749), .ZN(n5739) );
  INV_X1 U7395 ( .A(n7813), .ZN(n5733) );
  INV_X1 U7396 ( .A(n5731), .ZN(n5732) );
  OAI211_X1 U7397 ( .C1(n5733), .C2(n7811), .A(n8043), .B(n5732), .ZN(n5747)
         );
  NAND3_X1 U7398 ( .A1(n7699), .A2(n5788), .A3(n5789), .ZN(n5735) );
  INV_X1 U7399 ( .A(n5787), .ZN(n5734) );
  NAND2_X1 U7400 ( .A1(n7699), .A2(n5734), .ZN(n5741) );
  NAND3_X1 U7401 ( .A1(n7702), .A2(n5735), .A3(n5741), .ZN(n5736) );
  NAND3_X1 U7402 ( .A1(n5736), .A2(n5791), .A3(n9969), .ZN(n5737) );
  OR2_X1 U7403 ( .A1(n5747), .A2(n5737), .ZN(n5738) );
  OR3_X1 U7404 ( .A1(n5753), .A2(n5739), .A3(n5738), .ZN(n5832) );
  AND2_X1 U7405 ( .A1(n7702), .A2(n5742), .ZN(n5827) );
  AND2_X1 U7406 ( .A1(n5740), .A2(n5827), .ZN(n5754) );
  AND2_X1 U7407 ( .A1(n5743), .A2(n8202), .ZN(n8236) );
  AND2_X1 U7408 ( .A1(n7706), .A2(n7813), .ZN(n5748) );
  INV_X1 U7409 ( .A(n5744), .ZN(n5745) );
  OAI21_X1 U7410 ( .B1(n4991), .B2(n8043), .A(n5745), .ZN(n5746) );
  OAI21_X1 U7411 ( .B1(n5748), .B2(n5747), .A(n5746), .ZN(n5750) );
  NAND2_X1 U7412 ( .A1(n5750), .A2(n5749), .ZN(n5751) );
  AND2_X1 U7413 ( .A1(n8236), .A2(n5751), .ZN(n5752) );
  OR2_X1 U7414 ( .A1(n5753), .A2(n5752), .ZN(n5830) );
  OAI21_X1 U7415 ( .B1(n5832), .B2(n5754), .A(n5830), .ZN(n5766) );
  INV_X1 U7416 ( .A(n5755), .ZN(n5765) );
  INV_X1 U7417 ( .A(n5756), .ZN(n5761) );
  INV_X1 U7418 ( .A(n5757), .ZN(n5758) );
  NOR2_X1 U7419 ( .A1(n5759), .A2(n5758), .ZN(n5760) );
  NOR2_X1 U7420 ( .A1(n5761), .A2(n5760), .ZN(n5762) );
  OR2_X1 U7421 ( .A1(n5763), .A2(n5762), .ZN(n5764) );
  NAND4_X1 U7422 ( .A1(n8300), .A2(n5765), .A3(n8299), .A4(n5764), .ZN(n5837)
         );
  AOI21_X1 U7423 ( .B1(n5814), .B2(n5766), .A(n5837), .ZN(n5767) );
  AND2_X1 U7424 ( .A1(n8305), .A2(n8302), .ZN(n5838) );
  OAI211_X1 U7425 ( .C1(n5767), .C2(n5839), .A(n5777), .B(n5838), .ZN(n5768)
         );
  AND2_X1 U7426 ( .A1(n5842), .A2(n5768), .ZN(n5770) );
  NAND2_X1 U7427 ( .A1(n5774), .A2(n5775), .ZN(n5843) );
  OAI21_X1 U7428 ( .B1(n5770), .B2(n5843), .A(n5769), .ZN(n5772) );
  INV_X1 U7429 ( .A(n5813), .ZN(n5773) );
  NAND3_X1 U7430 ( .A1(n5773), .A2(n5868), .A3(n7754), .ZN(n5811) );
  INV_X1 U7431 ( .A(n9600), .ZN(n9593) );
  AND2_X1 U7432 ( .A1(n9755), .A2(n9476), .ZN(n8276) );
  INV_X1 U7433 ( .A(n9641), .ZN(n9634) );
  NAND2_X1 U7434 ( .A1(n5779), .A2(n8296), .ZN(n9664) );
  NAND2_X1 U7435 ( .A1(n8199), .A2(n5782), .ZN(n8047) );
  INV_X1 U7436 ( .A(n8047), .ZN(n8039) );
  NAND2_X1 U7437 ( .A1(n5785), .A2(n7707), .ZN(n7737) );
  INV_X1 U7438 ( .A(n7552), .ZN(n7636) );
  AND2_X1 U7439 ( .A1(n7217), .A2(n4966), .ZN(n5817) );
  NOR2_X1 U7440 ( .A1(n7653), .A2(n5817), .ZN(n7195) );
  NAND4_X1 U7441 ( .A1(n7632), .A2(n7195), .A3(n7636), .A4(n5786), .ZN(n5790)
         );
  INV_X1 U7442 ( .A(n10002), .ZN(n10013) );
  NOR3_X1 U7443 ( .A1(n5790), .A2(n10013), .A3(n10035), .ZN(n5793) );
  INV_X1 U7444 ( .A(n7563), .ZN(n9986) );
  NAND4_X1 U7445 ( .A1(n7688), .A2(n9968), .A3(n5793), .A4(n9986), .ZN(n5794)
         );
  NOR2_X1 U7446 ( .A1(n7737), .A2(n5794), .ZN(n5795) );
  NAND4_X1 U7447 ( .A1(n7978), .A2(n7708), .A3(n5795), .A4(n7818), .ZN(n5796)
         );
  NOR2_X1 U7448 ( .A1(n8044), .A2(n5796), .ZN(n5797) );
  NAND4_X1 U7449 ( .A1(n8229), .A2(n8039), .A3(n8209), .A4(n5797), .ZN(n5798)
         );
  NOR2_X1 U7450 ( .A1(n8238), .A2(n5798), .ZN(n5799) );
  NAND3_X1 U7451 ( .A1(n9695), .A2(n9714), .A3(n5799), .ZN(n5800) );
  NOR3_X1 U7452 ( .A1(n9664), .A2(n9681), .A3(n5800), .ZN(n5801) );
  NAND4_X1 U7453 ( .A1(n9623), .A2(n9634), .A3(n9655), .A4(n5801), .ZN(n5802)
         );
  NOR2_X1 U7454 ( .A1(n5802), .A2(n9610), .ZN(n5803) );
  AND4_X1 U7455 ( .A1(n8309), .A2(n8307), .A3(n9593), .A4(n5803), .ZN(n5804)
         );
  AND4_X1 U7456 ( .A1(n9549), .A2(n5850), .A3(n5846), .A4(n5804), .ZN(n5807)
         );
  INV_X1 U7457 ( .A(n5805), .ZN(n5849) );
  NAND3_X1 U7458 ( .A1(n5807), .A2(n5849), .A3(n5852), .ZN(n5812) );
  INV_X1 U7459 ( .A(n5808), .ZN(n5809) );
  NAND3_X1 U7460 ( .A1(n5812), .A2(n5809), .A3(n7913), .ZN(n5810) );
  NOR3_X1 U7461 ( .A1(n5813), .A2(n10011), .A3(n5812), .ZN(n5855) );
  INV_X1 U7462 ( .A(n5814), .ZN(n5835) );
  NAND2_X1 U7463 ( .A1(n5815), .A2(n5816), .ZN(n7637) );
  INV_X1 U7464 ( .A(n5817), .ZN(n5821) );
  NAND2_X1 U7465 ( .A1(n5818), .A2(n5819), .ZN(n5820) );
  NAND3_X1 U7466 ( .A1(n5821), .A2(n5868), .A3(n5820), .ZN(n5822) );
  NAND2_X1 U7467 ( .A1(n7634), .A2(n5822), .ZN(n5824) );
  OAI21_X1 U7468 ( .B1(n7637), .B2(n5824), .A(n5823), .ZN(n5826) );
  NAND2_X1 U7469 ( .A1(n5826), .A2(n5825), .ZN(n5828) );
  AND3_X1 U7470 ( .A1(n5829), .A2(n5828), .A3(n5827), .ZN(n5831) );
  OAI21_X1 U7471 ( .B1(n5832), .B2(n5831), .A(n5830), .ZN(n5833) );
  INV_X1 U7472 ( .A(n5833), .ZN(n5834) );
  NOR2_X1 U7473 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  NOR2_X1 U7474 ( .A1(n5837), .A2(n5836), .ZN(n5840) );
  OAI211_X1 U7475 ( .C1(n5840), .C2(n5839), .A(n8307), .B(n5838), .ZN(n5841)
         );
  NAND2_X1 U7476 ( .A1(n5842), .A2(n5841), .ZN(n5845) );
  INV_X1 U7477 ( .A(n5843), .ZN(n5844) );
  NAND2_X1 U7478 ( .A1(n5845), .A2(n5844), .ZN(n5848) );
  NAND3_X1 U7479 ( .A1(n5848), .A2(n5847), .A3(n5846), .ZN(n5851) );
  NAND3_X1 U7480 ( .A1(n5851), .A2(n5850), .A3(n5849), .ZN(n5853) );
  NAND2_X1 U7481 ( .A1(n5853), .A2(n5852), .ZN(n5864) );
  AOI21_X1 U7482 ( .B1(n5864), .B2(n10011), .A(n7573), .ZN(n5854) );
  INV_X1 U7483 ( .A(n6971), .ZN(n7021) );
  INV_X1 U7484 ( .A(n5875), .ZN(n5859) );
  NOR2_X1 U7485 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5873) );
  INV_X1 U7486 ( .A(n5873), .ZN(n5857) );
  NOR2_X1 U7487 ( .A1(n5857), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U7488 ( .A1(n5859), .A2(n5858), .ZN(n5861) );
  NAND2_X1 U7489 ( .A1(n5861), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5860) );
  MUX2_X1 U7490 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5860), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n5863) );
  NOR2_X1 U7491 ( .A1(n6999), .A2(P1_U3084), .ZN(n8017) );
  OAI21_X1 U7492 ( .B1(n5864), .B2(n7021), .A(n8017), .ZN(n5865) );
  INV_X1 U7493 ( .A(n5865), .ZN(n5866) );
  OR2_X1 U7494 ( .A1(n4537), .A2(n7006), .ZN(n7568) );
  INV_X1 U7495 ( .A(n7568), .ZN(n7193) );
  INV_X1 U7496 ( .A(n9926), .ZN(n9492) );
  INV_X1 U7497 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5871) );
  NAND3_X1 U7498 ( .A1(n5873), .A2(n5872), .A3(n5871), .ZN(n5874) );
  NAND2_X1 U7499 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  NAND2_X1 U7500 ( .A1(n5889), .A2(n6951), .ZN(n6715) );
  NAND3_X1 U7501 ( .A1(n7193), .A2(n9492), .A3(n7040), .ZN(n6986) );
  NAND2_X1 U7502 ( .A1(n6716), .A2(n8017), .ZN(n5891) );
  OAI211_X1 U7503 ( .C1(n6986), .C2(n9920), .A(P1_B_REG_SCAN_IN), .B(n5891), 
        .ZN(n5892) );
  NAND2_X1 U7504 ( .A1(n5893), .A2(n5892), .ZN(P1_U3240) );
  NOR2_X2 U7505 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5897) );
  NOR2_X2 U7506 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5896) );
  NOR2_X4 U7507 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5927) );
  NOR2_X1 U7508 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5900) );
  NOR2_X1 U7509 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n5904) );
  NOR2_X1 U7510 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5903) );
  NOR2_X1 U7511 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5902) );
  NAND4_X1 U7512 ( .A1(n6280), .A2(n5904), .A3(n5903), .A4(n5902), .ZN(n5915)
         );
  AND2_X2 U7513 ( .A1(n9034), .A2(n9038), .ZN(n5958) );
  NAND2_X1 U7514 ( .A1(n5958), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5911) );
  AND2_X2 U7515 ( .A1(n9034), .A2(n5906), .ZN(n5957) );
  NAND2_X1 U7516 ( .A1(n5957), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5910) );
  AND2_X4 U7517 ( .A1(n5907), .A2(n9038), .ZN(n5976) );
  NAND2_X1 U7518 ( .A1(n5976), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7519 ( .A1(n5994), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U7520 ( .A1(n4518), .A2(SI_0_), .ZN(n5912) );
  XNOR2_X1 U7521 ( .A(n5912), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9325) );
  INV_X1 U7522 ( .A(n5915), .ZN(n5916) );
  NAND2_X1 U7523 ( .A1(n5917), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5918) );
  INV_X1 U7524 ( .A(n5919), .ZN(n5920) );
  MUX2_X1 U7525 ( .A(n10173), .B(n9325), .S(n7284), .Z(n8124) );
  NAND2_X1 U7526 ( .A1(n5994), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U7527 ( .A1(n5958), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7528 ( .A1(n5957), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5922) );
  OR2_X1 U7529 ( .A1(n6177), .A2(n5307), .ZN(n5932) );
  NAND2_X1 U7530 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n10173), .ZN(n5926) );
  MUX2_X1 U7531 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5926), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5929) );
  INV_X1 U7532 ( .A(n5927), .ZN(n5928) );
  OR2_X1 U7533 ( .A1(n4385), .A2(n8538), .ZN(n5930) );
  AND3_X4 U7534 ( .A1(n5932), .A2(n5931), .A3(n5930), .ZN(n10194) );
  INV_X1 U7535 ( .A(n10194), .ZN(n7508) );
  NAND2_X1 U7536 ( .A1(n4376), .A2(n7508), .ZN(n5933) );
  NAND2_X1 U7537 ( .A1(n6571), .A2(n5933), .ZN(n5935) );
  OR2_X1 U7538 ( .A1(n4376), .A2(n7508), .ZN(n5934) );
  NAND2_X1 U7539 ( .A1(n5935), .A2(n5934), .ZN(n7836) );
  NAND2_X1 U7540 ( .A1(n5994), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U7541 ( .A1(n5958), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U7542 ( .A1(n5976), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U7543 ( .A1(n5957), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5936) );
  OR2_X1 U7544 ( .A1(n5954), .A2(n7046), .ZN(n5944) );
  OR2_X1 U7545 ( .A1(n6177), .A2(n5325), .ZN(n5943) );
  INV_X4 U7546 ( .A(n7284), .ZN(n7134) );
  NOR2_X1 U7547 ( .A1(n5927), .A2(n6283), .ZN(n5940) );
  MUX2_X1 U7548 ( .A(n6283), .B(n5940), .S(P2_IR_REG_2__SCAN_IN), .Z(n5941) );
  NAND2_X1 U7549 ( .A1(n7134), .A2(n7304), .ZN(n5942) );
  AND3_X2 U7550 ( .A1(n5944), .A2(n5943), .A3(n5942), .ZN(n6574) );
  NAND2_X1 U7551 ( .A1(n10146), .A2(n6574), .ZN(n6434) );
  NAND2_X1 U7552 ( .A1(n7836), .A2(n6546), .ZN(n5946) );
  OR2_X1 U7553 ( .A1(n10146), .A2(n10201), .ZN(n5945) );
  NAND2_X1 U7554 ( .A1(n5958), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U7555 ( .A1(n5976), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7556 ( .A1(n5957), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U7557 ( .A1(n5951), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5953) );
  INV_X1 U7558 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5952) );
  XNOR2_X1 U7559 ( .A(n5953), .B(n5952), .ZN(n7385) );
  INV_X1 U7560 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7031) );
  OR2_X1 U7561 ( .A1(n6177), .A2(n7031), .ZN(n5956) );
  NAND2_X1 U7562 ( .A1(n6404), .A2(n7030), .ZN(n5955) );
  NAND2_X1 U7563 ( .A1(n8535), .A2(n10212), .ZN(n6442) );
  NAND2_X1 U7564 ( .A1(n7796), .A2(n7802), .ZN(n7945) );
  NAND2_X1 U7565 ( .A1(n7957), .A2(n10212), .ZN(n7944) );
  NAND2_X1 U7566 ( .A1(n6396), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7567 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5973) );
  OAI21_X1 U7568 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5973), .ZN(n7950) );
  OR2_X1 U7569 ( .A1(n5975), .A2(n7950), .ZN(n5961) );
  INV_X2 U7570 ( .A(n5995), .ZN(n6356) );
  NAND2_X1 U7571 ( .A1(n6356), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U7572 ( .A1(n5976), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5959) );
  NAND4_X2 U7573 ( .A1(n5962), .A2(n5961), .A3(n5960), .A4(n5959), .ZN(n8534)
         );
  INV_X2 U7574 ( .A(n6177), .ZN(n5986) );
  OR2_X1 U7575 ( .A1(n5951), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7576 ( .A1(n5981), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5963) );
  XNOR2_X1 U7577 ( .A(n5963), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7321) );
  AOI22_X1 U7578 ( .A1(n5986), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7134), .B2(
        n7321), .ZN(n5965) );
  NAND2_X1 U7579 ( .A1(n7029), .A2(n6404), .ZN(n5964) );
  AND2_X2 U7580 ( .A1(n5965), .A2(n5964), .ZN(n10218) );
  NAND2_X1 U7581 ( .A1(n10144), .A2(n10218), .ZN(n5967) );
  AND2_X1 U7582 ( .A1(n7944), .A2(n5967), .ZN(n5966) );
  NAND2_X1 U7583 ( .A1(n7945), .A2(n5966), .ZN(n5970) );
  INV_X1 U7584 ( .A(n5967), .ZN(n5968) );
  INV_X1 U7585 ( .A(n10218), .ZN(n7959) );
  NAND2_X2 U7586 ( .A1(n6425), .A2(n6443), .ZN(n7954) );
  NAND2_X1 U7587 ( .A1(n5957), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5980) );
  INV_X1 U7588 ( .A(n5973), .ZN(n5971) );
  INV_X1 U7589 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7590 ( .A1(n5973), .A2(n5972), .ZN(n5974) );
  NAND2_X1 U7591 ( .A1(n6006), .A2(n5974), .ZN(n7855) );
  OR2_X1 U7592 ( .A1(n5975), .A2(n7855), .ZN(n5979) );
  NAND2_X1 U7593 ( .A1(n6356), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U7594 ( .A1(n5976), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5977) );
  NAND4_X1 U7595 ( .A1(n5980), .A2(n5979), .A3(n5978), .A4(n5977), .ZN(n8533)
         );
  INV_X1 U7596 ( .A(n5981), .ZN(n5983) );
  INV_X1 U7597 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7598 ( .A1(n5983), .A2(n5982), .ZN(n6015) );
  NAND2_X1 U7599 ( .A1(n6015), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5987) );
  XNOR2_X1 U7600 ( .A(n5987), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7336) );
  AOI22_X1 U7601 ( .A1(n5986), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7134), .B2(
        n7336), .ZN(n5984) );
  NAND2_X1 U7602 ( .A1(n6548), .A2(n7854), .ZN(n5985) );
  NAND2_X1 U7603 ( .A1(n7037), .A2(n6404), .ZN(n5993) );
  NAND2_X1 U7604 ( .A1(n5987), .A2(n9118), .ZN(n5988) );
  NAND2_X1 U7605 ( .A1(n5988), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5990) );
  INV_X1 U7606 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U7607 ( .A1(n5990), .A2(n5989), .ZN(n6001) );
  OR2_X1 U7608 ( .A1(n5990), .A2(n5989), .ZN(n5991) );
  AOI22_X1 U7609 ( .A1(n5986), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7134), .B2(
        n7360), .ZN(n5992) );
  NAND2_X1 U7610 ( .A1(n5993), .A2(n5992), .ZN(n7933) );
  NAND2_X1 U7611 ( .A1(n4375), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5999) );
  INV_X2 U7612 ( .A(n5994), .ZN(n6257) );
  INV_X1 U7613 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6005) );
  XNOR2_X1 U7614 ( .A(n6006), .B(n6005), .ZN(n7930) );
  OR2_X1 U7615 ( .A1(n6257), .A2(n7930), .ZN(n5998) );
  INV_X2 U7616 ( .A(n5995), .ZN(n6397) );
  NAND2_X1 U7617 ( .A1(n6397), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U7618 ( .A1(n5976), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7619 ( .A1(n7038), .A2(n6404), .ZN(n6004) );
  NAND2_X1 U7620 ( .A1(n6001), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6002) );
  XNOR2_X1 U7621 ( .A(n6002), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7409) );
  AOI22_X1 U7622 ( .A1(n5986), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7409), .B2(
        n7134), .ZN(n6003) );
  NAND2_X1 U7623 ( .A1(n6004), .A2(n6003), .ZN(n6602) );
  NAND2_X1 U7624 ( .A1(n4375), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6013) );
  OAI21_X1 U7625 ( .B1(n6006), .B2(n6005), .A(n7527), .ZN(n6009) );
  INV_X1 U7626 ( .A(n6006), .ZN(n6008) );
  NAND2_X1 U7627 ( .A1(n6009), .A2(n6025), .ZN(n7889) );
  OR2_X1 U7628 ( .A1(n6257), .A2(n7889), .ZN(n6012) );
  NAND2_X1 U7629 ( .A1(n6397), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7630 ( .A1(n5976), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6010) );
  NAND4_X1 U7631 ( .A1(n6013), .A2(n6012), .A3(n6011), .A4(n6010), .ZN(n8531)
         );
  INV_X1 U7632 ( .A(n8531), .ZN(n7939) );
  OR2_X1 U7633 ( .A1(n6602), .A2(n7939), .ZN(n8059) );
  NAND2_X1 U7634 ( .A1(n6602), .A2(n7939), .ZN(n6449) );
  NAND2_X1 U7635 ( .A1(n8059), .A2(n6449), .ZN(n7887) );
  OR2_X1 U7636 ( .A1(n6602), .A2(n8531), .ZN(n6014) );
  NAND2_X1 U7637 ( .A1(n7044), .A2(n6404), .ZN(n6022) );
  OR4_X2 U7638 ( .A1(n6015), .A2(P2_IR_REG_7__SCAN_IN), .A3(
        P2_IR_REG_5__SCAN_IN), .A4(P2_IR_REG_6__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7639 ( .A1(n6017), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6016) );
  MUX2_X1 U7640 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6016), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n6020) );
  INV_X1 U7641 ( .A(n6017), .ZN(n6019) );
  INV_X1 U7642 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7643 ( .A1(n6019), .A2(n6018), .ZN(n6042) );
  NAND2_X1 U7644 ( .A1(n6020), .A2(n6042), .ZN(n8556) );
  INV_X1 U7645 ( .A(n8556), .ZN(n7412) );
  AOI22_X1 U7646 ( .A1(n5986), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7134), .B2(
        n7412), .ZN(n6021) );
  NAND2_X1 U7647 ( .A1(n6022), .A2(n6021), .ZN(n10246) );
  NAND2_X1 U7648 ( .A1(n4374), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6030) );
  INV_X1 U7649 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7650 ( .A1(n6025), .A2(n6024), .ZN(n6026) );
  NAND2_X1 U7651 ( .A1(n6047), .A2(n6026), .ZN(n8069) );
  OR2_X1 U7652 ( .A1(n6257), .A2(n8069), .ZN(n6029) );
  NAND2_X1 U7653 ( .A1(n6397), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7654 ( .A1(n5976), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6027) );
  NAND4_X1 U7655 ( .A1(n6030), .A2(n6029), .A3(n6028), .A4(n6027), .ZN(n8530)
         );
  INV_X1 U7656 ( .A(n8530), .ZN(n7667) );
  OR2_X1 U7657 ( .A1(n10246), .A2(n7667), .ZN(n6452) );
  NAND2_X1 U7658 ( .A1(n4840), .A2(n7667), .ZN(n8104) );
  NAND2_X1 U7659 ( .A1(n10246), .A2(n8530), .ZN(n6031) );
  NAND2_X1 U7660 ( .A1(n6032), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6033) );
  XNOR2_X1 U7661 ( .A(n6033), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8587) );
  AOI22_X1 U7662 ( .A1(n5986), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7134), .B2(
        n8587), .ZN(n6034) );
  NAND2_X1 U7663 ( .A1(n6397), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6041) );
  INV_X1 U7664 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6046) );
  INV_X1 U7665 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6035) );
  OAI21_X1 U7666 ( .B1(n6047), .B2(n6046), .A(n6035), .ZN(n6037) );
  NAND2_X1 U7667 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n6036) );
  OR2_X2 U7668 ( .A1(n6047), .A2(n6036), .ZN(n6056) );
  NAND2_X1 U7669 ( .A1(n6037), .A2(n6056), .ZN(n8892) );
  OR2_X1 U7670 ( .A1(n6257), .A2(n8892), .ZN(n6040) );
  NAND2_X1 U7671 ( .A1(n5976), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7672 ( .A1(n4374), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6038) );
  NAND4_X1 U7673 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(n8528)
         );
  NAND2_X1 U7674 ( .A1(n10263), .A2(n7967), .ZN(n6457) );
  NAND2_X1 U7675 ( .A1(n9322), .A2(n6404), .ZN(n6045) );
  NAND2_X1 U7676 ( .A1(n6042), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6043) );
  XNOR2_X1 U7677 ( .A(n6043), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9319) );
  AOI22_X1 U7678 ( .A1(n5986), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7134), .B2(
        n9319), .ZN(n6044) );
  NAND2_X2 U7679 ( .A1(n6045), .A2(n6044), .ZN(n8114) );
  NAND2_X1 U7680 ( .A1(n6397), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6051) );
  XNOR2_X1 U7681 ( .A(n6047), .B(n6046), .ZN(n8115) );
  OR2_X1 U7682 ( .A1(n6257), .A2(n8115), .ZN(n6050) );
  NAND2_X1 U7683 ( .A1(n4375), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7684 ( .A1(n5976), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6048) );
  NAND4_X1 U7685 ( .A1(n6051), .A2(n6050), .A3(n6049), .A4(n6048), .ZN(n8529)
         );
  OR2_X1 U7686 ( .A1(n8114), .A2(n8529), .ZN(n8873) );
  INV_X1 U7687 ( .A(n8529), .ZN(n8883) );
  OR2_X1 U7688 ( .A1(n8114), .A2(n8883), .ZN(n6459) );
  NAND2_X1 U7689 ( .A1(n8114), .A2(n8883), .ZN(n8876) );
  NAND3_X1 U7690 ( .A1(n8879), .A2(n8102), .A3(n8873), .ZN(n6052) );
  NAND2_X1 U7691 ( .A1(n7062), .A2(n6404), .ZN(n6055) );
  OR2_X1 U7692 ( .A1(n6165), .A2(n6283), .ZN(n6053) );
  XNOR2_X1 U7693 ( .A(n6053), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7418) );
  AOI22_X1 U7694 ( .A1(n5986), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7134), .B2(
        n7418), .ZN(n6054) );
  NAND2_X1 U7695 ( .A1(n6055), .A2(n6054), .ZN(n7923) );
  NAND2_X1 U7696 ( .A1(n4374), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6061) );
  OR2_X2 U7697 ( .A1(n6056), .A2(n9161), .ZN(n6076) );
  NAND2_X1 U7698 ( .A1(n6056), .A2(n9161), .ZN(n6057) );
  NAND2_X1 U7699 ( .A1(n6076), .A2(n6057), .ZN(n7971) );
  OR2_X1 U7700 ( .A1(n6257), .A2(n7971), .ZN(n6060) );
  NAND2_X1 U7701 ( .A1(n6356), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7702 ( .A1(n5976), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6058) );
  NAND4_X1 U7703 ( .A1(n6061), .A2(n6060), .A3(n6059), .A4(n6058), .ZN(n8527)
         );
  OR2_X1 U7704 ( .A1(n7923), .A2(n8881), .ZN(n8137) );
  NAND2_X1 U7705 ( .A1(n7923), .A2(n8881), .ZN(n6545) );
  NAND2_X1 U7706 ( .A1(n8137), .A2(n6545), .ZN(n7964) );
  NAND2_X1 U7707 ( .A1(n7923), .A2(n8527), .ZN(n6062) );
  NAND2_X1 U7708 ( .A1(n7157), .A2(n6404), .ZN(n6065) );
  INV_X1 U7709 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7710 ( .A1(n6277), .A2(n6063), .ZN(n6119) );
  NAND2_X1 U7711 ( .A1(n6119), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6086) );
  XNOR2_X1 U7712 ( .A(n6086), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7486) );
  AOI22_X1 U7713 ( .A1(n5986), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7486), .B2(
        n7134), .ZN(n6064) );
  INV_X1 U7714 ( .A(n4375), .ZN(n6260) );
  INV_X1 U7715 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9215) );
  OR2_X1 U7716 ( .A1(n6260), .A2(n9215), .ZN(n6071) );
  NAND2_X1 U7717 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_13__SCAN_IN), 
        .ZN(n6066) );
  INV_X1 U7718 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6075) );
  INV_X1 U7719 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7470) );
  OAI21_X1 U7720 ( .B1(n6076), .B2(n6075), .A(n7470), .ZN(n6067) );
  NAND2_X1 U7721 ( .A1(n6091), .A2(n6067), .ZN(n8863) );
  OR2_X1 U7722 ( .A1(n6257), .A2(n8863), .ZN(n6070) );
  NAND2_X1 U7723 ( .A1(n6356), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7724 ( .A1(n5976), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6068) );
  NAND4_X1 U7725 ( .A1(n6071), .A2(n6070), .A3(n6069), .A4(n6068), .ZN(n8525)
         );
  OR2_X1 U7726 ( .A1(n9002), .A2(n8401), .ZN(n6474) );
  NAND2_X1 U7727 ( .A1(n9002), .A2(n8401), .ZN(n6473) );
  NAND2_X1 U7728 ( .A1(n6474), .A2(n6473), .ZN(n6343) );
  NAND2_X1 U7729 ( .A1(n7152), .A2(n6404), .ZN(n6074) );
  OR2_X1 U7730 ( .A1(n6277), .A2(n6283), .ZN(n6072) );
  XNOR2_X1 U7731 ( .A(n6072), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7463) );
  AOI22_X1 U7732 ( .A1(n5986), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7134), .B2(
        n7463), .ZN(n6073) );
  NAND2_X1 U7733 ( .A1(n6356), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6080) );
  XNOR2_X1 U7734 ( .A(n6076), .B(n6075), .ZN(n8132) );
  OR2_X1 U7735 ( .A1(n6257), .A2(n8132), .ZN(n6079) );
  NAND2_X1 U7736 ( .A1(n4374), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7737 ( .A1(n5976), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6077) );
  NAND4_X1 U7738 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n8526)
         );
  OR2_X1 U7739 ( .A1(n8134), .A2(n8526), .ZN(n8855) );
  NAND2_X1 U7740 ( .A1(n8127), .A2(n6081), .ZN(n6085) );
  OR2_X1 U7741 ( .A1(n8134), .A2(n8854), .ZN(n6463) );
  NAND2_X1 U7742 ( .A1(n8134), .A2(n8854), .ZN(n6552) );
  NAND2_X1 U7743 ( .A1(n6463), .A2(n6552), .ZN(n8128) );
  INV_X1 U7744 ( .A(n8855), .ZN(n6082) );
  NOR2_X1 U7745 ( .A1(n8128), .A2(n6082), .ZN(n6083) );
  AOI22_X1 U7746 ( .A1(n6343), .A2(n6083), .B1(n9002), .B2(n8525), .ZN(n6084)
         );
  NAND2_X1 U7747 ( .A1(n7164), .A2(n6404), .ZN(n6089) );
  NAND2_X1 U7748 ( .A1(n6086), .A2(n6116), .ZN(n6087) );
  NAND2_X1 U7749 ( .A1(n6087), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6100) );
  XNOR2_X1 U7750 ( .A(n6100), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7762) );
  AOI22_X1 U7751 ( .A1(n7762), .A2(n7134), .B1(n5986), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7752 ( .A1(n6356), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6096) );
  INV_X1 U7753 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9224) );
  NAND2_X1 U7754 ( .A1(n6091), .A2(n9224), .ZN(n6092) );
  NAND2_X1 U7755 ( .A1(n6107), .A2(n6092), .ZN(n8400) );
  OR2_X1 U7756 ( .A1(n6257), .A2(n8400), .ZN(n6095) );
  NAND2_X1 U7757 ( .A1(n4374), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7758 ( .A1(n5976), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6093) );
  NAND4_X1 U7759 ( .A1(n6096), .A2(n6095), .A3(n6094), .A4(n6093), .ZN(n8524)
         );
  OR2_X1 U7760 ( .A1(n8997), .A2(n8524), .ZN(n6099) );
  NAND2_X1 U7761 ( .A1(n8997), .A2(n8524), .ZN(n6097) );
  NAND2_X1 U7762 ( .A1(n6099), .A2(n6097), .ZN(n8077) );
  NAND2_X1 U7763 ( .A1(n7222), .A2(n6404), .ZN(n6104) );
  NAND2_X1 U7764 ( .A1(n6100), .A2(n6117), .ZN(n6101) );
  NAND2_X1 U7765 ( .A1(n6101), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6102) );
  XNOR2_X1 U7766 ( .A(n6102), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7783) );
  AOI22_X1 U7767 ( .A1(n7783), .A2(n7134), .B1(n5986), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7768 ( .A1(n4374), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7769 ( .A1(n6356), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6111) );
  INV_X1 U7770 ( .A(n6107), .ZN(n6105) );
  INV_X1 U7771 ( .A(n6123), .ZN(n6137) );
  INV_X1 U7772 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7773 ( .A1(n6107), .A2(n6106), .ZN(n6108) );
  AND2_X1 U7774 ( .A1(n6137), .A2(n6108), .ZN(n8834) );
  NAND2_X1 U7775 ( .A1(n5994), .A2(n8834), .ZN(n6110) );
  NAND2_X1 U7776 ( .A1(n5976), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6109) );
  NAND4_X1 U7777 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n8814)
         );
  INV_X1 U7778 ( .A(n8814), .ZN(n8453) );
  OR2_X1 U7779 ( .A1(n8992), .A2(n8453), .ZN(n6482) );
  NAND2_X1 U7780 ( .A1(n8992), .A2(n8453), .ZN(n6481) );
  NAND2_X1 U7781 ( .A1(n6482), .A2(n6481), .ZN(n8835) );
  OR2_X1 U7782 ( .A1(n8992), .A2(n8814), .ZN(n6113) );
  NAND2_X1 U7783 ( .A1(n6114), .A2(n6113), .ZN(n8801) );
  NAND2_X1 U7784 ( .A1(n7436), .A2(n6404), .ZN(n6122) );
  INV_X1 U7785 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6115) );
  NAND3_X1 U7786 ( .A1(n6117), .A2(n6116), .A3(n6115), .ZN(n6118) );
  OR2_X1 U7787 ( .A1(n6119), .A2(n6118), .ZN(n6132) );
  OAI21_X1 U7788 ( .B1(n6132), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6120) );
  XNOR2_X1 U7789 ( .A(n6120), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8598) );
  AOI22_X1 U7790 ( .A1(n8598), .A2(n7134), .B1(n5986), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n6121) );
  INV_X1 U7791 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n6131) );
  INV_X1 U7792 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6125) );
  NAND2_X1 U7793 ( .A1(n6139), .A2(n6125), .ZN(n6126) );
  NAND2_X1 U7794 ( .A1(n6157), .A2(n6126), .ZN(n8797) );
  OR2_X1 U7795 ( .A1(n8797), .A2(n6257), .ZN(n6130) );
  INV_X1 U7796 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9147) );
  OR2_X1 U7797 ( .A1(n6260), .A2(n9147), .ZN(n6128) );
  NAND2_X1 U7798 ( .A1(n6397), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6127) );
  AND2_X1 U7799 ( .A1(n6128), .A2(n6127), .ZN(n6129) );
  OAI211_X1 U7800 ( .C1(n6359), .C2(n6131), .A(n6130), .B(n6129), .ZN(n8817)
         );
  INV_X1 U7801 ( .A(n8817), .ZN(n8505) );
  NAND2_X1 U7802 ( .A1(n8980), .A2(n8505), .ZN(n6417) );
  NAND2_X1 U7803 ( .A1(n6418), .A2(n6417), .ZN(n8803) );
  NAND2_X1 U7804 ( .A1(n7277), .A2(n6404), .ZN(n6135) );
  NAND2_X1 U7805 ( .A1(n6132), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6133) );
  XNOR2_X1 U7806 ( .A(n6133), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8031) );
  AOI22_X1 U7807 ( .A1(n7134), .A2(n8031), .B1(n5986), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n6134) );
  INV_X1 U7808 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7809 ( .A1(n6137), .A2(n6136), .ZN(n6138) );
  NAND2_X1 U7810 ( .A1(n6139), .A2(n6138), .ZN(n8823) );
  INV_X1 U7811 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6140) );
  OAI22_X1 U7812 ( .A1(n8823), .A2(n6257), .B1(n6359), .B2(n6140), .ZN(n6143)
         );
  INV_X1 U7813 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8990) );
  NAND2_X1 U7814 ( .A1(n6397), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6141) );
  OAI21_X1 U7815 ( .B1(n6260), .B2(n8990), .A(n6141), .ZN(n6142) );
  NAND2_X1 U7816 ( .A1(n8984), .A2(n8523), .ZN(n8802) );
  NAND3_X1 U7817 ( .A1(n8801), .A2(n8803), .A3(n8802), .ZN(n6149) );
  INV_X1 U7818 ( .A(n8523), .ZN(n6144) );
  OR2_X1 U7819 ( .A1(n8984), .A2(n6144), .ZN(n6424) );
  NAND2_X1 U7820 ( .A1(n8984), .A2(n6144), .ZN(n6423) );
  NAND2_X1 U7821 ( .A1(n6424), .A2(n6423), .ZN(n8809) );
  INV_X1 U7822 ( .A(n8802), .ZN(n6145) );
  NOR2_X1 U7823 ( .A1(n8809), .A2(n6145), .ZN(n6147) );
  NOR2_X1 U7824 ( .A1(n8980), .A2(n8817), .ZN(n6146) );
  AOI21_X1 U7825 ( .B1(n8803), .B2(n6147), .A(n6146), .ZN(n6148) );
  NAND2_X1 U7826 ( .A1(n6149), .A2(n6148), .ZN(n8786) );
  NAND2_X1 U7827 ( .A1(n7683), .A2(n6404), .ZN(n6156) );
  NOR2_X1 U7828 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n6151) );
  NOR2_X1 U7829 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6150) );
  AND3_X1 U7830 ( .A1(n6152), .A2(n6151), .A3(n6150), .ZN(n6164) );
  NAND2_X1 U7831 ( .A1(n6277), .A2(n6164), .ZN(n6153) );
  NAND2_X1 U7832 ( .A1(n6153), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6154) );
  XNOR2_X1 U7833 ( .A(n6154), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8610) );
  AOI22_X1 U7834 ( .A1(n5986), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7134), .B2(
        n8610), .ZN(n6155) );
  NAND2_X1 U7835 ( .A1(n6157), .A2(n9173), .ZN(n6158) );
  NAND2_X1 U7836 ( .A1(n6171), .A2(n6158), .ZN(n8782) );
  AOI22_X1 U7837 ( .A1(n4375), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n6397), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7838 ( .A1(n5976), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6159) );
  OAI211_X1 U7839 ( .C1(n8782), .C2(n6257), .A(n6160), .B(n6159), .ZN(n8768)
         );
  NOR2_X1 U7840 ( .A1(n8974), .A2(n8768), .ZN(n6162) );
  NAND2_X1 U7841 ( .A1(n8974), .A2(n8768), .ZN(n6161) );
  NAND2_X1 U7842 ( .A1(n7753), .A2(n6404), .ZN(n6168) );
  NOR2_X1 U7843 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6163) );
  NAND3_X1 U7844 ( .A1(n6165), .A2(n6164), .A3(n6163), .ZN(n6166) );
  AOI22_X1 U7845 ( .A1(n5986), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8620), .B2(
        n7134), .ZN(n6167) );
  INV_X1 U7846 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6175) );
  INV_X1 U7847 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7848 ( .A1(n6171), .A2(n6170), .ZN(n6172) );
  NAND2_X1 U7849 ( .A1(n6180), .A2(n6172), .ZN(n8418) );
  OR2_X1 U7850 ( .A1(n8418), .A2(n6257), .ZN(n6174) );
  AOI22_X1 U7851 ( .A1(n4374), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n6397), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n6173) );
  OAI211_X1 U7852 ( .C1(n6359), .C2(n6175), .A(n6174), .B(n6173), .ZN(n8779)
         );
  AND2_X1 U7853 ( .A1(n8970), .A2(n8779), .ZN(n6176) );
  NAND2_X1 U7854 ( .A1(n7909), .A2(n6404), .ZN(n6179) );
  OR2_X1 U7855 ( .A1(n6406), .A2(n7918), .ZN(n6178) );
  NAND2_X2 U7856 ( .A1(n6179), .A2(n6178), .ZN(n8963) );
  INV_X1 U7857 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8482) );
  OR2_X2 U7858 ( .A1(n6180), .A2(n8482), .ZN(n6200) );
  NAND2_X1 U7859 ( .A1(n6180), .A2(n8482), .ZN(n6181) );
  AND2_X1 U7860 ( .A1(n6200), .A2(n6181), .ZN(n8755) );
  NAND2_X1 U7861 ( .A1(n8755), .A2(n5994), .ZN(n6187) );
  INV_X1 U7862 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7863 ( .A1(n6397), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7864 ( .A1(n4375), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6182) );
  OAI211_X1 U7865 ( .C1(n6359), .C2(n6184), .A(n6183), .B(n6182), .ZN(n6185)
         );
  INV_X1 U7866 ( .A(n6185), .ZN(n6186) );
  NAND2_X1 U7867 ( .A1(n6187), .A2(n6186), .ZN(n8769) );
  NAND2_X1 U7868 ( .A1(n8963), .A2(n8428), .ZN(n6502) );
  INV_X1 U7869 ( .A(n8963), .ZN(n8757) );
  NAND2_X1 U7870 ( .A1(n7912), .A2(n6404), .ZN(n6189) );
  OR2_X1 U7871 ( .A1(n6406), .A2(n7943), .ZN(n6188) );
  INV_X1 U7872 ( .A(n8741), .ZN(n8955) );
  XNOR2_X1 U7873 ( .A(n6200), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n8426) );
  NAND2_X1 U7874 ( .A1(n8426), .A2(n5994), .ZN(n6195) );
  INV_X1 U7875 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7876 ( .A1(n6397), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7877 ( .A1(n4375), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6190) );
  OAI211_X1 U7878 ( .C1(n6192), .C2(n6359), .A(n6191), .B(n6190), .ZN(n6193)
         );
  INV_X1 U7879 ( .A(n6193), .ZN(n6194) );
  NAND2_X1 U7880 ( .A1(n6195), .A2(n6194), .ZN(n8751) );
  INV_X1 U7881 ( .A(n8751), .ZN(n8497) );
  NAND2_X1 U7882 ( .A1(n8955), .A2(n8497), .ZN(n6197) );
  NAND2_X1 U7883 ( .A1(n7976), .A2(n6404), .ZN(n6199) );
  OR2_X1 U7884 ( .A1(n6406), .A2(n8244), .ZN(n6198) );
  INV_X1 U7885 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9133) );
  INV_X1 U7886 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8495) );
  OAI21_X1 U7887 ( .B1(n6200), .B2(n9133), .A(n8495), .ZN(n6203) );
  AND2_X1 U7888 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n6201) );
  NAND2_X1 U7889 ( .A1(n6203), .A2(n6213), .ZN(n8716) );
  OR2_X1 U7890 ( .A1(n8716), .A2(n6257), .ZN(n6209) );
  INV_X1 U7891 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7892 ( .A1(n4374), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7893 ( .A1(n5976), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6204) );
  OAI211_X1 U7894 ( .C1(n6228), .C2(n6206), .A(n6205), .B(n6204), .ZN(n6207)
         );
  INV_X1 U7895 ( .A(n6207), .ZN(n6208) );
  NAND2_X1 U7896 ( .A1(n8950), .A2(n8427), .ZN(n6488) );
  NAND2_X1 U7897 ( .A1(n8696), .A2(n6488), .ZN(n6350) );
  NAND2_X1 U7898 ( .A1(n8054), .A2(n6404), .ZN(n6211) );
  OR2_X1 U7899 ( .A1(n6406), .A2(n8057), .ZN(n6210) );
  INV_X1 U7900 ( .A(n6223), .ZN(n6224) );
  INV_X1 U7901 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U7902 ( .A1(n6213), .A2(n8409), .ZN(n6214) );
  NAND2_X1 U7903 ( .A1(n6224), .A2(n6214), .ZN(n8702) );
  OR2_X1 U7904 ( .A1(n8702), .A2(n6257), .ZN(n6220) );
  INV_X1 U7905 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7906 ( .A1(n6397), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7907 ( .A1(n4375), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6215) );
  OAI211_X1 U7908 ( .C1(n6217), .C2(n6359), .A(n6216), .B(n6215), .ZN(n6218)
         );
  INV_X1 U7909 ( .A(n6218), .ZN(n6219) );
  NAND2_X1 U7910 ( .A1(n6220), .A2(n6219), .ZN(n8726) );
  OR2_X1 U7911 ( .A1(n8945), .A2(n8496), .ZN(n6511) );
  NAND2_X1 U7912 ( .A1(n8945), .A2(n8496), .ZN(n6496) );
  INV_X1 U7913 ( .A(n8945), .ZN(n8705) );
  NAND2_X1 U7914 ( .A1(n8159), .A2(n6404), .ZN(n6222) );
  INV_X1 U7915 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n9291) );
  OR2_X1 U7916 ( .A1(n6406), .A2(n9291), .ZN(n6221) );
  INV_X1 U7917 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8474) );
  NAND2_X1 U7918 ( .A1(n6224), .A2(n8474), .ZN(n6225) );
  NAND2_X1 U7919 ( .A1(n6234), .A2(n6225), .ZN(n8681) );
  OR2_X1 U7920 ( .A1(n8681), .A2(n6257), .ZN(n6231) );
  INV_X1 U7921 ( .A(n6397), .ZN(n6228) );
  INV_X1 U7922 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9247) );
  NAND2_X1 U7923 ( .A1(n5976), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6227) );
  NAND2_X1 U7924 ( .A1(n4374), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6226) );
  OAI211_X1 U7925 ( .C1(n6228), .C2(n9247), .A(n6227), .B(n6226), .ZN(n6229)
         );
  INV_X1 U7926 ( .A(n6229), .ZN(n6230) );
  NAND2_X1 U7927 ( .A1(n6231), .A2(n6230), .ZN(n8699) );
  NAND2_X1 U7928 ( .A1(n8940), .A2(n8440), .ZN(n6516) );
  NAND2_X1 U7929 ( .A1(n8222), .A2(n6404), .ZN(n6233) );
  OR2_X1 U7930 ( .A1(n6406), .A2(n8227), .ZN(n6232) );
  INV_X1 U7931 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8437) );
  NAND2_X1 U7932 ( .A1(n6234), .A2(n8437), .ZN(n6235) );
  AND2_X1 U7933 ( .A1(n6246), .A2(n6235), .ZN(n8672) );
  NAND2_X1 U7934 ( .A1(n8672), .A2(n5994), .ZN(n6240) );
  INV_X1 U7935 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n9175) );
  NAND2_X1 U7936 ( .A1(n4374), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7937 ( .A1(n6397), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6236) );
  OAI211_X1 U7938 ( .C1(n9175), .C2(n6359), .A(n6237), .B(n6236), .ZN(n6238)
         );
  INV_X1 U7939 ( .A(n6238), .ZN(n6239) );
  NAND2_X1 U7940 ( .A1(n6240), .A2(n6239), .ZN(n8689) );
  INV_X1 U7941 ( .A(n8689), .ZN(n8475) );
  XNOR2_X1 U7942 ( .A(n8673), .B(n8475), .ZN(n8669) );
  NAND2_X1 U7943 ( .A1(n8670), .A2(n8669), .ZN(n8668) );
  NAND2_X1 U7944 ( .A1(n9042), .A2(n6404), .ZN(n6243) );
  OR2_X1 U7945 ( .A1(n6406), .A2(n9044), .ZN(n6242) );
  INV_X1 U7946 ( .A(n6246), .ZN(n6244) );
  INV_X1 U7947 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7948 ( .A1(n6246), .A2(n6245), .ZN(n6247) );
  NAND2_X1 U7949 ( .A1(n6255), .A2(n6247), .ZN(n8661) );
  OR2_X2 U7950 ( .A1(n8661), .A2(n6257), .ZN(n6252) );
  INV_X1 U7951 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9196) );
  NAND2_X1 U7952 ( .A1(n4375), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U7953 ( .A1(n5976), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6248) );
  OAI211_X1 U7954 ( .C1(n6228), .C2(n9196), .A(n6249), .B(n6248), .ZN(n6250)
         );
  INV_X1 U7955 ( .A(n6250), .ZN(n6251) );
  NAND2_X1 U7956 ( .A1(n8930), .A2(n8439), .ZN(n8632) );
  NAND2_X2 U7957 ( .A1(n6519), .A2(n8632), .ZN(n8651) );
  OR2_X1 U7958 ( .A1(n6406), .A2(n9041), .ZN(n6254) );
  INV_X1 U7959 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U7960 ( .A1(n6255), .A2(n6709), .ZN(n6256) );
  NAND2_X1 U7961 ( .A1(n6266), .A2(n6256), .ZN(n8640) );
  INV_X1 U7962 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9185) );
  NAND2_X1 U7963 ( .A1(n6356), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U7964 ( .A1(n5976), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6258) );
  OAI211_X1 U7965 ( .C1(n6260), .C2(n9185), .A(n6259), .B(n6258), .ZN(n6261)
         );
  INV_X1 U7966 ( .A(n6261), .ZN(n6262) );
  NAND2_X1 U7967 ( .A1(n8924), .A2(n8367), .ZN(n6522) );
  NAND2_X1 U7968 ( .A1(n8341), .A2(n6404), .ZN(n6265) );
  OR2_X1 U7969 ( .A1(n6406), .A2(n8342), .ZN(n6264) );
  INV_X1 U7970 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8365) );
  NAND2_X1 U7971 ( .A1(n6266), .A2(n8365), .ZN(n6267) );
  NAND2_X1 U7972 ( .A1(n8364), .A2(n5994), .ZN(n6273) );
  INV_X1 U7973 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7974 ( .A1(n4374), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U7975 ( .A1(n6356), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6268) );
  OAI211_X1 U7976 ( .C1(n6270), .C2(n6359), .A(n6269), .B(n6268), .ZN(n6271)
         );
  INV_X1 U7977 ( .A(n6271), .ZN(n6272) );
  NAND2_X1 U7978 ( .A1(n8919), .A2(n6710), .ZN(n6525) );
  OAI21_X1 U7979 ( .B1(n6274), .B2(n6385), .A(n8378), .ZN(n6275) );
  INV_X1 U7980 ( .A(n6275), .ZN(n8923) );
  NAND2_X1 U7981 ( .A1(n6280), .A2(n6316), .ZN(n6281) );
  NOR2_X1 U7982 ( .A1(n6285), .A2(n6283), .ZN(n6282) );
  MUX2_X1 U7983 ( .A(n6283), .B(n6282), .S(P2_IR_REG_25__SCAN_IN), .Z(n6287)
         );
  NAND2_X1 U7984 ( .A1(n6285), .A2(n6284), .ZN(n6293) );
  INV_X1 U7985 ( .A(n6293), .ZN(n6286) );
  NAND2_X1 U7986 ( .A1(n6317), .A2(n6316), .ZN(n6289) );
  XNOR2_X1 U7987 ( .A(n8160), .B(P2_B_REG_SCAN_IN), .ZN(n6292) );
  NAND2_X1 U7988 ( .A1(n8225), .A2(n6292), .ZN(n6295) );
  NAND2_X1 U7989 ( .A1(n6293), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6294) );
  INV_X1 U7990 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10184) );
  NOR2_X1 U7991 ( .A1(n6305), .A2(n6313), .ZN(n10185) );
  AOI21_X1 U7992 ( .B1(n10174), .B2(n10184), .A(n10185), .ZN(n8907) );
  NOR4_X1 U7993 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6299) );
  NOR4_X1 U7994 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6298) );
  NOR4_X1 U7995 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6297) );
  NOR4_X1 U7996 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6296) );
  NAND4_X1 U7997 ( .A1(n6299), .A2(n6298), .A3(n6297), .A4(n6296), .ZN(n6304)
         );
  NOR2_X1 U7998 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .ZN(
        n9056) );
  NOR4_X1 U7999 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6302) );
  NOR4_X1 U8000 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6301) );
  NOR4_X1 U8001 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6300) );
  NAND4_X1 U8002 ( .A1(n9056), .A2(n6302), .A3(n6301), .A4(n6300), .ZN(n6303)
         );
  OAI21_X1 U8003 ( .B1(n6304), .B2(n6303), .A(n10174), .ZN(n8905) );
  AND2_X1 U8004 ( .A1(n8907), .A2(n8905), .ZN(n6677) );
  INV_X1 U8005 ( .A(n8160), .ZN(n6306) );
  NAND2_X1 U8006 ( .A1(n6311), .A2(n6310), .ZN(n6680) );
  INV_X1 U8007 ( .A(n6313), .ZN(n9045) );
  INV_X1 U8008 ( .A(n10182), .ZN(n6315) );
  INV_X1 U8009 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10181) );
  NAND2_X1 U8010 ( .A1(n10174), .A2(n10181), .ZN(n6314) );
  NAND2_X1 U8011 ( .A1(n6321), .A2(n6320), .ZN(n6322) );
  NAND2_X1 U8012 ( .A1(n6322), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6324) );
  INV_X1 U8013 ( .A(n8902), .ZN(n6325) );
  NOR2_X1 U8014 ( .A1(n8908), .A2(n6325), .ZN(n6326) );
  NAND2_X1 U8015 ( .A1(n6684), .A2(n6326), .ZN(n6372) );
  AND2_X1 U8016 ( .A1(n7917), .A2(n8620), .ZN(n6327) );
  NAND2_X1 U8017 ( .A1(n6373), .A2(n6327), .ZN(n10269) );
  XNOR2_X1 U8018 ( .A(n6373), .B(n6569), .ZN(n6329) );
  OR2_X1 U8019 ( .A1(n6569), .A2(n4760), .ZN(n7795) );
  NAND2_X1 U8020 ( .A1(n8913), .A2(n7795), .ZN(n6330) );
  INV_X2 U8021 ( .A(n8124), .ZN(n10188) );
  OR2_X2 U8022 ( .A1(n8537), .A2(n10188), .ZN(n8147) );
  NAND2_X1 U8023 ( .A1(n4377), .A2(n10194), .ZN(n8145) );
  INV_X1 U8024 ( .A(n6546), .ZN(n7843) );
  NAND2_X1 U8025 ( .A1(n7842), .A2(n7843), .ZN(n7800) );
  NAND2_X1 U8026 ( .A1(n7800), .A2(n7801), .ZN(n6331) );
  INV_X1 U8027 ( .A(n7952), .ZN(n6332) );
  NOR2_X1 U8028 ( .A1(n7954), .A2(n6332), .ZN(n6333) );
  NAND2_X1 U8029 ( .A1(n7799), .A2(n6333), .ZN(n6334) );
  NAND2_X1 U8030 ( .A1(n6334), .A2(n6443), .ZN(n7848) );
  OR2_X1 U8031 ( .A1(n7528), .A2(n7933), .ZN(n6444) );
  NAND2_X1 U8032 ( .A1(n7933), .A2(n7528), .ZN(n7884) );
  INV_X1 U8033 ( .A(n7884), .ZN(n6336) );
  NOR2_X1 U8034 ( .A1(n7887), .A2(n6336), .ZN(n6337) );
  AND2_X1 U8035 ( .A1(n6452), .A2(n8059), .ZN(n6338) );
  INV_X1 U8036 ( .A(n8104), .ZN(n6339) );
  INV_X1 U8037 ( .A(n8876), .ZN(n6340) );
  AND2_X1 U8038 ( .A1(n6463), .A2(n8137), .ZN(n6553) );
  NAND2_X1 U8039 ( .A1(n6342), .A2(n6552), .ZN(n8852) );
  NAND2_X1 U8040 ( .A1(n8852), .A2(n8857), .ZN(n8851) );
  INV_X1 U8041 ( .A(n8524), .ZN(n8853) );
  INV_X1 U8042 ( .A(n6482), .ZN(n6344) );
  NAND2_X1 U8043 ( .A1(n8810), .A2(n8811), .ZN(n6345) );
  INV_X1 U8044 ( .A(n8768), .ZN(n8419) );
  NAND2_X1 U8045 ( .A1(n8974), .A2(n8419), .ZN(n6543) );
  INV_X1 U8046 ( .A(n8779), .ZN(n8504) );
  OR2_X1 U8047 ( .A1(n8970), .A2(n8504), .ZN(n6500) );
  NAND2_X1 U8048 ( .A1(n8970), .A2(n8504), .ZN(n8748) );
  NAND2_X1 U8049 ( .A1(n6500), .A2(n8748), .ZN(n8765) );
  INV_X1 U8050 ( .A(n8759), .ZN(n6347) );
  INV_X1 U8051 ( .A(n8748), .ZN(n6486) );
  NOR2_X1 U8052 ( .A1(n6347), .A2(n6486), .ZN(n6348) );
  INV_X1 U8053 ( .A(n6497), .ZN(n6349) );
  XNOR2_X1 U8054 ( .A(n8741), .B(n8751), .ZN(n8732) );
  NAND2_X1 U8055 ( .A1(n8741), .A2(n8497), .ZN(n8721) );
  INV_X1 U8056 ( .A(n8707), .ZN(n8695) );
  AND2_X1 U8057 ( .A1(n8695), .A2(n8696), .ZN(n6352) );
  NAND2_X1 U8058 ( .A1(n8685), .A2(n6353), .ZN(n8687) );
  INV_X1 U8059 ( .A(n8669), .ZN(n6556) );
  INV_X1 U8060 ( .A(n8651), .ZN(n8656) );
  NAND2_X1 U8061 ( .A1(n6561), .A2(n6328), .ZN(n6413) );
  INV_X1 U8062 ( .A(n6355), .ZN(n8387) );
  INV_X1 U8063 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U8064 ( .A1(n4375), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U8065 ( .A1(n6356), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6357) );
  OAI211_X1 U8066 ( .C1(n6360), .C2(n6359), .A(n6358), .B(n6357), .ZN(n6361)
         );
  AOI21_X1 U8067 ( .B1(n8387), .B2(n5994), .A(n6361), .ZN(n8368) );
  INV_X1 U8068 ( .A(n8368), .ZN(n8522) );
  INV_X1 U8069 ( .A(n6363), .ZN(n6364) );
  NAND2_X1 U8070 ( .A1(n8522), .A2(n8816), .ZN(n6366) );
  NAND2_X1 U8071 ( .A1(n8657), .A2(n8815), .ZN(n6365) );
  INV_X1 U8072 ( .A(n8970), .ZN(n8423) );
  NOR2_X2 U8073 ( .A1(n7853), .A2(n7933), .ZN(n7927) );
  INV_X1 U8074 ( .A(n6602), .ZN(n10239) );
  INV_X1 U8075 ( .A(n10246), .ZN(n8070) );
  INV_X1 U8076 ( .A(n7923), .ZN(n10274) );
  INV_X1 U8077 ( .A(n8134), .ZN(n10281) );
  NAND2_X1 U8078 ( .A1(n8130), .A2(n10281), .ZN(n8862) );
  OR2_X2 U8079 ( .A1(n8862), .A2(n9002), .ZN(n8080) );
  INV_X1 U8080 ( .A(n8992), .ZN(n8846) );
  INV_X1 U8081 ( .A(n8984), .ZN(n8826) );
  INV_X1 U8082 ( .A(n8919), .ZN(n6380) );
  INV_X1 U8083 ( .A(n8386), .ZN(n6371) );
  AOI21_X1 U8084 ( .B1(n8919), .B2(n4493), .A(n6371), .ZN(n8920) );
  INV_X1 U8085 ( .A(n6372), .ZN(n6377) );
  INV_X1 U8086 ( .A(n6567), .ZN(n6375) );
  NAND2_X1 U8087 ( .A1(n6375), .A2(n7917), .ZN(n7852) );
  INV_X1 U8088 ( .A(n7852), .ZN(n6376) );
  NOR2_X1 U8089 ( .A1(n6567), .A2(n7917), .ZN(n6378) );
  INV_X1 U8090 ( .A(n8891), .ZN(n8864) );
  AOI22_X1 U8091 ( .A1(n8364), .A2(n8864), .B1(n8866), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n6379) );
  OAI21_X1 U8092 ( .B1(n6380), .B2(n8893), .A(n6379), .ZN(n6381) );
  AOI21_X1 U8093 ( .B1(n8920), .B2(n8895), .A(n6381), .ZN(n6382) );
  OAI21_X1 U8094 ( .B1(n8922), .B2(n8872), .A(n6382), .ZN(n6383) );
  INV_X1 U8095 ( .A(n6383), .ZN(n6384) );
  INV_X1 U8096 ( .A(n6385), .ZN(n6557) );
  INV_X1 U8097 ( .A(n6526), .ZN(n6386) );
  NAND2_X1 U8098 ( .A1(n8329), .A2(n6404), .ZN(n6389) );
  OR2_X1 U8099 ( .A1(n6406), .A2(n9292), .ZN(n6388) );
  OR2_X1 U8100 ( .A1(n8914), .A2(n8368), .ZN(n6529) );
  NAND2_X1 U8101 ( .A1(n8914), .A2(n8368), .ZN(n6530) );
  NAND2_X1 U8102 ( .A1(n4374), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U8103 ( .A1(n5976), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U8104 ( .A1(n6397), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6390) );
  NAND3_X1 U8105 ( .A1(n6392), .A2(n6391), .A3(n6390), .ZN(n8623) );
  NOR2_X1 U8106 ( .A1(n8623), .A2(n6374), .ZN(n6401) );
  NAND2_X1 U8107 ( .A1(n8326), .A2(n6404), .ZN(n6394) );
  INV_X1 U8108 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9103) );
  OR2_X1 U8109 ( .A1(n6406), .A2(n9103), .ZN(n6393) );
  INV_X1 U8110 ( .A(n6530), .ZN(n6395) );
  AOI21_X1 U8111 ( .B1(n6401), .B2(n8627), .A(n6395), .ZN(n6403) );
  NAND2_X1 U8112 ( .A1(n4375), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U8113 ( .A1(n6397), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U8114 ( .A1(n5976), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6398) );
  NAND3_X1 U8115 ( .A1(n6400), .A2(n6399), .A3(n6398), .ZN(n8521) );
  INV_X1 U8116 ( .A(n8521), .ZN(n6409) );
  NOR2_X1 U8117 ( .A1(n8627), .A2(n6409), .ZN(n6528) );
  INV_X1 U8118 ( .A(n6401), .ZN(n6402) );
  NAND2_X1 U8119 ( .A1(n9030), .A2(n6404), .ZN(n6408) );
  INV_X1 U8120 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6405) );
  OR2_X1 U8121 ( .A1(n6406), .A2(n6405), .ZN(n6407) );
  INV_X1 U8122 ( .A(n8623), .ZN(n6410) );
  OR2_X1 U8123 ( .A1(n8899), .A2(n6410), .ZN(n6533) );
  NAND2_X1 U8124 ( .A1(n8627), .A2(n6409), .ZN(n6534) );
  NAND2_X1 U8125 ( .A1(n6533), .A2(n6534), .ZN(n6559) );
  NAND2_X1 U8126 ( .A1(n8899), .A2(n6410), .ZN(n6536) );
  OAI21_X1 U8127 ( .B1(n6411), .B2(n6559), .A(n6536), .ZN(n6412) );
  XNOR2_X1 U8128 ( .A(n6412), .B(n8620), .ZN(n6416) );
  NOR2_X1 U8129 ( .A1(n6680), .A2(P2_U3152), .ZN(n7280) );
  INV_X1 U8130 ( .A(n6413), .ZN(n6414) );
  OR2_X1 U8131 ( .A1(n7538), .A2(n6414), .ZN(n6415) );
  INV_X1 U8132 ( .A(n6417), .ZN(n6421) );
  NAND2_X1 U8133 ( .A1(n6544), .A2(n6418), .ZN(n6420) );
  AND2_X1 U8134 ( .A1(n6328), .A2(n8620), .ZN(n6419) );
  MUX2_X1 U8135 ( .A(n6421), .B(n6420), .S(n4382), .Z(n6422) );
  INV_X1 U8136 ( .A(n6422), .ZN(n6485) );
  MUX2_X1 U8137 ( .A(n6424), .B(n6423), .S(n4382), .Z(n6484) );
  INV_X1 U8138 ( .A(n8803), .ZN(n8790) );
  NAND2_X1 U8139 ( .A1(n6425), .A2(n6428), .ZN(n6427) );
  NAND2_X1 U8140 ( .A1(n6445), .A2(n6443), .ZN(n6426) );
  AND2_X1 U8141 ( .A1(n7952), .A2(n6425), .ZN(n6429) );
  OAI211_X1 U8142 ( .C1(n6447), .C2(n6429), .A(n6428), .B(n7884), .ZN(n6430)
         );
  NAND2_X1 U8143 ( .A1(n6430), .A2(n4382), .ZN(n6441) );
  NAND2_X1 U8144 ( .A1(n8537), .A2(n10188), .ZN(n8120) );
  AND2_X1 U8145 ( .A1(n8120), .A2(n6328), .ZN(n6431) );
  OAI211_X1 U8146 ( .C1(n6431), .C2(n8151), .A(n6434), .B(n8145), .ZN(n6432)
         );
  NAND2_X1 U8147 ( .A1(n6432), .A2(n7801), .ZN(n6437) );
  NAND2_X1 U8148 ( .A1(n8145), .A2(n8120), .ZN(n6433) );
  NAND3_X1 U8149 ( .A1(n6433), .A2(n7801), .A3(n8146), .ZN(n6435) );
  NAND2_X1 U8150 ( .A1(n6435), .A2(n6434), .ZN(n6436) );
  INV_X1 U8151 ( .A(n6447), .ZN(n6438) );
  NAND3_X1 U8152 ( .A1(n6439), .A2(n6438), .A3(n7797), .ZN(n6440) );
  AND2_X1 U8153 ( .A1(n6443), .A2(n6442), .ZN(n6446) );
  OAI211_X1 U8154 ( .C1(n6447), .C2(n6446), .A(n6445), .B(n6444), .ZN(n6448)
         );
  MUX2_X1 U8155 ( .A(n8059), .B(n6449), .S(n4382), .Z(n6450) );
  NAND3_X1 U8156 ( .A1(n6451), .A2(n8063), .A3(n6450), .ZN(n6454) );
  MUX2_X1 U8157 ( .A(n8104), .B(n6452), .S(n4382), .Z(n6453) );
  OR2_X1 U8158 ( .A1(n8876), .A2(n4400), .ZN(n6455) );
  OAI21_X1 U8159 ( .B1(n6459), .B2(n4382), .A(n6455), .ZN(n6456) );
  NOR2_X1 U8160 ( .A1(n8879), .A2(n6456), .ZN(n6461) );
  AND3_X1 U8161 ( .A1(n8137), .A2(n6458), .A3(n4382), .ZN(n6464) );
  INV_X1 U8162 ( .A(n6459), .ZN(n6460) );
  NAND2_X1 U8163 ( .A1(n6461), .A2(n6460), .ZN(n6462) );
  NAND2_X1 U8164 ( .A1(n8137), .A2(n8854), .ZN(n6465) );
  NAND3_X1 U8165 ( .A1(n10281), .A2(n4400), .A3(n6465), .ZN(n6471) );
  NAND2_X1 U8166 ( .A1(n6545), .A2(n8526), .ZN(n6466) );
  NAND3_X1 U8167 ( .A1(n8134), .A2(n6466), .A3(n4382), .ZN(n6470) );
  OR3_X1 U8168 ( .A1(n6545), .A2(n4400), .A3(n8526), .ZN(n6469) );
  INV_X1 U8169 ( .A(n8137), .ZN(n6467) );
  NAND3_X1 U8170 ( .A1(n6467), .A2(n4400), .A3(n8526), .ZN(n6468) );
  NAND2_X1 U8171 ( .A1(n8857), .A2(n6472), .ZN(n6476) );
  MUX2_X1 U8172 ( .A(n6474), .B(n6473), .S(n4382), .Z(n6475) );
  NAND3_X1 U8173 ( .A1(n6476), .A2(n8077), .A3(n6475), .ZN(n6480) );
  NAND2_X1 U8174 ( .A1(n8524), .A2(n4382), .ZN(n6478) );
  NAND2_X1 U8175 ( .A1(n8853), .A2(n4400), .ZN(n6477) );
  MUX2_X1 U8176 ( .A(n6478), .B(n6477), .S(n8997), .Z(n6479) );
  MUX2_X1 U8177 ( .A(n6482), .B(n6481), .S(n4382), .Z(n6483) );
  AOI21_X1 U8178 ( .B1(n6499), .B2(n6544), .A(n6486), .ZN(n6490) );
  NAND2_X1 U8179 ( .A1(n6497), .A2(n6500), .ZN(n6489) );
  AND3_X1 U8180 ( .A1(n8721), .A2(n4400), .A3(n6502), .ZN(n6487) );
  OAI211_X1 U8181 ( .C1(n6490), .C2(n6489), .A(n6488), .B(n6487), .ZN(n6495)
         );
  NAND2_X1 U8182 ( .A1(n8751), .A2(n4400), .ZN(n6492) );
  OAI22_X1 U8183 ( .A1(n8741), .A2(n6492), .B1(n8427), .B2(n4382), .ZN(n6491)
         );
  NAND2_X1 U8184 ( .A1(n8719), .A2(n6491), .ZN(n6494) );
  OR3_X1 U8185 ( .A1(n8741), .A2(n8427), .A3(n6492), .ZN(n6493) );
  AND3_X1 U8186 ( .A1(n6495), .A2(n6494), .A3(n6493), .ZN(n6510) );
  INV_X1 U8187 ( .A(n6496), .ZN(n8686) );
  NOR2_X1 U8188 ( .A1(n8751), .A2(n4400), .ZN(n6506) );
  AOI22_X1 U8189 ( .A1(n8741), .A2(n6506), .B1(n8427), .B2(n4382), .ZN(n6509)
         );
  OAI211_X1 U8190 ( .C1(n8741), .C2(n8497), .A(n6497), .B(n4382), .ZN(n6498)
         );
  INV_X1 U8191 ( .A(n6498), .ZN(n6505) );
  NAND3_X1 U8192 ( .A1(n6499), .A2(n6543), .A3(n8748), .ZN(n6501) );
  NAND2_X1 U8193 ( .A1(n6501), .A2(n6500), .ZN(n6503) );
  NAND2_X1 U8194 ( .A1(n6503), .A2(n6502), .ZN(n6504) );
  NAND3_X1 U8195 ( .A1(n8696), .A2(n6505), .A3(n6504), .ZN(n6508) );
  NAND3_X1 U8196 ( .A1(n8741), .A2(n8427), .A3(n6506), .ZN(n6507) );
  NAND2_X1 U8197 ( .A1(n6512), .A2(n6511), .ZN(n6513) );
  NAND2_X1 U8198 ( .A1(n6513), .A2(n4400), .ZN(n6514) );
  NAND2_X1 U8199 ( .A1(n6515), .A2(n6514), .ZN(n6517) );
  AOI21_X1 U8200 ( .B1(n6519), .B2(n4420), .A(n4382), .ZN(n6518) );
  AOI21_X1 U8201 ( .B1(n6520), .B2(n6519), .A(n6518), .ZN(n6521) );
  MUX2_X1 U8202 ( .A(n6523), .B(n6522), .S(n4382), .Z(n6524) );
  MUX2_X1 U8203 ( .A(n6526), .B(n6525), .S(n4400), .Z(n6527) );
  INV_X1 U8204 ( .A(n6528), .ZN(n6535) );
  AND2_X1 U8205 ( .A1(n6535), .A2(n6534), .ZN(n6532) );
  MUX2_X1 U8206 ( .A(n6530), .B(n6529), .S(n4400), .Z(n6531) );
  NAND2_X1 U8207 ( .A1(n6536), .A2(n6535), .ZN(n6558) );
  INV_X1 U8208 ( .A(n6558), .ZN(n6537) );
  AND2_X1 U8209 ( .A1(n8623), .A2(n4382), .ZN(n6539) );
  OAI21_X1 U8210 ( .B1(n8623), .B2(n4382), .A(n8899), .ZN(n6538) );
  OAI21_X1 U8211 ( .B1(n6539), .B2(n8899), .A(n6538), .ZN(n6540) );
  INV_X1 U8212 ( .A(n7280), .ZN(n8055) );
  INV_X1 U8213 ( .A(n9040), .ZN(n8383) );
  NAND4_X1 U8214 ( .A1(n8904), .A2(n8383), .A3(n8815), .A4(n6686), .ZN(n6541)
         );
  OAI211_X1 U8215 ( .C1(n6354), .C2(n8055), .A(n6541), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6566) );
  NAND2_X1 U8216 ( .A1(n6544), .A2(n6543), .ZN(n8785) );
  INV_X1 U8217 ( .A(n6545), .ZN(n6551) );
  INV_X1 U8218 ( .A(n8102), .ZN(n8105) );
  NOR2_X1 U8219 ( .A1(n8151), .A2(n6546), .ZN(n6547) );
  NAND4_X1 U8220 ( .A1(n6547), .A2(n6561), .A3(n8120), .A4(n8145), .ZN(n6549)
         );
  NOR4_X1 U8221 ( .A1(n6549), .A2(n7851), .A3(n7954), .A4(n7802), .ZN(n6550)
         );
  NOR4_X1 U8222 ( .A1(n8765), .A2(n8785), .A3(n8803), .A4(n6554), .ZN(n6555)
         );
  XNOR2_X1 U8223 ( .A(n6560), .B(n8620), .ZN(n6562) );
  OAI22_X1 U8224 ( .A1(n6562), .A2(n6328), .B1(n6561), .B2(n6568), .ZN(n6564)
         );
  NAND3_X1 U8225 ( .A1(n6564), .A2(n7280), .A3(n6563), .ZN(n6565) );
  BUF_X4 U8226 ( .A(n6589), .Z(n8352) );
  XNOR2_X1 U8227 ( .A(n8940), .B(n6673), .ZN(n8470) );
  NAND2_X1 U8228 ( .A1(n8726), .A2(n4383), .ZN(n8468) );
  AOI21_X1 U8229 ( .B1(n8470), .B2(n8440), .A(n8468), .ZN(n6667) );
  XNOR2_X1 U8230 ( .A(n8945), .B(n8352), .ZN(n6663) );
  NAND2_X1 U8231 ( .A1(n4377), .A2(n4383), .ZN(n7249) );
  NOR2_X1 U8232 ( .A1(n7250), .A2(n7249), .ZN(n6575) );
  INV_X1 U8233 ( .A(n6571), .ZN(n6572) );
  OR2_X1 U8234 ( .A1(n6589), .A2(n8124), .ZN(n6573) );
  NAND2_X1 U8235 ( .A1(n7541), .A2(n6573), .ZN(n7251) );
  NAND2_X1 U8236 ( .A1(n7250), .A2(n7249), .ZN(n7252) );
  NAND2_X1 U8237 ( .A1(n10146), .A2(n4384), .ZN(n6576) );
  NAND2_X1 U8238 ( .A1(n6577), .A2(n6576), .ZN(n7253) );
  OAI211_X1 U8239 ( .C1(n6575), .C2(n7251), .A(n7252), .B(n7253), .ZN(n6580)
         );
  INV_X1 U8240 ( .A(n6576), .ZN(n6579) );
  INV_X1 U8241 ( .A(n6577), .ZN(n6578) );
  NAND2_X1 U8242 ( .A1(n6579), .A2(n6578), .ZN(n7254) );
  NAND2_X1 U8243 ( .A1(n6580), .A2(n7254), .ZN(n10154) );
  AND2_X1 U8244 ( .A1(n8535), .A2(n4383), .ZN(n6581) );
  NAND2_X1 U8245 ( .A1(n6581), .A2(n6582), .ZN(n6586) );
  INV_X1 U8246 ( .A(n6581), .ZN(n6584) );
  INV_X1 U8247 ( .A(n6582), .ZN(n6583) );
  AND2_X1 U8248 ( .A1(n6586), .A2(n6585), .ZN(n10155) );
  NAND2_X1 U8249 ( .A1(n10154), .A2(n10155), .ZN(n10152) );
  NAND2_X1 U8250 ( .A1(n10152), .A2(n6586), .ZN(n7497) );
  INV_X1 U8251 ( .A(n7497), .ZN(n6588) );
  XNOR2_X1 U8252 ( .A(n6589), .B(n10218), .ZN(n6594) );
  NAND2_X1 U8253 ( .A1(n8534), .A2(n8351), .ZN(n6593) );
  XNOR2_X1 U8254 ( .A(n6594), .B(n6593), .ZN(n7498) );
  INV_X1 U8255 ( .A(n7498), .ZN(n6587) );
  NAND2_X1 U8256 ( .A1(n6588), .A2(n6587), .ZN(n7438) );
  XNOR2_X1 U8257 ( .A(n7854), .B(n6589), .ZN(n6590) );
  NAND2_X1 U8258 ( .A1(n6590), .A2(n6591), .ZN(n6597) );
  NAND2_X1 U8259 ( .A1(n6597), .A2(n6592), .ZN(n7443) );
  NAND2_X1 U8260 ( .A1(n6594), .A2(n6593), .ZN(n7439) );
  INV_X1 U8261 ( .A(n7439), .ZN(n6595) );
  XNOR2_X1 U8262 ( .A(n7933), .B(n8352), .ZN(n6598) );
  NAND2_X1 U8263 ( .A1(n8532), .A2(n8351), .ZN(n6599) );
  XNOR2_X1 U8264 ( .A(n6598), .B(n6599), .ZN(n7518) );
  INV_X1 U8265 ( .A(n6598), .ZN(n6600) );
  NAND2_X1 U8266 ( .A1(n6600), .A2(n6599), .ZN(n6601) );
  XNOR2_X1 U8267 ( .A(n6602), .B(n8352), .ZN(n6603) );
  AND2_X1 U8268 ( .A1(n8531), .A2(n8351), .ZN(n6604) );
  NAND2_X1 U8269 ( .A1(n6603), .A2(n6604), .ZN(n6608) );
  INV_X1 U8270 ( .A(n6603), .ZN(n6606) );
  INV_X1 U8271 ( .A(n6604), .ZN(n6605) );
  NAND2_X1 U8272 ( .A1(n6606), .A2(n6605), .ZN(n6607) );
  AND2_X1 U8273 ( .A1(n6608), .A2(n6607), .ZN(n7533) );
  NAND2_X1 U8274 ( .A1(n7534), .A2(n7533), .ZN(n7532) );
  XNOR2_X1 U8275 ( .A(n10246), .B(n8352), .ZN(n6611) );
  NAND2_X1 U8276 ( .A1(n8530), .A2(n8351), .ZN(n6609) );
  XNOR2_X1 U8277 ( .A(n6611), .B(n6609), .ZN(n7546) );
  INV_X1 U8278 ( .A(n6609), .ZN(n6610) );
  XNOR2_X1 U8279 ( .A(n8114), .B(n8352), .ZN(n6612) );
  AND2_X1 U8280 ( .A1(n8529), .A2(n8351), .ZN(n6613) );
  AND2_X1 U8281 ( .A1(n6612), .A2(n6613), .ZN(n7664) );
  INV_X1 U8282 ( .A(n6612), .ZN(n6615) );
  INV_X1 U8283 ( .A(n6613), .ZN(n6614) );
  XNOR2_X1 U8284 ( .A(n10263), .B(n6673), .ZN(n6617) );
  NAND2_X1 U8285 ( .A1(n8528), .A2(n8351), .ZN(n6616) );
  XNOR2_X1 U8286 ( .A(n6617), .B(n6616), .ZN(n7831) );
  OAI22_X2 U8287 ( .A1(n7830), .A2(n7831), .B1(n6617), .B2(n6616), .ZN(n7920)
         );
  XNOR2_X1 U8288 ( .A(n7923), .B(n8352), .ZN(n6620) );
  NAND2_X1 U8289 ( .A1(n8527), .A2(n8351), .ZN(n6618) );
  XNOR2_X1 U8290 ( .A(n6620), .B(n6618), .ZN(n7919) );
  INV_X1 U8291 ( .A(n6618), .ZN(n6619) );
  NAND2_X1 U8292 ( .A1(n6620), .A2(n6619), .ZN(n8006) );
  XNOR2_X1 U8293 ( .A(n8134), .B(n6673), .ZN(n6621) );
  NAND2_X1 U8294 ( .A1(n8526), .A2(n8351), .ZN(n6622) );
  NAND2_X1 U8295 ( .A1(n6621), .A2(n6622), .ZN(n6628) );
  INV_X1 U8296 ( .A(n6621), .ZN(n6624) );
  INV_X1 U8297 ( .A(n6622), .ZN(n6623) );
  NAND2_X1 U8298 ( .A1(n6624), .A2(n6623), .ZN(n6625) );
  NAND2_X1 U8299 ( .A1(n6628), .A2(n6625), .ZN(n8010) );
  INV_X1 U8300 ( .A(n8010), .ZN(n6626) );
  AND2_X1 U8301 ( .A1(n8006), .A2(n6626), .ZN(n6627) );
  XNOR2_X1 U8302 ( .A(n9002), .B(n6673), .ZN(n6629) );
  NAND2_X1 U8303 ( .A1(n8525), .A2(n8351), .ZN(n6630) );
  XNOR2_X1 U8304 ( .A(n6629), .B(n6630), .ZN(n8095) );
  INV_X1 U8305 ( .A(n6629), .ZN(n6632) );
  INV_X1 U8306 ( .A(n6630), .ZN(n6631) );
  XNOR2_X1 U8307 ( .A(n8997), .B(n6673), .ZN(n6633) );
  NAND2_X1 U8308 ( .A1(n8524), .A2(n8351), .ZN(n6634) );
  NAND2_X1 U8309 ( .A1(n6633), .A2(n6634), .ZN(n6638) );
  INV_X1 U8310 ( .A(n6633), .ZN(n6636) );
  INV_X1 U8311 ( .A(n6634), .ZN(n6635) );
  NAND2_X1 U8312 ( .A1(n6636), .A2(n6635), .ZN(n6637) );
  AND2_X1 U8313 ( .A1(n6638), .A2(n6637), .ZN(n8398) );
  NAND2_X1 U8314 ( .A1(n8396), .A2(n6638), .ZN(n8446) );
  XNOR2_X1 U8315 ( .A(n8992), .B(n6673), .ZN(n8445) );
  NAND2_X1 U8316 ( .A1(n8814), .A2(n4384), .ZN(n6639) );
  AND2_X1 U8317 ( .A1(n8445), .A2(n6639), .ZN(n6642) );
  INV_X1 U8318 ( .A(n8445), .ZN(n6640) );
  INV_X1 U8319 ( .A(n6639), .ZN(n8512) );
  NAND2_X1 U8320 ( .A1(n6640), .A2(n8512), .ZN(n6641) );
  XNOR2_X1 U8321 ( .A(n8984), .B(n8352), .ZN(n6645) );
  NAND2_X1 U8322 ( .A1(n8523), .A2(n8351), .ZN(n6643) );
  XNOR2_X1 U8323 ( .A(n6645), .B(n6643), .ZN(n8448) );
  INV_X1 U8324 ( .A(n6643), .ZN(n6644) );
  NAND2_X1 U8325 ( .A1(n8817), .A2(n8351), .ZN(n6648) );
  XNOR2_X1 U8326 ( .A(n8980), .B(n8352), .ZN(n6647) );
  XOR2_X1 U8327 ( .A(n6648), .B(n6647), .Z(n8460) );
  XNOR2_X1 U8328 ( .A(n8974), .B(n8352), .ZN(n6650) );
  NAND2_X1 U8329 ( .A1(n8768), .A2(n4383), .ZN(n6649) );
  XNOR2_X1 U8330 ( .A(n6650), .B(n6649), .ZN(n8502) );
  INV_X1 U8331 ( .A(n6649), .ZN(n6651) );
  AND2_X1 U8332 ( .A1(n8779), .A2(n4384), .ZN(n6653) );
  XNOR2_X1 U8333 ( .A(n8970), .B(n8352), .ZN(n6652) );
  NAND2_X1 U8334 ( .A1(n8769), .A2(n4383), .ZN(n6655) );
  XNOR2_X1 U8335 ( .A(n8963), .B(n8352), .ZN(n6654) );
  XOR2_X1 U8336 ( .A(n6655), .B(n6654), .Z(n8480) );
  INV_X1 U8337 ( .A(n6654), .ZN(n6656) );
  XNOR2_X1 U8338 ( .A(n8741), .B(n8352), .ZN(n6660) );
  NAND2_X1 U8339 ( .A1(n8751), .A2(n8351), .ZN(n6658) );
  XNOR2_X1 U8340 ( .A(n6660), .B(n6658), .ZN(n8424) );
  XNOR2_X1 U8341 ( .A(n8950), .B(n8352), .ZN(n8491) );
  NOR2_X1 U8342 ( .A1(n8427), .A2(n7538), .ZN(n8492) );
  NOR2_X1 U8343 ( .A1(n8491), .A2(n8492), .ZN(n6662) );
  INV_X1 U8344 ( .A(n6660), .ZN(n6657) );
  NOR2_X1 U8345 ( .A1(n6657), .A2(n6658), .ZN(n8488) );
  OAI21_X1 U8346 ( .B1(n8488), .B2(n8492), .A(n8491), .ZN(n6661) );
  INV_X1 U8347 ( .A(n6658), .ZN(n6659) );
  NAND2_X1 U8348 ( .A1(n8699), .A2(n4384), .ZN(n8471) );
  NOR2_X1 U8349 ( .A1(n8470), .A2(n8471), .ZN(n6666) );
  XNOR2_X1 U8350 ( .A(n8673), .B(n8352), .ZN(n6670) );
  NAND2_X1 U8351 ( .A1(n8689), .A2(n4383), .ZN(n8433) );
  INV_X1 U8352 ( .A(n6670), .ZN(n8434) );
  AND2_X1 U8353 ( .A1(n8436), .A2(n8434), .ZN(n6671) );
  XNOR2_X1 U8354 ( .A(n8930), .B(n6673), .ZN(n6675) );
  NAND2_X1 U8355 ( .A1(n8666), .A2(n8351), .ZN(n6674) );
  NOR2_X1 U8356 ( .A1(n6675), .A2(n6674), .ZN(n6699) );
  AOI21_X1 U8357 ( .B1(n6675), .B2(n6674), .A(n6699), .ZN(n6702) );
  NAND2_X1 U8358 ( .A1(n6707), .A2(n6702), .ZN(n6701) );
  AND2_X1 U8359 ( .A1(n10280), .A2(n7279), .ZN(n6676) );
  OAI211_X1 U8360 ( .C1(n6707), .C2(n6702), .A(n6701), .B(n10153), .ZN(n6694)
         );
  INV_X1 U8361 ( .A(n8930), .ZN(n6691) );
  NAND2_X1 U8362 ( .A1(n6677), .A2(n8908), .ZN(n6678) );
  NAND2_X1 U8363 ( .A1(n6678), .A2(n8903), .ZN(n7257) );
  NOR2_X1 U8364 ( .A1(n10175), .A2(n10280), .ZN(n6679) );
  NAND2_X1 U8365 ( .A1(n8902), .A2(n6680), .ZN(n6681) );
  NOR2_X1 U8366 ( .A1(n7281), .A2(n6681), .ZN(n6682) );
  NAND2_X1 U8367 ( .A1(n7257), .A2(n6682), .ZN(n6683) );
  NOR2_X1 U8368 ( .A1(n10161), .A2(n8661), .ZN(n6689) );
  INV_X1 U8369 ( .A(n6684), .ZN(n6685) );
  NOR2_X1 U8370 ( .A1(n6685), .A2(n9007), .ZN(n6687) );
  NAND2_X1 U8371 ( .A1(n6687), .A2(n6686), .ZN(n8516) );
  OAI22_X1 U8372 ( .A1(n8367), .A2(n10145), .B1(n10148), .B2(n8475), .ZN(n6688) );
  AOI211_X1 U8373 ( .C1(P2_REG3_REG_26__SCAN_IN), .C2(P2_U3152), .A(n6689), 
        .B(n6688), .ZN(n6690) );
  XNOR2_X1 U8374 ( .A(n8924), .B(n8352), .ZN(n6696) );
  INV_X1 U8375 ( .A(n6696), .ZN(n6698) );
  AND2_X1 U8376 ( .A1(n8657), .A2(n8351), .ZN(n6695) );
  INV_X1 U8377 ( .A(n6695), .ZN(n6697) );
  AOI21_X1 U8378 ( .B1(n6698), .B2(n6697), .A(n8371), .ZN(n6703) );
  INV_X1 U8379 ( .A(n6699), .ZN(n6704) );
  NAND2_X1 U8380 ( .A1(n6701), .A2(n6700), .ZN(n6708) );
  AND2_X1 U8381 ( .A1(n6702), .A2(n6703), .ZN(n6706) );
  INV_X1 U8382 ( .A(n6703), .ZN(n6705) );
  AOI21_X2 U8383 ( .B1(n6707), .B2(n6706), .A(n5031), .ZN(n8376) );
  NAND3_X1 U8384 ( .A1(n6708), .A2(n10153), .A3(n8376), .ZN(n6714) );
  OAI22_X1 U8385 ( .A1(n10161), .A2(n8640), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6709), .ZN(n6712) );
  OAI22_X1 U8386 ( .A1(n6710), .A2(n10145), .B1(n8439), .B2(n10148), .ZN(n6711) );
  AOI211_X1 U8387 ( .C1(n8924), .C2(n10151), .A(n6712), .B(n6711), .ZN(n6713)
         );
  NAND2_X1 U8388 ( .A1(n6714), .A2(n6713), .ZN(P2_U3216) );
  INV_X1 U8389 ( .A(n7007), .ZN(n6717) );
  AND2_X1 U8390 ( .A1(n6929), .A2(n9657), .ZN(n6718) );
  AOI21_X1 U8391 ( .B1(n9758), .B2(n6758), .A(n6718), .ZN(n9339) );
  NAND2_X1 U8392 ( .A1(n9755), .A2(n4380), .ZN(n6720) );
  NAND2_X1 U8393 ( .A1(n9476), .A2(n6947), .ZN(n6719) );
  NAND2_X1 U8394 ( .A1(n6720), .A2(n6719), .ZN(n6721) );
  INV_X4 U8395 ( .A(n6733), .ZN(n6945) );
  XNOR2_X1 U8396 ( .A(n6721), .B(n6945), .ZN(n6726) );
  INV_X1 U8397 ( .A(n6726), .ZN(n6724) );
  AND2_X1 U8398 ( .A1(n6929), .A2(n9476), .ZN(n6722) );
  AOI21_X1 U8399 ( .B1(n9755), .B2(n6758), .A(n6722), .ZN(n6725) );
  INV_X1 U8400 ( .A(n6725), .ZN(n6723) );
  NAND2_X1 U8401 ( .A1(n6724), .A2(n6723), .ZN(n9370) );
  AOI21_X1 U8402 ( .B1(n9339), .B2(n9370), .A(n9372), .ZN(n6923) );
  AND2_X1 U8403 ( .A1(n6729), .A2(n6728), .ZN(n7168) );
  INV_X1 U8404 ( .A(n6908), .ZN(n6736) );
  NAND2_X1 U8405 ( .A1(n7217), .A2(n6758), .ZN(n6731) );
  INV_X1 U8406 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6730) );
  NAND3_X1 U8407 ( .A1(n6732), .A2(n6731), .A3(n5034), .ZN(n7167) );
  INV_X1 U8408 ( .A(n7167), .ZN(n6734) );
  NAND2_X1 U8409 ( .A1(n6734), .A2(n4387), .ZN(n6735) );
  NAND2_X1 U8410 ( .A1(n7166), .A2(n6735), .ZN(n6742) );
  NAND2_X1 U8411 ( .A1(n5818), .A2(n6758), .ZN(n6738) );
  NAND2_X1 U8412 ( .A1(n4997), .A2(n6736), .ZN(n6737) );
  XNOR2_X1 U8413 ( .A(n6739), .B(n6945), .ZN(n6741) );
  INV_X1 U8414 ( .A(n6741), .ZN(n6740) );
  AOI22_X1 U8415 ( .A1(n6929), .A2(n5818), .B1(n4997), .B2(n6758), .ZN(n7215)
         );
  NAND2_X1 U8416 ( .A1(n6742), .A2(n6741), .ZN(n7213) );
  NAND2_X1 U8417 ( .A1(n9490), .A2(n6758), .ZN(n6744) );
  NAND2_X1 U8418 ( .A1(n6736), .A2(n7553), .ZN(n6743) );
  NAND2_X1 U8419 ( .A1(n6744), .A2(n6743), .ZN(n6745) );
  XNOR2_X1 U8420 ( .A(n6745), .B(n6945), .ZN(n6747) );
  AND2_X1 U8421 ( .A1(n6758), .A2(n7553), .ZN(n6746) );
  AOI21_X1 U8422 ( .B1(n6929), .B2(n9490), .A(n6746), .ZN(n6748) );
  NAND2_X1 U8423 ( .A1(n6747), .A2(n6748), .ZN(n6752) );
  INV_X1 U8424 ( .A(n6747), .ZN(n6750) );
  INV_X1 U8425 ( .A(n6748), .ZN(n6749) );
  NAND2_X1 U8426 ( .A1(n6750), .A2(n6749), .ZN(n6751) );
  AND2_X1 U8427 ( .A1(n6752), .A2(n6751), .ZN(n8335) );
  NAND2_X1 U8428 ( .A1(n8333), .A2(n6752), .ZN(n7205) );
  OAI22_X1 U8429 ( .A1(n10041), .A2(n6917), .B1(n10076), .B2(n6908), .ZN(n6753) );
  XNOR2_X1 U8430 ( .A(n6753), .B(n4387), .ZN(n7204) );
  INV_X1 U8431 ( .A(n7204), .ZN(n6757) );
  INV_X2 U8432 ( .A(n6754), .ZN(n6942) );
  OR2_X1 U8433 ( .A1(n10041), .A2(n6942), .ZN(n6756) );
  NAND2_X1 U8434 ( .A1(n6947), .A2(n7647), .ZN(n6755) );
  NAND2_X1 U8435 ( .A1(n6756), .A2(n6755), .ZN(n6762) );
  INV_X1 U8436 ( .A(n6762), .ZN(n7203) );
  NAND2_X1 U8437 ( .A1(n6757), .A2(n7203), .ZN(n7580) );
  OR2_X1 U8438 ( .A1(n10016), .A2(n6942), .ZN(n6761) );
  NAND2_X1 U8439 ( .A1(n5365), .A2(n6758), .ZN(n6760) );
  NAND2_X1 U8440 ( .A1(n6761), .A2(n6760), .ZN(n6764) );
  INV_X1 U8441 ( .A(n6764), .ZN(n7582) );
  NAND2_X1 U8442 ( .A1(n7583), .A2(n7582), .ZN(n6763) );
  NAND2_X1 U8443 ( .A1(n7580), .A2(n6763), .ZN(n6774) );
  NAND3_X1 U8444 ( .A1(n6763), .A2(n7204), .A3(n6762), .ZN(n6766) );
  INV_X1 U8445 ( .A(n7583), .ZN(n6765) );
  NAND2_X1 U8446 ( .A1(n6765), .A2(n6764), .ZN(n7584) );
  AND2_X1 U8447 ( .A1(n6766), .A2(n7584), .ZN(n6773) );
  NAND2_X1 U8448 ( .A1(n10038), .A2(n6758), .ZN(n6768) );
  NAND2_X1 U8449 ( .A1(n10006), .A2(n4380), .ZN(n6767) );
  NAND2_X1 U8450 ( .A1(n6768), .A2(n6767), .ZN(n6769) );
  XNOR2_X1 U8451 ( .A(n6769), .B(n4387), .ZN(n6779) );
  NAND2_X1 U8452 ( .A1(n6929), .A2(n10038), .ZN(n6771) );
  NAND2_X1 U8453 ( .A1(n10006), .A2(n6947), .ZN(n6770) );
  NAND2_X1 U8454 ( .A1(n6771), .A2(n6770), .ZN(n7588) );
  NAND2_X1 U8455 ( .A1(n6779), .A2(n7588), .ZN(n6772) );
  OAI211_X1 U8456 ( .C1(n7205), .C2(n6774), .A(n6773), .B(n6772), .ZN(n6782)
         );
  NAND2_X1 U8457 ( .A1(n9994), .A2(n4380), .ZN(n6775) );
  OAI21_X1 U8458 ( .B1(n10017), .B2(n6917), .A(n6775), .ZN(n6776) );
  XNOR2_X1 U8459 ( .A(n6776), .B(n6945), .ZN(n6783) );
  OR2_X1 U8460 ( .A1(n10017), .A2(n6942), .ZN(n6778) );
  NAND2_X1 U8461 ( .A1(n9994), .A2(n6947), .ZN(n6777) );
  AND2_X1 U8462 ( .A1(n6778), .A2(n6777), .ZN(n6784) );
  NAND2_X1 U8463 ( .A1(n6783), .A2(n6784), .ZN(n7720) );
  INV_X1 U8464 ( .A(n6779), .ZN(n7585) );
  INV_X1 U8465 ( .A(n7588), .ZN(n6780) );
  NAND2_X1 U8466 ( .A1(n7585), .A2(n6780), .ZN(n6781) );
  INV_X1 U8467 ( .A(n6783), .ZN(n6786) );
  INV_X1 U8468 ( .A(n6784), .ZN(n6785) );
  NAND2_X1 U8469 ( .A1(n6786), .A2(n6785), .ZN(n7721) );
  NAND2_X1 U8470 ( .A1(n10105), .A2(n6947), .ZN(n6789) );
  OR2_X1 U8471 ( .A1(n9988), .A2(n6942), .ZN(n6788) );
  NAND2_X1 U8472 ( .A1(n6789), .A2(n6788), .ZN(n7240) );
  NAND2_X1 U8473 ( .A1(n10105), .A2(n4380), .ZN(n6791) );
  OR2_X1 U8474 ( .A1(n9988), .A2(n6917), .ZN(n6790) );
  NAND2_X1 U8475 ( .A1(n6791), .A2(n6790), .ZN(n6792) );
  XNOR2_X1 U8476 ( .A(n6792), .B(n4387), .ZN(n7239) );
  NAND2_X1 U8477 ( .A1(n7242), .A2(n7240), .ZN(n6793) );
  NAND2_X1 U8478 ( .A1(n9976), .A2(n4380), .ZN(n6795) );
  OR2_X1 U8479 ( .A1(n7739), .A2(n6917), .ZN(n6794) );
  NAND2_X1 U8480 ( .A1(n6795), .A2(n6794), .ZN(n6796) );
  XNOR2_X1 U8481 ( .A(n6796), .B(n4387), .ZN(n7598) );
  NAND2_X1 U8482 ( .A1(n9976), .A2(n6947), .ZN(n6798) );
  OR2_X1 U8483 ( .A1(n7739), .A2(n6942), .ZN(n6797) );
  NAND2_X1 U8484 ( .A1(n6798), .A2(n6797), .ZN(n7599) );
  NAND2_X1 U8485 ( .A1(n7747), .A2(n4380), .ZN(n6800) );
  NAND2_X1 U8486 ( .A1(n9487), .A2(n6947), .ZN(n6799) );
  NAND2_X1 U8487 ( .A1(n6800), .A2(n6799), .ZN(n6801) );
  XNOR2_X1 U8488 ( .A(n6801), .B(n4387), .ZN(n6807) );
  NAND2_X1 U8489 ( .A1(n7747), .A2(n6947), .ZN(n6803) );
  NAND2_X1 U8490 ( .A1(n6929), .A2(n9487), .ZN(n6802) );
  NAND2_X1 U8491 ( .A1(n6803), .A2(n6802), .ZN(n6808) );
  AND2_X1 U8492 ( .A1(n6807), .A2(n6808), .ZN(n7596) );
  INV_X1 U8493 ( .A(n7596), .ZN(n6804) );
  INV_X1 U8494 ( .A(n7598), .ZN(n6805) );
  INV_X1 U8495 ( .A(n7599), .ZN(n7602) );
  NAND2_X1 U8496 ( .A1(n6805), .A2(n7602), .ZN(n6806) );
  INV_X1 U8497 ( .A(n6807), .ZN(n6810) );
  INV_X1 U8498 ( .A(n6808), .ZN(n6809) );
  NAND2_X1 U8499 ( .A1(n6810), .A2(n6809), .ZN(n7597) );
  NAND2_X1 U8500 ( .A1(n7815), .A2(n4380), .ZN(n6813) );
  OR2_X1 U8501 ( .A1(n7814), .A2(n6917), .ZN(n6812) );
  NAND2_X1 U8502 ( .A1(n6813), .A2(n6812), .ZN(n6814) );
  XNOR2_X1 U8503 ( .A(n6814), .B(n4387), .ZN(n6817) );
  NAND2_X1 U8504 ( .A1(n7815), .A2(n6947), .ZN(n6816) );
  OR2_X1 U8505 ( .A1(n7814), .A2(n6942), .ZN(n6815) );
  NAND2_X1 U8506 ( .A1(n6816), .A2(n6815), .ZN(n6818) );
  NAND2_X1 U8507 ( .A1(n6817), .A2(n6818), .ZN(n7614) );
  NAND2_X1 U8508 ( .A1(n7612), .A2(n7614), .ZN(n6821) );
  INV_X1 U8509 ( .A(n6817), .ZN(n6820) );
  INV_X1 U8510 ( .A(n6818), .ZN(n6819) );
  NAND2_X1 U8511 ( .A1(n6820), .A2(n6819), .ZN(n7613) );
  NAND2_X1 U8512 ( .A1(n9819), .A2(n4380), .ZN(n6823) );
  NAND2_X1 U8513 ( .A1(n9485), .A2(n6947), .ZN(n6822) );
  NAND2_X1 U8514 ( .A1(n6823), .A2(n6822), .ZN(n6824) );
  XNOR2_X1 U8515 ( .A(n6824), .B(n6945), .ZN(n6826) );
  AND2_X1 U8516 ( .A1(n6929), .A2(n9485), .ZN(n6825) );
  AOI21_X1 U8517 ( .B1(n9819), .B2(n6947), .A(n6825), .ZN(n6827) );
  XNOR2_X1 U8518 ( .A(n6826), .B(n6827), .ZN(n7787) );
  INV_X1 U8519 ( .A(n6826), .ZN(n6829) );
  INV_X1 U8520 ( .A(n6827), .ZN(n6828) );
  NAND2_X1 U8521 ( .A1(n9816), .A2(n4380), .ZN(n6831) );
  OR2_X1 U8522 ( .A1(n9483), .A2(n6917), .ZN(n6830) );
  NAND2_X1 U8523 ( .A1(n6831), .A2(n6830), .ZN(n6832) );
  XNOR2_X1 U8524 ( .A(n6832), .B(n4387), .ZN(n6834) );
  NOR2_X1 U8525 ( .A1(n9483), .A2(n6942), .ZN(n6833) );
  AOI21_X1 U8526 ( .B1(n9816), .B2(n6947), .A(n6833), .ZN(n6835) );
  XNOR2_X1 U8527 ( .A(n6834), .B(n6835), .ZN(n7996) );
  INV_X1 U8528 ( .A(n6834), .ZN(n6836) );
  NAND2_X1 U8529 ( .A1(n6836), .A2(n6835), .ZN(n6837) );
  AND2_X2 U8530 ( .A1(n7995), .A2(n6837), .ZN(n8087) );
  OAI22_X1 U8531 ( .A1(n9809), .A2(n6908), .B1(n8048), .B2(n6917), .ZN(n6838)
         );
  XNOR2_X1 U8532 ( .A(n6838), .B(n6945), .ZN(n8085) );
  OR2_X1 U8533 ( .A1(n9809), .A2(n6917), .ZN(n6840) );
  OR2_X1 U8534 ( .A1(n8048), .A2(n6942), .ZN(n6839) );
  AND2_X1 U8535 ( .A1(n6840), .A2(n6839), .ZN(n6842) );
  NAND2_X1 U8536 ( .A1(n8085), .A2(n6842), .ZN(n6841) );
  INV_X1 U8537 ( .A(n8085), .ZN(n6843) );
  INV_X1 U8538 ( .A(n6842), .ZN(n8084) );
  NAND2_X1 U8539 ( .A1(n6843), .A2(n8084), .ZN(n6844) );
  OAI22_X1 U8540 ( .A1(n8188), .A2(n6908), .B1(n8189), .B2(n6917), .ZN(n6845)
         );
  XNOR2_X1 U8541 ( .A(n6845), .B(n6945), .ZN(n8179) );
  OR2_X1 U8542 ( .A1(n8188), .A2(n6917), .ZN(n6847) );
  OR2_X1 U8543 ( .A1(n8189), .A2(n6942), .ZN(n6846) );
  AND2_X1 U8544 ( .A1(n6847), .A2(n6846), .ZN(n6849) );
  NAND2_X1 U8545 ( .A1(n8179), .A2(n6849), .ZN(n6854) );
  OAI22_X1 U8546 ( .A1(n8216), .A2(n6908), .B1(n9384), .B2(n6917), .ZN(n6848)
         );
  XNOR2_X1 U8547 ( .A(n6848), .B(n6945), .ZN(n6853) );
  INV_X1 U8548 ( .A(n8179), .ZN(n6850) );
  INV_X1 U8549 ( .A(n6849), .ZN(n8178) );
  NAND2_X1 U8550 ( .A1(n6850), .A2(n8178), .ZN(n6852) );
  AND2_X1 U8551 ( .A1(n6853), .A2(n6852), .ZN(n6851) );
  OAI22_X1 U8552 ( .A1(n8216), .A2(n6917), .B1(n9384), .B2(n6942), .ZN(n9460)
         );
  NAND2_X1 U8553 ( .A1(n9457), .A2(n9460), .ZN(n6858) );
  INV_X1 U8554 ( .A(n6852), .ZN(n6857) );
  INV_X1 U8555 ( .A(n6853), .ZN(n6855) );
  AND2_X1 U8556 ( .A1(n6855), .A2(n6854), .ZN(n6856) );
  OAI21_X2 U8557 ( .B1(n8177), .B2(n6857), .A(n6856), .ZN(n9458) );
  OAI22_X1 U8558 ( .A1(n8228), .A2(n6908), .B1(n9468), .B2(n6917), .ZN(n6859)
         );
  XNOR2_X1 U8559 ( .A(n6859), .B(n4387), .ZN(n6860) );
  OAI22_X1 U8560 ( .A1(n8228), .A2(n6917), .B1(n9468), .B2(n6942), .ZN(n6861)
         );
  AND2_X1 U8561 ( .A1(n6860), .A2(n6861), .ZN(n9380) );
  INV_X1 U8562 ( .A(n6860), .ZN(n6863) );
  INV_X1 U8563 ( .A(n6861), .ZN(n6862) );
  NAND2_X1 U8564 ( .A1(n6863), .A2(n6862), .ZN(n9379) );
  NAND2_X1 U8565 ( .A1(n9790), .A2(n4380), .ZN(n6865) );
  NAND2_X1 U8566 ( .A1(n9716), .A2(n6947), .ZN(n6864) );
  NAND2_X1 U8567 ( .A1(n6865), .A2(n6864), .ZN(n6866) );
  XNOR2_X1 U8568 ( .A(n6866), .B(n4387), .ZN(n6868) );
  AND2_X1 U8569 ( .A1(n9716), .A2(n6929), .ZN(n6867) );
  AOI21_X1 U8570 ( .B1(n9790), .B2(n6947), .A(n6867), .ZN(n6869) );
  XNOR2_X1 U8571 ( .A(n6868), .B(n6869), .ZN(n9391) );
  INV_X1 U8572 ( .A(n6868), .ZN(n6870) );
  NAND2_X1 U8573 ( .A1(n6870), .A2(n6869), .ZN(n6871) );
  NAND2_X1 U8574 ( .A1(n9783), .A2(n4380), .ZN(n6873) );
  NAND2_X1 U8575 ( .A1(n9696), .A2(n6947), .ZN(n6872) );
  NAND2_X1 U8576 ( .A1(n6873), .A2(n6872), .ZN(n6874) );
  XNOR2_X1 U8577 ( .A(n6874), .B(n6945), .ZN(n6877) );
  NAND2_X1 U8578 ( .A1(n9783), .A2(n6947), .ZN(n6876) );
  NAND2_X1 U8579 ( .A1(n9696), .A2(n6929), .ZN(n6875) );
  NAND2_X1 U8580 ( .A1(n6876), .A2(n6875), .ZN(n9429) );
  NAND2_X1 U8581 ( .A1(n9773), .A2(n4380), .ZN(n6880) );
  NAND2_X1 U8582 ( .A1(n9697), .A2(n6758), .ZN(n6879) );
  NAND2_X1 U8583 ( .A1(n6880), .A2(n6879), .ZN(n6881) );
  XNOR2_X1 U8584 ( .A(n6881), .B(n4387), .ZN(n6891) );
  NAND2_X1 U8585 ( .A1(n9773), .A2(n6758), .ZN(n6883) );
  NAND2_X1 U8586 ( .A1(n9697), .A2(n6929), .ZN(n6882) );
  NAND2_X1 U8587 ( .A1(n6883), .A2(n6882), .ZN(n6892) );
  NAND2_X1 U8588 ( .A1(n6891), .A2(n6892), .ZN(n9360) );
  NAND2_X1 U8589 ( .A1(n9778), .A2(n4380), .ZN(n6885) );
  NAND2_X1 U8590 ( .A1(n9717), .A2(n6947), .ZN(n6884) );
  NAND2_X1 U8591 ( .A1(n6885), .A2(n6884), .ZN(n6886) );
  XNOR2_X1 U8592 ( .A(n6886), .B(n6945), .ZN(n9358) );
  INV_X1 U8593 ( .A(n9358), .ZN(n9355) );
  NAND2_X1 U8594 ( .A1(n9778), .A2(n6947), .ZN(n6888) );
  NAND2_X1 U8595 ( .A1(n9717), .A2(n6929), .ZN(n6887) );
  AND2_X1 U8596 ( .A1(n6888), .A2(n6887), .ZN(n6890) );
  INV_X1 U8597 ( .A(n6890), .ZN(n9354) );
  NAND2_X1 U8598 ( .A1(n9355), .A2(n9354), .ZN(n6889) );
  NAND2_X1 U8599 ( .A1(n9360), .A2(n6889), .ZN(n6897) );
  INV_X1 U8600 ( .A(n6891), .ZN(n6894) );
  INV_X1 U8601 ( .A(n6892), .ZN(n6893) );
  NAND2_X1 U8602 ( .A1(n6894), .A2(n6893), .ZN(n9361) );
  NAND2_X1 U8603 ( .A1(n9770), .A2(n4380), .ZN(n6899) );
  OR2_X1 U8604 ( .A1(n9478), .A2(n6917), .ZN(n6898) );
  NAND2_X1 U8605 ( .A1(n6899), .A2(n6898), .ZN(n6900) );
  XNOR2_X1 U8606 ( .A(n6900), .B(n4387), .ZN(n6902) );
  NOR2_X1 U8607 ( .A1(n9478), .A2(n6942), .ZN(n6901) );
  AOI21_X1 U8608 ( .B1(n9770), .B2(n6947), .A(n6901), .ZN(n6903) );
  XNOR2_X1 U8609 ( .A(n6902), .B(n6903), .ZN(n9362) );
  INV_X1 U8610 ( .A(n6902), .ZN(n6904) );
  NAND2_X1 U8611 ( .A1(n6904), .A2(n6903), .ZN(n6905) );
  OR2_X1 U8612 ( .A1(n9654), .A2(n6917), .ZN(n6907) );
  OR2_X1 U8613 ( .A1(n9667), .A2(n6942), .ZN(n6906) );
  OAI22_X1 U8614 ( .A1(n9654), .A2(n6908), .B1(n9667), .B2(n6917), .ZN(n6909)
         );
  XNOR2_X1 U8615 ( .A(n6909), .B(n4387), .ZN(n9421) );
  NAND2_X1 U8616 ( .A1(n9758), .A2(n4380), .ZN(n6911) );
  NAND2_X1 U8617 ( .A1(n9657), .A2(n6947), .ZN(n6910) );
  NAND2_X1 U8618 ( .A1(n6911), .A2(n6910), .ZN(n6912) );
  XNOR2_X1 U8619 ( .A(n6912), .B(n6945), .ZN(n9337) );
  NAND2_X1 U8620 ( .A1(n9750), .A2(n4380), .ZN(n6919) );
  OR2_X1 U8621 ( .A1(n9625), .A2(n6917), .ZN(n6918) );
  NAND2_X1 U8622 ( .A1(n6919), .A2(n6918), .ZN(n6920) );
  XNOR2_X1 U8623 ( .A(n6920), .B(n6945), .ZN(n6925) );
  NOR2_X1 U8624 ( .A1(n9625), .A2(n6942), .ZN(n6921) );
  AOI21_X1 U8625 ( .B1(n9750), .B2(n6947), .A(n6921), .ZN(n6924) );
  AND2_X1 U8626 ( .A1(n6925), .A2(n6924), .ZN(n9445) );
  NAND2_X1 U8627 ( .A1(n9743), .A2(n4380), .ZN(n6927) );
  NAND2_X1 U8628 ( .A1(n9474), .A2(n6947), .ZN(n6926) );
  NAND2_X1 U8629 ( .A1(n6927), .A2(n6926), .ZN(n6928) );
  XNOR2_X1 U8630 ( .A(n6928), .B(n6945), .ZN(n6937) );
  AND2_X1 U8631 ( .A1(n6929), .A2(n9474), .ZN(n6930) );
  AOI21_X1 U8632 ( .B1(n9743), .B2(n6947), .A(n6930), .ZN(n6938) );
  XNOR2_X1 U8633 ( .A(n6937), .B(n6938), .ZN(n9444) );
  NAND2_X1 U8634 ( .A1(n9739), .A2(n4380), .ZN(n6932) );
  OR2_X1 U8635 ( .A1(n9602), .A2(n6917), .ZN(n6931) );
  NAND2_X1 U8636 ( .A1(n6932), .A2(n6931), .ZN(n6933) );
  XNOR2_X1 U8637 ( .A(n6933), .B(n6945), .ZN(n6936) );
  NOR2_X1 U8638 ( .A1(n9602), .A2(n6942), .ZN(n6934) );
  AOI21_X1 U8639 ( .B1(n9739), .B2(n6947), .A(n6934), .ZN(n6935) );
  NAND2_X1 U8640 ( .A1(n6936), .A2(n6935), .ZN(n6968) );
  OAI21_X1 U8641 ( .B1(n6936), .B2(n6935), .A(n6968), .ZN(n9326) );
  INV_X1 U8642 ( .A(n6937), .ZN(n6940) );
  INV_X1 U8643 ( .A(n6938), .ZN(n6939) );
  NOR2_X2 U8644 ( .A1(n9443), .A2(n6941), .ZN(n9330) );
  NAND2_X1 U8645 ( .A1(n9570), .A2(n6758), .ZN(n6944) );
  OR2_X1 U8646 ( .A1(n9582), .A2(n6942), .ZN(n6943) );
  NAND2_X1 U8647 ( .A1(n6944), .A2(n6943), .ZN(n6946) );
  XNOR2_X1 U8648 ( .A(n6946), .B(n6945), .ZN(n6949) );
  INV_X1 U8649 ( .A(n9582), .ZN(n9553) );
  AOI22_X1 U8650 ( .A1(n9570), .A2(n4380), .B1(n6947), .B2(n9553), .ZN(n6948)
         );
  XNOR2_X1 U8651 ( .A(n6949), .B(n6948), .ZN(n6966) );
  INV_X1 U8652 ( .A(n6966), .ZN(n6970) );
  NAND3_X1 U8653 ( .A1(n8163), .A2(P1_B_REG_SCAN_IN), .A3(n8223), .ZN(n6950)
         );
  INV_X1 U8654 ( .A(n7188), .ZN(n6953) );
  INV_X1 U8655 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6952) );
  INV_X1 U8656 ( .A(n6951), .ZN(n9857) );
  AND2_X1 U8657 ( .A1(n7199), .A2(n7040), .ZN(n6982) );
  NOR4_X1 U8658 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6957) );
  NOR4_X1 U8659 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6956) );
  NOR4_X1 U8660 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6955) );
  NOR4_X1 U8661 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n6954) );
  NAND4_X1 U8662 ( .A1(n6957), .A2(n6956), .A3(n6955), .A4(n6954), .ZN(n6962)
         );
  NOR2_X1 U8663 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .ZN(
        n9055) );
  NOR4_X1 U8664 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6960) );
  NOR4_X1 U8665 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6959) );
  NOR4_X1 U8666 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6958) );
  NAND4_X1 U8667 ( .A1(n9055), .A2(n6960), .A3(n6959), .A4(n6958), .ZN(n6961)
         );
  NOR2_X1 U8668 ( .A1(n6962), .A2(n6961), .ZN(n7189) );
  AND2_X1 U8669 ( .A1(n7189), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6963) );
  NAND2_X1 U8670 ( .A1(n9857), .A2(n8223), .ZN(n7186) );
  OAI21_X1 U8671 ( .B1(n7188), .B2(n6963), .A(n7186), .ZN(n7015) );
  INV_X1 U8672 ( .A(n7010), .ZN(n7011) );
  OR2_X1 U8673 ( .A1(n7015), .A2(n7011), .ZN(n6964) );
  NOR2_X1 U8674 ( .A1(n10106), .A2(n6964), .ZN(n6965) );
  NAND3_X1 U8675 ( .A1(n6966), .A2(n9448), .A3(n6968), .ZN(n6967) );
  NOR2_X1 U8676 ( .A1(n9330), .A2(n6967), .ZN(n6994) );
  INV_X1 U8677 ( .A(n6968), .ZN(n6969) );
  NAND3_X1 U8678 ( .A1(n6970), .A2(n9448), .A3(n6969), .ZN(n6993) );
  NOR2_X1 U8679 ( .A1(n9824), .A2(n5868), .ZN(n6973) );
  INV_X1 U8680 ( .A(n7191), .ZN(n6974) );
  INV_X1 U8681 ( .A(n7015), .ZN(n6981) );
  NAND2_X1 U8682 ( .A1(n6981), .A2(n7199), .ZN(n6985) );
  NAND2_X1 U8683 ( .A1(n6974), .A2(n6985), .ZN(n6980) );
  INV_X1 U8684 ( .A(n7016), .ZN(n6975) );
  NAND2_X1 U8685 ( .A1(n6977), .A2(n6976), .ZN(n6978) );
  NAND2_X1 U8686 ( .A1(n6978), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6979) );
  NAND3_X1 U8687 ( .A1(n6981), .A2(n7193), .A3(n9926), .ZN(n6984) );
  INV_X1 U8688 ( .A(n6982), .ZN(n6983) );
  NOR2_X1 U8689 ( .A1(n9467), .A2(n8313), .ZN(n6989) );
  OAI22_X1 U8690 ( .A1(n9451), .A2(n9602), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6987), .ZN(n6988) );
  AOI211_X1 U8691 ( .C1(n9569), .C2(n9462), .A(n6989), .B(n6988), .ZN(n6990)
         );
  NOR2_X1 U8692 ( .A1(n6994), .A2(n5027), .ZN(n6995) );
  NAND2_X1 U8693 ( .A1(n6996), .A2(n6995), .ZN(P1_U3218) );
  NAND2_X1 U8694 ( .A1(n7010), .A2(n7001), .ZN(n6997) );
  NAND2_X1 U8695 ( .A1(n6997), .A2(n6999), .ZN(n9496) );
  NAND2_X1 U8696 ( .A1(n9496), .A2(n9493), .ZN(n6998) );
  NAND2_X1 U8697 ( .A1(n6998), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8698 ( .A(n6999), .ZN(n7000) );
  NAND2_X1 U8699 ( .A1(n5869), .A2(n10011), .ZN(n7003) );
  XNOR2_X1 U8700 ( .A(n7637), .B(n7552), .ZN(n7014) );
  NAND2_X1 U8701 ( .A1(n7650), .A2(n7652), .ZN(n7651) );
  NAND2_X1 U8702 ( .A1(n5818), .A2(n4997), .ZN(n7004) );
  NAND2_X1 U8703 ( .A1(n7651), .A2(n7004), .ZN(n7559) );
  AND2_X1 U8704 ( .A1(n7559), .A2(n7636), .ZN(n7005) );
  NOR2_X1 U8705 ( .A1(n7559), .A2(n7636), .ZN(n7631) );
  OR2_X1 U8706 ( .A1(n7005), .A2(n7631), .ZN(n10073) );
  OR2_X1 U8707 ( .A1(n7006), .A2(n7017), .ZN(n7009) );
  OR2_X1 U8708 ( .A1(n7007), .A2(n7913), .ZN(n7008) );
  NAND2_X1 U8709 ( .A1(n10073), .A2(n10034), .ZN(n7013) );
  AOI22_X1 U8710 ( .A1(n7554), .A2(n10037), .B1(n9715), .B2(n5818), .ZN(n7012)
         );
  OAI211_X1 U8711 ( .C1(n10014), .C2(n7014), .A(n7013), .B(n7012), .ZN(n10071)
         );
  MUX2_X1 U8712 ( .A(n10071), .B(P1_REG2_REG_2__SCAN_IN), .S(n10047), .Z(n7028) );
  AND2_X1 U8713 ( .A1(n7017), .A2(n10011), .ZN(n7018) );
  NAND2_X1 U8714 ( .A1(n10033), .A2(n7018), .ZN(n8218) );
  INV_X1 U8715 ( .A(n8218), .ZN(n10029) );
  NAND2_X1 U8716 ( .A1(n10073), .A2(n10029), .ZN(n7026) );
  NOR2_X1 U8717 ( .A1(n7574), .A2(n7910), .ZN(n10007) );
  INV_X1 U8718 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7020) );
  OAI22_X1 U8719 ( .A1(n9710), .A2(n10069), .B1(n10031), .B2(n7020), .ZN(n7024) );
  NOR2_X1 U8720 ( .A1(n7574), .A2(n7021), .ZN(n7022) );
  NAND2_X1 U8721 ( .A1(n10033), .A2(n7022), .ZN(n9573) );
  OAI21_X1 U8722 ( .B1(n7659), .B2(n10069), .A(n7643), .ZN(n10070) );
  NOR2_X1 U8723 ( .A1(n9573), .A2(n10070), .ZN(n7023) );
  NOR2_X1 U8724 ( .A1(n7024), .A2(n7023), .ZN(n7025) );
  NAND2_X1 U8725 ( .A1(n7026), .A2(n7025), .ZN(n7027) );
  OR2_X1 U8726 ( .A1(n7028), .A2(n7027), .ZN(P1_U3289) );
  INV_X1 U8727 ( .A(n7304), .ZN(n7399) );
  AND2_X1 U8728 ( .A1(n4518), .A2(P2_U3152), .ZN(n9321) );
  NOR2_X1 U8729 ( .A1(n4518), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9320) );
  INV_X2 U8730 ( .A(n9320), .ZN(n9043) );
  OAI222_X1 U8731 ( .A1(n7399), .A2(P2_U3152), .B1(n9036), .B2(n7046), .C1(
        n5325), .C2(n9043), .ZN(P2_U3356) );
  INV_X1 U8732 ( .A(n7029), .ZN(n7050) );
  INV_X1 U8733 ( .A(n7321), .ZN(n7335) );
  OAI222_X1 U8734 ( .A1(n9043), .A2(n5080), .B1(n9036), .B2(n7050), .C1(
        P2_U3152), .C2(n7335), .ZN(P2_U3354) );
  INV_X2 U8735 ( .A(n9321), .ZN(n9036) );
  INV_X1 U8736 ( .A(n7030), .ZN(n7035) );
  OAI222_X1 U8737 ( .A1(n9043), .A2(n7031), .B1(n9036), .B2(n7035), .C1(
        P2_U3152), .C2(n7385), .ZN(P2_U3355) );
  OAI222_X1 U8738 ( .A1(n8538), .A2(P2_U3152), .B1(n9036), .B2(n7056), .C1(
        n5307), .C2(n9043), .ZN(P2_U3357) );
  INV_X1 U8739 ( .A(n7115), .ZN(n7034) );
  OAI222_X1 U8740 ( .A1(n8332), .A2(n5061), .B1(n7914), .B2(n7035), .C1(
        P1_U3084), .C2(n7034), .ZN(P1_U3350) );
  INV_X1 U8741 ( .A(n7036), .ZN(n7053) );
  INV_X1 U8742 ( .A(n7336), .ZN(n7351) );
  OAI222_X1 U8743 ( .A1(n9043), .A2(n5085), .B1(n9036), .B2(n7053), .C1(
        P2_U3152), .C2(n7351), .ZN(P2_U3353) );
  INV_X1 U8744 ( .A(n7037), .ZN(n7051) );
  INV_X1 U8745 ( .A(n7360), .ZN(n7320) );
  OAI222_X1 U8746 ( .A1(n9043), .A2(n5087), .B1(n9036), .B2(n7051), .C1(
        P2_U3152), .C2(n7320), .ZN(P2_U3352) );
  INV_X1 U8747 ( .A(n7038), .ZN(n7048) );
  INV_X1 U8748 ( .A(n7409), .ZN(n7371) );
  OAI222_X1 U8749 ( .A1(n9043), .A2(n5096), .B1(n9036), .B2(n7048), .C1(
        P2_U3152), .C2(n7371), .ZN(P2_U3351) );
  INV_X1 U8750 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n7041) );
  INV_X1 U8751 ( .A(n7186), .ZN(n7039) );
  AOI22_X1 U8752 ( .A1(n10062), .A2(n7041), .B1(n7040), .B2(n7039), .ZN(
        P1_U3441) );
  NAND2_X1 U8753 ( .A1(n10062), .A2(P1_D_REG_0__SCAN_IN), .ZN(n7042) );
  OAI21_X1 U8754 ( .B1(n10062), .B2(n7043), .A(n7042), .ZN(P1_U3440) );
  INV_X1 U8755 ( .A(n7044), .ZN(n7045) );
  OAI222_X1 U8756 ( .A1(n8332), .A2(n9049), .B1(n7914), .B2(n7045), .C1(
        P1_U3084), .C2(n7176), .ZN(P1_U3345) );
  OAI222_X1 U8757 ( .A1(n9043), .A2(n9052), .B1(n9036), .B2(n7045), .C1(
        P2_U3152), .C2(n8556), .ZN(P2_U3350) );
  INV_X1 U8758 ( .A(n9910), .ZN(n7047) );
  OAI222_X1 U8759 ( .A1(n7047), .A2(P1_U3084), .B1(n7914), .B2(n7046), .C1(
        n9048), .C2(n8332), .ZN(P1_U3351) );
  INV_X1 U8760 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7049) );
  INV_X1 U8761 ( .A(n7138), .ZN(n7144) );
  OAI222_X1 U8762 ( .A1(n8332), .A2(n7049), .B1(n7914), .B2(n7048), .C1(
        P1_U3084), .C2(n7144), .ZN(P1_U3346) );
  OAI222_X1 U8763 ( .A1(n8332), .A2(n5078), .B1(n7914), .B2(n7050), .C1(
        P1_U3084), .C2(n9935), .ZN(P1_U3349) );
  INV_X1 U8764 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7052) );
  INV_X1 U8765 ( .A(n7130), .ZN(n7095) );
  OAI222_X1 U8766 ( .A1(n8332), .A2(n7052), .B1(n7914), .B2(n7051), .C1(
        P1_U3084), .C2(n7095), .ZN(P1_U3347) );
  INV_X1 U8767 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7054) );
  INV_X1 U8768 ( .A(n7101), .ZN(n7092) );
  OAI222_X1 U8769 ( .A1(n8332), .A2(n7054), .B1(n7914), .B2(n7053), .C1(
        P1_U3084), .C2(n7092), .ZN(P1_U3348) );
  INV_X1 U8770 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7055) );
  OAI222_X1 U8771 ( .A1(n7079), .A2(P1_U3084), .B1(n7914), .B2(n7056), .C1(
        n7055), .C2(n8332), .ZN(P1_U3352) );
  INV_X1 U8772 ( .A(n9322), .ZN(n7057) );
  INV_X1 U8773 ( .A(n7232), .ZN(n7227) );
  OAI222_X1 U8774 ( .A1(n8332), .A2(n9046), .B1(n7914), .B2(n7057), .C1(n7227), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U8775 ( .A(n7058), .ZN(n7064) );
  AOI22_X1 U8776 ( .A1(n8587), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n9320), .ZN(n7059) );
  OAI21_X1 U8777 ( .B1(n7064), .B2(n9036), .A(n7059), .ZN(P2_U3348) );
  INV_X1 U8778 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7061) );
  NAND2_X1 U8779 ( .A1(n8623), .A2(P2_U3966), .ZN(n7060) );
  OAI21_X1 U8780 ( .B1(n7061), .B2(P2_U3966), .A(n7060), .ZN(P2_U3583) );
  INV_X1 U8781 ( .A(n7062), .ZN(n7063) );
  OAI222_X1 U8782 ( .A1(n8332), .A2(n9107), .B1(n7914), .B2(n7063), .C1(n7268), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U8783 ( .A(n7418), .ZN(n7454) );
  OAI222_X1 U8784 ( .A1(P2_U3152), .A2(n7454), .B1(n9036), .B2(n7063), .C1(
        n9060), .C2(n9043), .ZN(P2_U3347) );
  INV_X1 U8785 ( .A(n7267), .ZN(n7264) );
  OAI222_X1 U8786 ( .A1(n8332), .A2(n7065), .B1(n7914), .B2(n7064), .C1(n7264), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U8787 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7090) );
  NOR2_X1 U8788 ( .A1(n9920), .A2(P1_U3084), .ZN(n9851) );
  NAND2_X1 U8789 ( .A1(n9496), .A2(n9851), .ZN(n8263) );
  INV_X1 U8790 ( .A(n8263), .ZN(n7085) );
  NAND2_X1 U8791 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3084), .ZN(n7589) );
  INV_X1 U8792 ( .A(n7589), .ZN(n7076) );
  INV_X1 U8793 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7070) );
  INV_X1 U8794 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10132) );
  MUX2_X1 U8795 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10132), .S(n9910), .Z(n9914)
         );
  INV_X1 U8796 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10130) );
  MUX2_X1 U8797 ( .A(n10130), .B(P1_REG1_REG_1__SCAN_IN), .S(n7079), .Z(n9894)
         );
  AND2_X1 U8798 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9893) );
  NAND2_X1 U8799 ( .A1(n9894), .A2(n9893), .ZN(n9892) );
  NAND2_X1 U8800 ( .A1(n9891), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7067) );
  NAND2_X1 U8801 ( .A1(n9892), .A2(n7067), .ZN(n9913) );
  NAND2_X1 U8802 ( .A1(n9914), .A2(n9913), .ZN(n9912) );
  NAND2_X1 U8803 ( .A1(n9910), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7068) );
  NAND2_X1 U8804 ( .A1(n9912), .A2(n7068), .ZN(n7110) );
  INV_X1 U8805 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7069) );
  XNOR2_X1 U8806 ( .A(n7115), .B(n7069), .ZN(n7111) );
  XNOR2_X1 U8807 ( .A(n9935), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9936) );
  NAND2_X1 U8808 ( .A1(n7115), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9937) );
  XOR2_X1 U8809 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7101), .Z(n7072) );
  NOR2_X1 U8810 ( .A1(n9926), .A2(P1_U3084), .ZN(n9848) );
  AND2_X1 U8811 ( .A1(n9848), .A2(n9920), .ZN(n7071) );
  OAI211_X1 U8812 ( .C1(n7073), .C2(n7072), .A(n7091), .B(n9962), .ZN(n7074)
         );
  INV_X1 U8813 ( .A(n7074), .ZN(n7075) );
  AOI211_X1 U8814 ( .C1(n9957), .C2(n7101), .A(n7076), .B(n7075), .ZN(n7089)
         );
  INV_X1 U8815 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9904) );
  INV_X1 U8816 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7077) );
  AND2_X1 U8817 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9919) );
  NAND2_X1 U8818 ( .A1(n9891), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9905) );
  NAND2_X1 U8819 ( .A1(n9910), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7117) );
  INV_X1 U8820 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7642) );
  MUX2_X1 U8821 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n7642), .S(n7115), .Z(n7080)
         );
  NAND2_X1 U8822 ( .A1(n7115), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7082) );
  AND2_X1 U8823 ( .A1(n7119), .A2(n7082), .ZN(n9931) );
  MUX2_X1 U8824 ( .A(n5353), .B(P1_REG2_REG_4__SCAN_IN), .S(n9935), .Z(n9930)
         );
  AND2_X1 U8825 ( .A1(n9935), .A2(n5353), .ZN(n7083) );
  INV_X1 U8826 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10022) );
  MUX2_X1 U8827 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10022), .S(n7101), .Z(n7084)
         );
  INV_X1 U8828 ( .A(n7100), .ZN(n7087) );
  NOR3_X1 U8829 ( .A1(n9934), .A2(n7084), .A3(n7083), .ZN(n7086) );
  OAI21_X1 U8830 ( .B1(n7087), .B2(n7086), .A(n9932), .ZN(n7088) );
  OAI211_X1 U8831 ( .C1(n7090), .C2(n9947), .A(n7089), .B(n7088), .ZN(P1_U3246) );
  INV_X1 U8832 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7094) );
  INV_X1 U8833 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7093) );
  OAI21_X1 U8834 ( .B1(n7093), .B2(n7092), .A(n7091), .ZN(n7124) );
  MUX2_X1 U8835 ( .A(n7094), .B(P1_REG1_REG_6__SCAN_IN), .S(n7130), .Z(n7125)
         );
  NOR2_X1 U8836 ( .A1(n7124), .A2(n7125), .ZN(n7123) );
  XNOR2_X1 U8837 ( .A(n7138), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n7096) );
  AOI21_X1 U8838 ( .B1(n7097), .B2(n7096), .A(n7143), .ZN(n7109) );
  NAND2_X1 U8839 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3084), .ZN(n7243) );
  INV_X1 U8840 ( .A(n7243), .ZN(n7099) );
  NOR2_X1 U8841 ( .A1(n9947), .A2(n4527), .ZN(n7098) );
  AOI211_X1 U8842 ( .C1(n9957), .C2(n7138), .A(n7099), .B(n7098), .ZN(n7108)
         );
  INV_X1 U8843 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7102) );
  MUX2_X1 U8844 ( .A(n7102), .B(P1_REG2_REG_6__SCAN_IN), .S(n7130), .Z(n7127)
         );
  INV_X1 U8845 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7103) );
  MUX2_X1 U8846 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7103), .S(n7138), .Z(n7104)
         );
  OAI21_X1 U8847 ( .B1(n7105), .B2(n7104), .A(n7140), .ZN(n7106) );
  NAND2_X1 U8848 ( .A1(n7106), .A2(n9932), .ZN(n7107) );
  OAI211_X1 U8849 ( .C1(n7109), .C2(n9533), .A(n7108), .B(n7107), .ZN(P1_U3248) );
  INV_X1 U8850 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7122) );
  OAI211_X1 U8851 ( .C1(n7111), .C2(n7110), .A(n9962), .B(n9938), .ZN(n7113)
         );
  NAND2_X1 U8852 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7112) );
  NAND2_X1 U8853 ( .A1(n7113), .A2(n7112), .ZN(n7114) );
  AOI21_X1 U8854 ( .B1(n7115), .B2(n9957), .A(n7114), .ZN(n7121) );
  MUX2_X1 U8855 ( .A(n7642), .B(P1_REG2_REG_3__SCAN_IN), .S(n7115), .Z(n7116)
         );
  NAND3_X1 U8856 ( .A1(n9909), .A2(n7117), .A3(n7116), .ZN(n7118) );
  NAND3_X1 U8857 ( .A1(n9932), .A2(n7119), .A3(n7118), .ZN(n7120) );
  OAI211_X1 U8858 ( .C1(n7122), .C2(n9947), .A(n7121), .B(n7120), .ZN(P1_U3244) );
  AOI21_X1 U8859 ( .B1(n7125), .B2(n7124), .A(n7123), .ZN(n7133) );
  AOI211_X1 U8860 ( .C1(n7128), .C2(n7127), .A(n9950), .B(n7126), .ZN(n7129)
         );
  AOI21_X1 U8861 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n9961), .A(n7129), .ZN(
        n7132) );
  AND2_X1 U8862 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7727) );
  AOI21_X1 U8863 ( .B1(n9957), .B2(n7130), .A(n7727), .ZN(n7131) );
  OAI211_X1 U8864 ( .C1(n7133), .C2(n9533), .A(n7132), .B(n7131), .ZN(P1_U3247) );
  NAND2_X1 U8865 ( .A1(n10175), .A2(n8055), .ZN(n7135) );
  NAND2_X1 U8866 ( .A1(n7135), .A2(n7134), .ZN(n7137) );
  OR2_X1 U8867 ( .A1(n10175), .A2(n7279), .ZN(n7136) );
  NOR2_X1 U8868 ( .A1(n10164), .A2(P2_U3966), .ZN(P2_U3151) );
  XNOR2_X1 U8869 ( .A(n7177), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n7141) );
  NAND2_X1 U8870 ( .A1(n7141), .A2(n9492), .ZN(n7142) );
  XNOR2_X1 U8871 ( .A(n7142), .B(n7176), .ZN(n7151) );
  INV_X1 U8872 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7145) );
  XNOR2_X1 U8873 ( .A(n7176), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n7146) );
  OAI211_X1 U8874 ( .C1(n7147), .C2(n7146), .A(n7171), .B(n9962), .ZN(n7150)
         );
  NAND2_X1 U8875 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3084), .ZN(n7430) );
  INV_X1 U8876 ( .A(n7430), .ZN(n7148) );
  AOI21_X1 U8877 ( .B1(n9961), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n7148), .ZN(
        n7149) );
  OAI211_X1 U8878 ( .C1(n7151), .C2(n8263), .A(n7150), .B(n7149), .ZN(P1_U3249) );
  INV_X1 U8879 ( .A(n7152), .ZN(n7154) );
  INV_X1 U8880 ( .A(n7463), .ZN(n7473) );
  OAI222_X1 U8881 ( .A1(n9043), .A2(n7153), .B1(n9036), .B2(n7154), .C1(
        P2_U3152), .C2(n7473), .ZN(P2_U3346) );
  INV_X1 U8882 ( .A(n7866), .ZN(n7861) );
  OAI222_X1 U8883 ( .A1(n8332), .A2(n7155), .B1(n7914), .B2(n7154), .C1(
        P1_U3084), .C2(n7861), .ZN(P1_U3341) );
  NAND2_X1 U8884 ( .A1(n8322), .A2(P1_U4006), .ZN(n7156) );
  OAI21_X1 U8885 ( .B1(P1_U4006), .B2(n6405), .A(n7156), .ZN(P1_U3586) );
  INV_X1 U8886 ( .A(n7486), .ZN(n7159) );
  INV_X1 U8887 ( .A(n7157), .ZN(n7161) );
  OAI222_X1 U8888 ( .A1(P2_U3152), .A2(n7159), .B1(n9036), .B2(n7161), .C1(
        n7158), .C2(n9043), .ZN(P2_U3345) );
  INV_X1 U8889 ( .A(n8167), .ZN(n7160) );
  OAI222_X1 U8890 ( .A1(n8332), .A2(n9300), .B1(n7914), .B2(n7161), .C1(n7160), 
        .C2(P1_U3084), .ZN(P1_U3340) );
  INV_X1 U8891 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n7163) );
  NAND2_X1 U8892 ( .A1(n7217), .A2(P1_U4006), .ZN(n7162) );
  OAI21_X1 U8893 ( .B1(P1_U4006), .B2(n7163), .A(n7162), .ZN(P1_U3555) );
  INV_X1 U8894 ( .A(n7164), .ZN(n7185) );
  AOI22_X1 U8895 ( .A1(n7762), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n9320), .ZN(n7165) );
  OAI21_X1 U8896 ( .B1(n7185), .B2(n9036), .A(n7165), .ZN(P2_U3344) );
  OAI21_X1 U8897 ( .B1(n7168), .B2(n7167), .A(n7166), .ZN(n9921) );
  INV_X1 U8898 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7623) );
  OAI22_X1 U8899 ( .A1(n7731), .A2(n7623), .B1(n5313), .B2(n9467), .ZN(n7169)
         );
  AOI21_X1 U8900 ( .B1(n9448), .B2(n9921), .A(n7169), .ZN(n7170) );
  OAI21_X1 U8901 ( .B1(n4966), .B2(n9456), .A(n7170), .ZN(P1_U3230) );
  XNOR2_X1 U8902 ( .A(n7232), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n7173) );
  OAI21_X1 U8903 ( .B1(n10139), .B2(n7176), .A(n7171), .ZN(n7172) );
  NOR2_X1 U8904 ( .A1(n7172), .A2(n7173), .ZN(n7225) );
  AOI21_X1 U8905 ( .B1(n7173), .B2(n7172), .A(n7225), .ZN(n7184) );
  NAND2_X1 U8906 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3084), .ZN(n7606) );
  INV_X1 U8907 ( .A(n7606), .ZN(n7174) );
  AOI21_X1 U8908 ( .B1(n9957), .B2(n7232), .A(n7174), .ZN(n7175) );
  INV_X1 U8909 ( .A(n7175), .ZN(n7182) );
  XNOR2_X1 U8910 ( .A(n7232), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n7180) );
  INV_X1 U8911 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9210) );
  AOI211_X1 U8912 ( .C1(n7180), .C2(n7179), .A(n9950), .B(n4471), .ZN(n7181)
         );
  AOI211_X1 U8913 ( .C1(n9961), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7182), .B(
        n7181), .ZN(n7183) );
  OAI21_X1 U8914 ( .B1(n7184), .B2(n9533), .A(n7183), .ZN(P1_U3250) );
  INV_X1 U8915 ( .A(n8256), .ZN(n8172) );
  OAI222_X1 U8916 ( .A1(n8332), .A2(n9137), .B1(n7914), .B2(n7185), .C1(n8172), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  OAI21_X1 U8917 ( .B1(n7188), .B2(P1_D_REG_1__SCAN_IN), .A(n7186), .ZN(n7187)
         );
  OAI21_X1 U8918 ( .B1(n7189), .B2(n7188), .A(n7187), .ZN(n7190) );
  INV_X1 U8919 ( .A(n7199), .ZN(n7192) );
  INV_X1 U8920 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7198) );
  INV_X1 U8921 ( .A(n7574), .ZN(n7194) );
  NOR3_X1 U8922 ( .A1(n7195), .A2(n7194), .A3(n7193), .ZN(n7196) );
  AOI21_X1 U8923 ( .B1(n10037), .B2(n5818), .A(n7196), .ZN(n7629) );
  OAI21_X1 U8924 ( .B1(n4966), .B2(n7574), .A(n7629), .ZN(n7201) );
  NAND2_X1 U8925 ( .A1(n7201), .A2(n10129), .ZN(n7197) );
  OAI21_X1 U8926 ( .B1(n10129), .B2(n7198), .A(n7197), .ZN(P1_U3454) );
  NAND2_X1 U8927 ( .A1(n7201), .A2(n10143), .ZN(n7202) );
  OAI21_X1 U8928 ( .B1(n10143), .B2(n6730), .A(n7202), .ZN(P1_U3523) );
  XNOR2_X1 U8929 ( .A(n7204), .B(n7203), .ZN(n7207) );
  NAND2_X1 U8930 ( .A1(n7206), .A2(n7207), .ZN(n7581) );
  OAI21_X1 U8931 ( .B1(n7207), .B2(n7206), .A(n7581), .ZN(n7211) );
  AOI22_X1 U8932 ( .A1(n9464), .A2(n9490), .B1(n9440), .B2(n5364), .ZN(n7209)
         );
  MUX2_X1 U8933 ( .A(n9437), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n7208) );
  OAI211_X1 U8934 ( .C1(n9456), .C2(n10076), .A(n7209), .B(n7208), .ZN(n7210)
         );
  AOI21_X1 U8935 ( .B1(n7211), .B2(n9448), .A(n7210), .ZN(n7212) );
  INV_X1 U8936 ( .A(n7212), .ZN(P1_U3216) );
  NAND2_X1 U8937 ( .A1(n7214), .A2(n7213), .ZN(n7216) );
  XNOR2_X1 U8938 ( .A(n7216), .B(n7215), .ZN(n7221) );
  INV_X1 U8939 ( .A(n7731), .ZN(n8338) );
  INV_X1 U8940 ( .A(n7217), .ZN(n7654) );
  OAI22_X1 U8941 ( .A1(n7654), .A2(n9451), .B1(n9467), .B2(n7655), .ZN(n7219)
         );
  NOR2_X1 U8942 ( .A1(n9456), .A2(n5819), .ZN(n7218) );
  AOI211_X1 U8943 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n8338), .A(n7219), .B(
        n7218), .ZN(n7220) );
  OAI21_X1 U8944 ( .B1(n7221), .B2(n9472), .A(n7220), .ZN(P1_U3220) );
  INV_X1 U8945 ( .A(n7222), .ZN(n7223) );
  OAI222_X1 U8946 ( .A1(n8332), .A2(n9159), .B1(n7914), .B2(n7223), .C1(
        P1_U3084), .C2(n9505), .ZN(P1_U3338) );
  INV_X1 U8947 ( .A(n7783), .ZN(n7758) );
  OAI222_X1 U8948 ( .A1(n9043), .A2(n7224), .B1(n9036), .B2(n7223), .C1(
        P2_U3152), .C2(n7758), .ZN(P2_U3343) );
  INV_X1 U8949 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7226) );
  AOI21_X1 U8950 ( .B1(n7227), .B2(n7226), .A(n7225), .ZN(n7229) );
  XNOR2_X1 U8951 ( .A(n7267), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n7228) );
  NOR2_X1 U8952 ( .A1(n7229), .A2(n7228), .ZN(n7263) );
  AOI21_X1 U8953 ( .B1(n7229), .B2(n7228), .A(n7263), .ZN(n7238) );
  NAND2_X1 U8954 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3084), .ZN(n7617) );
  INV_X1 U8955 ( .A(n7617), .ZN(n7230) );
  AOI21_X1 U8956 ( .B1(n9957), .B2(n7267), .A(n7230), .ZN(n7231) );
  INV_X1 U8957 ( .A(n7231), .ZN(n7236) );
  XNOR2_X1 U8958 ( .A(n7267), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7233) );
  AOI211_X1 U8959 ( .C1(n7234), .C2(n7233), .A(n9950), .B(n7266), .ZN(n7235)
         );
  AOI211_X1 U8960 ( .C1(n9961), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n7236), .B(
        n7235), .ZN(n7237) );
  OAI21_X1 U8961 ( .B1(n7238), .B2(n9533), .A(n7237), .ZN(P1_U3251) );
  XOR2_X1 U8962 ( .A(n7240), .B(n7239), .Z(n7241) );
  XNOR2_X1 U8963 ( .A(n7242), .B(n7241), .ZN(n7248) );
  INV_X1 U8964 ( .A(n7739), .ZN(n9488) );
  OAI21_X1 U8965 ( .B1(n9451), .B2(n10017), .A(n7243), .ZN(n7244) );
  AOI21_X1 U8966 ( .B1(n9440), .B2(n9488), .A(n7244), .ZN(n7245) );
  OAI21_X1 U8967 ( .B1(n9437), .B2(n7576), .A(n7245), .ZN(n7246) );
  AOI21_X1 U8968 ( .B1(n9470), .B2(n10105), .A(n7246), .ZN(n7247) );
  OAI21_X1 U8969 ( .B1(n7248), .B2(n9472), .A(n7247), .ZN(P1_U3211) );
  XOR2_X1 U8970 ( .A(n7250), .B(n7249), .Z(n7511) );
  INV_X1 U8971 ( .A(n7251), .ZN(n7510) );
  NAND2_X1 U8972 ( .A1(n7511), .A2(n7510), .ZN(n7509) );
  NAND2_X1 U8973 ( .A1(n7509), .A2(n7252), .ZN(n7256) );
  NAND2_X1 U8974 ( .A1(n7254), .A2(n7253), .ZN(n7255) );
  XNOR2_X1 U8975 ( .A(n7256), .B(n7255), .ZN(n7262) );
  INV_X1 U8976 ( .A(n10148), .ZN(n7260) );
  NAND3_X1 U8977 ( .A1(n7257), .A2(n8904), .A3(n8902), .ZN(n7537) );
  AOI22_X1 U8978 ( .A1(n10151), .A2(n10201), .B1(n7537), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7258) );
  OAI21_X1 U8979 ( .B1(n10145), .B2(n7957), .A(n7258), .ZN(n7259) );
  AOI21_X1 U8980 ( .B1(n7260), .B2(n4377), .A(n7259), .ZN(n7261) );
  OAI21_X1 U8981 ( .B1(n8519), .B2(n7262), .A(n7261), .ZN(P2_U3239) );
  XNOR2_X1 U8982 ( .A(n7676), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n7672) );
  XOR2_X1 U8983 ( .A(n7672), .B(n7673), .Z(n7276) );
  NOR2_X1 U8984 ( .A1(n9268), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7790) );
  NOR2_X1 U8985 ( .A1(n4632), .A2(n7268), .ZN(n7265) );
  AOI211_X1 U8986 ( .C1(n9961), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n7790), .B(
        n7265), .ZN(n7275) );
  INV_X1 U8987 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7269) );
  MUX2_X1 U8988 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n7269), .S(n7268), .Z(n7270)
         );
  INV_X1 U8989 ( .A(n7270), .ZN(n7271) );
  OAI21_X1 U8990 ( .B1(n7272), .B2(n7271), .A(n7675), .ZN(n7273) );
  NAND2_X1 U8991 ( .A1(n7273), .A2(n9932), .ZN(n7274) );
  OAI211_X1 U8992 ( .C1(n7276), .C2(n9533), .A(n7275), .B(n7274), .ZN(P1_U3252) );
  INV_X1 U8993 ( .A(n7277), .ZN(n7386) );
  INV_X1 U8994 ( .A(n8332), .ZN(n9852) );
  AOI22_X1 U8995 ( .A1(n9522), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9852), .ZN(n7278) );
  OAI21_X1 U8996 ( .B1(n7386), .B2(n7914), .A(n7278), .ZN(P1_U3337) );
  INV_X1 U8997 ( .A(n7279), .ZN(n7283) );
  AOI21_X1 U8998 ( .B1(n7281), .B2(P2_STATE_REG_SCAN_IN), .A(n7280), .ZN(n7282) );
  OAI21_X1 U8999 ( .B1(n10175), .B2(n7283), .A(n7282), .ZN(n7285) );
  NAND2_X1 U9000 ( .A1(n7285), .A2(n4385), .ZN(n7302) );
  NAND2_X1 U9001 ( .A1(n7302), .A2(n8536), .ZN(n7286) );
  NAND2_X1 U9002 ( .A1(n7286), .A2(n8383), .ZN(n8618) );
  INV_X1 U9003 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7845) );
  INV_X1 U9004 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9163) );
  MUX2_X1 U9005 ( .A(n9163), .B(P2_REG2_REG_1__SCAN_IN), .S(n8538), .Z(n7287)
         );
  AND2_X1 U9006 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n10173), .ZN(n8542) );
  NAND2_X1 U9007 ( .A1(n7287), .A2(n8542), .ZN(n8540) );
  OAI21_X1 U9008 ( .B1(n9163), .B2(n8538), .A(n8540), .ZN(n7389) );
  NAND2_X1 U9009 ( .A1(n7304), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7373) );
  INV_X1 U9010 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7290) );
  MUX2_X1 U9011 ( .A(n7290), .B(P2_REG2_REG_3__SCAN_IN), .S(n7385), .Z(n7288)
         );
  NAND2_X1 U9012 ( .A1(n7289), .A2(n7288), .ZN(n7375) );
  OR2_X1 U9013 ( .A1(n7385), .A2(n7290), .ZN(n7324) );
  NAND2_X1 U9014 ( .A1(n7375), .A2(n7324), .ZN(n7292) );
  INV_X1 U9015 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7322) );
  MUX2_X1 U9016 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7322), .S(n7321), .Z(n7291)
         );
  NAND2_X1 U9017 ( .A1(n7292), .A2(n7291), .ZN(n7339) );
  NAND2_X1 U9018 ( .A1(n7321), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7338) );
  NAND2_X1 U9019 ( .A1(n7339), .A2(n7338), .ZN(n7295) );
  INV_X1 U9020 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7293) );
  MUX2_X1 U9021 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7293), .S(n7336), .Z(n7294)
         );
  NAND2_X1 U9022 ( .A1(n7295), .A2(n7294), .ZN(n7341) );
  NAND2_X1 U9023 ( .A1(n7336), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7300) );
  NAND2_X1 U9024 ( .A1(n7341), .A2(n7300), .ZN(n7298) );
  INV_X1 U9025 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7296) );
  MUX2_X1 U9026 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7296), .S(n7360), .Z(n7297)
         );
  NAND2_X1 U9027 ( .A1(n7298), .A2(n7297), .ZN(n7357) );
  MUX2_X1 U9028 ( .A(n7296), .B(P2_REG2_REG_6__SCAN_IN), .S(n7360), .Z(n7299)
         );
  NAND3_X1 U9029 ( .A1(n7341), .A2(n7300), .A3(n7299), .ZN(n7301) );
  NAND3_X1 U9030 ( .A1(n10163), .A2(n7357), .A3(n7301), .ZN(n7319) );
  INV_X1 U9031 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10300) );
  MUX2_X1 U9032 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10300), .S(n7360), .Z(n7313)
         );
  INV_X1 U9033 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10295) );
  MUX2_X1 U9034 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10295), .S(n7304), .Z(n7393)
         );
  INV_X1 U9035 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10293) );
  MUX2_X1 U9036 ( .A(n10293), .B(P2_REG1_REG_1__SCAN_IN), .S(n8538), .Z(n8546)
         );
  AND2_X1 U9037 ( .A1(n10173), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U9038 ( .A1(n8546), .A2(n8545), .ZN(n8544) );
  INV_X1 U9039 ( .A(n8538), .ZN(n8543) );
  NAND2_X1 U9040 ( .A1(n8543), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7303) );
  NAND2_X1 U9041 ( .A1(n8544), .A2(n7303), .ZN(n7392) );
  NAND2_X1 U9042 ( .A1(n7393), .A2(n7392), .ZN(n7391) );
  NAND2_X1 U9043 ( .A1(n7304), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7305) );
  NAND2_X1 U9044 ( .A1(n7391), .A2(n7305), .ZN(n7377) );
  XNOR2_X1 U9045 ( .A(n7385), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n7378) );
  NAND2_X1 U9046 ( .A1(n7377), .A2(n7378), .ZN(n7376) );
  INV_X1 U9047 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7306) );
  OR2_X1 U9048 ( .A1(n7385), .A2(n7306), .ZN(n7307) );
  NAND2_X1 U9049 ( .A1(n7376), .A2(n7307), .ZN(n7327) );
  INV_X1 U9050 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7308) );
  XNOR2_X1 U9051 ( .A(n7321), .B(n7308), .ZN(n7328) );
  NAND2_X1 U9052 ( .A1(n7327), .A2(n7328), .ZN(n7326) );
  NAND2_X1 U9053 ( .A1(n7321), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7309) );
  NAND2_X1 U9054 ( .A1(n7326), .A2(n7309), .ZN(n7343) );
  INV_X1 U9055 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7310) );
  XNOR2_X1 U9056 ( .A(n7336), .B(n7310), .ZN(n7344) );
  NAND2_X1 U9057 ( .A1(n7343), .A2(n7344), .ZN(n7342) );
  NAND2_X1 U9058 ( .A1(n7336), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7311) );
  NAND2_X1 U9059 ( .A1(n7342), .A2(n7311), .ZN(n7312) );
  NAND2_X1 U9060 ( .A1(n7312), .A2(n7313), .ZN(n7362) );
  OAI21_X1 U9061 ( .B1(n7313), .B2(n7312), .A(n7362), .ZN(n7316) );
  NAND2_X1 U9062 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7520) );
  INV_X1 U9063 ( .A(n7520), .ZN(n7314) );
  AOI21_X1 U9064 ( .B1(n10164), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7314), .ZN(
        n7315) );
  OAI21_X1 U9065 ( .B1(n10167), .B2(n7316), .A(n7315), .ZN(n7317) );
  INV_X1 U9066 ( .A(n7317), .ZN(n7318) );
  OAI211_X1 U9067 ( .C1(n10166), .C2(n7320), .A(n7319), .B(n7318), .ZN(
        P2_U3251) );
  MUX2_X1 U9068 ( .A(n7322), .B(P2_REG2_REG_4__SCAN_IN), .S(n7321), .Z(n7323)
         );
  NAND3_X1 U9069 ( .A1(n7375), .A2(n7324), .A3(n7323), .ZN(n7325) );
  NAND3_X1 U9070 ( .A1(n10163), .A2(n7339), .A3(n7325), .ZN(n7334) );
  OAI21_X1 U9071 ( .B1(n7328), .B2(n7327), .A(n7326), .ZN(n7331) );
  NAND2_X1 U9072 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7502) );
  INV_X1 U9073 ( .A(n7502), .ZN(n7329) );
  AOI21_X1 U9074 ( .B1(n10164), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n7329), .ZN(
        n7330) );
  OAI21_X1 U9075 ( .B1(n10167), .B2(n7331), .A(n7330), .ZN(n7332) );
  INV_X1 U9076 ( .A(n7332), .ZN(n7333) );
  OAI211_X1 U9077 ( .C1(n10166), .C2(n7335), .A(n7334), .B(n7333), .ZN(
        P2_U3249) );
  MUX2_X1 U9078 ( .A(n7293), .B(P2_REG2_REG_5__SCAN_IN), .S(n7336), .Z(n7337)
         );
  NAND3_X1 U9079 ( .A1(n7339), .A2(n7338), .A3(n7337), .ZN(n7340) );
  NAND3_X1 U9080 ( .A1(n10163), .A2(n7341), .A3(n7340), .ZN(n7350) );
  OAI21_X1 U9081 ( .B1(n7344), .B2(n7343), .A(n7342), .ZN(n7347) );
  NAND2_X1 U9082 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7445) );
  INV_X1 U9083 ( .A(n7445), .ZN(n7345) );
  AOI21_X1 U9084 ( .B1(n10164), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7345), .ZN(
        n7346) );
  OAI21_X1 U9085 ( .B1(n10167), .B2(n7347), .A(n7346), .ZN(n7348) );
  INV_X1 U9086 ( .A(n7348), .ZN(n7349) );
  OAI211_X1 U9087 ( .C1(n10166), .C2(n7351), .A(n7350), .B(n7349), .ZN(
        P2_U3250) );
  NAND2_X1 U9088 ( .A1(n7360), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7356) );
  NAND2_X1 U9089 ( .A1(n7357), .A2(n7356), .ZN(n7354) );
  INV_X1 U9090 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7352) );
  MUX2_X1 U9091 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7352), .S(n7409), .Z(n7353)
         );
  NAND2_X1 U9092 ( .A1(n7354), .A2(n7353), .ZN(n8559) );
  MUX2_X1 U9093 ( .A(n7352), .B(P2_REG2_REG_7__SCAN_IN), .S(n7409), .Z(n7355)
         );
  NAND3_X1 U9094 ( .A1(n7357), .A2(n7356), .A3(n7355), .ZN(n7358) );
  NAND3_X1 U9095 ( .A1(n10163), .A2(n8559), .A3(n7358), .ZN(n7370) );
  INV_X1 U9096 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7359) );
  XNOR2_X1 U9097 ( .A(n7409), .B(n7359), .ZN(n7364) );
  NAND2_X1 U9098 ( .A1(n7360), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7361) );
  NAND2_X1 U9099 ( .A1(n7362), .A2(n7361), .ZN(n7363) );
  NAND2_X1 U9100 ( .A1(n7363), .A2(n7364), .ZN(n7401) );
  OAI21_X1 U9101 ( .B1(n7364), .B2(n7363), .A(n7401), .ZN(n7367) );
  INV_X1 U9102 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7527) );
  NOR2_X1 U9103 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7527), .ZN(n7365) );
  AOI21_X1 U9104 ( .B1(n10164), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7365), .ZN(
        n7366) );
  OAI21_X1 U9105 ( .B1(n10167), .B2(n7367), .A(n7366), .ZN(n7368) );
  INV_X1 U9106 ( .A(n7368), .ZN(n7369) );
  OAI211_X1 U9107 ( .C1(n10166), .C2(n7371), .A(n7370), .B(n7369), .ZN(
        P2_U3252) );
  MUX2_X1 U9108 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7290), .S(n7385), .Z(n7372)
         );
  NAND3_X1 U9109 ( .A1(n7388), .A2(n7373), .A3(n7372), .ZN(n7374) );
  NAND3_X1 U9110 ( .A1(n10163), .A2(n7375), .A3(n7374), .ZN(n7384) );
  OAI21_X1 U9111 ( .B1(n7378), .B2(n7377), .A(n7376), .ZN(n7381) );
  INV_X1 U9112 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7379) );
  NOR2_X1 U9113 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7379), .ZN(n10149) );
  AOI21_X1 U9114 ( .B1(n10164), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n10149), .ZN(
        n7380) );
  OAI21_X1 U9115 ( .B1(n10167), .B2(n7381), .A(n7380), .ZN(n7382) );
  INV_X1 U9116 ( .A(n7382), .ZN(n7383) );
  OAI211_X1 U9117 ( .C1(n10166), .C2(n7385), .A(n7384), .B(n7383), .ZN(
        P2_U3248) );
  INV_X1 U9118 ( .A(n8031), .ZN(n7770) );
  OAI222_X1 U9119 ( .A1(n9043), .A2(n7387), .B1(n9036), .B2(n7386), .C1(n7770), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  OAI211_X1 U9120 ( .C1(n7390), .C2(n7389), .A(n10163), .B(n7388), .ZN(n7398)
         );
  OAI21_X1 U9121 ( .B1(n7393), .B2(n7392), .A(n7391), .ZN(n7395) );
  AOI22_X1 U9122 ( .A1(n10164), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n7394) );
  OAI21_X1 U9123 ( .B1(n10167), .B2(n7395), .A(n7394), .ZN(n7396) );
  INV_X1 U9124 ( .A(n7396), .ZN(n7397) );
  OAI211_X1 U9125 ( .C1(n10166), .C2(n7399), .A(n7398), .B(n7397), .ZN(
        P2_U3247) );
  INV_X1 U9126 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10312) );
  MUX2_X1 U9127 ( .A(n10312), .B(P2_REG1_REG_12__SCAN_IN), .S(n7463), .Z(n7408) );
  NAND2_X1 U9128 ( .A1(n7409), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7400) );
  NAND2_X1 U9129 ( .A1(n7401), .A2(n7400), .ZN(n8554) );
  XNOR2_X1 U9130 ( .A(n8556), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n8555) );
  NAND2_X1 U9131 ( .A1(n8554), .A2(n8555), .ZN(n8553) );
  NAND2_X1 U9132 ( .A1(n7412), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7402) );
  NAND2_X1 U9133 ( .A1(n8553), .A2(n7402), .ZN(n8571) );
  INV_X1 U9134 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10305) );
  MUX2_X1 U9135 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10305), .S(n9319), .Z(n8572)
         );
  NAND2_X1 U9136 ( .A1(n8571), .A2(n8572), .ZN(n8570) );
  NAND2_X1 U9137 ( .A1(n9319), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7403) );
  NAND2_X1 U9138 ( .A1(n8570), .A2(n7403), .ZN(n8585) );
  INV_X1 U9139 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10307) );
  MUX2_X1 U9140 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n10307), .S(n8587), .Z(n8586) );
  NAND2_X1 U9141 ( .A1(n8585), .A2(n8586), .ZN(n8584) );
  NAND2_X1 U9142 ( .A1(n8587), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7404) );
  NAND2_X1 U9143 ( .A1(n8584), .A2(n7404), .ZN(n7459) );
  INV_X1 U9144 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10309) );
  MUX2_X1 U9145 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10309), .S(n7418), .Z(n7458) );
  NAND2_X1 U9146 ( .A1(n7459), .A2(n7458), .ZN(n7457) );
  NAND2_X1 U9147 ( .A1(n7418), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7405) );
  NAND2_X1 U9148 ( .A1(n7457), .A2(n7405), .ZN(n7407) );
  INV_X1 U9149 ( .A(n7475), .ZN(n7406) );
  AOI21_X1 U9150 ( .B1(n7408), .B2(n7407), .A(n7406), .ZN(n7427) );
  NAND2_X1 U9151 ( .A1(n7409), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U9152 ( .A1(n8559), .A2(n8558), .ZN(n7411) );
  INV_X1 U9153 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8067) );
  MUX2_X1 U9154 ( .A(n8067), .B(P2_REG2_REG_8__SCAN_IN), .S(n8556), .Z(n7410)
         );
  NAND2_X1 U9155 ( .A1(n7412), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8565) );
  INV_X1 U9156 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7413) );
  MUX2_X1 U9157 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7413), .S(n9319), .Z(n7414)
         );
  NAND2_X1 U9158 ( .A1(n9319), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8578) );
  INV_X1 U9159 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8888) );
  MUX2_X1 U9160 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n8888), .S(n8587), .Z(n7415)
         );
  NAND2_X1 U9161 ( .A1(n7416), .A2(n7415), .ZN(n8581) );
  NAND2_X1 U9162 ( .A1(n8587), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7417) );
  NAND2_X1 U9163 ( .A1(n8581), .A2(n7417), .ZN(n7453) );
  INV_X1 U9164 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7969) );
  MUX2_X1 U9165 ( .A(n7969), .B(P2_REG2_REG_11__SCAN_IN), .S(n7418), .Z(n7452)
         );
  NAND2_X1 U9166 ( .A1(n7454), .A2(n7969), .ZN(n7419) );
  NAND2_X1 U9167 ( .A1(n7450), .A2(n7419), .ZN(n7421) );
  INV_X1 U9168 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n9212) );
  MUX2_X1 U9169 ( .A(n9212), .B(P2_REG2_REG_12__SCAN_IN), .S(n7463), .Z(n7420)
         );
  AOI21_X1 U9170 ( .B1(n7421), .B2(n7420), .A(n10165), .ZN(n7425) );
  NAND2_X1 U9171 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n8012) );
  INV_X1 U9172 ( .A(n8012), .ZN(n7422) );
  AOI21_X1 U9173 ( .B1(n10164), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7422), .ZN(
        n7423) );
  OAI21_X1 U9174 ( .B1(n10166), .B2(n7473), .A(n7423), .ZN(n7424) );
  AOI21_X1 U9175 ( .B1(n7425), .B2(n7465), .A(n7424), .ZN(n7426) );
  OAI21_X1 U9176 ( .B1(n7427), .B2(n10167), .A(n7426), .ZN(P2_U3257) );
  XNOR2_X1 U9177 ( .A(n7598), .B(n7602), .ZN(n7429) );
  XNOR2_X1 U9178 ( .A(n7600), .B(n7429), .ZN(n7435) );
  NAND2_X1 U9179 ( .A1(n9440), .A2(n9487), .ZN(n7431) );
  OAI211_X1 U9180 ( .C1(n9988), .C2(n9451), .A(n7431), .B(n7430), .ZN(n7432)
         );
  AOI21_X1 U9181 ( .B1(n9975), .B2(n9462), .A(n7432), .ZN(n7434) );
  NAND2_X1 U9182 ( .A1(n9470), .A2(n9976), .ZN(n7433) );
  OAI211_X1 U9183 ( .C1(n7435), .C2(n9472), .A(n7434), .B(n7433), .ZN(P1_U3219) );
  INV_X1 U9184 ( .A(n7436), .ZN(n7515) );
  AOI22_X1 U9185 ( .A1(n9532), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9852), .ZN(n7437) );
  OAI21_X1 U9186 ( .B1(n7515), .B2(n7914), .A(n7437), .ZN(P1_U3336) );
  NAND2_X1 U9187 ( .A1(n7500), .A2(n7439), .ZN(n7442) );
  INV_X1 U9188 ( .A(n7440), .ZN(n7441) );
  AOI211_X1 U9189 ( .C1(n7443), .C2(n7442), .A(n7441), .B(n8519), .ZN(n7448)
         );
  NAND2_X1 U9190 ( .A1(n10151), .A2(n7854), .ZN(n7444) );
  OAI211_X1 U9191 ( .C1(n10161), .C2(n7855), .A(n7445), .B(n7444), .ZN(n7447)
         );
  OAI22_X1 U9192 ( .A1(n10144), .A2(n10148), .B1(n10145), .B2(n7528), .ZN(
        n7446) );
  OR3_X1 U9193 ( .A1(n7448), .A2(n7447), .A3(n7446), .ZN(P2_U3229) );
  INV_X1 U9194 ( .A(P1_U4006), .ZN(n7526) );
  NAND2_X1 U9195 ( .A1(n7526), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7449) );
  OAI21_X1 U9196 ( .B1(n8313), .B2(n7526), .A(n7449), .ZN(P1_U3584) );
  INV_X1 U9197 ( .A(n7450), .ZN(n7451) );
  AOI21_X1 U9198 ( .B1(n7453), .B2(n7452), .A(n7451), .ZN(n7462) );
  NOR2_X1 U9199 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9161), .ZN(n7456) );
  NOR2_X1 U9200 ( .A1(n10166), .A2(n7454), .ZN(n7455) );
  AOI211_X1 U9201 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n10164), .A(n7456), .B(
        n7455), .ZN(n7461) );
  OAI211_X1 U9202 ( .C1(n7459), .C2(n7458), .A(n7457), .B(n10162), .ZN(n7460)
         );
  OAI211_X1 U9203 ( .C1(n7462), .C2(n10165), .A(n7461), .B(n7460), .ZN(
        P2_U3256) );
  NAND2_X1 U9204 ( .A1(n7463), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7464) );
  INV_X1 U9205 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7466) );
  MUX2_X1 U9206 ( .A(n7466), .B(P2_REG2_REG_13__SCAN_IN), .S(n7486), .Z(n7468)
         );
  INV_X1 U9207 ( .A(n7491), .ZN(n7467) );
  AOI21_X1 U9208 ( .B1(n7469), .B2(n7468), .A(n7467), .ZN(n7481) );
  INV_X1 U9209 ( .A(n10164), .ZN(n7777) );
  INV_X1 U9210 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7471) );
  OAI22_X1 U9211 ( .A1(n7777), .A2(n7471), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7470), .ZN(n7472) );
  AOI21_X1 U9212 ( .B1(n8588), .B2(n7486), .A(n7472), .ZN(n7480) );
  XNOR2_X1 U9213 ( .A(n7486), .B(n9215), .ZN(n7477) );
  NAND2_X1 U9214 ( .A1(n7473), .A2(n10312), .ZN(n7474) );
  NAND2_X1 U9215 ( .A1(n7475), .A2(n7474), .ZN(n7476) );
  NAND2_X1 U9216 ( .A1(n7476), .A2(n7477), .ZN(n7484) );
  OAI21_X1 U9217 ( .B1(n7477), .B2(n7476), .A(n7484), .ZN(n7478) );
  NAND2_X1 U9218 ( .A1(n7478), .A2(n10162), .ZN(n7479) );
  OAI211_X1 U9219 ( .C1(n7481), .C2(n10165), .A(n7480), .B(n7479), .ZN(
        P2_U3258) );
  INV_X1 U9220 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7482) );
  XNOR2_X1 U9221 ( .A(n7762), .B(n7482), .ZN(n7764) );
  OR2_X1 U9222 ( .A1(n7486), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7483) );
  XOR2_X1 U9223 ( .A(n7764), .B(n7765), .Z(n7496) );
  INV_X1 U9224 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9241) );
  AND2_X1 U9225 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8403) );
  INV_X1 U9226 ( .A(n8403), .ZN(n7485) );
  OAI21_X1 U9227 ( .B1(n7777), .B2(n9241), .A(n7485), .ZN(n7494) );
  OR2_X1 U9228 ( .A1(n7486), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7489) );
  INV_X1 U9229 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9240) );
  MUX2_X1 U9230 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n9240), .S(n7762), .Z(n7488)
         );
  NAND2_X1 U9231 ( .A1(n7487), .A2(n7488), .ZN(n7757) );
  INV_X1 U9232 ( .A(n7488), .ZN(n7490) );
  NAND3_X1 U9233 ( .A1(n7491), .A2(n7490), .A3(n7489), .ZN(n7492) );
  AOI21_X1 U9234 ( .B1(n7757), .B2(n7492), .A(n10165), .ZN(n7493) );
  AOI211_X1 U9235 ( .C1(n8588), .C2(n7762), .A(n7494), .B(n7493), .ZN(n7495)
         );
  OAI21_X1 U9236 ( .B1(n10167), .B2(n7496), .A(n7495), .ZN(P2_U3259) );
  OAI22_X1 U9237 ( .A1(n7957), .A2(n10148), .B1(n10145), .B2(n7958), .ZN(n7505) );
  NAND2_X1 U9238 ( .A1(n7497), .A2(n7498), .ZN(n7499) );
  AOI21_X1 U9239 ( .B1(n7500), .B2(n7499), .A(n8519), .ZN(n7504) );
  NAND2_X1 U9240 ( .A1(n10151), .A2(n7959), .ZN(n7501) );
  OAI211_X1 U9241 ( .C1(n10161), .C2(n7950), .A(n7502), .B(n7501), .ZN(n7503)
         );
  OR3_X1 U9242 ( .A1(n7505), .A2(n7504), .A3(n7503), .ZN(P2_U3232) );
  NAND2_X1 U9243 ( .A1(n8537), .A2(n8815), .ZN(n7507) );
  NAND2_X1 U9244 ( .A1(n10146), .A2(n8816), .ZN(n7506) );
  AND2_X1 U9245 ( .A1(n7507), .A2(n7506), .ZN(n8152) );
  AOI22_X1 U9246 ( .A1(n10151), .A2(n7508), .B1(n7537), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7514) );
  OAI21_X1 U9247 ( .B1(n7511), .B2(n7510), .A(n7509), .ZN(n7512) );
  NAND2_X1 U9248 ( .A1(n10153), .A2(n7512), .ZN(n7513) );
  OAI211_X1 U9249 ( .C1(n8152), .C2(n8516), .A(n7514), .B(n7513), .ZN(P2_U3224) );
  INV_X1 U9250 ( .A(n8598), .ZN(n8029) );
  OAI222_X1 U9251 ( .A1(n9043), .A2(n7516), .B1(n9036), .B2(n7515), .C1(n8029), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  OAI21_X1 U9252 ( .B1(n4474), .B2(n7518), .A(n7517), .ZN(n7523) );
  NAND2_X1 U9253 ( .A1(n10151), .A2(n7933), .ZN(n7519) );
  OAI211_X1 U9254 ( .C1(n10161), .C2(n7930), .A(n7520), .B(n7519), .ZN(n7522)
         );
  OAI22_X1 U9255 ( .A1(n7958), .A2(n10148), .B1(n10145), .B2(n7939), .ZN(n7521) );
  AOI211_X1 U9256 ( .C1(n10153), .C2(n7523), .A(n7522), .B(n7521), .ZN(n7524)
         );
  INV_X1 U9257 ( .A(n7524), .ZN(P2_U3241) );
  NAND2_X1 U9258 ( .A1(n7526), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7525) );
  OAI21_X1 U9259 ( .B1(n9602), .B2(n7526), .A(n7525), .ZN(P1_U3582) );
  INV_X1 U9260 ( .A(n7889), .ZN(n7531) );
  INV_X1 U9261 ( .A(n10161), .ZN(n8513) );
  OAI22_X1 U9262 ( .A1(n8459), .A2(n10239), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7527), .ZN(n7530) );
  OAI22_X1 U9263 ( .A1(n7528), .A2(n10148), .B1(n10145), .B2(n7667), .ZN(n7529) );
  AOI211_X1 U9264 ( .C1(n7531), .C2(n8513), .A(n7530), .B(n7529), .ZN(n7536)
         );
  OAI211_X1 U9265 ( .C1(n7534), .C2(n7533), .A(n7532), .B(n10153), .ZN(n7535)
         );
  NAND2_X1 U9266 ( .A1(n7536), .A2(n7535), .ZN(P2_U3215) );
  INV_X1 U9267 ( .A(n4376), .ZN(n7544) );
  AOI22_X1 U9268 ( .A1(n8124), .A2(n10151), .B1(n7537), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n7543) );
  INV_X1 U9269 ( .A(n8537), .ZN(n7539) );
  OAI21_X1 U9270 ( .B1(n7539), .B2(n7538), .A(n10188), .ZN(n7540) );
  NAND3_X1 U9271 ( .A1(n10153), .A2(n7541), .A3(n7540), .ZN(n7542) );
  OAI211_X1 U9272 ( .C1(n10145), .C2(n7544), .A(n7543), .B(n7542), .ZN(
        P2_U3234) );
  OAI211_X1 U9273 ( .C1(n7547), .C2(n7546), .A(n7545), .B(n10153), .ZN(n7551)
         );
  INV_X1 U9274 ( .A(n8516), .ZN(n7549) );
  OAI22_X1 U9275 ( .A1(n7939), .A2(n8882), .B1(n8883), .B2(n8880), .ZN(n8065)
         );
  AND2_X1 U9276 ( .A1(P2_U3152), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8552) );
  OAI22_X1 U9277 ( .A1(n8459), .A2(n8070), .B1(n10161), .B2(n8069), .ZN(n7548)
         );
  AOI211_X1 U9278 ( .C1(n7549), .C2(n8065), .A(n8552), .B(n7548), .ZN(n7550)
         );
  NAND2_X1 U9279 ( .A1(n7551), .A2(n7550), .ZN(P2_U3223) );
  NAND2_X1 U9280 ( .A1(n7552), .A2(n7556), .ZN(n7558) );
  NOR2_X1 U9281 ( .A1(n9490), .A2(n7553), .ZN(n7630) );
  NOR2_X1 U9282 ( .A1(n7554), .A2(n7647), .ZN(n7555) );
  AOI21_X1 U9283 ( .B1(n7556), .B2(n7630), .A(n7555), .ZN(n7557) );
  OAI21_X1 U9284 ( .B1(n7559), .B2(n7558), .A(n7557), .ZN(n10023) );
  NAND2_X1 U9285 ( .A1(n10023), .A2(n10035), .ZN(n7561) );
  NAND2_X1 U9286 ( .A1(n10016), .A2(n10082), .ZN(n7560) );
  NAND2_X1 U9287 ( .A1(n10038), .A2(n10006), .ZN(n9985) );
  AND2_X1 U9288 ( .A1(n7563), .A2(n9985), .ZN(n7562) );
  INV_X1 U9289 ( .A(n9994), .ZN(n9996) );
  NAND2_X1 U9290 ( .A1(n9996), .A2(n10017), .ZN(n7564) );
  INV_X1 U9291 ( .A(n7689), .ZN(n7566) );
  NAND2_X1 U9292 ( .A1(n7686), .A2(n7566), .ZN(n7567) );
  XNOR2_X1 U9293 ( .A(n7567), .B(n7688), .ZN(n10109) );
  INV_X1 U9294 ( .A(n7569), .ZN(n7570) );
  NOR2_X1 U9295 ( .A1(n9990), .A2(n7570), .ZN(n7571) );
  NAND2_X1 U9296 ( .A1(n7571), .A2(n7688), .ZN(n9970) );
  OAI21_X1 U9297 ( .B1(n7688), .B2(n7571), .A(n9970), .ZN(n7572) );
  INV_X1 U9298 ( .A(n10017), .ZN(n9489) );
  AOI222_X1 U9299 ( .A1(n10043), .A2(n7572), .B1(n9488), .B2(n10037), .C1(
        n9489), .C2(n9715), .ZN(n10108) );
  MUX2_X1 U9300 ( .A(n7103), .B(n10108), .S(n10033), .Z(n7579) );
  NAND2_X1 U9301 ( .A1(n10003), .A2(n9996), .ZN(n9995) );
  AOI211_X1 U9302 ( .C1(n10105), .C2(n9995), .A(n10121), .B(n4979), .ZN(n10104) );
  NOR2_X1 U9303 ( .A1(n7575), .A2(n10011), .ZN(n9616) );
  OAI22_X1 U9304 ( .A1(n5407), .A2(n9710), .B1(n7576), .B2(n10031), .ZN(n7577)
         );
  AOI21_X1 U9305 ( .B1(n10104), .B2(n9616), .A(n7577), .ZN(n7578) );
  OAI211_X1 U9306 ( .C1(n10109), .C2(n9722), .A(n7579), .B(n7578), .ZN(
        P1_U3284) );
  NAND2_X1 U9307 ( .A1(n7581), .A2(n7580), .ZN(n8344) );
  XNOR2_X1 U9308 ( .A(n7583), .B(n7582), .ZN(n8343) );
  OR2_X1 U9309 ( .A1(n8344), .A2(n8343), .ZN(n8345) );
  AND2_X1 U9310 ( .A1(n8345), .A2(n7584), .ZN(n7586) );
  NAND2_X1 U9311 ( .A1(n7586), .A2(n7585), .ZN(n7722) );
  OAI21_X1 U9312 ( .B1(n7586), .B2(n7585), .A(n7722), .ZN(n7587) );
  NOR2_X1 U9313 ( .A1(n7587), .A2(n7588), .ZN(n7724) );
  AOI21_X1 U9314 ( .B1(n7588), .B2(n7587), .A(n7724), .ZN(n7595) );
  NAND2_X1 U9315 ( .A1(n9464), .A2(n5364), .ZN(n7590) );
  OAI211_X1 U9316 ( .C1(n10017), .C2(n9467), .A(n7590), .B(n7589), .ZN(n7593)
         );
  NOR2_X1 U9317 ( .A1(n9437), .A2(n7591), .ZN(n7592) );
  AOI211_X1 U9318 ( .C1(n9470), .C2(n10006), .A(n7593), .B(n7592), .ZN(n7594)
         );
  OAI21_X1 U9319 ( .B1(n7595), .B2(n9472), .A(n7594), .ZN(P1_U3225) );
  NAND2_X1 U9320 ( .A1(n6804), .A2(n7597), .ZN(n7605) );
  INV_X1 U9321 ( .A(n7600), .ZN(n7603) );
  OAI21_X1 U9322 ( .B1(n7600), .B2(n7599), .A(n7598), .ZN(n7601) );
  OAI21_X1 U9323 ( .B1(n7603), .B2(n7602), .A(n7601), .ZN(n7604) );
  XOR2_X1 U9324 ( .A(n7605), .B(n7604), .Z(n7611) );
  INV_X1 U9325 ( .A(n7814), .ZN(n9486) );
  NAND2_X1 U9326 ( .A1(n9440), .A2(n9486), .ZN(n7607) );
  OAI211_X1 U9327 ( .C1(n7739), .C2(n9451), .A(n7607), .B(n7606), .ZN(n7609)
         );
  INV_X1 U9328 ( .A(n7747), .ZN(n10120) );
  NOR2_X1 U9329 ( .A1(n10120), .A2(n9456), .ZN(n7608) );
  AOI211_X1 U9330 ( .C1(n7746), .C2(n9462), .A(n7609), .B(n7608), .ZN(n7610)
         );
  OAI21_X1 U9331 ( .B1(n7611), .B2(n9472), .A(n7610), .ZN(P1_U3229) );
  NAND2_X1 U9332 ( .A1(n7614), .A2(n7613), .ZN(n7615) );
  XNOR2_X1 U9333 ( .A(n7616), .B(n7615), .ZN(n7622) );
  NAND2_X1 U9334 ( .A1(n9440), .A2(n9485), .ZN(n7618) );
  OAI211_X1 U9335 ( .C1(n9967), .C2(n9451), .A(n7618), .B(n7617), .ZN(n7620)
         );
  INV_X1 U9336 ( .A(n7815), .ZN(n7876) );
  NOR2_X1 U9337 ( .A1(n7876), .A2(n9456), .ZN(n7619) );
  AOI211_X1 U9338 ( .C1(n7714), .C2(n9462), .A(n7620), .B(n7619), .ZN(n7621)
         );
  OAI21_X1 U9339 ( .B1(n7622), .B2(n9472), .A(n7621), .ZN(P1_U3215) );
  INV_X1 U9340 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7624) );
  OAI22_X1 U9341 ( .A1(n10033), .A2(n7624), .B1(n7623), .B2(n10031), .ZN(n7625) );
  INV_X1 U9342 ( .A(n7625), .ZN(n7628) );
  OAI21_X1 U9343 ( .B1(n10050), .B2(n10028), .A(n7626), .ZN(n7627) );
  OAI211_X1 U9344 ( .C1(n7629), .C2(n10047), .A(n7628), .B(n7627), .ZN(
        P1_U3291) );
  NOR2_X1 U9345 ( .A1(n7631), .A2(n7630), .ZN(n7633) );
  XNOR2_X1 U9346 ( .A(n7633), .B(n7556), .ZN(n10075) );
  INV_X1 U9347 ( .A(n10034), .ZN(n7819) );
  INV_X1 U9348 ( .A(n7634), .ZN(n7635) );
  AOI21_X1 U9349 ( .B1(n7637), .B2(n7636), .A(n7635), .ZN(n7638) );
  XNOR2_X1 U9350 ( .A(n7638), .B(n7556), .ZN(n7640) );
  OAI22_X1 U9351 ( .A1(n7655), .A2(n10040), .B1(n10016), .B2(n10018), .ZN(
        n7639) );
  AOI21_X1 U9352 ( .B1(n7640), .B2(n10043), .A(n7639), .ZN(n7641) );
  OAI21_X1 U9353 ( .B1(n10075), .B2(n7819), .A(n7641), .ZN(n10078) );
  NAND2_X1 U9354 ( .A1(n10078), .A2(n10033), .ZN(n7649) );
  OAI22_X1 U9355 ( .A1(n10033), .A2(n7642), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10031), .ZN(n7646) );
  NAND2_X1 U9356 ( .A1(n7643), .A2(n7647), .ZN(n7644) );
  NAND2_X1 U9357 ( .A1(n10024), .A2(n7644), .ZN(n10077) );
  NOR2_X1 U9358 ( .A1(n9573), .A2(n10077), .ZN(n7645) );
  AOI211_X1 U9359 ( .C1(n10050), .C2(n7647), .A(n7646), .B(n7645), .ZN(n7648)
         );
  OAI211_X1 U9360 ( .C1(n10075), .C2(n8218), .A(n7649), .B(n7648), .ZN(
        P1_U3288) );
  OAI21_X1 U9361 ( .B1(n7650), .B2(n7652), .A(n7651), .ZN(n10063) );
  OAI21_X1 U9362 ( .B1(n5786), .B2(n7653), .A(n5815), .ZN(n7657) );
  OAI22_X1 U9363 ( .A1(n7655), .A2(n10018), .B1(n7654), .B2(n10040), .ZN(n7656) );
  AOI21_X1 U9364 ( .B1(n7657), .B2(n10043), .A(n7656), .ZN(n7658) );
  OAI21_X1 U9365 ( .B1(n7819), .B2(n10063), .A(n7658), .ZN(n10065) );
  OAI211_X1 U9366 ( .C1(n5819), .C2(n4966), .A(n4933), .B(n10004), .ZN(n10064)
         );
  INV_X1 U9367 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7660) );
  OAI22_X1 U9368 ( .A1(n10064), .A2(n10011), .B1(n10031), .B2(n7660), .ZN(
        n7661) );
  OAI21_X1 U9369 ( .B1(n10065), .B2(n7661), .A(n10033), .ZN(n7663) );
  AOI22_X1 U9370 ( .A1(n10050), .A2(n4997), .B1(n10047), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7662) );
  OAI211_X1 U9371 ( .C1(n10063), .C2(n8218), .A(n7663), .B(n7662), .ZN(
        P1_U3290) );
  NOR2_X1 U9372 ( .A1(n4470), .A2(n7664), .ZN(n7665) );
  XNOR2_X1 U9373 ( .A(n7666), .B(n7665), .ZN(n7671) );
  NAND2_X1 U9374 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8568) );
  OAI21_X1 U9375 ( .B1(n10161), .B2(n8115), .A(n8568), .ZN(n7669) );
  OAI22_X1 U9376 ( .A1(n7667), .A2(n10148), .B1(n10145), .B2(n7967), .ZN(n7668) );
  AOI211_X1 U9377 ( .C1(n10151), .C2(n8114), .A(n7669), .B(n7668), .ZN(n7670)
         );
  OAI21_X1 U9378 ( .B1(n7671), .B2(n8519), .A(n7670), .ZN(P2_U3233) );
  XOR2_X1 U9379 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7866), .Z(n7862) );
  XOR2_X1 U9380 ( .A(n7862), .B(n7863), .Z(n7682) );
  NAND2_X1 U9381 ( .A1(n9957), .A2(n7866), .ZN(n7674) );
  NAND2_X1 U9382 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7998) );
  NAND2_X1 U9383 ( .A1(n7674), .A2(n7998), .ZN(n7680) );
  XNOR2_X1 U9384 ( .A(n7866), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7678) );
  AOI211_X1 U9385 ( .C1(n7678), .C2(n7677), .A(n9950), .B(n7865), .ZN(n7679)
         );
  AOI211_X1 U9386 ( .C1(n9961), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n7680), .B(
        n7679), .ZN(n7681) );
  OAI21_X1 U9387 ( .B1(n9533), .B2(n7682), .A(n7681), .ZN(P1_U3253) );
  INV_X1 U9388 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7684) );
  INV_X1 U9389 ( .A(n7683), .ZN(n7685) );
  INV_X1 U9390 ( .A(n9956), .ZN(n8254) );
  OAI222_X1 U9391 ( .A1(n8332), .A2(n7684), .B1(n7914), .B2(n7685), .C1(
        P1_U3084), .C2(n8254), .ZN(P1_U3335) );
  INV_X1 U9392 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n9235) );
  INV_X1 U9393 ( .A(n8610), .ZN(n8603) );
  OAI222_X1 U9394 ( .A1(n9043), .A2(n9235), .B1(n9036), .B2(n7685), .C1(
        P2_U3152), .C2(n8603), .ZN(P2_U3340) );
  INV_X1 U9395 ( .A(n7688), .ZN(n7687) );
  NAND2_X1 U9396 ( .A1(n9976), .A2(n9488), .ZN(n7692) );
  OR2_X1 U9397 ( .A1(n7747), .A2(n9487), .ZN(n7693) );
  NAND2_X1 U9398 ( .A1(n7747), .A2(n9487), .ZN(n7694) );
  INV_X1 U9399 ( .A(n7817), .ZN(n7697) );
  AOI21_X1 U9400 ( .B1(n7708), .B2(n7695), .A(n7697), .ZN(n7874) );
  AOI22_X1 U9401 ( .A1(n9715), .A2(n9487), .B1(n9485), .B2(n10037), .ZN(n7712)
         );
  INV_X1 U9402 ( .A(n7699), .ZN(n7701) );
  INV_X1 U9403 ( .A(n9969), .ZN(n7700) );
  NAND2_X1 U9404 ( .A1(n7812), .A2(n7707), .ZN(n7709) );
  XNOR2_X1 U9405 ( .A(n7709), .B(n7708), .ZN(n7710) );
  NAND2_X1 U9406 ( .A1(n7710), .A2(n10043), .ZN(n7711) );
  OAI211_X1 U9407 ( .C1(n7874), .C2(n7819), .A(n7712), .B(n7711), .ZN(n7877)
         );
  NAND2_X1 U9408 ( .A1(n7877), .A2(n10033), .ZN(n7719) );
  OAI211_X1 U9409 ( .C1(n7745), .C2(n7876), .A(n10004), .B(n7823), .ZN(n7875)
         );
  INV_X1 U9410 ( .A(n7875), .ZN(n7717) );
  INV_X1 U9411 ( .A(n10031), .ZN(n10009) );
  AOI22_X1 U9412 ( .A1(n10047), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7714), .B2(
        n10009), .ZN(n7715) );
  OAI21_X1 U9413 ( .B1(n7876), .B2(n9710), .A(n7715), .ZN(n7716) );
  AOI21_X1 U9414 ( .B1(n7717), .B2(n9616), .A(n7716), .ZN(n7718) );
  OAI211_X1 U9415 ( .C1(n7874), .C2(n8218), .A(n7719), .B(n7718), .ZN(P1_U3281) );
  NAND2_X1 U9416 ( .A1(n7721), .A2(n7720), .ZN(n7726) );
  INV_X1 U9417 ( .A(n7722), .ZN(n7723) );
  NOR2_X1 U9418 ( .A1(n7724), .A2(n7723), .ZN(n7725) );
  XOR2_X1 U9419 ( .A(n7726), .B(n7725), .Z(n7733) );
  AND2_X1 U9420 ( .A1(n9994), .A2(n10106), .ZN(n10096) );
  NAND2_X1 U9421 ( .A1(n9462), .A2(n9993), .ZN(n7729) );
  AOI21_X1 U9422 ( .B1(n9464), .B2(n10038), .A(n7727), .ZN(n7728) );
  OAI211_X1 U9423 ( .C1(n9988), .C2(n9467), .A(n7729), .B(n7728), .ZN(n7730)
         );
  AOI21_X1 U9424 ( .B1(n7731), .B2(n10096), .A(n7730), .ZN(n7732) );
  OAI21_X1 U9425 ( .B1(n7733), .B2(n9472), .A(n7732), .ZN(P1_U3237) );
  XNOR2_X1 U9426 ( .A(n7734), .B(n7737), .ZN(n7743) );
  NAND2_X1 U9427 ( .A1(n7735), .A2(n7736), .ZN(n7738) );
  XNOR2_X1 U9428 ( .A(n7738), .B(n7737), .ZN(n7741) );
  OAI22_X1 U9429 ( .A1(n7739), .A2(n10040), .B1(n7814), .B2(n10018), .ZN(n7740) );
  AOI21_X1 U9430 ( .B1(n7741), .B2(n10043), .A(n7740), .ZN(n7742) );
  OAI21_X1 U9431 ( .B1(n7743), .B2(n7819), .A(n7742), .ZN(n10123) );
  INV_X1 U9432 ( .A(n10123), .ZN(n7752) );
  INV_X1 U9433 ( .A(n7743), .ZN(n10125) );
  NOR2_X1 U9434 ( .A1(n9977), .A2(n10120), .ZN(n7744) );
  OR2_X1 U9435 ( .A1(n7745), .A2(n7744), .ZN(n10122) );
  AOI22_X1 U9436 ( .A1(n10047), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7746), .B2(
        n10009), .ZN(n7749) );
  NAND2_X1 U9437 ( .A1(n7747), .A2(n10050), .ZN(n7748) );
  OAI211_X1 U9438 ( .C1(n10122), .C2(n9573), .A(n7749), .B(n7748), .ZN(n7750)
         );
  AOI21_X1 U9439 ( .B1(n10125), .B2(n10029), .A(n7750), .ZN(n7751) );
  OAI21_X1 U9440 ( .B1(n7752), .B2(n10047), .A(n7751), .ZN(P1_U3282) );
  INV_X1 U9441 ( .A(n7753), .ZN(n7755) );
  OAI222_X1 U9442 ( .A1(n8332), .A2(n9250), .B1(n7914), .B2(n7755), .C1(
        P1_U3084), .C2(n7754), .ZN(P1_U3334) );
  OAI222_X1 U9443 ( .A1(n9043), .A2(n9077), .B1(n9036), .B2(n7755), .C1(n4760), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OR2_X1 U9444 ( .A1(n7762), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U9445 ( .A1(n7757), .A2(n7756), .ZN(n7759) );
  NAND2_X1 U9446 ( .A1(n7759), .A2(n7758), .ZN(n7761) );
  OR2_X1 U9447 ( .A1(n7759), .A2(n7758), .ZN(n7760) );
  NAND2_X1 U9448 ( .A1(n7761), .A2(n7760), .ZN(n7778) );
  MUX2_X1 U9449 ( .A(n6140), .B(P2_REG2_REG_16__SCAN_IN), .S(n8031), .Z(n8020)
         );
  XNOR2_X1 U9450 ( .A(n8021), .B(n8020), .ZN(n7774) );
  XNOR2_X1 U9451 ( .A(n8031), .B(n8990), .ZN(n7768) );
  NOR2_X1 U9452 ( .A1(n7762), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7763) );
  AOI21_X1 U9453 ( .B1(n7765), .B2(n7764), .A(n7763), .ZN(n7766) );
  XOR2_X1 U9454 ( .A(n7783), .B(n7766), .Z(n7775) );
  AOI21_X1 U9455 ( .B1(n7766), .B2(n7783), .A(n7785), .ZN(n7767) );
  NAND2_X1 U9456 ( .A1(n7767), .A2(n7768), .ZN(n8030) );
  OAI21_X1 U9457 ( .B1(n7768), .B2(n7767), .A(n8030), .ZN(n7769) );
  NAND2_X1 U9458 ( .A1(n7769), .A2(n10162), .ZN(n7773) );
  AND2_X1 U9459 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8455) );
  NOR2_X1 U9460 ( .A1(n10166), .A2(n7770), .ZN(n7771) );
  AOI211_X1 U9461 ( .C1(P2_ADDR_REG_16__SCAN_IN), .C2(n10164), .A(n8455), .B(
        n7771), .ZN(n7772) );
  OAI211_X1 U9462 ( .C1(n7774), .C2(n10165), .A(n7773), .B(n7772), .ZN(
        P2_U3261) );
  OAI21_X1 U9463 ( .B1(n7775), .B2(P2_REG1_REG_15__SCAN_IN), .A(n10162), .ZN(
        n7786) );
  INV_X1 U9464 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7776) );
  NAND2_X1 U9465 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8514) );
  OAI21_X1 U9466 ( .B1(n7777), .B2(n7776), .A(n8514), .ZN(n7782) );
  NAND2_X1 U9467 ( .A1(n7778), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7779) );
  AOI21_X1 U9468 ( .B1(n7780), .B2(n7779), .A(n10165), .ZN(n7781) );
  AOI211_X1 U9469 ( .C1(n8588), .C2(n7783), .A(n7782), .B(n7781), .ZN(n7784)
         );
  OAI21_X1 U9470 ( .B1(n7786), .B2(n7785), .A(n7784), .ZN(P2_U3260) );
  INV_X1 U9471 ( .A(n9819), .ZN(n7826) );
  AOI21_X1 U9472 ( .B1(n7788), .B2(n7787), .A(n9472), .ZN(n7789) );
  NAND2_X1 U9473 ( .A1(n7789), .A2(n4924), .ZN(n7794) );
  AOI21_X1 U9474 ( .B1(n9464), .B2(n9486), .A(n7790), .ZN(n7791) );
  OAI21_X1 U9475 ( .B1(n9483), .B2(n9467), .A(n7791), .ZN(n7792) );
  AOI21_X1 U9476 ( .B1(n5037), .B2(n9462), .A(n7792), .ZN(n7793) );
  OAI211_X1 U9477 ( .C1(n7826), .C2(n9456), .A(n7794), .B(n7793), .ZN(P1_U3234) );
  OR2_X1 U9478 ( .A1(n8872), .A2(n7795), .ZN(n8898) );
  XNOR2_X1 U9479 ( .A(n7797), .B(n7796), .ZN(n10209) );
  OAI22_X1 U9480 ( .A1(n8898), .A2(n10209), .B1(n8893), .B2(n10212), .ZN(n7810) );
  XNOR2_X1 U9481 ( .A(n7838), .B(n10212), .ZN(n10210) );
  NOR2_X1 U9482 ( .A1(n8891), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7798) );
  AOI21_X1 U9483 ( .B1(n8895), .B2(n10210), .A(n7798), .ZN(n7808) );
  NAND3_X1 U9484 ( .A1(n7841), .A2(n7802), .A3(n7801), .ZN(n7803) );
  NAND2_X1 U9485 ( .A1(n7953), .A2(n7803), .ZN(n7804) );
  NAND2_X1 U9486 ( .A1(n7804), .A2(n8886), .ZN(n7806) );
  AOI22_X1 U9487 ( .A1(n8815), .A2(n10146), .B1(n8534), .B2(n8816), .ZN(n7805)
         );
  OAI211_X1 U9488 ( .C1(n10209), .C2(n8913), .A(n7806), .B(n7805), .ZN(n10213)
         );
  NAND2_X1 U9489 ( .A1(n8393), .A2(n10213), .ZN(n7807) );
  OAI211_X1 U9490 ( .C1(n7290), .C2(n8393), .A(n7808), .B(n7807), .ZN(n7809)
         );
  OR2_X1 U9491 ( .A1(n7810), .A2(n7809), .ZN(P2_U3293) );
  XOR2_X1 U9492 ( .A(n7902), .B(n7818), .Z(n7822) );
  OAI22_X1 U9493 ( .A1(n7814), .A2(n10040), .B1(n9483), .B2(n10018), .ZN(n7821) );
  OR2_X1 U9494 ( .A1(n7815), .A2(n9486), .ZN(n7816) );
  NAND2_X1 U9495 ( .A1(n7817), .A2(n7816), .ZN(n7898) );
  XNOR2_X1 U9496 ( .A(n7898), .B(n7818), .ZN(n9823) );
  NOR2_X1 U9497 ( .A1(n9823), .A2(n7819), .ZN(n7820) );
  AOI211_X1 U9498 ( .C1(n7822), .C2(n10043), .A(n7821), .B(n7820), .ZN(n9822)
         );
  INV_X1 U9499 ( .A(n7904), .ZN(n7824) );
  AOI21_X1 U9500 ( .B1(n9819), .B2(n7823), .A(n7824), .ZN(n9820) );
  AOI22_X1 U9501 ( .A1(n10047), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n5037), .B2(
        n10009), .ZN(n7825) );
  OAI21_X1 U9502 ( .B1(n7826), .B2(n9710), .A(n7825), .ZN(n7828) );
  NOR2_X1 U9503 ( .A1(n9823), .A2(n8218), .ZN(n7827) );
  AOI211_X1 U9504 ( .C1(n9820), .C2(n10028), .A(n7828), .B(n7827), .ZN(n7829)
         );
  OAI21_X1 U9505 ( .B1(n9822), .B2(n10047), .A(n7829), .ZN(P1_U3280) );
  XNOR2_X1 U9506 ( .A(n7830), .B(n7831), .ZN(n7835) );
  NAND2_X1 U9507 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n8582) );
  OAI21_X1 U9508 ( .B1(n10161), .B2(n8892), .A(n8582), .ZN(n7833) );
  OAI22_X1 U9509 ( .A1(n8883), .A2(n10148), .B1(n10145), .B2(n8881), .ZN(n7832) );
  AOI211_X1 U9510 ( .C1(n10151), .C2(n10263), .A(n7833), .B(n7832), .ZN(n7834)
         );
  OAI21_X1 U9511 ( .B1(n7835), .B2(n8519), .A(n7834), .ZN(P2_U3219) );
  XNOR2_X1 U9512 ( .A(n7836), .B(n7843), .ZN(n10205) );
  NAND2_X1 U9513 ( .A1(n8144), .A2(n10201), .ZN(n7837) );
  AND2_X1 U9514 ( .A1(n7838), .A2(n7837), .ZN(n10202) );
  AOI22_X1 U9515 ( .A1(n8895), .A2(n10202), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n8864), .ZN(n7839) );
  OAI21_X1 U9516 ( .B1(n10205), .B2(n8850), .A(n7839), .ZN(n7840) );
  AOI21_X1 U9517 ( .B1(n8825), .B2(n10201), .A(n7840), .ZN(n7847) );
  OAI21_X1 U9518 ( .B1(n7843), .B2(n7842), .A(n7841), .ZN(n7844) );
  AOI222_X1 U9519 ( .A1(n8886), .A2(n7844), .B1(n8535), .B2(n8816), .C1(n4377), 
        .C2(n8815), .ZN(n10204) );
  MUX2_X1 U9520 ( .A(n10204), .B(n7845), .S(n8872), .Z(n7846) );
  NAND2_X1 U9521 ( .A1(n7847), .A2(n7846), .ZN(P2_U3294) );
  XNOR2_X1 U9522 ( .A(n7848), .B(n7851), .ZN(n7849) );
  AOI222_X1 U9523 ( .A1(n8886), .A2(n7849), .B1(n8532), .B2(n8816), .C1(n8534), 
        .C2(n8815), .ZN(n10227) );
  INV_X1 U9524 ( .A(n8850), .ZN(n8761) );
  XNOR2_X1 U9525 ( .A(n7851), .B(n7850), .ZN(n10230) );
  OR2_X1 U9526 ( .A1(n8872), .A2(n8620), .ZN(n8676) );
  INV_X1 U9527 ( .A(n8676), .ZN(n8807) );
  INV_X1 U9528 ( .A(n7853), .ZN(n7929) );
  AOI211_X1 U9529 ( .C1(n7854), .C2(n7949), .A(n10282), .B(n7929), .ZN(n10224)
         );
  OAI22_X1 U9530 ( .A1(n8393), .A2(n7293), .B1(n7855), .B2(n8891), .ZN(n7856)
         );
  AOI21_X1 U9531 ( .B1(n8807), .B2(n10224), .A(n7856), .ZN(n7857) );
  OAI21_X1 U9532 ( .B1(n10226), .B2(n8893), .A(n7857), .ZN(n7858) );
  AOI21_X1 U9533 ( .B1(n8761), .B2(n10230), .A(n7858), .ZN(n7859) );
  OAI21_X1 U9534 ( .B1(n8872), .B2(n10227), .A(n7859), .ZN(P2_U3291) );
  XNOR2_X1 U9535 ( .A(n8167), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n8164) );
  INV_X1 U9536 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7860) );
  XOR2_X1 U9537 ( .A(n8164), .B(n8165), .Z(n7873) );
  NAND2_X1 U9538 ( .A1(n9957), .A2(n8167), .ZN(n7864) );
  NAND2_X1 U9539 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8088) );
  NAND2_X1 U9540 ( .A1(n7864), .A2(n8088), .ZN(n7871) );
  NAND2_X1 U9541 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n8167), .ZN(n7867) );
  OAI21_X1 U9542 ( .B1(n8167), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7867), .ZN(
        n7868) );
  AOI211_X1 U9543 ( .C1(n7869), .C2(n7868), .A(n9950), .B(n8166), .ZN(n7870)
         );
  AOI211_X1 U9544 ( .C1(n9961), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n7871), .B(
        n7870), .ZN(n7872) );
  OAI21_X1 U9545 ( .B1(n9533), .B2(n7873), .A(n7872), .ZN(P1_U3254) );
  INV_X1 U9546 ( .A(n7874), .ZN(n7879) );
  OAI21_X1 U9547 ( .B1(n7876), .B2(n10119), .A(n7875), .ZN(n7878) );
  AOI211_X1 U9548 ( .C1(n10126), .C2(n7879), .A(n7878), .B(n7877), .ZN(n7882)
         );
  NAND2_X1 U9549 ( .A1(n10127), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7880) );
  OAI21_X1 U9550 ( .B1(n7882), .B2(n10127), .A(n7880), .ZN(P1_U3484) );
  NAND2_X1 U9551 ( .A1(n10141), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7881) );
  OAI21_X1 U9552 ( .B1(n7882), .B2(n10141), .A(n7881), .ZN(P1_U3533) );
  NAND2_X1 U9553 ( .A1(n7934), .A2(n7884), .ZN(n7885) );
  XNOR2_X1 U9554 ( .A(n7885), .B(n4381), .ZN(n7886) );
  AOI222_X1 U9555 ( .A1(n8886), .A2(n7886), .B1(n8530), .B2(n8816), .C1(n8532), 
        .C2(n8815), .ZN(n10241) );
  XNOR2_X1 U9556 ( .A(n7888), .B(n7887), .ZN(n10244) );
  NOR2_X1 U9557 ( .A1(n8891), .A2(n7889), .ZN(n7890) );
  AOI21_X1 U9558 ( .B1(n8872), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7890), .ZN(
        n7894) );
  NOR2_X1 U9559 ( .A1(n7927), .A2(n10239), .ZN(n7891) );
  OR2_X1 U9560 ( .A1(n8068), .A2(n7891), .ZN(n10240) );
  INV_X1 U9561 ( .A(n10240), .ZN(n7892) );
  NAND2_X1 U9562 ( .A1(n8895), .A2(n7892), .ZN(n7893) );
  OAI211_X1 U9563 ( .C1(n10239), .C2(n8893), .A(n7894), .B(n7893), .ZN(n7895)
         );
  AOI21_X1 U9564 ( .B1(n8761), .B2(n10244), .A(n7895), .ZN(n7896) );
  OAI21_X1 U9565 ( .B1(n10241), .B2(n8872), .A(n7896), .ZN(P2_U3289) );
  NAND2_X1 U9566 ( .A1(n7898), .A2(n7897), .ZN(n7900) );
  NAND2_X1 U9567 ( .A1(n7900), .A2(n7899), .ZN(n7979) );
  XNOR2_X1 U9568 ( .A(n7979), .B(n7978), .ZN(n9818) );
  OAI222_X1 U9569 ( .A1(n10040), .A2(n8000), .B1(n10018), .B2(n8048), .C1(
        n10014), .C2(n7903), .ZN(n9814) );
  INV_X1 U9570 ( .A(n9816), .ZN(n8005) );
  AOI211_X1 U9571 ( .C1(n9816), .C2(n7904), .A(n10121), .B(n7988), .ZN(n9815)
         );
  NAND2_X1 U9572 ( .A1(n9815), .A2(n9616), .ZN(n7906) );
  AOI22_X1 U9573 ( .A1(n10047), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8002), .B2(
        n10009), .ZN(n7905) );
  OAI211_X1 U9574 ( .C1(n8005), .C2(n9710), .A(n7906), .B(n7905), .ZN(n7907)
         );
  AOI21_X1 U9575 ( .B1(n9814), .B2(n10033), .A(n7907), .ZN(n7908) );
  OAI21_X1 U9576 ( .B1(n9818), .B2(n9722), .A(n7908), .ZN(P1_U3279) );
  INV_X1 U9577 ( .A(n7909), .ZN(n7916) );
  OAI222_X1 U9578 ( .A1(n8332), .A2(n7911), .B1(n7914), .B2(n7916), .C1(n7910), 
        .C2(P1_U3084), .ZN(P1_U3333) );
  INV_X1 U9579 ( .A(n7912), .ZN(n7942) );
  OAI222_X1 U9580 ( .A1(n8332), .A2(n7915), .B1(n7914), .B2(n7942), .C1(n7913), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  OAI222_X1 U9581 ( .A1(n9043), .A2(n7918), .B1(P2_U3152), .B2(n7917), .C1(
        n9036), .C2(n7916), .ZN(P2_U3338) );
  XNOR2_X1 U9582 ( .A(n7920), .B(n7919), .ZN(n7925) );
  OAI22_X1 U9583 ( .A1(n10161), .A2(n7971), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9161), .ZN(n7922) );
  OAI22_X1 U9584 ( .A1(n8854), .A2(n10145), .B1(n10148), .B2(n7967), .ZN(n7921) );
  AOI211_X1 U9585 ( .C1(n10151), .C2(n7923), .A(n7922), .B(n7921), .ZN(n7924)
         );
  OAI21_X1 U9586 ( .B1(n7925), .B2(n8519), .A(n7924), .ZN(P2_U3238) );
  XNOR2_X1 U9587 ( .A(n7926), .B(n7937), .ZN(n10232) );
  NOR2_X1 U9588 ( .A1(n8393), .A2(n7296), .ZN(n7932) );
  INV_X1 U9589 ( .A(n8895), .ZN(n8743) );
  INV_X1 U9590 ( .A(n7933), .ZN(n10233) );
  INV_X1 U9591 ( .A(n7927), .ZN(n7928) );
  OAI21_X1 U9592 ( .B1(n10233), .B2(n7929), .A(n7928), .ZN(n10234) );
  OAI22_X1 U9593 ( .A1(n8743), .A2(n10234), .B1(n7930), .B2(n8891), .ZN(n7931)
         );
  AOI211_X1 U9594 ( .C1(n8825), .C2(n7933), .A(n7932), .B(n7931), .ZN(n7941)
         );
  INV_X1 U9595 ( .A(n7934), .ZN(n7935) );
  AOI21_X1 U9596 ( .B1(n7937), .B2(n7936), .A(n7935), .ZN(n7938) );
  OAI222_X1 U9597 ( .A1(n8880), .A2(n7939), .B1(n8882), .B2(n7958), .C1(n8821), 
        .C2(n7938), .ZN(n10235) );
  NAND2_X1 U9598 ( .A1(n10235), .A2(n8393), .ZN(n7940) );
  OAI211_X1 U9599 ( .C1(n10232), .C2(n8850), .A(n7941), .B(n7940), .ZN(
        P2_U3290) );
  OAI222_X1 U9600 ( .A1(n9043), .A2(n7943), .B1(P2_U3152), .B2(n6374), .C1(
        n9036), .C2(n7942), .ZN(P2_U3337) );
  NAND2_X1 U9601 ( .A1(n7945), .A2(n7944), .ZN(n7946) );
  XOR2_X1 U9602 ( .A(n7954), .B(n7946), .Z(n10217) );
  OR2_X1 U9603 ( .A1(n7947), .A2(n10218), .ZN(n7948) );
  NAND2_X1 U9604 ( .A1(n7949), .A2(n7948), .ZN(n10219) );
  OAI22_X1 U9605 ( .A1(n8743), .A2(n10219), .B1(n7950), .B2(n8891), .ZN(n7951)
         );
  AOI21_X1 U9606 ( .B1(n8866), .B2(P2_REG2_REG_4__SCAN_IN), .A(n7951), .ZN(
        n7961) );
  NAND2_X1 U9607 ( .A1(n7953), .A2(n7952), .ZN(n7955) );
  XNOR2_X1 U9608 ( .A(n7955), .B(n7954), .ZN(n7956) );
  OAI222_X1 U9609 ( .A1(n8880), .A2(n7958), .B1(n8882), .B2(n7957), .C1(n7956), 
        .C2(n8821), .ZN(n10220) );
  AOI22_X1 U9610 ( .A1(n8825), .A2(n7959), .B1(n8393), .B2(n10220), .ZN(n7960)
         );
  OAI211_X1 U9611 ( .C1(n10217), .C2(n8850), .A(n7961), .B(n7960), .ZN(
        P2_U3292) );
  OAI21_X1 U9612 ( .B1(n7963), .B2(n7964), .A(n7962), .ZN(n10273) );
  XOR2_X1 U9613 ( .A(n7965), .B(n7964), .Z(n7966) );
  OAI222_X1 U9614 ( .A1(n8882), .A2(n7967), .B1(n8880), .B2(n8854), .C1(n8821), 
        .C2(n7966), .ZN(n10276) );
  INV_X1 U9615 ( .A(n10276), .ZN(n7968) );
  MUX2_X1 U9616 ( .A(n7969), .B(n7968), .S(n8393), .Z(n7975) );
  NOR2_X1 U9617 ( .A1(n8889), .A2(n10274), .ZN(n7970) );
  OR2_X1 U9618 ( .A1(n8130), .A2(n7970), .ZN(n10275) );
  INV_X1 U9619 ( .A(n10275), .ZN(n7973) );
  OAI22_X1 U9620 ( .A1(n8893), .A2(n10274), .B1(n8891), .B2(n7971), .ZN(n7972)
         );
  AOI21_X1 U9621 ( .B1(n7973), .B2(n8895), .A(n7972), .ZN(n7974) );
  OAI211_X1 U9622 ( .C1(n8850), .C2(n10273), .A(n7975), .B(n7974), .ZN(
        P2_U3285) );
  INV_X1 U9623 ( .A(n7976), .ZN(n8243) );
  OAI222_X1 U9624 ( .A1(n8332), .A2(n7977), .B1(n7914), .B2(n8243), .C1(
        P1_U3084), .C2(n6716), .ZN(P1_U3331) );
  INV_X1 U9625 ( .A(n8044), .ZN(n7980) );
  XNOR2_X1 U9626 ( .A(n8038), .B(n7980), .ZN(n9808) );
  NAND2_X1 U9627 ( .A1(n9808), .A2(n10034), .ZN(n7987) );
  INV_X1 U9628 ( .A(n7981), .ZN(n7982) );
  XNOR2_X1 U9629 ( .A(n8045), .B(n8044), .ZN(n7985) );
  OAI22_X1 U9630 ( .A1(n9483), .A2(n10040), .B1(n8189), .B2(n10018), .ZN(n7984) );
  AOI21_X1 U9631 ( .B1(n7985), .B2(n10043), .A(n7984), .ZN(n7986) );
  NAND2_X1 U9632 ( .A1(n7987), .A2(n7986), .ZN(n9812) );
  INV_X1 U9633 ( .A(n9812), .ZN(n7994) );
  NOR2_X1 U9634 ( .A1(n7988), .A2(n9809), .ZN(n7989) );
  OR2_X1 U9635 ( .A1(n8040), .A2(n7989), .ZN(n9810) );
  AOI22_X1 U9636 ( .A1(n10047), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8092), .B2(
        n10009), .ZN(n7991) );
  NAND2_X1 U9637 ( .A1(n8036), .A2(n10050), .ZN(n7990) );
  OAI211_X1 U9638 ( .C1(n9810), .C2(n9573), .A(n7991), .B(n7990), .ZN(n7992)
         );
  AOI21_X1 U9639 ( .B1(n9808), .B2(n10029), .A(n7992), .ZN(n7993) );
  OAI21_X1 U9640 ( .B1(n7994), .B2(n10047), .A(n7993), .ZN(P1_U3278) );
  OAI21_X1 U9641 ( .B1(n7996), .B2(n4469), .A(n7995), .ZN(n7997) );
  NAND2_X1 U9642 ( .A1(n7997), .A2(n9448), .ZN(n8004) );
  INV_X1 U9643 ( .A(n8048), .ZN(n9482) );
  NAND2_X1 U9644 ( .A1(n9440), .A2(n9482), .ZN(n7999) );
  OAI211_X1 U9645 ( .C1(n8000), .C2(n9451), .A(n7999), .B(n7998), .ZN(n8001)
         );
  AOI21_X1 U9646 ( .B1(n8002), .B2(n9462), .A(n8001), .ZN(n8003) );
  OAI211_X1 U9647 ( .C1(n8005), .C2(n9456), .A(n8004), .B(n8003), .ZN(P1_U3222) );
  NAND2_X1 U9648 ( .A1(n4506), .A2(n8006), .ZN(n8011) );
  INV_X1 U9649 ( .A(n8008), .ZN(n8009) );
  AOI21_X1 U9650 ( .B1(n8011), .B2(n8010), .A(n8009), .ZN(n8016) );
  OAI21_X1 U9651 ( .B1(n10161), .B2(n8132), .A(n8012), .ZN(n8014) );
  OAI22_X1 U9652 ( .A1(n8401), .A2(n10145), .B1(n10148), .B2(n8881), .ZN(n8013) );
  AOI211_X1 U9653 ( .C1(n10151), .C2(n8134), .A(n8014), .B(n8013), .ZN(n8015)
         );
  OAI21_X1 U9654 ( .B1(n8016), .B2(n8519), .A(n8015), .ZN(P2_U3226) );
  INV_X1 U9655 ( .A(n8054), .ZN(n8019) );
  AOI21_X1 U9656 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9852), .A(n8017), .ZN(
        n8018) );
  OAI21_X1 U9657 ( .B1(n8019), .B2(n7914), .A(n8018), .ZN(P1_U3330) );
  NAND2_X1 U9658 ( .A1(n8031), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8022) );
  MUX2_X1 U9659 ( .A(n6131), .B(P2_REG2_REG_17__SCAN_IN), .S(n8598), .Z(n8023)
         );
  INV_X1 U9660 ( .A(n8023), .ZN(n8024) );
  OAI211_X1 U9661 ( .C1(n8025), .C2(n8024), .A(n10163), .B(n8593), .ZN(n8028)
         );
  NAND2_X1 U9662 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8462) );
  INV_X1 U9663 ( .A(n8462), .ZN(n8026) );
  AOI21_X1 U9664 ( .B1(n10164), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8026), .ZN(
        n8027) );
  OAI211_X1 U9665 ( .C1(n10166), .C2(n8029), .A(n8028), .B(n8027), .ZN(n8035)
         );
  OAI21_X1 U9666 ( .B1(n8031), .B2(P2_REG1_REG_16__SCAN_IN), .A(n8030), .ZN(
        n8033) );
  XNOR2_X1 U9667 ( .A(n8598), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8032) );
  NOR2_X1 U9668 ( .A1(n8032), .A2(n8033), .ZN(n8597) );
  AOI211_X1 U9669 ( .C1(n8033), .C2(n8032), .A(n8597), .B(n10167), .ZN(n8034)
         );
  OR2_X1 U9670 ( .A1(n8035), .A2(n8034), .ZN(P2_U3262) );
  NAND2_X1 U9671 ( .A1(n9809), .A2(n8048), .ZN(n8037) );
  XNOR2_X1 U9672 ( .A(n8191), .B(n8039), .ZN(n9807) );
  INV_X1 U9673 ( .A(n8040), .ZN(n8041) );
  AOI211_X1 U9674 ( .C1(n9804), .C2(n8041), .A(n10121), .B(n4969), .ZN(n9803)
         );
  AOI22_X1 U9675 ( .A1(n10047), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8181), .B2(
        n10009), .ZN(n8042) );
  OAI21_X1 U9676 ( .B1(n8188), .B2(n9710), .A(n8042), .ZN(n8052) );
  AOI21_X1 U9677 ( .B1(n8046), .B2(n8047), .A(n10014), .ZN(n8050) );
  OAI22_X1 U9678 ( .A1(n8048), .A2(n10040), .B1(n9384), .B2(n10018), .ZN(n8049) );
  AOI21_X1 U9679 ( .B1(n8050), .B2(n8200), .A(n8049), .ZN(n9806) );
  NOR2_X1 U9680 ( .A1(n9806), .A2(n10047), .ZN(n8051) );
  AOI211_X1 U9681 ( .C1(n9803), .C2(n9616), .A(n8052), .B(n8051), .ZN(n8053)
         );
  OAI21_X1 U9682 ( .B1(n9722), .B2(n9807), .A(n8053), .ZN(P1_U3277) );
  NAND2_X1 U9683 ( .A1(n8054), .A2(n9321), .ZN(n8056) );
  OAI211_X1 U9684 ( .C1(n8057), .C2(n9043), .A(n8056), .B(n8055), .ZN(P2_U3335) );
  XNOR2_X1 U9685 ( .A(n8058), .B(n8063), .ZN(n10250) );
  NAND2_X1 U9686 ( .A1(n8060), .A2(n8059), .ZN(n8062) );
  INV_X1 U9687 ( .A(n8062), .ZN(n8064) );
  INV_X1 U9688 ( .A(n8063), .ZN(n8061) );
  OR2_X1 U9689 ( .A1(n8062), .A2(n8061), .ZN(n8106) );
  OAI21_X1 U9690 ( .B1(n8064), .B2(n8063), .A(n8106), .ZN(n8066) );
  AOI21_X1 U9691 ( .B1(n8066), .B2(n8886), .A(n8065), .ZN(n10249) );
  MUX2_X1 U9692 ( .A(n10249), .B(n8067), .S(n8866), .Z(n8073) );
  XNOR2_X1 U9693 ( .A(n8068), .B(n4840), .ZN(n10247) );
  OAI22_X1 U9694 ( .A1(n8893), .A2(n8070), .B1(n8891), .B2(n8069), .ZN(n8071)
         );
  AOI21_X1 U9695 ( .B1(n8895), .B2(n10247), .A(n8071), .ZN(n8072) );
  OAI211_X1 U9696 ( .C1(n10250), .C2(n8850), .A(n8073), .B(n8072), .ZN(
        P2_U3288) );
  INV_X1 U9697 ( .A(n8074), .ZN(n8075) );
  AOI21_X1 U9698 ( .B1(n8077), .B2(n8076), .A(n8075), .ZN(n9001) );
  XNOR2_X1 U9699 ( .A(n8078), .B(n8077), .ZN(n8079) );
  AOI222_X1 U9700 ( .A1(n8886), .A2(n8079), .B1(n8814), .B2(n8816), .C1(n8525), 
        .C2(n8815), .ZN(n9000) );
  MUX2_X1 U9701 ( .A(n9240), .B(n9000), .S(n8393), .Z(n8083) );
  AOI21_X1 U9702 ( .B1(n8997), .B2(n8080), .A(n8842), .ZN(n8998) );
  INV_X1 U9703 ( .A(n8997), .ZN(n8407) );
  OAI22_X1 U9704 ( .A1(n8407), .A2(n8893), .B1(n8400), .B2(n8891), .ZN(n8081)
         );
  AOI21_X1 U9705 ( .B1(n8998), .B2(n8895), .A(n8081), .ZN(n8082) );
  OAI211_X1 U9706 ( .C1(n9001), .C2(n8850), .A(n8083), .B(n8082), .ZN(P2_U3282) );
  XNOR2_X1 U9707 ( .A(n8085), .B(n8084), .ZN(n8086) );
  XNOR2_X1 U9708 ( .A(n8087), .B(n8086), .ZN(n8094) );
  INV_X1 U9709 ( .A(n8189), .ZN(n9481) );
  NAND2_X1 U9710 ( .A1(n9440), .A2(n9481), .ZN(n8089) );
  OAI211_X1 U9711 ( .C1(n9483), .C2(n9451), .A(n8089), .B(n8088), .ZN(n8091)
         );
  NOR2_X1 U9712 ( .A1(n9809), .A2(n9456), .ZN(n8090) );
  AOI211_X1 U9713 ( .C1(n8092), .C2(n9462), .A(n8091), .B(n8090), .ZN(n8093)
         );
  OAI21_X1 U9714 ( .B1(n8094), .B2(n9472), .A(n8093), .ZN(P1_U3232) );
  XNOR2_X1 U9715 ( .A(n8096), .B(n8095), .ZN(n8100) );
  OAI22_X1 U9716 ( .A1(n10161), .A2(n8863), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7470), .ZN(n8098) );
  OAI22_X1 U9717 ( .A1(n8854), .A2(n10148), .B1(n10145), .B2(n8853), .ZN(n8097) );
  AOI211_X1 U9718 ( .C1(n10151), .C2(n9002), .A(n8098), .B(n8097), .ZN(n8099)
         );
  OAI21_X1 U9719 ( .B1(n8100), .B2(n8519), .A(n8099), .ZN(P2_U3236) );
  OR2_X1 U9720 ( .A1(n8101), .A2(n8102), .ZN(n8874) );
  NAND2_X1 U9721 ( .A1(n8101), .A2(n8102), .ZN(n8103) );
  NAND2_X1 U9722 ( .A1(n8874), .A2(n8103), .ZN(n10260) );
  INV_X1 U9723 ( .A(n10260), .ZN(n8119) );
  NAND3_X1 U9724 ( .A1(n8106), .A2(n8105), .A3(n8104), .ZN(n8107) );
  AND2_X1 U9725 ( .A1(n8877), .A2(n8107), .ZN(n8110) );
  INV_X1 U9726 ( .A(n8913), .ZN(n10253) );
  NAND2_X1 U9727 ( .A1(n10260), .A2(n10253), .ZN(n8109) );
  AOI22_X1 U9728 ( .A1(n8815), .A2(n8530), .B1(n8528), .B2(n8816), .ZN(n8108)
         );
  OAI211_X1 U9729 ( .C1(n8821), .C2(n8110), .A(n8109), .B(n8108), .ZN(n10258)
         );
  MUX2_X1 U9730 ( .A(n10258), .B(P2_REG2_REG_9__SCAN_IN), .S(n8866), .Z(n8111)
         );
  INV_X1 U9731 ( .A(n8111), .ZN(n8118) );
  INV_X1 U9732 ( .A(n8890), .ZN(n8112) );
  AOI21_X1 U9733 ( .B1(n8114), .B2(n8113), .A(n8112), .ZN(n10255) );
  INV_X1 U9734 ( .A(n8114), .ZN(n10256) );
  OAI22_X1 U9735 ( .A1(n8893), .A2(n10256), .B1(n8891), .B2(n8115), .ZN(n8116)
         );
  AOI21_X1 U9736 ( .B1(n8895), .B2(n10255), .A(n8116), .ZN(n8117) );
  OAI211_X1 U9737 ( .C1(n8119), .C2(n8898), .A(n8118), .B(n8117), .ZN(P2_U3287) );
  NAND2_X1 U9738 ( .A1(n8147), .A2(n8120), .ZN(n8121) );
  INV_X1 U9739 ( .A(n8121), .ZN(n10189) );
  AOI22_X1 U9740 ( .A1(n8121), .A2(n8886), .B1(n8816), .B2(n4376), .ZN(n10187)
         );
  INV_X1 U9741 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n8122) );
  OAI22_X1 U9742 ( .A1(n8866), .A2(n10187), .B1(n8122), .B2(n8891), .ZN(n8123)
         );
  AOI21_X1 U9743 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n8872), .A(n8123), .ZN(
        n8126) );
  OAI21_X1 U9744 ( .B1(n8825), .B2(n8895), .A(n8124), .ZN(n8125) );
  OAI211_X1 U9745 ( .C1(n10189), .C2(n8850), .A(n8126), .B(n8125), .ZN(
        P2_U3296) );
  INV_X1 U9746 ( .A(n8127), .ZN(n8129) );
  INV_X1 U9747 ( .A(n8128), .ZN(n8138) );
  OAI21_X1 U9748 ( .B1(n8129), .B2(n8128), .A(n8856), .ZN(n10286) );
  OR2_X1 U9749 ( .A1(n8130), .A2(n10281), .ZN(n8131) );
  NAND2_X1 U9750 ( .A1(n8862), .A2(n8131), .ZN(n10283) );
  INV_X1 U9751 ( .A(n8132), .ZN(n8133) );
  AOI22_X1 U9752 ( .A1(n8825), .A2(n8134), .B1(n8864), .B2(n8133), .ZN(n8135)
         );
  OAI21_X1 U9753 ( .B1(n10283), .B2(n8743), .A(n8135), .ZN(n8142) );
  NAND2_X1 U9754 ( .A1(n8136), .A2(n8137), .ZN(n8139) );
  XNOR2_X1 U9755 ( .A(n8139), .B(n8138), .ZN(n8140) );
  OAI222_X1 U9756 ( .A1(n8882), .A2(n8881), .B1(n8880), .B2(n8401), .C1(n8821), 
        .C2(n8140), .ZN(n10284) );
  MUX2_X1 U9757 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n10284), .S(n8393), .Z(n8141) );
  AOI211_X1 U9758 ( .C1(n8761), .C2(n10286), .A(n8142), .B(n8141), .ZN(n8143)
         );
  INV_X1 U9759 ( .A(n8143), .ZN(P2_U3284) );
  OAI21_X1 U9760 ( .B1(n10188), .B2(n10194), .A(n8144), .ZN(n10195) );
  INV_X1 U9761 ( .A(n8145), .ZN(n8150) );
  NAND2_X1 U9762 ( .A1(n8146), .A2(n8145), .ZN(n8156) );
  INV_X1 U9763 ( .A(n8147), .ZN(n8148) );
  NAND2_X1 U9764 ( .A1(n8156), .A2(n8148), .ZN(n8149) );
  OAI211_X1 U9765 ( .C1(n8151), .C2(n8150), .A(n8886), .B(n8149), .ZN(n8153)
         );
  AND2_X1 U9766 ( .A1(n8153), .A2(n8152), .ZN(n10196) );
  MUX2_X1 U9767 ( .A(n10196), .B(n9163), .S(n8866), .Z(n8155) );
  INV_X1 U9768 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9225) );
  NAND2_X1 U9769 ( .A1(n8864), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8154) );
  OAI211_X1 U9770 ( .C1(n8743), .C2(n10195), .A(n8155), .B(n8154), .ZN(n8158)
         );
  XOR2_X1 U9771 ( .A(n6571), .B(n8156), .Z(n10193) );
  OAI22_X1 U9772 ( .A1(n10194), .A2(n8893), .B1(n8850), .B2(n10193), .ZN(n8157) );
  OR2_X1 U9773 ( .A1(n8158), .A2(n8157), .ZN(P2_U3295) );
  INV_X1 U9774 ( .A(n8159), .ZN(n8162) );
  OAI222_X1 U9775 ( .A1(P2_U3152), .A2(n8160), .B1(n9036), .B2(n8162), .C1(
        n9291), .C2(n9043), .ZN(P2_U3334) );
  INV_X1 U9776 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8161) );
  OAI222_X1 U9777 ( .A1(P1_U3084), .A2(n8163), .B1(n7914), .B2(n8162), .C1(
        n8161), .C2(n8332), .ZN(P1_U3329) );
  XNOR2_X1 U9778 ( .A(n8256), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n8257) );
  XNOR2_X1 U9779 ( .A(n8255), .B(n8257), .ZN(n8176) );
  INV_X1 U9780 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8170) );
  AOI211_X1 U9781 ( .C1(n8170), .C2(n8169), .A(n9950), .B(n8245), .ZN(n8171)
         );
  INV_X1 U9782 ( .A(n8171), .ZN(n8175) );
  INV_X1 U9783 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9134) );
  NOR2_X1 U9784 ( .A1(n9134), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8182) );
  NOR2_X1 U9785 ( .A1(n4632), .A2(n8172), .ZN(n8173) );
  AOI211_X1 U9786 ( .C1(n9961), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n8182), .B(
        n8173), .ZN(n8174) );
  OAI211_X1 U9787 ( .C1(n9533), .C2(n8176), .A(n8175), .B(n8174), .ZN(P1_U3255) );
  XNOR2_X1 U9788 ( .A(n8179), .B(n8178), .ZN(n8180) );
  XNOR2_X1 U9789 ( .A(n8177), .B(n8180), .ZN(n8187) );
  NAND2_X1 U9790 ( .A1(n9462), .A2(n8181), .ZN(n8184) );
  AOI21_X1 U9791 ( .B1(n9464), .B2(n9482), .A(n8182), .ZN(n8183) );
  OAI211_X1 U9792 ( .C1(n9384), .C2(n9467), .A(n8184), .B(n8183), .ZN(n8185)
         );
  AOI21_X1 U9793 ( .B1(n9804), .B2(n9470), .A(n8185), .ZN(n8186) );
  OAI21_X1 U9794 ( .B1(n8187), .B2(n9472), .A(n8186), .ZN(P1_U3213) );
  INV_X1 U9795 ( .A(n9384), .ZN(n9480) );
  NAND2_X1 U9796 ( .A1(n9804), .A2(n9481), .ZN(n8190) );
  XNOR2_X1 U9797 ( .A(n8230), .B(n8229), .ZN(n9797) );
  NAND2_X1 U9798 ( .A1(n9795), .A2(n8213), .ZN(n8195) );
  NOR2_X1 U9799 ( .A1(n8228), .A2(n9710), .ZN(n8198) );
  INV_X1 U9800 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8196) );
  OAI22_X1 U9801 ( .A1(n10033), .A2(n8196), .B1(n9387), .B2(n10031), .ZN(n8197) );
  AOI211_X1 U9802 ( .C1(n9794), .C2(n9616), .A(n8198), .B(n8197), .ZN(n8206)
         );
  NAND2_X1 U9803 ( .A1(n8237), .A2(n8202), .ZN(n8203) );
  XNOR2_X1 U9804 ( .A(n8203), .B(n8229), .ZN(n8204) );
  OAI222_X1 U9805 ( .A1(n10040), .A2(n9384), .B1(n10018), .B2(n9436), .C1(
        n10014), .C2(n8204), .ZN(n9793) );
  NAND2_X1 U9806 ( .A1(n9793), .A2(n10033), .ZN(n8205) );
  OAI211_X1 U9807 ( .C1(n9797), .C2(n9722), .A(n8206), .B(n8205), .ZN(P1_U3275) );
  XOR2_X1 U9808 ( .A(n8207), .B(n8209), .Z(n8217) );
  XNOR2_X1 U9809 ( .A(n8208), .B(n8209), .ZN(n8211) );
  AOI22_X1 U9810 ( .A1(n9481), .A2(n9715), .B1(n10037), .B2(n9479), .ZN(n8210)
         );
  OAI21_X1 U9811 ( .B1(n8211), .B2(n10014), .A(n8210), .ZN(n8212) );
  AOI21_X1 U9812 ( .B1(n8217), .B2(n10034), .A(n8212), .ZN(n9801) );
  AOI21_X1 U9813 ( .B1(n9798), .B2(n8214), .A(n8194), .ZN(n9799) );
  AOI22_X1 U9814 ( .A1(n10047), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9461), .B2(
        n10009), .ZN(n8215) );
  OAI21_X1 U9815 ( .B1(n8216), .B2(n9710), .A(n8215), .ZN(n8220) );
  INV_X1 U9816 ( .A(n8217), .ZN(n9802) );
  NOR2_X1 U9817 ( .A1(n9802), .A2(n8218), .ZN(n8219) );
  AOI211_X1 U9818 ( .C1(n9799), .C2(n10028), .A(n8220), .B(n8219), .ZN(n8221)
         );
  OAI21_X1 U9819 ( .B1(n10047), .B2(n9801), .A(n8221), .ZN(P1_U3276) );
  INV_X1 U9820 ( .A(n8222), .ZN(n8226) );
  OAI222_X1 U9821 ( .A1(n8332), .A2(n8224), .B1(n7914), .B2(n8226), .C1(
        P1_U3084), .C2(n8223), .ZN(P1_U3328) );
  OAI222_X1 U9822 ( .A1(n9043), .A2(n8227), .B1(n9036), .B2(n8226), .C1(
        P2_U3152), .C2(n8225), .ZN(P2_U3333) );
  XNOR2_X1 U9823 ( .A(n8267), .B(n8238), .ZN(n9792) );
  AOI211_X1 U9824 ( .C1(n9790), .C2(n8231), .A(n10121), .B(n8287), .ZN(n9789)
         );
  INV_X1 U9825 ( .A(n9790), .ZN(n8268) );
  NOR2_X1 U9826 ( .A1(n8268), .A2(n9710), .ZN(n8234) );
  INV_X1 U9827 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8232) );
  OAI22_X1 U9828 ( .A1(n10033), .A2(n8232), .B1(n9395), .B2(n10031), .ZN(n8233) );
  AOI211_X1 U9829 ( .C1(n9789), .C2(n9616), .A(n8234), .B(n8233), .ZN(n8242)
         );
  AOI21_X1 U9830 ( .B1(n8237), .B2(n8236), .A(n8235), .ZN(n8291) );
  XOR2_X1 U9831 ( .A(n8238), .B(n8291), .Z(n8239) );
  OAI222_X1 U9832 ( .A1(n10018), .A2(n8240), .B1(n10040), .B2(n9468), .C1(
        n8239), .C2(n10014), .ZN(n9788) );
  NAND2_X1 U9833 ( .A1(n9788), .A2(n10033), .ZN(n8241) );
  OAI211_X1 U9834 ( .C1(n9792), .C2(n9722), .A(n8242), .B(n8241), .ZN(P1_U3274) );
  OAI222_X1 U9835 ( .A1(n9043), .A2(n8244), .B1(n9036), .B2(n8243), .C1(n6373), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  NOR2_X1 U9836 ( .A1(n8247), .A2(n9505), .ZN(n8248) );
  XNOR2_X1 U9837 ( .A(n8247), .B(n9505), .ZN(n9508) );
  INV_X1 U9838 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9507) );
  NOR2_X1 U9839 ( .A1(n9508), .A2(n9507), .ZN(n9506) );
  NAND2_X1 U9840 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9522), .ZN(n8249) );
  OAI21_X1 U9841 ( .B1(n9522), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8249), .ZN(
        n9516) );
  NAND2_X1 U9842 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9532), .ZN(n8250) );
  OAI21_X1 U9843 ( .B1(n9532), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8250), .ZN(
        n9528) );
  AND2_X1 U9844 ( .A1(n9532), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8251) );
  NAND2_X1 U9845 ( .A1(n9956), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8252) );
  OAI21_X1 U9846 ( .B1(n9956), .B2(P1_REG2_REG_18__SCAN_IN), .A(n8252), .ZN(
        n9952) );
  XNOR2_X1 U9847 ( .A(n8253), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n8264) );
  INV_X1 U9848 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9237) );
  AOI22_X1 U9849 ( .A1(n9956), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9237), .B2(
        n8254), .ZN(n9960) );
  INV_X1 U9850 ( .A(n8255), .ZN(n8258) );
  NOR2_X1 U9851 ( .A1(n9505), .A2(n8259), .ZN(n8260) );
  INV_X1 U9852 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9279) );
  XNOR2_X1 U9853 ( .A(n8259), .B(n9505), .ZN(n9501) );
  NOR2_X1 U9854 ( .A1(n9279), .A2(n9501), .ZN(n9502) );
  NOR2_X1 U9855 ( .A1(n8260), .A2(n9502), .ZN(n9520) );
  XNOR2_X1 U9856 ( .A(n9522), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9519) );
  XNOR2_X1 U9857 ( .A(n9532), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9535) );
  NAND2_X1 U9858 ( .A1(n9960), .A2(n9959), .ZN(n9958) );
  OAI21_X1 U9859 ( .B1(n9956), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9958), .ZN(
        n8261) );
  XNOR2_X1 U9860 ( .A(n8261), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8262) );
  AOI22_X1 U9861 ( .A1(n8264), .A2(n9932), .B1(n9962), .B2(n8262), .ZN(n8265)
         );
  NAND2_X1 U9862 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9348) );
  NOR2_X1 U9863 ( .A1(n9790), .A2(n9716), .ZN(n8269) );
  INV_X1 U9864 ( .A(n9778), .ZN(n9692) );
  NAND2_X1 U9865 ( .A1(n9662), .A2(n9664), .ZN(n8274) );
  NOR2_X1 U9866 ( .A1(n9654), .A2(n9667), .ZN(n8275) );
  INV_X1 U9867 ( .A(n9667), .ZN(n9477) );
  INV_X1 U9868 ( .A(n9625), .ZN(n9475) );
  NAND2_X1 U9869 ( .A1(n8277), .A2(n9625), .ZN(n8278) );
  NOR2_X1 U9870 ( .A1(n9743), .A2(n9474), .ZN(n8280) );
  INV_X1 U9871 ( .A(n9743), .ZN(n9598) );
  NOR2_X1 U9872 ( .A1(n9590), .A2(n8307), .ZN(n8282) );
  NAND2_X1 U9873 ( .A1(n9587), .A2(n9602), .ZN(n8283) );
  INV_X1 U9874 ( .A(n8283), .ZN(n8281) );
  NOR2_X1 U9875 ( .A1(n8282), .A2(n8281), .ZN(n8286) );
  INV_X1 U9876 ( .A(n9783), .ZN(n9711) );
  OAI21_X1 U9877 ( .B1(n4972), .B2(n4391), .A(n5035), .ZN(n9574) );
  OAI22_X1 U9878 ( .A1(n9574), .A2(n10121), .B1(n4972), .B2(n10119), .ZN(n8288) );
  INV_X1 U9879 ( .A(n8288), .ZN(n8318) );
  NAND2_X1 U9880 ( .A1(n9713), .A2(n9714), .ZN(n9712) );
  NAND2_X1 U9881 ( .A1(n9712), .A2(n8292), .ZN(n9694) );
  INV_X1 U9882 ( .A(n8302), .ZN(n8304) );
  INV_X1 U9883 ( .A(n8305), .ZN(n8306) );
  OR2_X1 U9884 ( .A1(n8310), .A2(n8309), .ZN(n8311) );
  NAND2_X1 U9885 ( .A1(n9551), .A2(n8311), .ZN(n8312) );
  NAND2_X1 U9886 ( .A1(n8312), .A2(n10043), .ZN(n8316) );
  OR2_X1 U9887 ( .A1(n9602), .A2(n10040), .ZN(n8314) );
  AND2_X1 U9888 ( .A1(n8314), .A2(n5029), .ZN(n8315) );
  NAND2_X1 U9889 ( .A1(n8316), .A2(n8315), .ZN(n9567) );
  INV_X1 U9890 ( .A(n9567), .ZN(n8317) );
  MUX2_X1 U9891 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n8319), .S(n10129), .Z(
        P1_U3519) );
  MUX2_X1 U9892 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n8319), .S(n10143), .Z(
        P1_U3551) );
  NAND2_X1 U9893 ( .A1(n9542), .A2(n9560), .ZN(n9541) );
  INV_X1 U9894 ( .A(n9920), .ZN(n8320) );
  AND2_X1 U9895 ( .A1(n8320), .A2(P1_B_REG_SCAN_IN), .ZN(n8321) );
  NOR2_X1 U9896 ( .A1(n10018), .A2(n8321), .ZN(n9555) );
  NAND2_X1 U9897 ( .A1(n9555), .A2(n8322), .ZN(n9728) );
  NOR2_X1 U9898 ( .A1(n10047), .A2(n9728), .ZN(n9544) );
  NOR2_X1 U9899 ( .A1(n8323), .A2(n9710), .ZN(n8324) );
  AOI211_X1 U9900 ( .C1(n10047), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9544), .B(
        n8324), .ZN(n8325) );
  OAI21_X1 U9901 ( .B1(n9725), .B2(n9573), .A(n8325), .ZN(P1_U3261) );
  INV_X1 U9902 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8328) );
  INV_X1 U9903 ( .A(n8326), .ZN(n9035) );
  OAI222_X1 U9904 ( .A1(n8332), .A2(n8328), .B1(n7914), .B2(n9035), .C1(n8327), 
        .C2(P1_U3084), .ZN(P1_U3323) );
  INV_X1 U9905 ( .A(n8329), .ZN(n9037) );
  OAI222_X1 U9906 ( .A1(n8332), .A2(n8331), .B1(n7914), .B2(n9037), .C1(n8330), 
        .C2(P1_U3084), .ZN(P1_U3324) );
  OAI21_X1 U9907 ( .B1(n8335), .B2(n8334), .A(n8333), .ZN(n8336) );
  NAND2_X1 U9908 ( .A1(n8336), .A2(n9448), .ZN(n8340) );
  OAI22_X1 U9909 ( .A1(n5313), .A2(n9451), .B1(n9467), .B2(n10041), .ZN(n8337)
         );
  AOI21_X1 U9910 ( .B1(n8338), .B2(P1_REG3_REG_2__SCAN_IN), .A(n8337), .ZN(
        n8339) );
  OAI211_X1 U9911 ( .C1(n10069), .C2(n9456), .A(n8340), .B(n8339), .ZN(
        P1_U3235) );
  INV_X1 U9912 ( .A(n8341), .ZN(n9850) );
  OAI222_X1 U9913 ( .A1(n9043), .A2(n8342), .B1(P2_U3152), .B2(n6363), .C1(
        n9036), .C2(n9850), .ZN(P2_U3330) );
  AOI21_X1 U9914 ( .B1(n8344), .B2(n8343), .A(n9472), .ZN(n8346) );
  NAND2_X1 U9915 ( .A1(n8346), .A2(n8345), .ZN(n8350) );
  NAND2_X1 U9916 ( .A1(n9440), .A2(n10038), .ZN(n8347) );
  NAND2_X1 U9917 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9942) );
  OAI211_X1 U9918 ( .C1(n10041), .C2(n9451), .A(n8347), .B(n9942), .ZN(n8348)
         );
  AOI21_X1 U9919 ( .B1(n10030), .B2(n9462), .A(n8348), .ZN(n8349) );
  OAI211_X1 U9920 ( .C1(n10082), .C2(n9456), .A(n8350), .B(n8349), .ZN(
        P1_U3228) );
  NAND2_X1 U9921 ( .A1(n8919), .A2(n10280), .ZN(n8357) );
  NAND2_X1 U9922 ( .A1(n8635), .A2(n4384), .ZN(n8353) );
  XNOR2_X1 U9923 ( .A(n8353), .B(n8352), .ZN(n8356) );
  MUX2_X1 U9924 ( .A(n8919), .B(n8357), .S(n8356), .Z(n8355) );
  NAND2_X1 U9925 ( .A1(n8919), .A2(n10151), .ZN(n8354) );
  NAND2_X1 U9926 ( .A1(n8354), .A2(n8519), .ZN(n8359) );
  INV_X1 U9927 ( .A(n8372), .ZN(n8375) );
  MUX2_X1 U9928 ( .A(n8357), .B(n8919), .S(n8356), .Z(n8358) );
  INV_X1 U9929 ( .A(n8358), .ZN(n8362) );
  INV_X1 U9930 ( .A(n8371), .ZN(n8360) );
  NAND2_X1 U9931 ( .A1(n8360), .A2(n8359), .ZN(n8361) );
  INV_X1 U9932 ( .A(n8364), .ZN(n8366) );
  OAI22_X1 U9933 ( .A1(n8366), .A2(n10161), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8365), .ZN(n8370) );
  OAI22_X1 U9934 ( .A1(n8368), .A2(n10145), .B1(n8367), .B2(n10148), .ZN(n8369) );
  AOI211_X1 U9935 ( .C1(n8372), .C2(n8371), .A(n8370), .B(n8369), .ZN(n8373)
         );
  OAI211_X1 U9936 ( .C1(n8376), .C2(n8375), .A(n8374), .B(n8373), .ZN(P2_U3222) );
  OR2_X1 U9937 ( .A1(n8380), .A2(n4452), .ZN(n8382) );
  AOI21_X1 U9938 ( .B1(n8383), .B2(P2_B_REG_SCAN_IN), .A(n8880), .ZN(n8624) );
  AOI21_X1 U9939 ( .B1(n8914), .B2(n8386), .A(n8628), .ZN(n8915) );
  INV_X1 U9940 ( .A(n8914), .ZN(n8389) );
  AOI22_X1 U9941 ( .A1(P2_REG2_REG_29__SCAN_IN), .A2(n8866), .B1(n8387), .B2(
        n8864), .ZN(n8388) );
  OAI21_X1 U9942 ( .B1(n8389), .B2(n8893), .A(n8388), .ZN(n8390) );
  OAI21_X1 U9943 ( .B1(n8918), .B2(n8850), .A(n8395), .ZN(P2_U3267) );
  OAI21_X1 U9944 ( .B1(n8398), .B2(n8397), .A(n8396), .ZN(n8399) );
  NAND2_X1 U9945 ( .A1(n8399), .A2(n10153), .ZN(n8406) );
  INV_X1 U9946 ( .A(n8400), .ZN(n8404) );
  OAI22_X1 U9947 ( .A1(n8401), .A2(n10148), .B1(n10145), .B2(n8453), .ZN(n8402) );
  AOI211_X1 U9948 ( .C1(n8513), .C2(n8404), .A(n8403), .B(n8402), .ZN(n8405)
         );
  OAI211_X1 U9949 ( .C1(n8407), .C2(n8459), .A(n8406), .B(n8405), .ZN(P2_U3217) );
  INV_X1 U9950 ( .A(n8408), .ZN(n8469) );
  XNOR2_X1 U9951 ( .A(n8469), .B(n8468), .ZN(n8413) );
  OAI22_X1 U9952 ( .A1(n10161), .A2(n8702), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8409), .ZN(n8411) );
  OAI22_X1 U9953 ( .A1(n8427), .A2(n10148), .B1(n10145), .B2(n8440), .ZN(n8410) );
  AOI211_X1 U9954 ( .C1(n8945), .C2(n10151), .A(n8411), .B(n8410), .ZN(n8412)
         );
  OAI21_X1 U9955 ( .B1(n8413), .B2(n8519), .A(n8412), .ZN(P2_U3218) );
  OAI21_X1 U9956 ( .B1(n8416), .B2(n8415), .A(n8414), .ZN(n8417) );
  NAND2_X1 U9957 ( .A1(n8417), .A2(n10153), .ZN(n8422) );
  INV_X1 U9958 ( .A(n8418), .ZN(n8773) );
  AND2_X1 U9959 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8621) );
  OAI22_X1 U9960 ( .A1(n8419), .A2(n10148), .B1(n10145), .B2(n8428), .ZN(n8420) );
  AOI211_X1 U9961 ( .C1(n8513), .C2(n8773), .A(n8621), .B(n8420), .ZN(n8421)
         );
  OAI211_X1 U9962 ( .C1(n8423), .C2(n8459), .A(n8422), .B(n8421), .ZN(P2_U3221) );
  XNOR2_X1 U9963 ( .A(n8425), .B(n8424), .ZN(n8432) );
  INV_X1 U9964 ( .A(n8426), .ZN(n8739) );
  OAI22_X1 U9965 ( .A1(n10161), .A2(n8739), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9133), .ZN(n8430) );
  OAI22_X1 U9966 ( .A1(n8428), .A2(n10148), .B1(n10145), .B2(n8427), .ZN(n8429) );
  AOI211_X1 U9967 ( .C1(n8741), .C2(n10151), .A(n8430), .B(n8429), .ZN(n8431)
         );
  OAI21_X1 U9968 ( .B1(n8432), .B2(n8519), .A(n8431), .ZN(P2_U3225) );
  XNOR2_X1 U9969 ( .A(n8434), .B(n8433), .ZN(n8435) );
  XNOR2_X1 U9970 ( .A(n8436), .B(n8435), .ZN(n8444) );
  INV_X1 U9971 ( .A(n8672), .ZN(n8438) );
  OAI22_X1 U9972 ( .A1(n10161), .A2(n8438), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8437), .ZN(n8442) );
  OAI22_X1 U9973 ( .A1(n8440), .A2(n10148), .B1(n10145), .B2(n8439), .ZN(n8441) );
  AOI211_X1 U9974 ( .C1(n8673), .C2(n10151), .A(n8442), .B(n8441), .ZN(n8443)
         );
  OAI21_X1 U9975 ( .B1(n8444), .B2(n8519), .A(n8443), .ZN(P2_U3227) );
  NAND2_X1 U9976 ( .A1(n8446), .A2(n8445), .ZN(n8447) );
  OAI21_X1 U9977 ( .B1(n8446), .B2(n8445), .A(n8447), .ZN(n8511) );
  NOR2_X1 U9978 ( .A1(n8511), .A2(n8512), .ZN(n8510) );
  INV_X1 U9979 ( .A(n8447), .ZN(n8449) );
  NOR3_X1 U9980 ( .A1(n8510), .A2(n8449), .A3(n8448), .ZN(n8452) );
  INV_X1 U9981 ( .A(n8450), .ZN(n8451) );
  OAI21_X1 U9982 ( .B1(n8452), .B2(n8451), .A(n10153), .ZN(n8458) );
  INV_X1 U9983 ( .A(n8823), .ZN(n8456) );
  OAI22_X1 U9984 ( .A1(n8453), .A2(n10148), .B1(n10145), .B2(n8505), .ZN(n8454) );
  AOI211_X1 U9985 ( .C1(n8513), .C2(n8456), .A(n8455), .B(n8454), .ZN(n8457)
         );
  OAI211_X1 U9986 ( .C1(n8826), .C2(n8459), .A(n8458), .B(n8457), .ZN(P2_U3228) );
  XNOR2_X1 U9987 ( .A(n4513), .B(n8460), .ZN(n8466) );
  NOR2_X1 U9988 ( .A1(n10161), .A2(n8797), .ZN(n8464) );
  AOI22_X1 U9989 ( .A1(n8768), .A2(n8816), .B1(n8815), .B2(n8523), .ZN(n8792)
         );
  OAI21_X1 U9990 ( .B1(n8516), .B2(n8792), .A(n8462), .ZN(n8463) );
  AOI211_X1 U9991 ( .C1(n8980), .C2(n10151), .A(n8464), .B(n8463), .ZN(n8465)
         );
  OAI21_X1 U9992 ( .B1(n8466), .B2(n8519), .A(n8465), .ZN(P2_U3230) );
  OAI21_X1 U9993 ( .B1(n8469), .B2(n8468), .A(n8467), .ZN(n8473) );
  XOR2_X1 U9994 ( .A(n8471), .B(n8470), .Z(n8472) );
  XNOR2_X1 U9995 ( .A(n8473), .B(n8472), .ZN(n8479) );
  OAI22_X1 U9996 ( .A1(n10161), .A2(n8681), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8474), .ZN(n8477) );
  OAI22_X1 U9997 ( .A1(n8496), .A2(n10148), .B1(n10145), .B2(n8475), .ZN(n8476) );
  AOI211_X1 U9998 ( .C1(n8940), .C2(n10151), .A(n8477), .B(n8476), .ZN(n8478)
         );
  OAI21_X1 U9999 ( .B1(n8479), .B2(n8519), .A(n8478), .ZN(P2_U3231) );
  XNOR2_X1 U10000 ( .A(n8481), .B(n8480), .ZN(n8487) );
  INV_X1 U10001 ( .A(n8755), .ZN(n8483) );
  OAI22_X1 U10002 ( .A1(n10161), .A2(n8483), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8482), .ZN(n8485) );
  OAI22_X1 U10003 ( .A1(n8497), .A2(n10145), .B1(n10148), .B2(n8504), .ZN(
        n8484) );
  AOI211_X1 U10004 ( .C1(n8963), .C2(n10151), .A(n8485), .B(n8484), .ZN(n8486)
         );
  OAI21_X1 U10005 ( .B1(n8487), .B2(n8519), .A(n8486), .ZN(P2_U3235) );
  INV_X1 U10006 ( .A(n8488), .ZN(n8489) );
  NAND2_X1 U10007 ( .A1(n8490), .A2(n8489), .ZN(n8494) );
  XOR2_X1 U10008 ( .A(n8492), .B(n8491), .Z(n8493) );
  XNOR2_X1 U10009 ( .A(n8494), .B(n8493), .ZN(n8501) );
  OAI22_X1 U10010 ( .A1(n10161), .A2(n8716), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8495), .ZN(n8499) );
  OAI22_X1 U10011 ( .A1(n8497), .A2(n10148), .B1(n10145), .B2(n8496), .ZN(
        n8498) );
  AOI211_X1 U10012 ( .C1(n8950), .C2(n10151), .A(n8499), .B(n8498), .ZN(n8500)
         );
  OAI21_X1 U10013 ( .B1(n8501), .B2(n8519), .A(n8500), .ZN(P2_U3237) );
  XNOR2_X1 U10014 ( .A(n8503), .B(n8502), .ZN(n8509) );
  NAND2_X1 U10015 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8599) );
  OAI21_X1 U10016 ( .B1(n10161), .B2(n8782), .A(n8599), .ZN(n8507) );
  OAI22_X1 U10017 ( .A1(n8505), .A2(n10148), .B1(n10145), .B2(n8504), .ZN(
        n8506) );
  AOI211_X1 U10018 ( .C1(n8974), .C2(n10151), .A(n8507), .B(n8506), .ZN(n8508)
         );
  OAI21_X1 U10019 ( .B1(n8509), .B2(n8519), .A(n8508), .ZN(P2_U3240) );
  AOI21_X1 U10020 ( .B1(n8512), .B2(n8511), .A(n8510), .ZN(n8520) );
  AOI22_X1 U10021 ( .A1(n8816), .A2(n8523), .B1(n8524), .B2(n8815), .ZN(n8837)
         );
  NAND2_X1 U10022 ( .A1(n8513), .A2(n8834), .ZN(n8515) );
  OAI211_X1 U10023 ( .C1(n8837), .C2(n8516), .A(n8515), .B(n8514), .ZN(n8517)
         );
  AOI21_X1 U10024 ( .B1(n8992), .B2(n10151), .A(n8517), .ZN(n8518) );
  OAI21_X1 U10025 ( .B1(n8520), .B2(n8519), .A(n8518), .ZN(P2_U3243) );
  MUX2_X1 U10026 ( .A(n8521), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8536), .Z(
        P2_U3582) );
  MUX2_X1 U10027 ( .A(n8522), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8536), .Z(
        P2_U3581) );
  MUX2_X1 U10028 ( .A(n8635), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8536), .Z(
        P2_U3580) );
  MUX2_X1 U10029 ( .A(n8657), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8536), .Z(
        P2_U3579) );
  MUX2_X1 U10030 ( .A(n8666), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8536), .Z(
        P2_U3578) );
  MUX2_X1 U10031 ( .A(n8689), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8536), .Z(
        P2_U3577) );
  MUX2_X1 U10032 ( .A(n8699), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8536), .Z(
        P2_U3576) );
  MUX2_X1 U10033 ( .A(n8726), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8536), .Z(
        P2_U3575) );
  MUX2_X1 U10034 ( .A(n8734), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8536), .Z(
        P2_U3574) );
  MUX2_X1 U10035 ( .A(n8751), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8536), .Z(
        P2_U3573) );
  MUX2_X1 U10036 ( .A(n8769), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8536), .Z(
        P2_U3572) );
  MUX2_X1 U10037 ( .A(n8779), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8536), .Z(
        P2_U3571) );
  MUX2_X1 U10038 ( .A(n8768), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8536), .Z(
        P2_U3570) );
  MUX2_X1 U10039 ( .A(n8817), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8536), .Z(
        P2_U3569) );
  MUX2_X1 U10040 ( .A(n8523), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8536), .Z(
        P2_U3568) );
  MUX2_X1 U10041 ( .A(n8814), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8536), .Z(
        P2_U3567) );
  MUX2_X1 U10042 ( .A(n8524), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8536), .Z(
        P2_U3566) );
  MUX2_X1 U10043 ( .A(n8525), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8536), .Z(
        P2_U3565) );
  MUX2_X1 U10044 ( .A(n8526), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8536), .Z(
        P2_U3564) );
  MUX2_X1 U10045 ( .A(n8527), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8536), .Z(
        P2_U3563) );
  MUX2_X1 U10046 ( .A(n8528), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8536), .Z(
        P2_U3562) );
  MUX2_X1 U10047 ( .A(n8529), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8536), .Z(
        P2_U3561) );
  MUX2_X1 U10048 ( .A(n8530), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8536), .Z(
        P2_U3560) );
  MUX2_X1 U10049 ( .A(n8531), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8536), .Z(
        P2_U3559) );
  MUX2_X1 U10050 ( .A(n8532), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8536), .Z(
        P2_U3558) );
  MUX2_X1 U10051 ( .A(n8533), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8536), .Z(
        P2_U3557) );
  MUX2_X1 U10052 ( .A(n8534), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8536), .Z(
        P2_U3556) );
  MUX2_X1 U10053 ( .A(n8535), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8536), .Z(
        P2_U3555) );
  MUX2_X1 U10054 ( .A(n10146), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8536), .Z(
        P2_U3554) );
  MUX2_X1 U10055 ( .A(n4377), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8536), .Z(
        P2_U3553) );
  MUX2_X1 U10056 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8537), .S(P2_U3966), .Z(
        P2_U3552) );
  MUX2_X1 U10057 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n9163), .S(n8538), .Z(n8539)
         );
  INV_X1 U10058 ( .A(n8539), .ZN(n8541) );
  OAI211_X1 U10059 ( .C1(n8542), .C2(n8541), .A(n10163), .B(n8540), .ZN(n8550)
         );
  AOI22_X1 U10060 ( .A1(n10164), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n8549) );
  NAND2_X1 U10061 ( .A1(n8588), .A2(n8543), .ZN(n8548) );
  OAI211_X1 U10062 ( .C1(n8546), .C2(n8545), .A(n10162), .B(n8544), .ZN(n8547)
         );
  NAND4_X1 U10063 ( .A1(n8550), .A2(n8549), .A3(n8548), .A4(n8547), .ZN(
        P2_U3246) );
  NOR2_X1 U10064 ( .A1(n10166), .A2(n8556), .ZN(n8551) );
  AOI211_X1 U10065 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n10164), .A(n8552), .B(
        n8551), .ZN(n8563) );
  OAI211_X1 U10066 ( .C1(n8555), .C2(n8554), .A(n10162), .B(n8553), .ZN(n8562)
         );
  MUX2_X1 U10067 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n8067), .S(n8556), .Z(n8557)
         );
  NAND3_X1 U10068 ( .A1(n8559), .A2(n8558), .A3(n8557), .ZN(n8560) );
  NAND3_X1 U10069 ( .A1(n10163), .A2(n8566), .A3(n8560), .ZN(n8561) );
  NAND3_X1 U10070 ( .A1(n8563), .A2(n8562), .A3(n8561), .ZN(P2_U3253) );
  MUX2_X1 U10071 ( .A(n7413), .B(P2_REG2_REG_9__SCAN_IN), .S(n9319), .Z(n8564)
         );
  NAND3_X1 U10072 ( .A1(n8566), .A2(n8565), .A3(n8564), .ZN(n8567) );
  NAND3_X1 U10073 ( .A1(n10163), .A2(n8579), .A3(n8567), .ZN(n8576) );
  INV_X1 U10074 ( .A(n8568), .ZN(n8569) );
  AOI21_X1 U10075 ( .B1(n10164), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8569), .ZN(
        n8575) );
  OAI211_X1 U10076 ( .C1(n8572), .C2(n8571), .A(n10162), .B(n8570), .ZN(n8574)
         );
  NAND2_X1 U10077 ( .A1(n8588), .A2(n9319), .ZN(n8573) );
  NAND4_X1 U10078 ( .A1(n8576), .A2(n8575), .A3(n8574), .A4(n8573), .ZN(
        P2_U3254) );
  MUX2_X1 U10079 ( .A(n8888), .B(P2_REG2_REG_10__SCAN_IN), .S(n8587), .Z(n8577) );
  NAND3_X1 U10080 ( .A1(n8579), .A2(n8578), .A3(n8577), .ZN(n8580) );
  NAND3_X1 U10081 ( .A1(n10163), .A2(n8581), .A3(n8580), .ZN(n8592) );
  INV_X1 U10082 ( .A(n8582), .ZN(n8583) );
  AOI21_X1 U10083 ( .B1(n10164), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n8583), .ZN(
        n8591) );
  OAI211_X1 U10084 ( .C1(n8586), .C2(n8585), .A(n10162), .B(n8584), .ZN(n8590)
         );
  NAND2_X1 U10085 ( .A1(n8588), .A2(n8587), .ZN(n8589) );
  NAND4_X1 U10086 ( .A1(n8592), .A2(n8591), .A3(n8590), .A4(n8589), .ZN(
        P2_U3255) );
  NAND2_X1 U10087 ( .A1(n8598), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U10088 ( .A1(n8594), .A2(n8593), .ZN(n8595) );
  AOI21_X1 U10089 ( .B1(n8596), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8607), .ZN(
        n8606) );
  INV_X1 U10090 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9119) );
  XNOR2_X1 U10091 ( .A(n8610), .B(n9119), .ZN(n8613) );
  XNOR2_X1 U10092 ( .A(n8613), .B(n8612), .ZN(n8602) );
  NAND2_X1 U10093 ( .A1(n10164), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n8600) );
  NAND2_X1 U10094 ( .A1(n8600), .A2(n8599), .ZN(n8601) );
  AOI21_X1 U10095 ( .B1(n10162), .B2(n8602), .A(n8601), .ZN(n8605) );
  OR2_X1 U10096 ( .A1(n10166), .A2(n8603), .ZN(n8604) );
  OAI211_X1 U10097 ( .C1(n8606), .C2(n10165), .A(n8605), .B(n8604), .ZN(
        P2_U3263) );
  NOR2_X1 U10098 ( .A1(n8608), .A2(n8607), .ZN(n8609) );
  XOR2_X1 U10099 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8609), .Z(n8619) );
  INV_X1 U10100 ( .A(n8619), .ZN(n8615) );
  NOR2_X1 U10101 ( .A1(n8610), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8611) );
  AOI21_X1 U10102 ( .B1(n8613), .B2(n8612), .A(n8611), .ZN(n8614) );
  XNOR2_X1 U10103 ( .A(n8614), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U10104 ( .A1(n10162), .A2(n8616), .ZN(n8617) );
  NAND2_X1 U10105 ( .A1(n8912), .A2(n8628), .ZN(n8622) );
  NAND2_X1 U10106 ( .A1(n8624), .A2(n8623), .ZN(n8910) );
  NOR2_X1 U10107 ( .A1(n8866), .A2(n8910), .ZN(n8629) );
  AOI21_X1 U10108 ( .B1(n8866), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8629), .ZN(
        n8626) );
  NAND2_X1 U10109 ( .A1(n8899), .A2(n8825), .ZN(n8625) );
  OAI211_X1 U10110 ( .C1(n8901), .C2(n8743), .A(n8626), .B(n8625), .ZN(
        P2_U3265) );
  XNOR2_X1 U10111 ( .A(n8628), .B(n8627), .ZN(n8909) );
  NAND2_X1 U10112 ( .A1(n8909), .A2(n8895), .ZN(n8631) );
  AOI21_X1 U10113 ( .B1(n8872), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8629), .ZN(
        n8630) );
  OAI211_X1 U10114 ( .C1(n8912), .C2(n8893), .A(n8631), .B(n8630), .ZN(
        P2_U3266) );
  NAND2_X1 U10115 ( .A1(n8654), .A2(n8632), .ZN(n8634) );
  AOI21_X2 U10116 ( .B1(n8638), .B2(n8886), .A(n8637), .ZN(n8927) );
  AOI21_X1 U10117 ( .B1(n8924), .B2(n8658), .A(n8639), .ZN(n8925) );
  INV_X1 U10118 ( .A(n8640), .ZN(n8641) );
  AOI22_X1 U10119 ( .A1(P2_REG2_REG_27__SCAN_IN), .A2(n8866), .B1(n8641), .B2(
        n8864), .ZN(n8642) );
  OAI21_X1 U10120 ( .B1(n4674), .B2(n8893), .A(n8642), .ZN(n8648) );
  OAI21_X1 U10121 ( .B1(n8645), .B2(n8644), .A(n8643), .ZN(n8646) );
  INV_X1 U10122 ( .A(n8646), .ZN(n8928) );
  NOR2_X1 U10123 ( .A1(n8928), .A2(n8850), .ZN(n8647) );
  AOI211_X1 U10124 ( .C1(n8925), .C2(n8895), .A(n8648), .B(n8647), .ZN(n8649)
         );
  OAI21_X1 U10125 ( .B1(n8866), .B2(n8927), .A(n8649), .ZN(P2_U3269) );
  OAI21_X1 U10126 ( .B1(n8652), .B2(n8651), .A(n8650), .ZN(n8653) );
  INV_X1 U10127 ( .A(n8653), .ZN(n8933) );
  AOI21_X1 U10128 ( .B1(n8671), .B2(n8930), .A(n10282), .ZN(n8659) );
  AND2_X1 U10129 ( .A1(n8659), .A2(n8658), .ZN(n8929) );
  NAND2_X1 U10130 ( .A1(n8929), .A2(n4760), .ZN(n8660) );
  OAI211_X1 U10131 ( .C1(n8891), .C2(n8661), .A(n8932), .B(n8660), .ZN(n8662)
         );
  NAND2_X1 U10132 ( .A1(n8662), .A2(n8393), .ZN(n8664) );
  AOI22_X1 U10133 ( .A1(n8930), .A2(n8825), .B1(n8872), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8663) );
  OAI211_X1 U10134 ( .C1(n8933), .C2(n8850), .A(n8664), .B(n8663), .ZN(
        P2_U3270) );
  XNOR2_X1 U10135 ( .A(n8665), .B(n8669), .ZN(n8667) );
  AOI222_X1 U10136 ( .A1(n8886), .A2(n8667), .B1(n8666), .B2(n8816), .C1(n8699), .C2(n8815), .ZN(n8939) );
  OAI21_X1 U10137 ( .B1(n8670), .B2(n8669), .A(n8668), .ZN(n8937) );
  OAI211_X1 U10138 ( .C1(n8935), .C2(n8680), .A(n10265), .B(n8671), .ZN(n8934)
         );
  AOI22_X1 U10139 ( .A1(n8866), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8672), .B2(
        n8864), .ZN(n8675) );
  NAND2_X1 U10140 ( .A1(n8673), .A2(n8825), .ZN(n8674) );
  OAI211_X1 U10141 ( .C1(n8934), .C2(n8676), .A(n8675), .B(n8674), .ZN(n8677)
         );
  AOI21_X1 U10142 ( .B1(n8937), .B2(n8761), .A(n8677), .ZN(n8678) );
  OAI21_X1 U10143 ( .B1(n8939), .B2(n8872), .A(n8678), .ZN(P2_U3271) );
  XNOR2_X1 U10144 ( .A(n8679), .B(n4643), .ZN(n8944) );
  AOI21_X1 U10145 ( .B1(n8940), .B2(n8701), .A(n8680), .ZN(n8941) );
  INV_X1 U10146 ( .A(n8940), .ZN(n8684) );
  INV_X1 U10147 ( .A(n8681), .ZN(n8682) );
  AOI22_X1 U10148 ( .A1(n8866), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8682), .B2(
        n8864), .ZN(n8683) );
  OAI21_X1 U10149 ( .B1(n8684), .B2(n8893), .A(n8683), .ZN(n8693) );
  INV_X1 U10150 ( .A(n8685), .ZN(n8698) );
  OAI21_X1 U10151 ( .B1(n8698), .B2(n8686), .A(n4643), .ZN(n8688) );
  NAND3_X1 U10152 ( .A1(n8688), .A2(n8886), .A3(n8687), .ZN(n8691) );
  AOI22_X1 U10153 ( .A1(n8689), .A2(n8816), .B1(n8815), .B2(n8726), .ZN(n8690)
         );
  NOR2_X1 U10154 ( .A1(n8943), .A2(n8872), .ZN(n8692) );
  AOI211_X1 U10155 ( .C1(n8941), .C2(n8895), .A(n8693), .B(n8692), .ZN(n8694)
         );
  OAI21_X1 U10156 ( .B1(n8850), .B2(n8944), .A(n8694), .ZN(P2_U3272) );
  AOI21_X1 U10157 ( .B1(n8720), .B2(n8696), .A(n8695), .ZN(n8697) );
  AOI222_X1 U10158 ( .A1(n8886), .A2(n8700), .B1(n8699), .B2(n8816), .C1(n8734), .C2(n8815), .ZN(n8948) );
  AOI21_X1 U10159 ( .B1(n8945), .B2(n8713), .A(n6370), .ZN(n8946) );
  NOR2_X1 U10160 ( .A1(n8891), .A2(n8702), .ZN(n8703) );
  AOI21_X1 U10161 ( .B1(n8866), .B2(P2_REG2_REG_23__SCAN_IN), .A(n8703), .ZN(
        n8704) );
  OAI21_X1 U10162 ( .B1(n8705), .B2(n8893), .A(n8704), .ZN(n8710) );
  OAI21_X1 U10163 ( .B1(n8708), .B2(n8707), .A(n8706), .ZN(n8949) );
  NOR2_X1 U10164 ( .A1(n8949), .A2(n8850), .ZN(n8709) );
  AOI211_X1 U10165 ( .C1(n8946), .C2(n8895), .A(n8710), .B(n8709), .ZN(n8711)
         );
  OAI21_X1 U10166 ( .B1(n8872), .B2(n4386), .A(n8711), .ZN(P2_U3273) );
  XNOR2_X1 U10167 ( .A(n8712), .B(n4645), .ZN(n8954) );
  INV_X1 U10168 ( .A(n8736), .ZN(n8715) );
  INV_X1 U10169 ( .A(n8713), .ZN(n8714) );
  AOI21_X1 U10170 ( .B1(n8950), .B2(n8715), .A(n8714), .ZN(n8951) );
  INV_X1 U10171 ( .A(n8716), .ZN(n8717) );
  AOI22_X1 U10172 ( .A1(n8866), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8717), .B2(
        n8864), .ZN(n8718) );
  OAI21_X1 U10173 ( .B1(n8719), .B2(n8893), .A(n8718), .ZN(n8728) );
  AND2_X1 U10174 ( .A1(n8751), .A2(n8815), .ZN(n8725) );
  INV_X1 U10175 ( .A(n8720), .ZN(n8723) );
  AOI21_X1 U10176 ( .B1(n8731), .B2(n8721), .A(n4645), .ZN(n8722) );
  NOR3_X1 U10177 ( .A1(n8723), .A2(n8722), .A3(n8821), .ZN(n8724) );
  AOI211_X1 U10178 ( .C1(n8816), .C2(n8726), .A(n8725), .B(n8724), .ZN(n8953)
         );
  NOR2_X1 U10179 ( .A1(n8953), .A2(n8872), .ZN(n8727) );
  AOI211_X1 U10180 ( .C1(n8951), .C2(n8895), .A(n8728), .B(n8727), .ZN(n8729)
         );
  OAI21_X1 U10181 ( .B1(n8850), .B2(n8954), .A(n8729), .ZN(P2_U3274) );
  XOR2_X1 U10182 ( .A(n8732), .B(n8730), .Z(n8960) );
  OAI21_X1 U10183 ( .B1(n8733), .B2(n8732), .A(n8731), .ZN(n8735) );
  AOI222_X1 U10184 ( .A1(n8886), .A2(n8735), .B1(n8734), .B2(n8816), .C1(n8769), .C2(n8815), .ZN(n8959) );
  INV_X1 U10185 ( .A(n8959), .ZN(n8745) );
  AND2_X1 U10186 ( .A1(n8741), .A2(n5022), .ZN(n8737) );
  OR2_X1 U10187 ( .A1(n8737), .A2(n8736), .ZN(n8956) );
  NAND2_X1 U10188 ( .A1(n8866), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8738) );
  OAI21_X1 U10189 ( .B1(n8891), .B2(n8739), .A(n8738), .ZN(n8740) );
  AOI21_X1 U10190 ( .B1(n8741), .B2(n8825), .A(n8740), .ZN(n8742) );
  OAI21_X1 U10191 ( .B1(n8956), .B2(n8743), .A(n8742), .ZN(n8744) );
  AOI21_X1 U10192 ( .B1(n8745), .B2(n8393), .A(n8744), .ZN(n8746) );
  OAI21_X1 U10193 ( .B1(n8960), .B2(n8850), .A(n8746), .ZN(P2_U3275) );
  AOI21_X1 U10194 ( .B1(n8766), .B2(n8748), .A(n8759), .ZN(n8749) );
  AOI22_X1 U10195 ( .A1(n8751), .A2(n8816), .B1(n8815), .B2(n8779), .ZN(n8752)
         );
  NAND2_X1 U10196 ( .A1(n8771), .A2(n8963), .ZN(n8754) );
  AND2_X1 U10197 ( .A1(n5022), .A2(n8754), .ZN(n8964) );
  AOI22_X1 U10198 ( .A1(n8866), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8755), .B2(
        n8864), .ZN(n8756) );
  OAI21_X1 U10199 ( .B1(n8757), .B2(n8893), .A(n8756), .ZN(n8758) );
  AOI21_X1 U10200 ( .B1(n8895), .B2(n8964), .A(n8758), .ZN(n8763) );
  NAND2_X1 U10201 ( .A1(n8760), .A2(n8759), .ZN(n8961) );
  NAND3_X1 U10202 ( .A1(n8962), .A2(n8961), .A3(n8761), .ZN(n8762) );
  OAI211_X1 U10203 ( .C1(n8968), .C2(n8872), .A(n8763), .B(n8762), .ZN(
        P2_U3276) );
  XNOR2_X1 U10204 ( .A(n8764), .B(n8765), .ZN(n8973) );
  OAI21_X1 U10205 ( .B1(n8767), .B2(n6346), .A(n8766), .ZN(n8770) );
  AOI222_X1 U10206 ( .A1(n8886), .A2(n8770), .B1(n8769), .B2(n8816), .C1(n8768), .C2(n8815), .ZN(n8972) );
  INV_X1 U10207 ( .A(n8771), .ZN(n8772) );
  AOI211_X1 U10208 ( .C1(n8970), .C2(n4837), .A(n10282), .B(n8772), .ZN(n8969)
         );
  AOI22_X1 U10209 ( .A1(n8969), .A2(n4760), .B1(n8864), .B2(n8773), .ZN(n8774)
         );
  AOI21_X1 U10210 ( .B1(n8972), .B2(n8774), .A(n8866), .ZN(n8775) );
  INV_X1 U10211 ( .A(n8775), .ZN(n8777) );
  AOI22_X1 U10212 ( .A1(n8970), .A2(n8825), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n8872), .ZN(n8776) );
  OAI211_X1 U10213 ( .C1(n8973), .C2(n8850), .A(n8777), .B(n8776), .ZN(
        P2_U3277) );
  XNOR2_X1 U10214 ( .A(n8778), .B(n8785), .ZN(n8780) );
  AOI222_X1 U10215 ( .A1(n8886), .A2(n8780), .B1(n8779), .B2(n8816), .C1(n8817), .C2(n8815), .ZN(n8977) );
  AOI21_X1 U10216 ( .B1(n8974), .B2(n8795), .A(n8781), .ZN(n8975) );
  INV_X1 U10217 ( .A(n8782), .ZN(n8783) );
  AOI22_X1 U10218 ( .A1(n8866), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8783), .B2(
        n8864), .ZN(n8784) );
  OAI21_X1 U10219 ( .B1(n4835), .B2(n8893), .A(n8784), .ZN(n8788) );
  XOR2_X1 U10220 ( .A(n8786), .B(n8785), .Z(n8978) );
  NOR2_X1 U10221 ( .A1(n8978), .A2(n8850), .ZN(n8787) );
  AOI211_X1 U10222 ( .C1(n8975), .C2(n8895), .A(n8788), .B(n8787), .ZN(n8789)
         );
  OAI21_X1 U10223 ( .B1(n8866), .B2(n8977), .A(n8789), .ZN(P2_U3278) );
  XNOR2_X1 U10224 ( .A(n8791), .B(n8790), .ZN(n8794) );
  INV_X1 U10225 ( .A(n8792), .ZN(n8793) );
  AOI21_X1 U10226 ( .B1(n8794), .B2(n8886), .A(n8793), .ZN(n8982) );
  INV_X1 U10227 ( .A(n8795), .ZN(n8796) );
  AOI211_X1 U10228 ( .C1(n8980), .C2(n8828), .A(n10282), .B(n8796), .ZN(n8979)
         );
  INV_X1 U10229 ( .A(n8980), .ZN(n8800) );
  INV_X1 U10230 ( .A(n8797), .ZN(n8798) );
  AOI22_X1 U10231 ( .A1(n8866), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8798), .B2(
        n8864), .ZN(n8799) );
  OAI21_X1 U10232 ( .B1(n8800), .B2(n8893), .A(n8799), .ZN(n8806) );
  NAND2_X1 U10233 ( .A1(n8813), .A2(n8802), .ZN(n8804) );
  XNOR2_X1 U10234 ( .A(n8804), .B(n8803), .ZN(n8983) );
  NOR2_X1 U10235 ( .A1(n8983), .A2(n8850), .ZN(n8805) );
  AOI211_X1 U10236 ( .C1(n8979), .C2(n8807), .A(n8806), .B(n8805), .ZN(n8808)
         );
  OAI21_X1 U10237 ( .B1(n8872), .B2(n8982), .A(n8808), .ZN(P2_U3279) );
  XNOR2_X1 U10238 ( .A(n8810), .B(n8809), .ZN(n8820) );
  NAND2_X1 U10239 ( .A1(n8801), .A2(n8811), .ZN(n8812) );
  NAND2_X1 U10240 ( .A1(n8813), .A2(n8812), .ZN(n8987) );
  OR2_X1 U10241 ( .A1(n8987), .A2(n8913), .ZN(n8819) );
  AOI22_X1 U10242 ( .A1(n8817), .A2(n8816), .B1(n8815), .B2(n8814), .ZN(n8818)
         );
  OAI211_X1 U10243 ( .C1(n8821), .C2(n8820), .A(n8819), .B(n8818), .ZN(n8989)
         );
  NAND2_X1 U10244 ( .A1(n8866), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8822) );
  OAI21_X1 U10245 ( .B1(n8891), .B2(n8823), .A(n8822), .ZN(n8824) );
  AOI21_X1 U10246 ( .B1(n8984), .B2(n8825), .A(n8824), .ZN(n8830) );
  OR2_X1 U10247 ( .A1(n8843), .A2(n8826), .ZN(n8827) );
  AND2_X1 U10248 ( .A1(n8828), .A2(n8827), .ZN(n8985) );
  NAND2_X1 U10249 ( .A1(n8985), .A2(n8895), .ZN(n8829) );
  OAI211_X1 U10250 ( .C1(n8987), .C2(n8898), .A(n8830), .B(n8829), .ZN(n8831)
         );
  AOI21_X1 U10251 ( .B1(n8393), .B2(n8989), .A(n8831), .ZN(n8832) );
  INV_X1 U10252 ( .A(n8832), .ZN(P2_U3280) );
  XNOR2_X1 U10253 ( .A(n8833), .B(n4802), .ZN(n8996) );
  INV_X1 U10254 ( .A(n8834), .ZN(n8840) );
  XNOR2_X1 U10255 ( .A(n8836), .B(n8835), .ZN(n8839) );
  INV_X1 U10256 ( .A(n8837), .ZN(n8838) );
  AOI21_X1 U10257 ( .B1(n8839), .B2(n8886), .A(n8838), .ZN(n8995) );
  OAI21_X1 U10258 ( .B1(n8840), .B2(n8891), .A(n8995), .ZN(n8841) );
  NAND2_X1 U10259 ( .A1(n8841), .A2(n8393), .ZN(n8849) );
  INV_X1 U10260 ( .A(n8842), .ZN(n8844) );
  AOI21_X1 U10261 ( .B1(n8992), .B2(n8844), .A(n8843), .ZN(n8993) );
  INV_X1 U10262 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8845) );
  OAI22_X1 U10263 ( .A1(n8846), .A2(n8893), .B1(n8393), .B2(n8845), .ZN(n8847)
         );
  AOI21_X1 U10264 ( .B1(n8993), .B2(n8895), .A(n8847), .ZN(n8848) );
  OAI211_X1 U10265 ( .C1(n8996), .C2(n8850), .A(n8849), .B(n8848), .ZN(
        P2_U3281) );
  OAI21_X1 U10266 ( .B1(n8857), .B2(n8852), .A(n8851), .ZN(n8861) );
  OAI22_X1 U10267 ( .A1(n8854), .A2(n8882), .B1(n8853), .B2(n8880), .ZN(n8860)
         );
  NAND2_X1 U10268 ( .A1(n8856), .A2(n8855), .ZN(n8858) );
  XNOR2_X1 U10269 ( .A(n8858), .B(n8857), .ZN(n9006) );
  NOR2_X1 U10270 ( .A1(n9006), .A2(n8913), .ZN(n8859) );
  AOI211_X1 U10271 ( .C1(n8886), .C2(n8861), .A(n8860), .B(n8859), .ZN(n9005)
         );
  XOR2_X1 U10272 ( .A(n8862), .B(n9002), .Z(n9003) );
  INV_X1 U10273 ( .A(n9002), .ZN(n8868) );
  INV_X1 U10274 ( .A(n8863), .ZN(n8865) );
  AOI22_X1 U10275 ( .A1(n8866), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8865), .B2(
        n8864), .ZN(n8867) );
  OAI21_X1 U10276 ( .B1(n8868), .B2(n8893), .A(n8867), .ZN(n8870) );
  NOR2_X1 U10277 ( .A1(n9006), .A2(n8898), .ZN(n8869) );
  AOI211_X1 U10278 ( .C1(n9003), .C2(n8895), .A(n8870), .B(n8869), .ZN(n8871)
         );
  OAI21_X1 U10279 ( .B1(n9005), .B2(n8872), .A(n8871), .ZN(P2_U3283) );
  NAND2_X1 U10280 ( .A1(n8874), .A2(n8873), .ZN(n8875) );
  XOR2_X1 U10281 ( .A(n8879), .B(n8875), .Z(n10270) );
  NAND2_X1 U10282 ( .A1(n8877), .A2(n8876), .ZN(n8878) );
  XOR2_X1 U10283 ( .A(n8879), .B(n8878), .Z(n8887) );
  OAI22_X1 U10284 ( .A1(n8883), .A2(n8882), .B1(n8881), .B2(n8880), .ZN(n8885)
         );
  NOR2_X1 U10285 ( .A1(n10270), .A2(n8913), .ZN(n8884) );
  AOI211_X1 U10286 ( .C1(n8887), .C2(n8886), .A(n8885), .B(n8884), .ZN(n10268)
         );
  MUX2_X1 U10287 ( .A(n8888), .B(n10268), .S(n8393), .Z(n8897) );
  AOI21_X1 U10288 ( .B1(n10263), .B2(n8890), .A(n8889), .ZN(n10266) );
  OAI22_X1 U10289 ( .A1(n8893), .A2(n4838), .B1(n8892), .B2(n8891), .ZN(n8894)
         );
  AOI21_X1 U10290 ( .B1(n10266), .B2(n8895), .A(n8894), .ZN(n8896) );
  OAI211_X1 U10291 ( .C1(n10270), .C2(n8898), .A(n8897), .B(n8896), .ZN(
        P2_U3286) );
  NAND2_X1 U10292 ( .A1(n8899), .A2(n10264), .ZN(n8900) );
  OAI211_X1 U10293 ( .C1(n8901), .C2(n10282), .A(n8900), .B(n8910), .ZN(n9009)
         );
  NAND4_X1 U10294 ( .A1(n8905), .A2(n8904), .A3(n8903), .A4(n8902), .ZN(n8906)
         );
  MUX2_X1 U10295 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9009), .S(n10314), .Z(
        P2_U3551) );
  NAND2_X1 U10296 ( .A1(n8909), .A2(n10265), .ZN(n8911) );
  OAI211_X1 U10297 ( .C1(n8912), .C2(n10280), .A(n8911), .B(n8910), .ZN(n9010)
         );
  MUX2_X1 U10298 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9010), .S(n10314), .Z(
        P2_U3550) );
  AOI22_X1 U10299 ( .A1(n8915), .A2(n10265), .B1(n10264), .B2(n8914), .ZN(
        n8916) );
  MUX2_X1 U10300 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9011), .S(n10314), .Z(
        P2_U3549) );
  AOI22_X1 U10301 ( .A1(n8920), .A2(n10265), .B1(n10264), .B2(n8919), .ZN(
        n8921) );
  OAI211_X1 U10302 ( .C1(n8923), .C2(n10206), .A(n8922), .B(n8921), .ZN(n9012)
         );
  MUX2_X1 U10303 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9012), .S(n10314), .Z(
        P2_U3548) );
  AOI22_X1 U10304 ( .A1(n8925), .A2(n10265), .B1(n10264), .B2(n8924), .ZN(
        n8926) );
  OAI211_X1 U10305 ( .C1(n8928), .C2(n10206), .A(n8927), .B(n8926), .ZN(n9013)
         );
  MUX2_X1 U10306 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9013), .S(n10314), .Z(
        P2_U3547) );
  AOI21_X1 U10307 ( .B1(n10264), .B2(n8930), .A(n8929), .ZN(n8931) );
  OAI211_X1 U10308 ( .C1(n8933), .C2(n10206), .A(n8932), .B(n8931), .ZN(n9014)
         );
  MUX2_X1 U10309 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9014), .S(n10314), .Z(
        P2_U3546) );
  OAI21_X1 U10310 ( .B1(n8935), .B2(n10280), .A(n8934), .ZN(n8936) );
  AOI21_X1 U10311 ( .B1(n8937), .B2(n10287), .A(n8936), .ZN(n8938) );
  NAND2_X1 U10312 ( .A1(n8939), .A2(n8938), .ZN(n9015) );
  MUX2_X1 U10313 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9015), .S(n10314), .Z(
        P2_U3545) );
  AOI22_X1 U10314 ( .A1(n8941), .A2(n10265), .B1(n10264), .B2(n8940), .ZN(
        n8942) );
  OAI211_X1 U10315 ( .C1(n8944), .C2(n10206), .A(n8943), .B(n8942), .ZN(n9016)
         );
  MUX2_X1 U10316 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9016), .S(n10314), .Z(
        P2_U3544) );
  AOI22_X1 U10317 ( .A1(n8946), .A2(n10265), .B1(n10264), .B2(n8945), .ZN(
        n8947) );
  OAI211_X1 U10318 ( .C1(n10206), .C2(n8949), .A(n4386), .B(n8947), .ZN(n9017)
         );
  MUX2_X1 U10319 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9017), .S(n10314), .Z(
        P2_U3543) );
  AOI22_X1 U10320 ( .A1(n8951), .A2(n10265), .B1(n10264), .B2(n8950), .ZN(
        n8952) );
  OAI211_X1 U10321 ( .C1(n10206), .C2(n8954), .A(n8953), .B(n8952), .ZN(n9018)
         );
  MUX2_X1 U10322 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9018), .S(n10314), .Z(
        P2_U3542) );
  OAI22_X1 U10323 ( .A1(n8956), .A2(n10282), .B1(n8955), .B2(n10280), .ZN(
        n8957) );
  INV_X1 U10324 ( .A(n8957), .ZN(n8958) );
  OAI211_X1 U10325 ( .C1(n10206), .C2(n8960), .A(n8959), .B(n8958), .ZN(n9019)
         );
  MUX2_X1 U10326 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9019), .S(n10314), .Z(
        P2_U3541) );
  NAND3_X1 U10327 ( .A1(n8962), .A2(n8961), .A3(n10287), .ZN(n8966) );
  AOI22_X1 U10328 ( .A1(n8964), .A2(n10265), .B1(n10264), .B2(n8963), .ZN(
        n8965) );
  AND2_X1 U10329 ( .A1(n8966), .A2(n8965), .ZN(n8967) );
  NAND2_X1 U10330 ( .A1(n8968), .A2(n8967), .ZN(n9020) );
  MUX2_X1 U10331 ( .A(n9020), .B(P2_REG1_REG_20__SCAN_IN), .S(n10311), .Z(
        P2_U3540) );
  AOI21_X1 U10332 ( .B1(n10264), .B2(n8970), .A(n8969), .ZN(n8971) );
  OAI211_X1 U10333 ( .C1(n10206), .C2(n8973), .A(n8972), .B(n8971), .ZN(n9021)
         );
  MUX2_X1 U10334 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9021), .S(n10314), .Z(
        P2_U3539) );
  AOI22_X1 U10335 ( .A1(n8975), .A2(n10265), .B1(n10264), .B2(n8974), .ZN(
        n8976) );
  OAI211_X1 U10336 ( .C1(n10206), .C2(n8978), .A(n8977), .B(n8976), .ZN(n9022)
         );
  MUX2_X1 U10337 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9022), .S(n10314), .Z(
        P2_U3538) );
  AOI21_X1 U10338 ( .B1(n10264), .B2(n8980), .A(n8979), .ZN(n8981) );
  OAI211_X1 U10339 ( .C1(n8983), .C2(n10206), .A(n8982), .B(n8981), .ZN(n9023)
         );
  MUX2_X1 U10340 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9023), .S(n10314), .Z(
        P2_U3537) );
  AOI22_X1 U10341 ( .A1(n8985), .A2(n10265), .B1(n10264), .B2(n8984), .ZN(
        n8986) );
  OAI21_X1 U10342 ( .B1(n8987), .B2(n10269), .A(n8986), .ZN(n8988) );
  NOR2_X1 U10343 ( .A1(n8989), .A2(n8988), .ZN(n9024) );
  MUX2_X1 U10344 ( .A(n8990), .B(n9024), .S(n10314), .Z(n8991) );
  INV_X1 U10345 ( .A(n8991), .ZN(P2_U3536) );
  AOI22_X1 U10346 ( .A1(n8993), .A2(n10265), .B1(n10264), .B2(n8992), .ZN(
        n8994) );
  OAI211_X1 U10347 ( .C1(n8996), .C2(n10206), .A(n8995), .B(n8994), .ZN(n9027)
         );
  MUX2_X1 U10348 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9027), .S(n10314), .Z(
        P2_U3535) );
  AOI22_X1 U10349 ( .A1(n8998), .A2(n10265), .B1(n10264), .B2(n8997), .ZN(
        n8999) );
  OAI211_X1 U10350 ( .C1(n9001), .C2(n10206), .A(n9000), .B(n8999), .ZN(n9028)
         );
  MUX2_X1 U10351 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9028), .S(n10314), .Z(
        P2_U3534) );
  AOI22_X1 U10352 ( .A1(n9003), .A2(n10265), .B1(n10264), .B2(n9002), .ZN(
        n9004) );
  OAI211_X1 U10353 ( .C1(n9006), .C2(n10269), .A(n9005), .B(n9004), .ZN(n9029)
         );
  MUX2_X1 U10354 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9029), .S(n10314), .Z(
        P2_U3533) );
  MUX2_X1 U10355 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9009), .S(n10290), .Z(
        P2_U3519) );
  MUX2_X1 U10356 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9010), .S(n10290), .Z(
        P2_U3518) );
  MUX2_X1 U10357 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9012), .S(n10290), .Z(
        P2_U3516) );
  MUX2_X1 U10358 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9013), .S(n10290), .Z(
        P2_U3515) );
  MUX2_X1 U10359 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9014), .S(n10290), .Z(
        P2_U3514) );
  MUX2_X1 U10360 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9015), .S(n10290), .Z(
        P2_U3513) );
  MUX2_X1 U10361 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9016), .S(n10290), .Z(
        P2_U3512) );
  MUX2_X1 U10362 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9017), .S(n10290), .Z(
        P2_U3511) );
  MUX2_X1 U10363 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9018), .S(n10290), .Z(
        P2_U3510) );
  MUX2_X1 U10364 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9019), .S(n10290), .Z(
        P2_U3509) );
  MUX2_X1 U10365 ( .A(n9020), .B(P2_REG0_REG_20__SCAN_IN), .S(n10288), .Z(
        P2_U3508) );
  MUX2_X1 U10366 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9021), .S(n10290), .Z(
        P2_U3507) );
  MUX2_X1 U10367 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9022), .S(n10290), .Z(
        P2_U3505) );
  MUX2_X1 U10368 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9023), .S(n10290), .Z(
        P2_U3502) );
  INV_X1 U10369 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9025) );
  MUX2_X1 U10370 ( .A(n9025), .B(n9024), .S(n10290), .Z(n9026) );
  INV_X1 U10371 ( .A(n9026), .ZN(P2_U3499) );
  MUX2_X1 U10372 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9027), .S(n10290), .Z(
        P2_U3496) );
  MUX2_X1 U10373 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9028), .S(n10290), .Z(
        P2_U3493) );
  MUX2_X1 U10374 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9029), .S(n10290), .Z(
        P2_U3490) );
  INV_X1 U10375 ( .A(n9030), .ZN(n9847) );
  NOR4_X1 U10376 ( .A1(n9031), .A2(P2_IR_REG_30__SCAN_IN), .A3(n6283), .A4(
        P2_U3152), .ZN(n9032) );
  AOI21_X1 U10377 ( .B1(n9320), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9032), .ZN(
        n9033) );
  OAI21_X1 U10378 ( .B1(n9847), .B2(n9036), .A(n9033), .ZN(P2_U3327) );
  OAI222_X1 U10379 ( .A1(n9043), .A2(n9103), .B1(n9036), .B2(n9035), .C1(n9034), .C2(P2_U3152), .ZN(P2_U3328) );
  OAI222_X1 U10380 ( .A1(P2_U3152), .A2(n9038), .B1(n9036), .B2(n9037), .C1(
        n9292), .C2(n9043), .ZN(P2_U3329) );
  INV_X1 U10381 ( .A(n9039), .ZN(n9854) );
  OAI222_X1 U10382 ( .A1(n9043), .A2(n9041), .B1(P2_U3152), .B2(n9040), .C1(
        n9036), .C2(n9854), .ZN(P2_U3331) );
  INV_X1 U10383 ( .A(n9042), .ZN(n9856) );
  OAI222_X1 U10384 ( .A1(P2_U3152), .A2(n9045), .B1(n9036), .B2(n9856), .C1(
        n9044), .C2(n9043), .ZN(P2_U3332) );
  INV_X1 U10385 ( .A(SI_6_), .ZN(n9047) );
  NAND4_X1 U10386 ( .A1(n9049), .A2(n9048), .A3(n9047), .A4(n9046), .ZN(n9054)
         );
  AND4_X1 U10387 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(P1_REG1_REG_11__SCAN_IN), 
        .A3(P1_REG1_REG_3__SCAN_IN), .A4(P2_REG2_REG_29__SCAN_IN), .ZN(n9050)
         );
  INV_X1 U10388 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n9286) );
  AND4_X1 U10389 ( .A1(n9050), .A2(n7471), .A3(n5049), .A4(n9286), .ZN(n9051)
         );
  NAND4_X1 U10390 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .A3(
        P2_RD_REG_SCAN_IN), .A4(n9051), .ZN(n9053) );
  NOR4_X1 U10391 ( .A1(n9054), .A2(n9053), .A3(n9052), .A4(n5085), .ZN(n9101)
         );
  INV_X1 U10392 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10058) );
  INV_X1 U10393 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9266) );
  NAND4_X1 U10394 ( .A1(n9056), .A2(n9055), .A3(P1_ADDR_REG_3__SCAN_IN), .A4(
        n9266), .ZN(n9059) );
  NAND4_X1 U10395 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .A3(P2_ADDR_REG_15__SCAN_IN), .A4(P2_ADDR_REG_14__SCAN_IN), .ZN(n9058)
         );
  NAND4_X1 U10396 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .A3(P1_ADDR_REG_7__SCAN_IN), .A4(P1_ADDR_REG_8__SCAN_IN), .ZN(n9057)
         );
  NOR4_X1 U10397 ( .A1(n10058), .A2(n9059), .A3(n9058), .A4(n9057), .ZN(n9100)
         );
  INV_X1 U10398 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9122) );
  NOR4_X1 U10399 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(P1_REG1_REG_13__SCAN_IN), 
        .A3(n9122), .A4(n9103), .ZN(n9064) );
  INV_X1 U10400 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9108) );
  NOR4_X1 U10401 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P2_DATAO_REG_11__SCAN_IN), 
        .A3(n9060), .A4(n9108), .ZN(n9063) );
  INV_X1 U10402 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9138) );
  NOR4_X1 U10403 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_REG2_REG_16__SCAN_IN), 
        .A3(P2_REG3_REG_21__SCAN_IN), .A4(n9138), .ZN(n9062) );
  NOR4_X1 U10404 ( .A1(P1_REG0_REG_23__SCAN_IN), .A2(P2_REG2_REG_7__SCAN_IN), 
        .A3(n9131), .A4(n9119), .ZN(n9061) );
  AND4_X1 U10405 ( .A1(n9064), .A2(n9063), .A3(n9062), .A4(n9061), .ZN(n9070)
         );
  NAND4_X1 U10406 ( .A1(SI_22_), .A2(P1_REG3_REG_21__SCAN_IN), .A3(
        P2_IR_REG_21__SCAN_IN), .A4(P2_REG0_REG_24__SCAN_IN), .ZN(n9065) );
  NOR3_X1 U10407 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .A3(n9065), .ZN(n9069) );
  NAND4_X1 U10408 ( .A1(P1_D_REG_16__SCAN_IN), .A2(SI_26_), .A3(
        P1_REG3_REG_27__SCAN_IN), .A4(P2_REG1_REG_5__SCAN_IN), .ZN(n9067) );
  INV_X1 U10409 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9252) );
  NAND4_X1 U10410 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(P1_REG1_REG_18__SCAN_IN), .A3(n9252), .A4(n9240), .ZN(n9066) );
  NOR4_X1 U10411 ( .A1(n9067), .A2(P2_DATAO_REG_19__SCAN_IN), .A3(
        P1_IR_REG_26__SCAN_IN), .A4(n9066), .ZN(n9068) );
  AND3_X1 U10412 ( .A1(n9070), .A2(n9069), .A3(n9068), .ZN(n9099) );
  INV_X1 U10413 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10128) );
  INV_X1 U10414 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10068) );
  NOR4_X1 U10415 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(n10128), .A3(n10068), 
        .A4(n9279), .ZN(n9072) );
  INV_X1 U10416 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9071) );
  NAND3_X1 U10417 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9072), .A3(n9071), .ZN(
        n9083) );
  NOR4_X1 U10418 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(P1_REG2_REG_26__SCAN_IN), 
        .A3(P1_REG1_REG_31__SCAN_IN), .A4(n9292), .ZN(n9074) );
  INV_X1 U10419 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9226) );
  NOR4_X1 U10420 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .A3(
        n9226), .A4(n9225), .ZN(n9073) );
  NAND3_X1 U10421 ( .A1(n9075), .A2(n9074), .A3(n9073), .ZN(n9076) );
  INV_X1 U10422 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9923) );
  OR4_X1 U10423 ( .A1(n9076), .A2(n9300), .A3(n9923), .A4(P1_D_REG_7__SCAN_IN), 
        .ZN(n9082) );
  INV_X1 U10424 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9078) );
  NAND4_X1 U10425 ( .A1(n9078), .A2(n9077), .A3(P2_IR_REG_13__SCAN_IN), .A4(
        P2_REG3_REG_14__SCAN_IN), .ZN(n9081) );
  INV_X1 U10426 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9079) );
  NAND4_X1 U10427 ( .A1(n5877), .A2(n9079), .A3(P1_IR_REG_15__SCAN_IN), .A4(
        P1_REG3_REG_5__SCAN_IN), .ZN(n9080) );
  NOR4_X1 U10428 ( .A1(n9083), .A2(n9082), .A3(n9081), .A4(n9080), .ZN(n9086)
         );
  NAND4_X1 U10429 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P2_REG2_REG_12__SCAN_IN), 
        .A3(n9210), .A4(n9215), .ZN(n9084) );
  NOR3_X1 U10430 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(P2_REG0_REG_22__SCAN_IN), 
        .A3(n9084), .ZN(n9085) );
  NAND2_X1 U10431 ( .A1(n9086), .A2(n9085), .ZN(n9097) );
  NAND4_X1 U10432 ( .A1(P1_REG0_REG_10__SCAN_IN), .A2(P2_REG3_REG_13__SCAN_IN), 
        .A3(n9173), .A4(n6405), .ZN(n9096) );
  NAND4_X1 U10433 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P1_REG3_REG_22__SCAN_IN), 
        .A3(P2_REG3_REG_11__SCAN_IN), .A4(n9163), .ZN(n9095) );
  NOR4_X1 U10434 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P2_DATAO_REG_15__SCAN_IN), 
        .A3(P2_REG1_REG_17__SCAN_IN), .A4(P2_REG0_REG_1__SCAN_IN), .ZN(n9093)
         );
  INV_X1 U10435 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9145) );
  NOR4_X1 U10436 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(P1_REG2_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .A4(n9145), .ZN(n9092) );
  NAND4_X1 U10437 ( .A1(SI_24_), .A2(P2_IR_REG_14__SCAN_IN), .A3(
        P2_REG1_REG_27__SCAN_IN), .A4(n7077), .ZN(n9090) );
  INV_X1 U10438 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10208) );
  NAND4_X1 U10439 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P2_REG2_REG_25__SCAN_IN), 
        .A3(n10184), .A4(n10208), .ZN(n9089) );
  NAND4_X1 U10440 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), 
        .A3(n9196), .A4(n9200), .ZN(n9088) );
  NAND4_X1 U10441 ( .A1(P1_REG1_REG_14__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), 
        .A3(P2_REG3_REG_4__SCAN_IN), .A4(P2_REG0_REG_10__SCAN_IN), .ZN(n9087)
         );
  NOR4_X1 U10442 ( .A1(n9090), .A2(n9089), .A3(n9088), .A4(n9087), .ZN(n9091)
         );
  NAND3_X1 U10443 ( .A1(n9093), .A2(n9092), .A3(n9091), .ZN(n9094) );
  NOR4_X1 U10444 ( .A1(n9097), .A2(n9096), .A3(n9095), .A4(n9094), .ZN(n9098)
         );
  NAND4_X1 U10445 ( .A1(n9101), .A2(n9100), .A3(n9099), .A4(n9098), .ZN(n9318)
         );
  INV_X1 U10446 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10056) );
  AOI22_X1 U10447 ( .A1(n9103), .A2(keyinput82), .B1(n10056), .B2(keyinput64), 
        .ZN(n9102) );
  OAI221_X1 U10448 ( .B1(n9103), .B2(keyinput82), .C1(n10056), .C2(keyinput64), 
        .A(n9102), .ZN(n9114) );
  INV_X1 U10449 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9331) );
  AOI22_X1 U10450 ( .A1(n9105), .A2(keyinput48), .B1(keyinput31), .B2(n9331), 
        .ZN(n9104) );
  OAI221_X1 U10451 ( .B1(n9105), .B2(keyinput48), .C1(n9331), .C2(keyinput31), 
        .A(n9104), .ZN(n9113) );
  AOI22_X1 U10452 ( .A1(n9108), .A2(keyinput61), .B1(n9107), .B2(keyinput110), 
        .ZN(n9106) );
  OAI221_X1 U10453 ( .B1(n9108), .B2(keyinput61), .C1(n9107), .C2(keyinput110), 
        .A(n9106), .ZN(n9112) );
  XNOR2_X1 U10454 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(keyinput5), .ZN(n9110) );
  XNOR2_X1 U10455 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput70), .ZN(n9109) );
  NAND2_X1 U10456 ( .A1(n9110), .A2(n9109), .ZN(n9111) );
  NOR4_X1 U10457 ( .A1(n9114), .A2(n9113), .A3(n9112), .A4(n9111), .ZN(n9157)
         );
  INV_X1 U10458 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9116) );
  AOI22_X1 U10459 ( .A1(n9116), .A2(keyinput21), .B1(keyinput50), .B2(n7352), 
        .ZN(n9115) );
  OAI221_X1 U10460 ( .B1(n9116), .B2(keyinput21), .C1(n7352), .C2(keyinput50), 
        .A(n9115), .ZN(n9128) );
  INV_X1 U10461 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9118) );
  AOI22_X1 U10462 ( .A1(n9119), .A2(keyinput73), .B1(n9118), .B2(keyinput55), 
        .ZN(n9117) );
  OAI221_X1 U10463 ( .B1(n9119), .B2(keyinput73), .C1(n9118), .C2(keyinput55), 
        .A(n9117), .ZN(n9127) );
  INV_X1 U10464 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9121) );
  AOI22_X1 U10465 ( .A1(n9122), .A2(keyinput125), .B1(keyinput54), .B2(n9121), 
        .ZN(n9120) );
  OAI221_X1 U10466 ( .B1(n9122), .B2(keyinput125), .C1(n9121), .C2(keyinput54), 
        .A(n9120), .ZN(n9126) );
  XNOR2_X1 U10467 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(keyinput16), .ZN(n9124)
         );
  XNOR2_X1 U10468 ( .A(SI_6_), .B(keyinput44), .ZN(n9123) );
  NAND2_X1 U10469 ( .A1(n9124), .A2(n9123), .ZN(n9125) );
  NOR4_X1 U10470 ( .A1(n9128), .A2(n9127), .A3(n9126), .A4(n9125), .ZN(n9156)
         );
  INV_X1 U10471 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9130) );
  AOI22_X1 U10472 ( .A1(n9131), .A2(keyinput66), .B1(keyinput94), .B2(n9130), 
        .ZN(n9129) );
  OAI221_X1 U10473 ( .B1(n9131), .B2(keyinput66), .C1(n9130), .C2(keyinput94), 
        .A(n9129), .ZN(n9142) );
  AOI22_X1 U10474 ( .A1(n9134), .A2(keyinput9), .B1(keyinput117), .B2(n9133), 
        .ZN(n9132) );
  OAI221_X1 U10475 ( .B1(n9134), .B2(keyinput9), .C1(n9133), .C2(keyinput117), 
        .A(n9132), .ZN(n9141) );
  AOI22_X1 U10476 ( .A1(n8196), .A2(keyinput0), .B1(keyinput20), .B2(n4526), 
        .ZN(n9135) );
  OAI221_X1 U10477 ( .B1(n8196), .B2(keyinput0), .C1(n4526), .C2(keyinput20), 
        .A(n9135), .ZN(n9140) );
  AOI22_X1 U10478 ( .A1(n9138), .A2(keyinput116), .B1(n9137), .B2(keyinput58), 
        .ZN(n9136) );
  OAI221_X1 U10479 ( .B1(n9138), .B2(keyinput116), .C1(n9137), .C2(keyinput58), 
        .A(n9136), .ZN(n9139) );
  NOR4_X1 U10480 ( .A1(n9142), .A2(n9141), .A3(n9140), .A4(n9139), .ZN(n9155)
         );
  AOI22_X1 U10481 ( .A1(n7122), .A2(keyinput19), .B1(n7471), .B2(keyinput105), 
        .ZN(n9143) );
  OAI221_X1 U10482 ( .B1(n7122), .B2(keyinput19), .C1(n7471), .C2(keyinput105), 
        .A(n9143), .ZN(n9153) );
  INV_X1 U10483 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10059) );
  AOI22_X1 U10484 ( .A1(n9145), .A2(keyinput108), .B1(n10059), .B2(keyinput87), 
        .ZN(n9144) );
  OAI221_X1 U10485 ( .B1(n9145), .B2(keyinput108), .C1(n10059), .C2(keyinput87), .A(n9144), .ZN(n9152) );
  INV_X1 U10486 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10053) );
  AOI22_X1 U10487 ( .A1(n10053), .A2(keyinput22), .B1(keyinput74), .B2(n9147), 
        .ZN(n9146) );
  OAI221_X1 U10488 ( .B1(n10053), .B2(keyinput22), .C1(n9147), .C2(keyinput74), 
        .A(n9146), .ZN(n9151) );
  XNOR2_X1 U10489 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput11), .ZN(n9149) );
  XNOR2_X1 U10490 ( .A(keyinput127), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9148) );
  NAND2_X1 U10491 ( .A1(n9149), .A2(n9148), .ZN(n9150) );
  NOR4_X1 U10492 ( .A1(n9153), .A2(n9152), .A3(n9151), .A4(n9150), .ZN(n9154)
         );
  NAND4_X1 U10493 ( .A1(n9157), .A2(n9156), .A3(n9155), .A4(n9154), .ZN(n9316)
         );
  INV_X1 U10494 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10200) );
  AOI22_X1 U10495 ( .A1(n10200), .A2(keyinput49), .B1(n9159), .B2(keyinput3), 
        .ZN(n9158) );
  OAI221_X1 U10496 ( .B1(n10200), .B2(keyinput49), .C1(n9159), .C2(keyinput3), 
        .A(n9158), .ZN(n9169) );
  INV_X1 U10497 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9424) );
  AOI22_X1 U10498 ( .A1(n9161), .A2(keyinput101), .B1(n9424), .B2(keyinput107), 
        .ZN(n9160) );
  OAI221_X1 U10499 ( .B1(n9161), .B2(keyinput101), .C1(n9424), .C2(keyinput107), .A(n9160), .ZN(n9168) );
  INV_X1 U10500 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10179) );
  AOI22_X1 U10501 ( .A1(n10179), .A2(keyinput99), .B1(keyinput84), .B2(n9163), 
        .ZN(n9162) );
  OAI221_X1 U10502 ( .B1(n10179), .B2(keyinput99), .C1(n9163), .C2(keyinput84), 
        .A(n9162), .ZN(n9167) );
  INV_X1 U10503 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9165) );
  AOI22_X1 U10504 ( .A1(n7470), .A2(keyinput93), .B1(n9165), .B2(keyinput13), 
        .ZN(n9164) );
  OAI221_X1 U10505 ( .B1(n7470), .B2(keyinput93), .C1(n9165), .C2(keyinput13), 
        .A(n9164), .ZN(n9166) );
  NOR4_X1 U10506 ( .A1(n9169), .A2(n9168), .A3(n9167), .A4(n9166), .ZN(n9208)
         );
  INV_X1 U10507 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9171) );
  AOI22_X1 U10508 ( .A1(n10184), .A2(keyinput45), .B1(keyinput102), .B2(n9171), 
        .ZN(n9170) );
  OAI221_X1 U10509 ( .B1(n10184), .B2(keyinput45), .C1(n9171), .C2(keyinput102), .A(n9170), .ZN(n9181) );
  INV_X1 U10510 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U10511 ( .A1(n9173), .A2(keyinput72), .B1(keyinput106), .B2(n10317), 
        .ZN(n9172) );
  OAI221_X1 U10512 ( .B1(n9173), .B2(keyinput72), .C1(n10317), .C2(keyinput106), .A(n9172), .ZN(n9180) );
  AOI22_X1 U10513 ( .A1(n10208), .A2(keyinput17), .B1(n9175), .B2(keyinput124), 
        .ZN(n9174) );
  OAI221_X1 U10514 ( .B1(n10208), .B2(keyinput17), .C1(n9175), .C2(keyinput124), .A(n9174), .ZN(n9179) );
  XOR2_X1 U10515 ( .A(n6405), .B(keyinput14), .Z(n9177) );
  XNOR2_X1 U10516 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput97), .ZN(n9176) );
  NAND2_X1 U10517 ( .A1(n9177), .A2(n9176), .ZN(n9178) );
  NOR4_X1 U10518 ( .A1(n9181), .A2(n9180), .A3(n9179), .A4(n9178), .ZN(n9207)
         );
  INV_X1 U10519 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10178) );
  INV_X1 U10520 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9183) );
  AOI22_X1 U10521 ( .A1(n10178), .A2(keyinput103), .B1(n9183), .B2(keyinput76), 
        .ZN(n9182) );
  OAI221_X1 U10522 ( .B1(n10178), .B2(keyinput103), .C1(n9183), .C2(keyinput76), .A(n9182), .ZN(n9192) );
  AOI22_X1 U10523 ( .A1(n5446), .A2(keyinput118), .B1(keyinput25), .B2(n9185), 
        .ZN(n9184) );
  OAI221_X1 U10524 ( .B1(n5446), .B2(keyinput118), .C1(n9185), .C2(keyinput25), 
        .A(n9184), .ZN(n9191) );
  XOR2_X1 U10525 ( .A(n5178), .B(keyinput85), .Z(n9189) );
  XNOR2_X1 U10526 ( .A(keyinput100), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9188) );
  XNOR2_X1 U10527 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput80), .ZN(n9187) );
  XNOR2_X1 U10528 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput91), .ZN(n9186) );
  NAND4_X1 U10529 ( .A1(n9189), .A2(n9188), .A3(n9187), .A4(n9186), .ZN(n9190)
         );
  NOR3_X1 U10530 ( .A1(n9192), .A2(n9191), .A3(n9190), .ZN(n9206) );
  INV_X1 U10531 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9194) );
  INV_X1 U10532 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10272) );
  AOI22_X1 U10533 ( .A1(n9194), .A2(keyinput7), .B1(keyinput121), .B2(n10272), 
        .ZN(n9193) );
  OAI221_X1 U10534 ( .B1(n9194), .B2(keyinput7), .C1(n10272), .C2(keyinput121), 
        .A(n9193), .ZN(n9204) );
  INV_X1 U10535 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10055) );
  AOI22_X1 U10536 ( .A1(n10055), .A2(keyinput79), .B1(keyinput33), .B2(n9196), 
        .ZN(n9195) );
  OAI221_X1 U10537 ( .B1(n10055), .B2(keyinput79), .C1(n9196), .C2(keyinput33), 
        .A(n9195), .ZN(n9203) );
  INV_X1 U10538 ( .A(P2_RD_REG_SCAN_IN), .ZN(n9198) );
  AOI22_X1 U10539 ( .A1(n9198), .A2(keyinput123), .B1(keyinput83), .B2(n8365), 
        .ZN(n9197) );
  OAI221_X1 U10540 ( .B1(n9198), .B2(keyinput123), .C1(n8365), .C2(keyinput83), 
        .A(n9197), .ZN(n9202) );
  AOI22_X1 U10541 ( .A1(n9200), .A2(keyinput113), .B1(n10058), .B2(keyinput96), 
        .ZN(n9199) );
  OAI221_X1 U10542 ( .B1(n9200), .B2(keyinput113), .C1(n10058), .C2(keyinput96), .A(n9199), .ZN(n9201) );
  NOR4_X1 U10543 ( .A1(n9204), .A2(n9203), .A3(n9202), .A4(n9201), .ZN(n9205)
         );
  NAND4_X1 U10544 ( .A1(n9208), .A2(n9207), .A3(n9206), .A4(n9205), .ZN(n9315)
         );
  AOI22_X1 U10545 ( .A1(n7660), .A2(keyinput112), .B1(n9210), .B2(keyinput109), 
        .ZN(n9209) );
  OAI221_X1 U10546 ( .B1(n7660), .B2(keyinput112), .C1(n9210), .C2(keyinput109), .A(n9209), .ZN(n9221) );
  INV_X1 U10547 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10351) );
  AOI22_X1 U10548 ( .A1(n10351), .A2(keyinput71), .B1(n9212), .B2(keyinput12), 
        .ZN(n9211) );
  OAI221_X1 U10549 ( .B1(n10351), .B2(keyinput71), .C1(n9212), .C2(keyinput12), 
        .A(n9211), .ZN(n9220) );
  INV_X1 U10550 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9214) );
  AOI22_X1 U10551 ( .A1(n9215), .A2(keyinput1), .B1(n9214), .B2(keyinput47), 
        .ZN(n9213) );
  OAI221_X1 U10552 ( .B1(n9215), .B2(keyinput1), .C1(n9214), .C2(keyinput47), 
        .A(n9213), .ZN(n9219) );
  XNOR2_X1 U10553 ( .A(P2_REG0_REG_22__SCAN_IN), .B(keyinput78), .ZN(n9217) );
  XNOR2_X1 U10554 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput122), .ZN(n9216)
         );
  NAND2_X1 U10555 ( .A1(n9217), .A2(n9216), .ZN(n9218) );
  NOR4_X1 U10556 ( .A1(n9221), .A2(n9220), .A3(n9219), .A4(n9218), .ZN(n9263)
         );
  INV_X1 U10557 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10177) );
  AOI22_X1 U10558 ( .A1(n10177), .A2(keyinput60), .B1(keyinput38), .B2(n8122), 
        .ZN(n9222) );
  OAI221_X1 U10559 ( .B1(n10177), .B2(keyinput60), .C1(n8122), .C2(keyinput38), 
        .A(n9222), .ZN(n9233) );
  AOI22_X1 U10560 ( .A1(n9225), .A2(keyinput23), .B1(n9224), .B2(keyinput43), 
        .ZN(n9223) );
  OAI221_X1 U10561 ( .B1(n9225), .B2(keyinput23), .C1(n9224), .C2(keyinput43), 
        .A(n9223), .ZN(n9232) );
  XOR2_X1 U10562 ( .A(n9226), .B(keyinput57), .Z(n9230) );
  XNOR2_X1 U10563 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput15), .ZN(n9229) );
  XNOR2_X1 U10564 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput92), .ZN(n9228) );
  XNOR2_X1 U10565 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(keyinput2), .ZN(n9227) );
  NAND4_X1 U10566 ( .A1(n9230), .A2(n9229), .A3(n9228), .A4(n9227), .ZN(n9231)
         );
  NOR3_X1 U10567 ( .A1(n9233), .A2(n9232), .A3(n9231), .ZN(n9262) );
  AOI22_X1 U10568 ( .A1(n5898), .A2(keyinput29), .B1(n9235), .B2(keyinput42), 
        .ZN(n9234) );
  OAI221_X1 U10569 ( .B1(n5898), .B2(keyinput29), .C1(n9235), .C2(keyinput42), 
        .A(n9234), .ZN(n9245) );
  AOI22_X1 U10570 ( .A1(n4527), .A2(keyinput27), .B1(n9237), .B2(keyinput18), 
        .ZN(n9236) );
  OAI221_X1 U10571 ( .B1(n4527), .B2(keyinput27), .C1(n9237), .C2(keyinput18), 
        .A(n9236), .ZN(n9244) );
  INV_X1 U10572 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10057) );
  AOI22_X1 U10573 ( .A1(n7310), .A2(keyinput75), .B1(n10057), .B2(keyinput68), 
        .ZN(n9238) );
  OAI221_X1 U10574 ( .B1(n7310), .B2(keyinput75), .C1(n10057), .C2(keyinput68), 
        .A(n9238), .ZN(n9243) );
  AOI22_X1 U10575 ( .A1(n9241), .A2(keyinput39), .B1(n9240), .B2(keyinput67), 
        .ZN(n9239) );
  OAI221_X1 U10576 ( .B1(n9241), .B2(keyinput39), .C1(n9240), .C2(keyinput67), 
        .A(n9239), .ZN(n9242) );
  NOR4_X1 U10577 ( .A1(n9245), .A2(n9244), .A3(n9243), .A4(n9242), .ZN(n9261)
         );
  AOI22_X1 U10578 ( .A1(n6278), .A2(keyinput53), .B1(keyinput40), .B2(n9247), 
        .ZN(n9246) );
  OAI221_X1 U10579 ( .B1(n6278), .B2(keyinput53), .C1(n9247), .C2(keyinput40), 
        .A(n9246), .ZN(n9259) );
  AOI22_X1 U10580 ( .A1(n9250), .A2(keyinput111), .B1(keyinput41), .B2(n9249), 
        .ZN(n9248) );
  OAI221_X1 U10581 ( .B1(n9250), .B2(keyinput111), .C1(n9249), .C2(keyinput41), 
        .A(n9248), .ZN(n9258) );
  AOI22_X1 U10582 ( .A1(n9253), .A2(keyinput8), .B1(keyinput34), .B2(n9252), 
        .ZN(n9251) );
  OAI221_X1 U10583 ( .B1(n9253), .B2(keyinput8), .C1(n9252), .C2(keyinput34), 
        .A(n9251), .ZN(n9257) );
  XNOR2_X1 U10584 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput62), .ZN(n9255) );
  XNOR2_X1 U10585 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput126), .ZN(n9254) );
  NAND2_X1 U10586 ( .A1(n9255), .A2(n9254), .ZN(n9256) );
  NOR4_X1 U10587 ( .A1(n9259), .A2(n9258), .A3(n9257), .A4(n9256), .ZN(n9260)
         );
  NAND4_X1 U10588 ( .A1(n9263), .A2(n9262), .A3(n9261), .A4(n9260), .ZN(n9314)
         );
  INV_X1 U10589 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U10590 ( .A1(n10128), .A2(keyinput65), .B1(keyinput115), .B2(n10176), .ZN(n9264) );
  OAI221_X1 U10591 ( .B1(n10128), .B2(keyinput65), .C1(n10176), .C2(
        keyinput115), .A(n9264), .ZN(n9274) );
  INV_X1 U10592 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10054) );
  AOI22_X1 U10593 ( .A1(n10054), .A2(keyinput4), .B1(keyinput10), .B2(n9266), 
        .ZN(n9265) );
  OAI221_X1 U10594 ( .B1(n10054), .B2(keyinput4), .C1(n9266), .C2(keyinput10), 
        .A(n9265), .ZN(n9273) );
  AOI22_X1 U10595 ( .A1(n10068), .A2(keyinput81), .B1(n9268), .B2(keyinput104), 
        .ZN(n9267) );
  OAI221_X1 U10596 ( .B1(n10068), .B2(keyinput81), .C1(n9268), .C2(keyinput104), .A(n9267), .ZN(n9272) );
  XNOR2_X1 U10597 ( .A(P1_REG1_REG_26__SCAN_IN), .B(keyinput95), .ZN(n9270) );
  XNOR2_X1 U10598 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput56), .ZN(n9269) );
  NAND2_X1 U10599 ( .A1(n9270), .A2(n9269), .ZN(n9271) );
  NOR4_X1 U10600 ( .A1(n9274), .A2(n9273), .A3(n9272), .A4(n9271), .ZN(n9312)
         );
  INV_X1 U10601 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9276) );
  AOI22_X1 U10602 ( .A1(keyinput51), .A2(n9276), .B1(keyinput89), .B2(n5952), 
        .ZN(n9275) );
  OAI21_X1 U10603 ( .B1(n9276), .B2(keyinput51), .A(n9275), .ZN(n9284) );
  AOI22_X1 U10604 ( .A1(n5049), .A2(keyinput77), .B1(keyinput24), .B2(n7776), 
        .ZN(n9277) );
  OAI221_X1 U10605 ( .B1(n5049), .B2(keyinput77), .C1(n7776), .C2(keyinput24), 
        .A(n9277), .ZN(n9283) );
  AOI22_X1 U10606 ( .A1(n6360), .A2(keyinput52), .B1(n9279), .B2(keyinput86), 
        .ZN(n9278) );
  OAI221_X1 U10607 ( .B1(n6360), .B2(keyinput52), .C1(n9279), .C2(keyinput86), 
        .A(n9278), .ZN(n9282) );
  AOI22_X1 U10608 ( .A1(n7069), .A2(keyinput46), .B1(n9374), .B2(keyinput69), 
        .ZN(n9280) );
  OAI221_X1 U10609 ( .B1(n7069), .B2(keyinput46), .C1(n9374), .C2(keyinput69), 
        .A(n9280), .ZN(n9281) );
  NOR4_X1 U10610 ( .A1(n9284), .A2(n9283), .A3(n9282), .A4(n9281), .ZN(n9311)
         );
  AOI22_X1 U10611 ( .A1(n4619), .A2(keyinput37), .B1(keyinput36), .B2(n9286), 
        .ZN(n9285) );
  OAI221_X1 U10612 ( .B1(n4619), .B2(keyinput37), .C1(n9286), .C2(keyinput36), 
        .A(n9285), .ZN(n9298) );
  INV_X1 U10613 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9289) );
  INV_X1 U10614 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9288) );
  AOI22_X1 U10615 ( .A1(n9289), .A2(keyinput6), .B1(keyinput26), .B2(n9288), 
        .ZN(n9287) );
  OAI221_X1 U10616 ( .B1(n9289), .B2(keyinput6), .C1(n9288), .C2(keyinput26), 
        .A(n9287), .ZN(n9297) );
  AOI22_X1 U10617 ( .A1(n9292), .A2(keyinput119), .B1(n9291), .B2(keyinput88), 
        .ZN(n9290) );
  OAI221_X1 U10618 ( .B1(n9292), .B2(keyinput119), .C1(n9291), .C2(keyinput88), 
        .A(n9290), .ZN(n9296) );
  XNOR2_X1 U10619 ( .A(P2_REG0_REG_19__SCAN_IN), .B(keyinput28), .ZN(n9294) );
  XNOR2_X1 U10620 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput30), .ZN(n9293) );
  NAND2_X1 U10621 ( .A1(n9294), .A2(n9293), .ZN(n9295) );
  NOR4_X1 U10622 ( .A1(n9298), .A2(n9297), .A3(n9296), .A4(n9295), .ZN(n9310)
         );
  AOI22_X1 U10623 ( .A1(n9300), .A2(keyinput59), .B1(n5877), .B2(keyinput32), 
        .ZN(n9299) );
  OAI221_X1 U10624 ( .B1(n9300), .B2(keyinput59), .C1(n5877), .C2(keyinput32), 
        .A(n9299), .ZN(n9308) );
  INV_X1 U10625 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10060) );
  XNOR2_X1 U10626 ( .A(keyinput35), .B(n10060), .ZN(n9307) );
  XNOR2_X1 U10627 ( .A(keyinput90), .B(n9078), .ZN(n9306) );
  XNOR2_X1 U10628 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput114), .ZN(n9304) );
  XNOR2_X1 U10629 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput98), .ZN(n9303) );
  XNOR2_X1 U10630 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput63), .ZN(n9302) );
  XNOR2_X1 U10631 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput120), .ZN(n9301) );
  NAND4_X1 U10632 ( .A1(n9304), .A2(n9303), .A3(n9302), .A4(n9301), .ZN(n9305)
         );
  NOR4_X1 U10633 ( .A1(n9308), .A2(n9307), .A3(n9306), .A4(n9305), .ZN(n9309)
         );
  NAND4_X1 U10634 ( .A1(n9312), .A2(n9311), .A3(n9310), .A4(n9309), .ZN(n9313)
         );
  NOR4_X1 U10635 ( .A1(n9316), .A2(n9315), .A3(n9314), .A4(n9313), .ZN(n9317)
         );
  OAI221_X1 U10636 ( .B1(keyinput89), .B2(n5952), .C1(keyinput89), .C2(n9318), 
        .A(n9317), .ZN(n9324) );
  AOI222_X1 U10637 ( .A1(n9322), .A2(n9321), .B1(P1_DATAO_REG_9__SCAN_IN), 
        .B2(n9320), .C1(n9319), .C2(P2_STATE_REG_SCAN_IN), .ZN(n9323) );
  XOR2_X1 U10638 ( .A(n9324), .B(n9323), .Z(P2_U3349) );
  MUX2_X1 U10639 ( .A(n9325), .B(n10173), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3358) );
  INV_X1 U10640 ( .A(n9328), .ZN(n9329) );
  OAI21_X1 U10641 ( .B1(n9330), .B2(n9329), .A(n9448), .ZN(n9335) );
  NOR2_X1 U10642 ( .A1(n9467), .A2(n9582), .ZN(n9333) );
  OAI22_X1 U10643 ( .A1(n9451), .A2(n9612), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9331), .ZN(n9332) );
  AOI211_X1 U10644 ( .C1(n9585), .C2(n9462), .A(n9333), .B(n9332), .ZN(n9334)
         );
  INV_X1 U10645 ( .A(n9758), .ZN(n9639) );
  AND3_X1 U10646 ( .A1(n9336), .A2(n9337), .A3(n9420), .ZN(n9340) );
  INV_X1 U10647 ( .A(n9401), .ZN(n9342) );
  OAI21_X1 U10648 ( .B1(n9400), .B2(n9340), .A(n9339), .ZN(n9341) );
  OAI211_X1 U10649 ( .C1(n9342), .C2(n9400), .A(n9448), .B(n9341), .ZN(n9346)
         );
  AOI22_X1 U10650 ( .A1(n9464), .A2(n9477), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9343) );
  OAI21_X1 U10651 ( .B1(n9643), .B2(n9467), .A(n9343), .ZN(n9344) );
  AOI21_X1 U10652 ( .B1(n9637), .B2(n9462), .A(n9344), .ZN(n9345) );
  OAI211_X1 U10653 ( .C1(n9639), .C2(n9456), .A(n9346), .B(n9345), .ZN(
        P1_U3214) );
  XNOR2_X1 U10654 ( .A(n9358), .B(n9354), .ZN(n9347) );
  XNOR2_X1 U10655 ( .A(n9356), .B(n9347), .ZN(n9353) );
  NOR2_X1 U10656 ( .A1(n9437), .A2(n9689), .ZN(n9351) );
  NAND2_X1 U10657 ( .A1(n9696), .A2(n9464), .ZN(n9349) );
  OAI211_X1 U10658 ( .C1(n9666), .C2(n9467), .A(n9349), .B(n9348), .ZN(n9350)
         );
  OAI21_X1 U10659 ( .B1(n9353), .B2(n9472), .A(n9352), .ZN(P1_U3217) );
  INV_X1 U10660 ( .A(n9356), .ZN(n9359) );
  OAI21_X1 U10661 ( .B1(n9356), .B2(n9355), .A(n9354), .ZN(n9357) );
  OAI21_X1 U10662 ( .B1(n9359), .B2(n9358), .A(n9357), .ZN(n9412) );
  NAND2_X1 U10663 ( .A1(n9360), .A2(n9361), .ZN(n9413) );
  NOR2_X1 U10664 ( .A1(n9412), .A2(n9413), .ZN(n9411) );
  INV_X1 U10665 ( .A(n9361), .ZN(n9363) );
  NOR3_X1 U10666 ( .A1(n9411), .A2(n9363), .A3(n9362), .ZN(n9364) );
  OAI21_X1 U10667 ( .B1(n9364), .B2(n4444), .A(n9448), .ZN(n9368) );
  AOI22_X1 U10668 ( .A1(n9697), .A2(n9464), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9365) );
  OAI21_X1 U10669 ( .B1(n9667), .B2(n9467), .A(n9365), .ZN(n9366) );
  AOI21_X1 U10670 ( .B1(n9670), .B2(n9462), .A(n9366), .ZN(n9367) );
  OAI211_X1 U10671 ( .C1(n9369), .C2(n9456), .A(n9368), .B(n9367), .ZN(
        P1_U3221) );
  INV_X1 U10672 ( .A(n9370), .ZN(n9371) );
  OR2_X1 U10673 ( .A1(n9371), .A2(n9372), .ZN(n9399) );
  OAI21_X1 U10674 ( .B1(n9373), .B2(n9446), .A(n9448), .ZN(n9378) );
  NOR2_X1 U10675 ( .A1(n9467), .A2(n9612), .ZN(n9376) );
  OAI22_X1 U10676 ( .A1(n9451), .A2(n9643), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9374), .ZN(n9375) );
  AOI211_X1 U10677 ( .C1(n9617), .C2(n9462), .A(n9376), .B(n9375), .ZN(n9377)
         );
  OAI211_X1 U10678 ( .C1(n8277), .C2(n9456), .A(n9378), .B(n9377), .ZN(
        P1_U3223) );
  NOR2_X1 U10679 ( .A1(n4921), .A2(n9380), .ZN(n9381) );
  XNOR2_X1 U10680 ( .A(n9382), .B(n9381), .ZN(n9390) );
  NOR2_X1 U10681 ( .A1(n9383), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9521) );
  NOR2_X1 U10682 ( .A1(n9451), .A2(n9384), .ZN(n9385) );
  AOI211_X1 U10683 ( .C1(n9440), .C2(n9716), .A(n9521), .B(n9385), .ZN(n9386)
         );
  OAI21_X1 U10684 ( .B1(n9437), .B2(n9387), .A(n9386), .ZN(n9388) );
  AOI21_X1 U10685 ( .B1(n9795), .B2(n9470), .A(n9388), .ZN(n9389) );
  OAI21_X1 U10686 ( .B1(n9390), .B2(n9472), .A(n9389), .ZN(P1_U3224) );
  XOR2_X1 U10687 ( .A(n9392), .B(n9391), .Z(n9398) );
  NAND2_X1 U10688 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9527) );
  OAI21_X1 U10689 ( .B1(n9451), .B2(n9468), .A(n9527), .ZN(n9393) );
  AOI21_X1 U10690 ( .B1(n9440), .B2(n9696), .A(n9393), .ZN(n9394) );
  OAI21_X1 U10691 ( .B1(n9437), .B2(n9395), .A(n9394), .ZN(n9396) );
  AOI21_X1 U10692 ( .B1(n9790), .B2(n9470), .A(n9396), .ZN(n9397) );
  OAI21_X1 U10693 ( .B1(n9398), .B2(n9472), .A(n9397), .ZN(P1_U3226) );
  INV_X1 U10694 ( .A(n9755), .ZN(n9410) );
  OAI21_X1 U10695 ( .B1(n9401), .B2(n9400), .A(n9399), .ZN(n9402) );
  INV_X1 U10696 ( .A(n9402), .ZN(n9403) );
  OAI21_X1 U10697 ( .B1(n9404), .B2(n9403), .A(n9448), .ZN(n9409) );
  NOR2_X1 U10698 ( .A1(n9467), .A2(n9625), .ZN(n9407) );
  OAI22_X1 U10699 ( .A1(n9451), .A2(n9624), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9405), .ZN(n9406) );
  AOI211_X1 U10700 ( .C1(n9627), .C2(n9462), .A(n9407), .B(n9406), .ZN(n9408)
         );
  OAI211_X1 U10701 ( .C1(n9410), .C2(n9456), .A(n9409), .B(n9408), .ZN(
        P1_U3227) );
  AOI21_X1 U10702 ( .B1(n9413), .B2(n9412), .A(n9411), .ZN(n9418) );
  AOI22_X1 U10703 ( .A1(n9717), .A2(n9464), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9415) );
  NAND2_X1 U10704 ( .A1(n9462), .A2(n9678), .ZN(n9414) );
  OAI211_X1 U10705 ( .C1(n9478), .C2(n9467), .A(n9415), .B(n9414), .ZN(n9416)
         );
  AOI21_X1 U10706 ( .B1(n9773), .B2(n9470), .A(n9416), .ZN(n9417) );
  OAI21_X1 U10707 ( .B1(n9418), .B2(n9472), .A(n9417), .ZN(P1_U3231) );
  NAND2_X1 U10708 ( .A1(n9420), .A2(n9419), .ZN(n9422) );
  XNOR2_X1 U10709 ( .A(n9422), .B(n9421), .ZN(n9423) );
  NAND2_X1 U10710 ( .A1(n9423), .A2(n9448), .ZN(n9428) );
  NOR2_X1 U10711 ( .A1(n9467), .A2(n9624), .ZN(n9426) );
  OAI22_X1 U10712 ( .A1(n9478), .A2(n9451), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9424), .ZN(n9425) );
  AOI211_X1 U10713 ( .C1(n9652), .C2(n9462), .A(n9426), .B(n9425), .ZN(n9427)
         );
  OAI211_X1 U10714 ( .C1(n9654), .C2(n9456), .A(n9428), .B(n9427), .ZN(
        P1_U3233) );
  INV_X1 U10715 ( .A(n9431), .ZN(n9435) );
  AOI21_X1 U10716 ( .B1(n9431), .B2(n9430), .A(n9429), .ZN(n9432) );
  NOR2_X1 U10717 ( .A1(n9432), .A2(n9472), .ZN(n9433) );
  OAI21_X1 U10718 ( .B1(n9435), .B2(n9434), .A(n9433), .ZN(n9442) );
  NAND2_X1 U10719 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9949) );
  OAI21_X1 U10720 ( .B1(n9436), .B2(n9451), .A(n9949), .ZN(n9439) );
  NOR2_X1 U10721 ( .A1(n9437), .A2(n9707), .ZN(n9438) );
  AOI211_X1 U10722 ( .C1(n9440), .C2(n9717), .A(n9439), .B(n9438), .ZN(n9441)
         );
  OAI211_X1 U10723 ( .C1(n9711), .C2(n9456), .A(n9442), .B(n9441), .ZN(
        P1_U3236) );
  INV_X1 U10724 ( .A(n9443), .ZN(n9449) );
  OAI21_X1 U10725 ( .B1(n9446), .B2(n9445), .A(n9444), .ZN(n9447) );
  NAND3_X1 U10726 ( .A1(n9449), .A2(n9448), .A3(n9447), .ZN(n9455) );
  NOR2_X1 U10727 ( .A1(n9467), .A2(n9602), .ZN(n9453) );
  INV_X1 U10728 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9450) );
  OAI22_X1 U10729 ( .A1(n9451), .A2(n9625), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9450), .ZN(n9452) );
  AOI211_X1 U10730 ( .C1(n9596), .C2(n9462), .A(n9453), .B(n9452), .ZN(n9454)
         );
  OAI211_X1 U10731 ( .C1(n9598), .C2(n9456), .A(n9455), .B(n9454), .ZN(
        P1_U3238) );
  NAND2_X1 U10732 ( .A1(n9458), .A2(n9457), .ZN(n9459) );
  XOR2_X1 U10733 ( .A(n9460), .B(n9459), .Z(n9473) );
  NAND2_X1 U10734 ( .A1(n9462), .A2(n9461), .ZN(n9466) );
  NOR2_X1 U10735 ( .A1(n9463), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9510) );
  AOI21_X1 U10736 ( .B1(n9464), .B2(n9481), .A(n9510), .ZN(n9465) );
  OAI211_X1 U10737 ( .C1(n9468), .C2(n9467), .A(n9466), .B(n9465), .ZN(n9469)
         );
  AOI21_X1 U10738 ( .B1(n9798), .B2(n9470), .A(n9469), .ZN(n9471) );
  OAI21_X1 U10739 ( .B1(n9473), .B2(n9472), .A(n9471), .ZN(P1_U3239) );
  MUX2_X1 U10740 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9554), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10741 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9553), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10742 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9474), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10743 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9475), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10744 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9476), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10745 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9657), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10746 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9477), .S(P1_U4006), .Z(
        P1_U3577) );
  INV_X1 U10747 ( .A(n9478), .ZN(n9682) );
  MUX2_X1 U10748 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9682), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10749 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9697), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10750 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9717), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10751 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9696), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10752 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9716), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10753 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9479), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10754 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9480), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10755 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9481), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10756 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9482), .S(P1_U4006), .Z(
        P1_U3568) );
  INV_X1 U10757 ( .A(n9483), .ZN(n9484) );
  MUX2_X1 U10758 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9484), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10759 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9485), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10760 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9486), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10761 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9487), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10762 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9488), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10763 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n5406), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10764 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9489), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10765 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n10038), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10766 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n5364), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10767 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n7554), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10768 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9490), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10769 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n5818), .S(P1_U4006), .Z(
        P1_U3556) );
  NAND2_X1 U10770 ( .A1(n9961), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n9500) );
  NAND3_X1 U10771 ( .A1(n9962), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6730), .ZN(
        n9499) );
  OR2_X1 U10772 ( .A1(n9920), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9491) );
  NAND2_X1 U10773 ( .A1(n9492), .A2(n9491), .ZN(n9924) );
  XNOR2_X1 U10774 ( .A(n9924), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9495) );
  AOI21_X1 U10775 ( .B1(n9920), .B2(n6730), .A(P1_U3084), .ZN(n9494) );
  NAND4_X1 U10776 ( .A1(n9496), .A2(n9495), .A3(n9494), .A4(n9493), .ZN(n9498)
         );
  NAND2_X1 U10777 ( .A1(P1_U3084), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9497) );
  NAND4_X1 U10778 ( .A1(n9500), .A2(n9499), .A3(n9498), .A4(n9497), .ZN(
        P1_U3241) );
  INV_X1 U10779 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9514) );
  INV_X1 U10780 ( .A(n9501), .ZN(n9504) );
  INV_X1 U10781 ( .A(n9502), .ZN(n9503) );
  OAI211_X1 U10782 ( .C1(n9504), .C2(P1_REG1_REG_15__SCAN_IN), .A(n9962), .B(
        n9503), .ZN(n9513) );
  INV_X1 U10783 ( .A(n9505), .ZN(n9511) );
  AOI211_X1 U10784 ( .C1(n9508), .C2(n9507), .A(n9506), .B(n9950), .ZN(n9509)
         );
  AOI211_X1 U10785 ( .C1(n9957), .C2(n9511), .A(n9510), .B(n9509), .ZN(n9512)
         );
  OAI211_X1 U10786 ( .C1(n9947), .C2(n9514), .A(n9513), .B(n9512), .ZN(
        P1_U3256) );
  AOI211_X1 U10787 ( .C1(n9517), .C2(n9516), .A(n9515), .B(n9950), .ZN(n9526)
         );
  AOI211_X1 U10788 ( .C1(n9520), .C2(n9519), .A(n9518), .B(n9533), .ZN(n9525)
         );
  AOI21_X1 U10789 ( .B1(n9957), .B2(n9522), .A(n9521), .ZN(n9523) );
  OAI21_X1 U10790 ( .B1(n9947), .B2(n9171), .A(n9523), .ZN(n9524) );
  OR3_X1 U10791 ( .A1(n9526), .A2(n9525), .A3(n9524), .ZN(P1_U3257) );
  INV_X1 U10792 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9540) );
  INV_X1 U10793 ( .A(n9527), .ZN(n9531) );
  AOI211_X1 U10794 ( .C1(n9529), .C2(n9528), .A(n4461), .B(n9950), .ZN(n9530)
         );
  AOI211_X1 U10795 ( .C1(n9957), .C2(n9532), .A(n9531), .B(n9530), .ZN(n9539)
         );
  AOI211_X1 U10796 ( .C1(n9536), .C2(n9535), .A(n9534), .B(n9533), .ZN(n9537)
         );
  INV_X1 U10797 ( .A(n9537), .ZN(n9538) );
  OAI211_X1 U10798 ( .C1(n9947), .C2(n9540), .A(n9539), .B(n9538), .ZN(
        P1_U3258) );
  OAI21_X1 U10799 ( .B1(n9542), .B2(n9560), .A(n9541), .ZN(n9729) );
  NOR2_X1 U10800 ( .A1(n9542), .A2(n9710), .ZN(n9543) );
  AOI211_X1 U10801 ( .C1(n10047), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9544), .B(
        n9543), .ZN(n9545) );
  OAI21_X1 U10802 ( .B1(n9729), .B2(n9573), .A(n9545), .ZN(P1_U3262) );
  XNOR2_X1 U10803 ( .A(n9547), .B(n9549), .ZN(n9730) );
  INV_X1 U10804 ( .A(n9730), .ZN(n9566) );
  AOI22_X1 U10805 ( .A1(n9731), .A2(n10050), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n10047), .ZN(n9565) );
  INV_X1 U10806 ( .A(n9549), .ZN(n9548) );
  NAND4_X1 U10807 ( .A1(n9551), .A2(n9548), .A3(n9550), .A4(n10043), .ZN(n9558) );
  NAND3_X1 U10808 ( .A1(n9570), .A2(n9582), .A3(n10043), .ZN(n9552) );
  OR2_X1 U10809 ( .A1(n9548), .A2(n9552), .ZN(n9557) );
  AOI22_X1 U10810 ( .A1(n9555), .A2(n9554), .B1(n9553), .B2(n9715), .ZN(n9556)
         );
  NAND3_X1 U10811 ( .A1(n9559), .A2(n9558), .A3(n5023), .ZN(n9735) );
  AOI211_X1 U10812 ( .C1(n9731), .C2(n5035), .A(n10121), .B(n9560), .ZN(n9733)
         );
  INV_X1 U10813 ( .A(n9733), .ZN(n9562) );
  OAI22_X1 U10814 ( .A1(n9562), .A2(n10011), .B1(n10031), .B2(n9561), .ZN(
        n9563) );
  OAI21_X1 U10815 ( .B1(n9735), .B2(n9563), .A(n10033), .ZN(n9564) );
  OAI211_X1 U10816 ( .C1(n9566), .C2(n9722), .A(n9565), .B(n9564), .ZN(
        P1_U3355) );
  NAND2_X1 U10817 ( .A1(n9567), .A2(n10033), .ZN(n9579) );
  INV_X1 U10818 ( .A(n9568), .ZN(n9577) );
  INV_X1 U10819 ( .A(n9722), .ZN(n9576) );
  AOI22_X1 U10820 ( .A1(n10047), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9569), 
        .B2(n10009), .ZN(n9572) );
  NAND2_X1 U10821 ( .A1(n9570), .A2(n10050), .ZN(n9571) );
  OAI211_X1 U10822 ( .C1(n9574), .C2(n9573), .A(n9572), .B(n9571), .ZN(n9575)
         );
  AOI21_X1 U10823 ( .B1(n9577), .B2(n9576), .A(n9575), .ZN(n9578) );
  NAND2_X1 U10824 ( .A1(n9579), .A2(n9578), .ZN(P1_U3263) );
  AOI211_X1 U10825 ( .C1(n9581), .C2(n9589), .A(n10014), .B(n9580), .ZN(n9584)
         );
  OAI22_X1 U10826 ( .A1(n9612), .A2(n10040), .B1(n9582), .B2(n10018), .ZN(
        n9583) );
  AOI211_X1 U10827 ( .C1(n9739), .C2(n4976), .A(n10121), .B(n4391), .ZN(n9738)
         );
  AOI22_X1 U10828 ( .A1(n10047), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9585), 
        .B2(n10009), .ZN(n9586) );
  OAI21_X1 U10829 ( .B1(n9587), .B2(n9710), .A(n9586), .ZN(n9588) );
  AOI21_X1 U10830 ( .B1(n9738), .B2(n9616), .A(n9588), .ZN(n9592) );
  XNOR2_X1 U10831 ( .A(n9590), .B(n9589), .ZN(n9742) );
  OR2_X1 U10832 ( .A1(n9742), .A2(n9722), .ZN(n9591) );
  OAI211_X1 U10833 ( .C1(n9741), .C2(n10047), .A(n9592), .B(n9591), .ZN(
        P1_U3264) );
  XNOR2_X1 U10834 ( .A(n9594), .B(n9593), .ZN(n9747) );
  AOI21_X1 U10835 ( .B1(n9743), .B2(n9613), .A(n9595), .ZN(n9744) );
  AOI22_X1 U10836 ( .A1(n10047), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9596), 
        .B2(n10009), .ZN(n9597) );
  OAI21_X1 U10837 ( .B1(n9598), .B2(n9710), .A(n9597), .ZN(n9606) );
  AOI211_X1 U10838 ( .C1(n9601), .C2(n9600), .A(n10014), .B(n9599), .ZN(n9604)
         );
  OAI22_X1 U10839 ( .A1(n9625), .A2(n10040), .B1(n9602), .B2(n10018), .ZN(
        n9603) );
  NOR2_X1 U10840 ( .A1(n9604), .A2(n9603), .ZN(n9746) );
  NOR2_X1 U10841 ( .A1(n9746), .A2(n10047), .ZN(n9605) );
  AOI211_X1 U10842 ( .C1(n10028), .C2(n9744), .A(n9606), .B(n9605), .ZN(n9607)
         );
  OAI21_X1 U10843 ( .B1(n9747), .B2(n9722), .A(n9607), .ZN(P1_U3265) );
  XOR2_X1 U10844 ( .A(n9610), .B(n9608), .Z(n9752) );
  XOR2_X1 U10845 ( .A(n9610), .B(n9609), .Z(n9611) );
  OAI222_X1 U10846 ( .A1(n10018), .A2(n9612), .B1(n10040), .B2(n9643), .C1(
        n10014), .C2(n9611), .ZN(n9748) );
  INV_X1 U10847 ( .A(n9626), .ZN(n9615) );
  INV_X1 U10848 ( .A(n9613), .ZN(n9614) );
  AOI211_X1 U10849 ( .C1(n9750), .C2(n9615), .A(n10121), .B(n9614), .ZN(n9749)
         );
  NAND2_X1 U10850 ( .A1(n9749), .A2(n9616), .ZN(n9619) );
  AOI22_X1 U10851 ( .A1(n10047), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9617), 
        .B2(n10009), .ZN(n9618) );
  OAI211_X1 U10852 ( .C1(n8277), .C2(n9710), .A(n9619), .B(n9618), .ZN(n9620)
         );
  AOI21_X1 U10853 ( .B1(n9748), .B2(n10033), .A(n9620), .ZN(n9621) );
  OAI21_X1 U10854 ( .B1(n9752), .B2(n9722), .A(n9621), .ZN(P1_U3266) );
  XOR2_X1 U10855 ( .A(n9623), .B(n9622), .Z(n9757) );
  AOI22_X1 U10856 ( .A1(n9755), .A2(n10050), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10047), .ZN(n9632) );
  AOI211_X1 U10857 ( .C1(n9755), .C2(n9635), .A(n10121), .B(n9626), .ZN(n9754)
         );
  INV_X1 U10858 ( .A(n9754), .ZN(n9629) );
  INV_X1 U10859 ( .A(n9627), .ZN(n9628) );
  OAI22_X1 U10860 ( .A1(n9629), .A2(n10011), .B1(n10031), .B2(n9628), .ZN(
        n9630) );
  OAI21_X1 U10861 ( .B1(n9753), .B2(n9630), .A(n10033), .ZN(n9631) );
  OAI211_X1 U10862 ( .C1(n9757), .C2(n9722), .A(n9632), .B(n9631), .ZN(
        P1_U3267) );
  XNOR2_X1 U10863 ( .A(n9633), .B(n9634), .ZN(n9762) );
  INV_X1 U10864 ( .A(n9635), .ZN(n9636) );
  AOI21_X1 U10865 ( .B1(n9758), .B2(n9650), .A(n9636), .ZN(n9759) );
  AOI22_X1 U10866 ( .A1(n10047), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9637), 
        .B2(n10009), .ZN(n9638) );
  OAI21_X1 U10867 ( .B1(n9639), .B2(n9710), .A(n9638), .ZN(n9647) );
  AOI211_X1 U10868 ( .C1(n9642), .C2(n9641), .A(n10014), .B(n9640), .ZN(n9645)
         );
  OAI22_X1 U10869 ( .A1(n9643), .A2(n10018), .B1(n9667), .B2(n10040), .ZN(
        n9644) );
  NOR2_X1 U10870 ( .A1(n9645), .A2(n9644), .ZN(n9761) );
  NOR2_X1 U10871 ( .A1(n9761), .A2(n10047), .ZN(n9646) );
  AOI211_X1 U10872 ( .C1(n9759), .C2(n10028), .A(n9647), .B(n9646), .ZN(n9648)
         );
  OAI21_X1 U10873 ( .B1(n9762), .B2(n9722), .A(n9648), .ZN(P1_U3268) );
  XOR2_X1 U10874 ( .A(n9649), .B(n9655), .Z(n9767) );
  INV_X1 U10875 ( .A(n9668), .ZN(n9651) );
  AOI21_X1 U10876 ( .B1(n9763), .B2(n9651), .A(n4984), .ZN(n9764) );
  AOI22_X1 U10877 ( .A1(n10047), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9652), 
        .B2(n10009), .ZN(n9653) );
  OAI21_X1 U10878 ( .B1(n9654), .B2(n9710), .A(n9653), .ZN(n9660) );
  XNOR2_X1 U10879 ( .A(n9656), .B(n9655), .ZN(n9658) );
  AOI222_X1 U10880 ( .A1(n10043), .A2(n9658), .B1(n9657), .B2(n10037), .C1(
        n9682), .C2(n9715), .ZN(n9766) );
  NOR2_X1 U10881 ( .A1(n9766), .A2(n10047), .ZN(n9659) );
  AOI211_X1 U10882 ( .C1(n9764), .C2(n10028), .A(n9660), .B(n9659), .ZN(n9661)
         );
  OAI21_X1 U10883 ( .B1(n9767), .B2(n9722), .A(n9661), .ZN(P1_U3269) );
  XNOR2_X1 U10884 ( .A(n9662), .B(n9664), .ZN(n9772) );
  AOI22_X1 U10885 ( .A1(n9770), .A2(n10050), .B1(n10047), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9675) );
  XOR2_X1 U10886 ( .A(n9663), .B(n9664), .Z(n9665) );
  OAI222_X1 U10887 ( .A1(n10018), .A2(n9667), .B1(n10040), .B2(n9666), .C1(
        n10014), .C2(n9665), .ZN(n9768) );
  INV_X1 U10888 ( .A(n9677), .ZN(n9669) );
  AOI211_X1 U10889 ( .C1(n9770), .C2(n9669), .A(n10121), .B(n9668), .ZN(n9769)
         );
  INV_X1 U10890 ( .A(n9769), .ZN(n9672) );
  INV_X1 U10891 ( .A(n9670), .ZN(n9671) );
  OAI22_X1 U10892 ( .A1(n9672), .A2(n10011), .B1(n10031), .B2(n9671), .ZN(
        n9673) );
  OAI21_X1 U10893 ( .B1(n9768), .B2(n9673), .A(n10033), .ZN(n9674) );
  OAI211_X1 U10894 ( .C1(n9772), .C2(n9722), .A(n9675), .B(n9674), .ZN(
        P1_U3270) );
  XNOR2_X1 U10895 ( .A(n9676), .B(n9681), .ZN(n9777) );
  AOI21_X1 U10896 ( .B1(n9773), .B2(n9688), .A(n9677), .ZN(n9774) );
  AOI22_X1 U10897 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(n10047), .B1(n9678), 
        .B2(n10009), .ZN(n9679) );
  OAI21_X1 U10898 ( .B1(n4987), .B2(n9710), .A(n9679), .ZN(n9685) );
  XOR2_X1 U10899 ( .A(n9681), .B(n9680), .Z(n9683) );
  AOI222_X1 U10900 ( .A1(n10043), .A2(n9683), .B1(n9682), .B2(n10037), .C1(
        n9717), .C2(n9715), .ZN(n9776) );
  NOR2_X1 U10901 ( .A1(n9776), .A2(n10047), .ZN(n9684) );
  AOI211_X1 U10902 ( .C1(n9774), .C2(n10028), .A(n9685), .B(n9684), .ZN(n9686)
         );
  OAI21_X1 U10903 ( .B1(n9777), .B2(n9722), .A(n9686), .ZN(P1_U3271) );
  XNOR2_X1 U10904 ( .A(n9687), .B(n9695), .ZN(n9782) );
  AOI21_X1 U10905 ( .B1(n9778), .B2(n9704), .A(n4983), .ZN(n9779) );
  INV_X1 U10906 ( .A(n9689), .ZN(n9690) );
  AOI22_X1 U10907 ( .A1(n10047), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9690), 
        .B2(n10009), .ZN(n9691) );
  OAI21_X1 U10908 ( .B1(n9692), .B2(n9710), .A(n9691), .ZN(n9700) );
  OAI21_X1 U10909 ( .B1(n9695), .B2(n9694), .A(n9693), .ZN(n9698) );
  AOI222_X1 U10910 ( .A1(n10043), .A2(n9698), .B1(n9697), .B2(n10037), .C1(
        n9696), .C2(n9715), .ZN(n9781) );
  NOR2_X1 U10911 ( .A1(n9781), .A2(n10047), .ZN(n9699) );
  AOI211_X1 U10912 ( .C1(n9779), .C2(n10028), .A(n9700), .B(n9699), .ZN(n9701)
         );
  OAI21_X1 U10913 ( .B1(n9722), .B2(n9782), .A(n9701), .ZN(P1_U3272) );
  XNOR2_X1 U10914 ( .A(n9703), .B(n9702), .ZN(n9787) );
  INV_X1 U10915 ( .A(n8287), .ZN(n9706) );
  INV_X1 U10916 ( .A(n9704), .ZN(n9705) );
  AOI21_X1 U10917 ( .B1(n9783), .B2(n9706), .A(n9705), .ZN(n9784) );
  INV_X1 U10918 ( .A(n9707), .ZN(n9708) );
  AOI22_X1 U10919 ( .A1(n10047), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9708), 
        .B2(n10009), .ZN(n9709) );
  OAI21_X1 U10920 ( .B1(n9711), .B2(n9710), .A(n9709), .ZN(n9720) );
  OAI21_X1 U10921 ( .B1(n9714), .B2(n9713), .A(n9712), .ZN(n9718) );
  AOI222_X1 U10922 ( .A1(n10043), .A2(n9718), .B1(n9717), .B2(n10037), .C1(
        n9716), .C2(n9715), .ZN(n9786) );
  NOR2_X1 U10923 ( .A1(n9786), .A2(n10047), .ZN(n9719) );
  AOI211_X1 U10924 ( .C1(n9784), .C2(n10028), .A(n9720), .B(n9719), .ZN(n9721)
         );
  OAI21_X1 U10925 ( .B1(n9722), .B2(n9787), .A(n9721), .ZN(P1_U3273) );
  NAND2_X1 U10926 ( .A1(n9723), .A2(n10106), .ZN(n9724) );
  OAI211_X1 U10927 ( .C1(n9725), .C2(n10121), .A(n9728), .B(n9724), .ZN(n9825)
         );
  MUX2_X1 U10928 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9825), .S(n10143), .Z(
        P1_U3554) );
  NAND2_X1 U10929 ( .A1(n9726), .A2(n10106), .ZN(n9727) );
  OAI211_X1 U10930 ( .C1(n9729), .C2(n10121), .A(n9728), .B(n9727), .ZN(n9826)
         );
  MUX2_X1 U10931 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9826), .S(n10143), .Z(
        P1_U3553) );
  NAND2_X1 U10932 ( .A1(n9730), .A2(n10093), .ZN(n9737) );
  INV_X1 U10933 ( .A(n9731), .ZN(n9732) );
  NOR2_X1 U10934 ( .A1(n9732), .A2(n10119), .ZN(n9734) );
  NOR3_X1 U10935 ( .A1(n9735), .A2(n9734), .A3(n9733), .ZN(n9736) );
  NAND2_X1 U10936 ( .A1(n9737), .A2(n9736), .ZN(n9827) );
  MUX2_X1 U10937 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9827), .S(n10143), .Z(
        P1_U3552) );
  AOI21_X1 U10938 ( .B1(n10106), .B2(n9739), .A(n9738), .ZN(n9740) );
  MUX2_X1 U10939 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9828), .S(n10143), .Z(
        P1_U3550) );
  AOI22_X1 U10940 ( .A1(n9744), .A2(n10004), .B1(n10106), .B2(n9743), .ZN(
        n9745) );
  OAI211_X1 U10941 ( .C1(n9747), .C2(n10110), .A(n9746), .B(n9745), .ZN(n9829)
         );
  MUX2_X1 U10942 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9829), .S(n10143), .Z(
        P1_U3549) );
  OAI21_X1 U10943 ( .B1(n9752), .B2(n10110), .A(n9751), .ZN(n9830) );
  MUX2_X1 U10944 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9830), .S(n10143), .Z(
        P1_U3548) );
  AOI211_X1 U10945 ( .C1(n10106), .C2(n9755), .A(n9754), .B(n9753), .ZN(n9756)
         );
  AOI22_X1 U10946 ( .A1(n9759), .A2(n10004), .B1(n10106), .B2(n9758), .ZN(
        n9760) );
  OAI211_X1 U10947 ( .C1(n9762), .C2(n10110), .A(n9761), .B(n9760), .ZN(n9832)
         );
  MUX2_X1 U10948 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9832), .S(n10143), .Z(
        P1_U3546) );
  AOI22_X1 U10949 ( .A1(n9764), .A2(n10004), .B1(n10106), .B2(n9763), .ZN(
        n9765) );
  OAI211_X1 U10950 ( .C1(n9767), .C2(n10110), .A(n9766), .B(n9765), .ZN(n9833)
         );
  MUX2_X1 U10951 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9833), .S(n10143), .Z(
        P1_U3545) );
  AOI211_X1 U10952 ( .C1(n10106), .C2(n9770), .A(n9769), .B(n9768), .ZN(n9771)
         );
  OAI21_X1 U10953 ( .B1(n9772), .B2(n10110), .A(n9771), .ZN(n9834) );
  MUX2_X1 U10954 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9834), .S(n10143), .Z(
        P1_U3544) );
  AOI22_X1 U10955 ( .A1(n9774), .A2(n10004), .B1(n10106), .B2(n9773), .ZN(
        n9775) );
  OAI211_X1 U10956 ( .C1(n9777), .C2(n10110), .A(n9776), .B(n9775), .ZN(n9835)
         );
  MUX2_X1 U10957 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9835), .S(n10143), .Z(
        P1_U3543) );
  AOI22_X1 U10958 ( .A1(n9779), .A2(n10004), .B1(n10106), .B2(n9778), .ZN(
        n9780) );
  OAI211_X1 U10959 ( .C1(n9782), .C2(n10110), .A(n9781), .B(n9780), .ZN(n9836)
         );
  MUX2_X1 U10960 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9836), .S(n10143), .Z(
        P1_U3542) );
  AOI22_X1 U10961 ( .A1(n9784), .A2(n10004), .B1(n10106), .B2(n9783), .ZN(
        n9785) );
  OAI211_X1 U10962 ( .C1(n9787), .C2(n10110), .A(n9786), .B(n9785), .ZN(n9837)
         );
  MUX2_X1 U10963 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9837), .S(n10143), .Z(
        P1_U3541) );
  AOI211_X1 U10964 ( .C1(n10106), .C2(n9790), .A(n9789), .B(n9788), .ZN(n9791)
         );
  OAI21_X1 U10965 ( .B1(n9792), .B2(n10110), .A(n9791), .ZN(n9838) );
  MUX2_X1 U10966 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9838), .S(n10143), .Z(
        P1_U3540) );
  AOI211_X1 U10967 ( .C1(n10106), .C2(n9795), .A(n9794), .B(n9793), .ZN(n9796)
         );
  OAI21_X1 U10968 ( .B1(n9797), .B2(n10110), .A(n9796), .ZN(n9839) );
  MUX2_X1 U10969 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9839), .S(n10143), .Z(
        P1_U3539) );
  AOI22_X1 U10970 ( .A1(n9799), .A2(n10004), .B1(n10106), .B2(n9798), .ZN(
        n9800) );
  OAI211_X1 U10971 ( .C1(n9802), .C2(n9824), .A(n9801), .B(n9800), .ZN(n9840)
         );
  MUX2_X1 U10972 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9840), .S(n10143), .Z(
        P1_U3538) );
  AOI21_X1 U10973 ( .B1(n10106), .B2(n9804), .A(n9803), .ZN(n9805) );
  OAI211_X1 U10974 ( .C1(n9807), .C2(n10110), .A(n9806), .B(n9805), .ZN(n9841)
         );
  MUX2_X1 U10975 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9841), .S(n10143), .Z(
        P1_U3537) );
  AND2_X1 U10976 ( .A1(n9808), .A2(n10126), .ZN(n9813) );
  OAI22_X1 U10977 ( .A1(n9810), .A2(n10121), .B1(n9809), .B2(n10119), .ZN(
        n9811) );
  MUX2_X1 U10978 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9842), .S(n10143), .Z(
        P1_U3536) );
  AOI211_X1 U10979 ( .C1(n10106), .C2(n9816), .A(n9815), .B(n9814), .ZN(n9817)
         );
  OAI21_X1 U10980 ( .B1(n10110), .B2(n9818), .A(n9817), .ZN(n9843) );
  MUX2_X1 U10981 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9843), .S(n10143), .Z(
        P1_U3535) );
  AOI22_X1 U10982 ( .A1(n9820), .A2(n10004), .B1(n10106), .B2(n9819), .ZN(
        n9821) );
  OAI211_X1 U10983 ( .C1(n9824), .C2(n9823), .A(n9822), .B(n9821), .ZN(n9844)
         );
  MUX2_X1 U10984 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9844), .S(n10143), .Z(
        P1_U3534) );
  MUX2_X1 U10985 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9825), .S(n10129), .Z(
        P1_U3522) );
  MUX2_X1 U10986 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9826), .S(n10129), .Z(
        P1_U3521) );
  MUX2_X1 U10987 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9827), .S(n10129), .Z(
        P1_U3520) );
  MUX2_X1 U10988 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9828), .S(n10129), .Z(
        P1_U3518) );
  MUX2_X1 U10989 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9829), .S(n10129), .Z(
        P1_U3517) );
  MUX2_X1 U10990 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9830), .S(n10129), .Z(
        P1_U3516) );
  MUX2_X1 U10991 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9831), .S(n10129), .Z(
        P1_U3515) );
  MUX2_X1 U10992 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9832), .S(n10129), .Z(
        P1_U3514) );
  MUX2_X1 U10993 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9833), .S(n10129), .Z(
        P1_U3513) );
  MUX2_X1 U10994 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9834), .S(n10129), .Z(
        P1_U3512) );
  MUX2_X1 U10995 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9835), .S(n10129), .Z(
        P1_U3511) );
  MUX2_X1 U10996 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9836), .S(n10129), .Z(
        P1_U3510) );
  MUX2_X1 U10997 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9837), .S(n10129), .Z(
        P1_U3508) );
  MUX2_X1 U10998 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9838), .S(n10129), .Z(
        P1_U3505) );
  MUX2_X1 U10999 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9839), .S(n10129), .Z(
        P1_U3502) );
  MUX2_X1 U11000 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9840), .S(n10129), .Z(
        P1_U3499) );
  MUX2_X1 U11001 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9841), .S(n10129), .Z(
        P1_U3496) );
  MUX2_X1 U11002 ( .A(n9842), .B(P1_REG0_REG_13__SCAN_IN), .S(n10127), .Z(
        P1_U3493) );
  MUX2_X1 U11003 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9843), .S(n10129), .Z(
        P1_U3490) );
  MUX2_X1 U11004 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n9844), .S(n10129), .Z(
        P1_U3487) );
  NOR4_X1 U11005 ( .A1(n5243), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5050), .A4(
        P1_U3084), .ZN(n9845) );
  AOI21_X1 U11006 ( .B1(n9852), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9845), .ZN(
        n9846) );
  OAI21_X1 U11007 ( .B1(n9847), .B2(n7914), .A(n9846), .ZN(P1_U3322) );
  AOI21_X1 U11008 ( .B1(n9852), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n9848), .ZN(
        n9849) );
  OAI21_X1 U11009 ( .B1(n9850), .B2(n7914), .A(n9849), .ZN(P1_U3325) );
  AOI21_X1 U11010 ( .B1(n9852), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n9851), .ZN(
        n9853) );
  OAI21_X1 U11011 ( .B1(n9854), .B2(n7914), .A(n9853), .ZN(P1_U3326) );
  OAI222_X1 U11012 ( .A1(P1_U3084), .A2(n9857), .B1(n7914), .B2(n9856), .C1(
        n9855), .C2(n8332), .ZN(P1_U3327) );
  MUX2_X1 U11013 ( .A(n9858), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U11014 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9859) );
  AOI21_X1 U11015 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9859), .ZN(n10321) );
  NOR2_X1 U11016 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9860) );
  AOI21_X1 U11017 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9860), .ZN(n10324) );
  NOR2_X1 U11018 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9861) );
  AOI21_X1 U11019 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9861), .ZN(n10327) );
  NOR2_X1 U11020 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9862) );
  AOI21_X1 U11021 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9862), .ZN(n10330) );
  NOR2_X1 U11022 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9863) );
  AOI21_X1 U11023 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9863), .ZN(n10333) );
  NOR2_X1 U11024 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9871) );
  XNOR2_X1 U11025 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10361) );
  NAND2_X1 U11026 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9869) );
  XOR2_X1 U11027 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10359) );
  NAND2_X1 U11028 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9867) );
  AOI21_X1 U11029 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10315) );
  NAND2_X1 U11030 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n9864) );
  NOR2_X1 U11031 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10316), .ZN(n9865) );
  XOR2_X1 U11032 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10356) );
  NAND2_X1 U11033 ( .A1(n10357), .A2(n10356), .ZN(n9866) );
  NAND2_X1 U11034 ( .A1(n9867), .A2(n9866), .ZN(n10358) );
  NAND2_X1 U11035 ( .A1(n10359), .A2(n10358), .ZN(n9868) );
  NAND2_X1 U11036 ( .A1(n9869), .A2(n9868), .ZN(n10360) );
  NOR2_X1 U11037 ( .A1(n10361), .A2(n10360), .ZN(n9870) );
  NOR2_X1 U11038 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9872), .ZN(n10346) );
  NAND2_X1 U11039 ( .A1(n9874), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9876) );
  NAND2_X1 U11040 ( .A1(n10344), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9875) );
  NAND2_X1 U11041 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9877), .ZN(n9879) );
  NAND2_X1 U11042 ( .A1(n10343), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9878) );
  NAND2_X1 U11043 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9880), .ZN(n9882) );
  NAND2_X1 U11044 ( .A1(n10348), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9881) );
  NAND2_X1 U11045 ( .A1(n9882), .A2(n9881), .ZN(n9883) );
  INV_X1 U11046 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10355) );
  XNOR2_X1 U11047 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9883), .ZN(n10354) );
  NAND2_X1 U11048 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9885) );
  OAI21_X1 U11049 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9885), .ZN(n10341) );
  NAND2_X1 U11050 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9886) );
  OAI21_X1 U11051 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9886), .ZN(n10338) );
  NOR2_X1 U11052 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9887) );
  AOI21_X1 U11053 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9887), .ZN(n10335) );
  NAND2_X1 U11054 ( .A1(n10330), .A2(n10329), .ZN(n10328) );
  NAND2_X1 U11055 ( .A1(n10327), .A2(n10326), .ZN(n10325) );
  NAND2_X1 U11056 ( .A1(n10324), .A2(n10323), .ZN(n10322) );
  NAND2_X1 U11057 ( .A1(n10321), .A2(n10320), .ZN(n10319) );
  NOR2_X1 U11058 ( .A1(n10351), .A2(n10350), .ZN(n9888) );
  NAND2_X1 U11059 ( .A1(n10351), .A2(n10350), .ZN(n10349) );
  XOR2_X1 U11060 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n9889) );
  XNOR2_X1 U11061 ( .A(n9890), .B(n9889), .ZN(ADD_1071_U4) );
  XNOR2_X1 U11062 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11063 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  NAND2_X1 U11064 ( .A1(n9957), .A2(n9891), .ZN(n9898) );
  OAI21_X1 U11065 ( .B1(n9894), .B2(n9893), .A(n9892), .ZN(n9895) );
  INV_X1 U11066 ( .A(n9895), .ZN(n9896) );
  AOI22_X1 U11067 ( .A1(n9962), .A2(n9896), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        P1_U3084), .ZN(n9897) );
  OAI211_X1 U11068 ( .C1(n9947), .C2(n9899), .A(n9898), .B(n9897), .ZN(n9900)
         );
  INV_X1 U11069 ( .A(n9900), .ZN(n9903) );
  OAI211_X1 U11070 ( .C1(n9919), .C2(n9901), .A(n9932), .B(n9906), .ZN(n9902)
         );
  NAND2_X1 U11071 ( .A1(n9903), .A2(n9902), .ZN(P1_U3242) );
  INV_X1 U11072 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9929) );
  MUX2_X1 U11073 ( .A(n9904), .B(P1_REG2_REG_2__SCAN_IN), .S(n9910), .Z(n9907)
         );
  NAND3_X1 U11074 ( .A1(n9907), .A2(n9906), .A3(n9905), .ZN(n9908) );
  NAND3_X1 U11075 ( .A1(n9932), .A2(n9909), .A3(n9908), .ZN(n9918) );
  NAND2_X1 U11076 ( .A1(n9957), .A2(n9910), .ZN(n9917) );
  NAND2_X1 U11077 ( .A1(P1_U3084), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9916) );
  OAI211_X1 U11078 ( .C1(n9914), .C2(n9913), .A(n9962), .B(n9912), .ZN(n9915)
         );
  AND4_X1 U11079 ( .A1(n9918), .A2(n9917), .A3(n9916), .A4(n9915), .ZN(n9928)
         );
  INV_X1 U11080 ( .A(n9919), .ZN(n9922) );
  MUX2_X1 U11081 ( .A(n9922), .B(n9921), .S(n9920), .Z(n9927) );
  NAND2_X1 U11082 ( .A1(n9924), .A2(n9923), .ZN(n9925) );
  OAI211_X1 U11083 ( .C1(n9927), .C2(n9926), .A(P1_U4006), .B(n9925), .ZN(
        n9945) );
  OAI211_X1 U11084 ( .C1(n9929), .C2(n9947), .A(n9928), .B(n9945), .ZN(
        P1_U3243) );
  INV_X1 U11085 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9948) );
  NOR2_X1 U11086 ( .A1(n9931), .A2(n9930), .ZN(n9933) );
  OAI21_X1 U11087 ( .B1(n9934), .B2(n9933), .A(n9932), .ZN(n9944) );
  NAND2_X1 U11088 ( .A1(n9957), .A2(n4500), .ZN(n9943) );
  AOI21_X1 U11089 ( .B1(n9938), .B2(n9937), .A(n9936), .ZN(n9939) );
  OAI21_X1 U11090 ( .B1(n9940), .B2(n9939), .A(n9962), .ZN(n9941) );
  AND4_X1 U11091 ( .A1(n9944), .A2(n9943), .A3(n9942), .A4(n9941), .ZN(n9946)
         );
  OAI211_X1 U11092 ( .C1(n9948), .C2(n9947), .A(n9946), .B(n9945), .ZN(
        P1_U3245) );
  INV_X1 U11093 ( .A(n9949), .ZN(n9955) );
  AOI211_X1 U11094 ( .C1(n9953), .C2(n9952), .A(n9951), .B(n9950), .ZN(n9954)
         );
  AOI211_X1 U11095 ( .C1(n9957), .C2(n9956), .A(n9955), .B(n9954), .ZN(n9965)
         );
  OAI21_X1 U11096 ( .B1(n9960), .B2(n9959), .A(n9958), .ZN(n9963) );
  AOI22_X1 U11097 ( .A1(n9963), .A2(n9962), .B1(n9961), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U11098 ( .A1(n9965), .A2(n9964), .ZN(P1_U3259) );
  XOR2_X1 U11099 ( .A(n9968), .B(n9966), .Z(n10117) );
  OAI22_X1 U11100 ( .A1(n9967), .A2(n10018), .B1(n9988), .B2(n10040), .ZN(
        n9974) );
  AOI21_X1 U11101 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(n9972) );
  INV_X1 U11102 ( .A(n7735), .ZN(n9971) );
  NOR3_X1 U11103 ( .A1(n9972), .A2(n9971), .A3(n10014), .ZN(n9973) );
  AOI211_X1 U11104 ( .C1(n10034), .C2(n10117), .A(n9974), .B(n9973), .ZN(
        n10114) );
  AOI222_X1 U11105 ( .A1(n9976), .A2(n10050), .B1(P1_REG2_REG_8__SCAN_IN), 
        .B2(n10047), .C1(n10009), .C2(n9975), .ZN(n9981) );
  INV_X1 U11106 ( .A(n9977), .ZN(n9978) );
  OAI21_X1 U11107 ( .B1(n4981), .B2(n4979), .A(n9978), .ZN(n10113) );
  INV_X1 U11108 ( .A(n10113), .ZN(n9979) );
  AOI22_X1 U11109 ( .A1(n10117), .A2(n10029), .B1(n10028), .B2(n9979), .ZN(
        n9980) );
  OAI211_X1 U11110 ( .C1(n10047), .C2(n10114), .A(n9981), .B(n9980), .ZN(
        P1_U3283) );
  INV_X1 U11111 ( .A(n9983), .ZN(n9984) );
  NAND2_X1 U11112 ( .A1(n9984), .A2(n10013), .ZN(n10000) );
  NAND2_X1 U11113 ( .A1(n10000), .A2(n9985), .ZN(n9987) );
  XNOR2_X1 U11114 ( .A(n9987), .B(n9986), .ZN(n10102) );
  OAI22_X1 U11115 ( .A1(n9989), .A2(n10040), .B1(n9988), .B2(n10018), .ZN(
        n9992) );
  AOI211_X1 U11116 ( .C1(n7563), .C2(n7698), .A(n10014), .B(n9990), .ZN(n9991)
         );
  AOI211_X1 U11117 ( .C1(n10102), .C2(n10034), .A(n9992), .B(n9991), .ZN(
        n10099) );
  OAI21_X1 U11118 ( .B1(n10003), .B2(n9996), .A(n9995), .ZN(n10098) );
  INV_X1 U11119 ( .A(n10098), .ZN(n9997) );
  AOI22_X1 U11120 ( .A1(n10102), .A2(n10029), .B1(n10028), .B2(n9997), .ZN(
        n9998) );
  OAI211_X1 U11121 ( .C1(n10047), .C2(n10099), .A(n9999), .B(n9998), .ZN(
        P1_U3285) );
  INV_X1 U11122 ( .A(n10000), .ZN(n10001) );
  AOI21_X1 U11123 ( .B1(n10002), .B2(n9983), .A(n10001), .ZN(n10094) );
  INV_X1 U11124 ( .A(n10003), .ZN(n10005) );
  OAI211_X1 U11125 ( .C1(n10090), .C2(n10025), .A(n10005), .B(n10004), .ZN(
        n10089) );
  AOI22_X1 U11126 ( .A1(n10009), .A2(n10008), .B1(n10007), .B2(n10006), .ZN(
        n10010) );
  OAI21_X1 U11127 ( .B1(n10089), .B2(n10011), .A(n10010), .ZN(n10019) );
  XNOR2_X1 U11128 ( .A(n10012), .B(n10013), .ZN(n10015) );
  OAI222_X1 U11129 ( .A1(n10018), .A2(n10017), .B1(n10040), .B2(n10016), .C1(
        n10015), .C2(n10014), .ZN(n10091) );
  AOI211_X1 U11130 ( .C1(n10020), .C2(n10094), .A(n10019), .B(n10091), .ZN(
        n10021) );
  AOI22_X1 U11131 ( .A1(n10047), .A2(n10022), .B1(n10021), .B2(n10033), .ZN(
        P1_U3286) );
  XNOR2_X1 U11132 ( .A(n10023), .B(n10035), .ZN(n10085) );
  AND2_X1 U11133 ( .A1(n10024), .A2(n5365), .ZN(n10026) );
  OR2_X1 U11134 ( .A1(n10026), .A2(n10025), .ZN(n10083) );
  INV_X1 U11135 ( .A(n10083), .ZN(n10027) );
  AOI22_X1 U11136 ( .A1(n10085), .A2(n10029), .B1(n10028), .B2(n10027), .ZN(
        n10052) );
  INV_X1 U11137 ( .A(n10030), .ZN(n10032) );
  OAI22_X1 U11138 ( .A1(n10033), .A2(n5353), .B1(n10032), .B2(n10031), .ZN(
        n10049) );
  NAND2_X1 U11139 ( .A1(n10085), .A2(n10034), .ZN(n10046) );
  INV_X1 U11140 ( .A(n10035), .ZN(n10036) );
  XNOR2_X1 U11141 ( .A(n5740), .B(n10036), .ZN(n10044) );
  NAND2_X1 U11142 ( .A1(n10038), .A2(n10037), .ZN(n10039) );
  OAI21_X1 U11143 ( .B1(n10041), .B2(n10040), .A(n10039), .ZN(n10042) );
  AOI21_X1 U11144 ( .B1(n10044), .B2(n10043), .A(n10042), .ZN(n10045) );
  AND2_X1 U11145 ( .A1(n10046), .A2(n10045), .ZN(n10087) );
  NOR2_X1 U11146 ( .A1(n10087), .A2(n10047), .ZN(n10048) );
  AOI211_X1 U11147 ( .C1(n10050), .C2(n5365), .A(n10049), .B(n10048), .ZN(
        n10051) );
  NAND2_X1 U11148 ( .A1(n10052), .A2(n10051), .ZN(P1_U3287) );
  AND2_X1 U11149 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10062), .ZN(P1_U3292) );
  AND2_X1 U11150 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10062), .ZN(P1_U3293) );
  NOR2_X1 U11151 ( .A1(n10061), .A2(n10053), .ZN(P1_U3294) );
  AND2_X1 U11152 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10062), .ZN(P1_U3295) );
  AND2_X1 U11153 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10062), .ZN(P1_U3296) );
  AND2_X1 U11154 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10062), .ZN(P1_U3297) );
  AND2_X1 U11155 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10062), .ZN(P1_U3298) );
  NOR2_X1 U11156 ( .A1(n10061), .A2(n10054), .ZN(P1_U3299) );
  AND2_X1 U11157 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10062), .ZN(P1_U3300) );
  AND2_X1 U11158 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10062), .ZN(P1_U3301) );
  AND2_X1 U11159 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10062), .ZN(P1_U3302) );
  AND2_X1 U11160 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10062), .ZN(P1_U3303) );
  NOR2_X1 U11161 ( .A1(n10061), .A2(n10055), .ZN(P1_U3304) );
  AND2_X1 U11162 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10062), .ZN(P1_U3305) );
  NOR2_X1 U11163 ( .A1(n10061), .A2(n10056), .ZN(P1_U3306) );
  NOR2_X1 U11164 ( .A1(n10061), .A2(n10057), .ZN(P1_U3307) );
  AND2_X1 U11165 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10062), .ZN(P1_U3308) );
  AND2_X1 U11166 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10062), .ZN(P1_U3309) );
  NOR2_X1 U11167 ( .A1(n10061), .A2(n10058), .ZN(P1_U3310) );
  AND2_X1 U11168 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10062), .ZN(P1_U3311) );
  NOR2_X1 U11169 ( .A1(n10061), .A2(n10059), .ZN(P1_U3312) );
  AND2_X1 U11170 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10062), .ZN(P1_U3313) );
  AND2_X1 U11171 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10062), .ZN(P1_U3314) );
  AND2_X1 U11172 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10062), .ZN(P1_U3315) );
  NOR2_X1 U11173 ( .A1(n10061), .A2(n10060), .ZN(P1_U3316) );
  AND2_X1 U11174 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10062), .ZN(P1_U3317) );
  AND2_X1 U11175 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10062), .ZN(P1_U3318) );
  AND2_X1 U11176 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10062), .ZN(P1_U3319) );
  AND2_X1 U11177 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10062), .ZN(P1_U3320) );
  AND2_X1 U11178 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10062), .ZN(P1_U3321) );
  INV_X1 U11179 ( .A(n10063), .ZN(n10067) );
  OAI21_X1 U11180 ( .B1(n5819), .B2(n10119), .A(n10064), .ZN(n10066) );
  AOI211_X1 U11181 ( .C1(n10126), .C2(n10067), .A(n10066), .B(n10065), .ZN(
        n10131) );
  AOI22_X1 U11182 ( .A1(n10129), .A2(n10131), .B1(n10068), .B2(n10127), .ZN(
        P1_U3457) );
  OAI22_X1 U11183 ( .A1(n10070), .A2(n10121), .B1(n10069), .B2(n10119), .ZN(
        n10072) );
  AOI211_X1 U11184 ( .C1(n10126), .C2(n10073), .A(n10072), .B(n10071), .ZN(
        n10133) );
  INV_X1 U11185 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10074) );
  AOI22_X1 U11186 ( .A1(n10129), .A2(n10133), .B1(n10074), .B2(n10127), .ZN(
        P1_U3460) );
  INV_X1 U11187 ( .A(n10075), .ZN(n10080) );
  OAI22_X1 U11188 ( .A1(n10077), .A2(n10121), .B1(n10076), .B2(n10119), .ZN(
        n10079) );
  AOI211_X1 U11189 ( .C1(n10126), .C2(n10080), .A(n10079), .B(n10078), .ZN(
        n10134) );
  INV_X1 U11190 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10081) );
  AOI22_X1 U11191 ( .A1(n10129), .A2(n10134), .B1(n10081), .B2(n10127), .ZN(
        P1_U3463) );
  OAI22_X1 U11192 ( .A1(n10083), .A2(n10121), .B1(n10082), .B2(n10119), .ZN(
        n10084) );
  AOI21_X1 U11193 ( .B1(n10085), .B2(n10126), .A(n10084), .ZN(n10086) );
  AND2_X1 U11194 ( .A1(n10087), .A2(n10086), .ZN(n10135) );
  INV_X1 U11195 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10088) );
  AOI22_X1 U11196 ( .A1(n10129), .A2(n10135), .B1(n10088), .B2(n10127), .ZN(
        P1_U3466) );
  OAI21_X1 U11197 ( .B1(n10090), .B2(n10119), .A(n10089), .ZN(n10092) );
  AOI211_X1 U11198 ( .C1(n10094), .C2(n10093), .A(n10092), .B(n10091), .ZN(
        n10136) );
  INV_X1 U11199 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U11200 ( .A1(n10129), .A2(n10136), .B1(n10095), .B2(n10127), .ZN(
        P1_U3469) );
  INV_X1 U11201 ( .A(n10096), .ZN(n10097) );
  OAI21_X1 U11202 ( .B1(n10098), .B2(n10121), .A(n10097), .ZN(n10101) );
  INV_X1 U11203 ( .A(n10099), .ZN(n10100) );
  AOI211_X1 U11204 ( .C1(n10126), .C2(n10102), .A(n10101), .B(n10100), .ZN(
        n10137) );
  INV_X1 U11205 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10103) );
  AOI22_X1 U11206 ( .A1(n10129), .A2(n10137), .B1(n10103), .B2(n10127), .ZN(
        P1_U3472) );
  AOI21_X1 U11207 ( .B1(n10106), .B2(n10105), .A(n10104), .ZN(n10107) );
  OAI211_X1 U11208 ( .C1(n10110), .C2(n10109), .A(n10108), .B(n10107), .ZN(
        n10111) );
  INV_X1 U11209 ( .A(n10111), .ZN(n10138) );
  INV_X1 U11210 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U11211 ( .A1(n10129), .A2(n10138), .B1(n10112), .B2(n10127), .ZN(
        P1_U3475) );
  OAI22_X1 U11212 ( .A1(n10113), .A2(n10121), .B1(n4981), .B2(n10119), .ZN(
        n10116) );
  INV_X1 U11213 ( .A(n10114), .ZN(n10115) );
  AOI211_X1 U11214 ( .C1(n10126), .C2(n10117), .A(n10116), .B(n10115), .ZN(
        n10140) );
  INV_X1 U11215 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10118) );
  AOI22_X1 U11216 ( .A1(n10129), .A2(n10140), .B1(n10118), .B2(n10127), .ZN(
        P1_U3478) );
  OAI22_X1 U11217 ( .A1(n10122), .A2(n10121), .B1(n10120), .B2(n10119), .ZN(
        n10124) );
  AOI211_X1 U11218 ( .C1(n10126), .C2(n10125), .A(n10124), .B(n10123), .ZN(
        n10142) );
  AOI22_X1 U11219 ( .A1(n10129), .A2(n10142), .B1(n10128), .B2(n10127), .ZN(
        P1_U3481) );
  AOI22_X1 U11220 ( .A1(n10143), .A2(n10131), .B1(n10130), .B2(n10141), .ZN(
        P1_U3524) );
  AOI22_X1 U11221 ( .A1(n10143), .A2(n10133), .B1(n10132), .B2(n10141), .ZN(
        P1_U3525) );
  AOI22_X1 U11222 ( .A1(n10143), .A2(n10134), .B1(n7069), .B2(n10141), .ZN(
        P1_U3526) );
  AOI22_X1 U11223 ( .A1(n10143), .A2(n10135), .B1(n7070), .B2(n10141), .ZN(
        P1_U3527) );
  AOI22_X1 U11224 ( .A1(n10143), .A2(n10136), .B1(n7093), .B2(n10141), .ZN(
        P1_U3528) );
  AOI22_X1 U11225 ( .A1(n10143), .A2(n10137), .B1(n7094), .B2(n10141), .ZN(
        P1_U3529) );
  AOI22_X1 U11226 ( .A1(n10143), .A2(n10138), .B1(n7145), .B2(n10141), .ZN(
        P1_U3530) );
  INV_X1 U11227 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10139) );
  AOI22_X1 U11228 ( .A1(n10143), .A2(n10140), .B1(n10139), .B2(n10141), .ZN(
        P1_U3531) );
  AOI22_X1 U11229 ( .A1(n10143), .A2(n10142), .B1(n7226), .B2(n10141), .ZN(
        P1_U3532) );
  OR2_X1 U11230 ( .A1(n10145), .A2(n10144), .ZN(n10159) );
  INV_X1 U11231 ( .A(n10146), .ZN(n10147) );
  OR2_X1 U11232 ( .A1(n10148), .A2(n10147), .ZN(n10158) );
  AOI21_X1 U11233 ( .B1(n10151), .B2(n10150), .A(n10149), .ZN(n10157) );
  OAI211_X1 U11234 ( .C1(n10155), .C2(n10154), .A(n10153), .B(n10152), .ZN(
        n10156) );
  AND4_X1 U11235 ( .A1(n10159), .A2(n10158), .A3(n10157), .A4(n10156), .ZN(
        n10160) );
  OAI21_X1 U11236 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n10161), .A(n10160), .ZN(
        P2_U3220) );
  AOI22_X1 U11237 ( .A1(n10163), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10162), .ZN(n10172) );
  AOI22_X1 U11238 ( .A1(n10164), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10171) );
  NOR2_X1 U11239 ( .A1(n10165), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10169) );
  OAI21_X1 U11240 ( .B1(n10167), .B2(P2_REG1_REG_0__SCAN_IN), .A(n10166), .ZN(
        n10168) );
  OAI21_X1 U11241 ( .B1(n10169), .B2(n10168), .A(n10173), .ZN(n10170) );
  OAI211_X1 U11242 ( .C1(n10173), .C2(n10172), .A(n10171), .B(n10170), .ZN(
        P2_U3245) );
  AND2_X1 U11243 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10183), .ZN(P2_U3297) );
  AND2_X1 U11244 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10183), .ZN(P2_U3298) );
  AND2_X1 U11245 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10183), .ZN(P2_U3299) );
  AND2_X1 U11246 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10183), .ZN(P2_U3300) );
  AND2_X1 U11247 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10183), .ZN(P2_U3301) );
  NOR2_X1 U11248 ( .A1(n10180), .A2(n10176), .ZN(P2_U3302) );
  NOR2_X1 U11249 ( .A1(n10180), .A2(n10177), .ZN(P2_U3303) );
  AND2_X1 U11250 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10183), .ZN(P2_U3304) );
  AND2_X1 U11251 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10183), .ZN(P2_U3305) );
  NOR2_X1 U11252 ( .A1(n10180), .A2(n10178), .ZN(P2_U3306) );
  AND2_X1 U11253 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10183), .ZN(P2_U3307) );
  AND2_X1 U11254 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10183), .ZN(P2_U3308) );
  AND2_X1 U11255 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10183), .ZN(P2_U3309) );
  AND2_X1 U11256 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10183), .ZN(P2_U3310) );
  AND2_X1 U11257 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10183), .ZN(P2_U3311) );
  AND2_X1 U11258 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10183), .ZN(P2_U3312) );
  AND2_X1 U11259 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10183), .ZN(P2_U3313) );
  AND2_X1 U11260 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10183), .ZN(P2_U3314) );
  AND2_X1 U11261 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10183), .ZN(P2_U3315) );
  AND2_X1 U11262 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10183), .ZN(P2_U3316) );
  AND2_X1 U11263 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10183), .ZN(P2_U3317) );
  NOR2_X1 U11264 ( .A1(n10180), .A2(n10179), .ZN(P2_U3318) );
  AND2_X1 U11265 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10183), .ZN(P2_U3319) );
  AND2_X1 U11266 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10183), .ZN(P2_U3320) );
  AND2_X1 U11267 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10183), .ZN(P2_U3321) );
  AND2_X1 U11268 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10183), .ZN(P2_U3322) );
  AND2_X1 U11269 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10183), .ZN(P2_U3323) );
  AND2_X1 U11270 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10183), .ZN(P2_U3324) );
  AND2_X1 U11271 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10183), .ZN(P2_U3325) );
  AND2_X1 U11272 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10183), .ZN(P2_U3326) );
  AOI22_X1 U11273 ( .A1(n10186), .A2(n10182), .B1(n10181), .B2(n10183), .ZN(
        P2_U3437) );
  AOI22_X1 U11274 ( .A1(n10186), .A2(n10185), .B1(n10184), .B2(n10183), .ZN(
        P2_U3438) );
  INV_X1 U11275 ( .A(n10187), .ZN(n10191) );
  OAI22_X1 U11276 ( .A1(n10189), .A2(n10206), .B1(n6567), .B2(n10188), .ZN(
        n10190) );
  NOR2_X1 U11277 ( .A1(n10191), .A2(n10190), .ZN(n10292) );
  INV_X1 U11278 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10192) );
  AOI22_X1 U11279 ( .A1(n10290), .A2(n10292), .B1(n10192), .B2(n10288), .ZN(
        P2_U3451) );
  INV_X1 U11280 ( .A(n10193), .ZN(n10199) );
  OAI22_X1 U11281 ( .A1(n10195), .A2(n10282), .B1(n10194), .B2(n10280), .ZN(
        n10198) );
  INV_X1 U11282 ( .A(n10196), .ZN(n10197) );
  AOI211_X1 U11283 ( .C1(n10287), .C2(n10199), .A(n10198), .B(n10197), .ZN(
        n10294) );
  AOI22_X1 U11284 ( .A1(n10290), .A2(n10294), .B1(n10200), .B2(n10288), .ZN(
        P2_U3454) );
  AOI22_X1 U11285 ( .A1(n10202), .A2(n10265), .B1(n10264), .B2(n10201), .ZN(
        n10203) );
  OAI211_X1 U11286 ( .C1(n10206), .C2(n10205), .A(n10204), .B(n10203), .ZN(
        n10207) );
  INV_X1 U11287 ( .A(n10207), .ZN(n10296) );
  AOI22_X1 U11288 ( .A1(n10290), .A2(n10296), .B1(n10208), .B2(n10288), .ZN(
        P2_U3457) );
  INV_X1 U11289 ( .A(n10269), .ZN(n10261) );
  INV_X1 U11290 ( .A(n10209), .ZN(n10215) );
  NAND2_X1 U11291 ( .A1(n10210), .A2(n10265), .ZN(n10211) );
  OAI21_X1 U11292 ( .B1(n10212), .B2(n10280), .A(n10211), .ZN(n10214) );
  AOI211_X1 U11293 ( .C1(n10261), .C2(n10215), .A(n10214), .B(n10213), .ZN(
        n10297) );
  INV_X1 U11294 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10216) );
  AOI22_X1 U11295 ( .A1(n10290), .A2(n10297), .B1(n10216), .B2(n10288), .ZN(
        P2_U3460) );
  INV_X1 U11296 ( .A(n10217), .ZN(n10222) );
  OAI22_X1 U11297 ( .A1(n10219), .A2(n10282), .B1(n10218), .B2(n10280), .ZN(
        n10221) );
  AOI211_X1 U11298 ( .C1(n10287), .C2(n10222), .A(n10221), .B(n10220), .ZN(
        n10298) );
  INV_X1 U11299 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10223) );
  AOI22_X1 U11300 ( .A1(n10290), .A2(n10298), .B1(n10223), .B2(n10288), .ZN(
        P2_U3463) );
  INV_X1 U11301 ( .A(n10224), .ZN(n10225) );
  OAI21_X1 U11302 ( .B1(n10226), .B2(n10280), .A(n10225), .ZN(n10229) );
  INV_X1 U11303 ( .A(n10227), .ZN(n10228) );
  AOI211_X1 U11304 ( .C1(n10287), .C2(n10230), .A(n10229), .B(n10228), .ZN(
        n10299) );
  INV_X1 U11305 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10231) );
  AOI22_X1 U11306 ( .A1(n10290), .A2(n10299), .B1(n10231), .B2(n10288), .ZN(
        P2_U3466) );
  INV_X1 U11307 ( .A(n10232), .ZN(n10237) );
  OAI22_X1 U11308 ( .A1(n10234), .A2(n10282), .B1(n10233), .B2(n10280), .ZN(
        n10236) );
  AOI211_X1 U11309 ( .C1(n10237), .C2(n10287), .A(n10236), .B(n10235), .ZN(
        n10301) );
  INV_X1 U11310 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10238) );
  AOI22_X1 U11311 ( .A1(n10290), .A2(n10301), .B1(n10238), .B2(n10288), .ZN(
        P2_U3469) );
  OAI22_X1 U11312 ( .A1(n10240), .A2(n10282), .B1(n10239), .B2(n10280), .ZN(
        n10243) );
  INV_X1 U11313 ( .A(n10241), .ZN(n10242) );
  AOI211_X1 U11314 ( .C1(n10287), .C2(n10244), .A(n10243), .B(n10242), .ZN(
        n10302) );
  INV_X1 U11315 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10245) );
  AOI22_X1 U11316 ( .A1(n10290), .A2(n10302), .B1(n10245), .B2(n10288), .ZN(
        P2_U3472) );
  INV_X1 U11317 ( .A(n10250), .ZN(n10252) );
  AOI22_X1 U11318 ( .A1(n10247), .A2(n10265), .B1(n10264), .B2(n4840), .ZN(
        n10248) );
  OAI211_X1 U11319 ( .C1(n10250), .C2(n10269), .A(n10249), .B(n10248), .ZN(
        n10251) );
  AOI21_X1 U11320 ( .B1(n10253), .B2(n10252), .A(n10251), .ZN(n10304) );
  INV_X1 U11321 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U11322 ( .A1(n10290), .A2(n10304), .B1(n10254), .B2(n10288), .ZN(
        P2_U3475) );
  INV_X1 U11323 ( .A(n10255), .ZN(n10257) );
  OAI22_X1 U11324 ( .A1(n10257), .A2(n10282), .B1(n10256), .B2(n10280), .ZN(
        n10259) );
  AOI211_X1 U11325 ( .C1(n10261), .C2(n10260), .A(n10259), .B(n10258), .ZN(
        n10306) );
  INV_X1 U11326 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10262) );
  AOI22_X1 U11327 ( .A1(n10290), .A2(n10306), .B1(n10262), .B2(n10288), .ZN(
        P2_U3478) );
  AOI22_X1 U11328 ( .A1(n10266), .A2(n10265), .B1(n10264), .B2(n10263), .ZN(
        n10267) );
  OAI211_X1 U11329 ( .C1(n10270), .C2(n10269), .A(n10268), .B(n10267), .ZN(
        n10271) );
  INV_X1 U11330 ( .A(n10271), .ZN(n10308) );
  AOI22_X1 U11331 ( .A1(n10290), .A2(n10308), .B1(n10272), .B2(n10288), .ZN(
        P2_U3481) );
  INV_X1 U11332 ( .A(n10273), .ZN(n10278) );
  OAI22_X1 U11333 ( .A1(n10275), .A2(n10282), .B1(n10274), .B2(n10280), .ZN(
        n10277) );
  AOI211_X1 U11334 ( .C1(n10278), .C2(n10287), .A(n10277), .B(n10276), .ZN(
        n10310) );
  INV_X1 U11335 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10279) );
  AOI22_X1 U11336 ( .A1(n10290), .A2(n10310), .B1(n10279), .B2(n10288), .ZN(
        P2_U3484) );
  OAI22_X1 U11337 ( .A1(n10283), .A2(n10282), .B1(n10281), .B2(n10280), .ZN(
        n10285) );
  AOI211_X1 U11338 ( .C1(n10287), .C2(n10286), .A(n10285), .B(n10284), .ZN(
        n10313) );
  INV_X1 U11339 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U11340 ( .A1(n10290), .A2(n10313), .B1(n10289), .B2(n10288), .ZN(
        P2_U3487) );
  INV_X1 U11341 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10291) );
  AOI22_X1 U11342 ( .A1(n10314), .A2(n10292), .B1(n10291), .B2(n10311), .ZN(
        P2_U3520) );
  AOI22_X1 U11343 ( .A1(n10314), .A2(n10294), .B1(n10293), .B2(n10311), .ZN(
        P2_U3521) );
  AOI22_X1 U11344 ( .A1(n10314), .A2(n10296), .B1(n10295), .B2(n10311), .ZN(
        P2_U3522) );
  AOI22_X1 U11345 ( .A1(n10314), .A2(n10297), .B1(n7306), .B2(n10311), .ZN(
        P2_U3523) );
  AOI22_X1 U11346 ( .A1(n10314), .A2(n10298), .B1(n7308), .B2(n10311), .ZN(
        P2_U3524) );
  AOI22_X1 U11347 ( .A1(n10314), .A2(n10299), .B1(n7310), .B2(n10311), .ZN(
        P2_U3525) );
  AOI22_X1 U11348 ( .A1(n10314), .A2(n10301), .B1(n10300), .B2(n10311), .ZN(
        P2_U3526) );
  AOI22_X1 U11349 ( .A1(n10314), .A2(n10302), .B1(n7359), .B2(n10311), .ZN(
        P2_U3527) );
  INV_X1 U11350 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U11351 ( .A1(n10314), .A2(n10304), .B1(n10303), .B2(n10311), .ZN(
        P2_U3528) );
  AOI22_X1 U11352 ( .A1(n10314), .A2(n10306), .B1(n10305), .B2(n10311), .ZN(
        P2_U3529) );
  AOI22_X1 U11353 ( .A1(n10314), .A2(n10308), .B1(n10307), .B2(n10311), .ZN(
        P2_U3530) );
  AOI22_X1 U11354 ( .A1(n10314), .A2(n10310), .B1(n10309), .B2(n10311), .ZN(
        P2_U3531) );
  AOI22_X1 U11355 ( .A1(n10314), .A2(n10313), .B1(n10312), .B2(n10311), .ZN(
        P2_U3532) );
  NOR2_X1 U11356 ( .A1(n10316), .A2(n10315), .ZN(n10318) );
  XNOR2_X1 U11357 ( .A(n10318), .B(n10317), .ZN(ADD_1071_U5) );
  XOR2_X1 U11358 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11359 ( .B1(n10321), .B2(n10320), .A(n10319), .ZN(ADD_1071_U56) );
  OAI21_X1 U11360 ( .B1(n10324), .B2(n10323), .A(n10322), .ZN(ADD_1071_U57) );
  OAI21_X1 U11361 ( .B1(n10327), .B2(n10326), .A(n10325), .ZN(ADD_1071_U58) );
  OAI21_X1 U11362 ( .B1(n10330), .B2(n10329), .A(n10328), .ZN(ADD_1071_U59) );
  OAI21_X1 U11363 ( .B1(n10333), .B2(n10332), .A(n10331), .ZN(ADD_1071_U60) );
  OAI21_X1 U11364 ( .B1(n10336), .B2(n10335), .A(n10334), .ZN(ADD_1071_U61) );
  AOI21_X1 U11365 ( .B1(n10339), .B2(n10338), .A(n10337), .ZN(ADD_1071_U62) );
  AOI21_X1 U11366 ( .B1(n10342), .B2(n10341), .A(n10340), .ZN(ADD_1071_U63) );
  XOR2_X1 U11367 ( .A(n10343), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11368 ( .A(n10344), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11369 ( .A1(n10346), .A2(n10345), .ZN(n10347) );
  XOR2_X1 U11370 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10347), .Z(ADD_1071_U51) );
  XOR2_X1 U11371 ( .A(n10348), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  OAI21_X1 U11372 ( .B1(n10351), .B2(n10350), .A(n10349), .ZN(n10352) );
  XNOR2_X1 U11373 ( .A(n10352), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11374 ( .B1(n10355), .B2(n10354), .A(n10353), .ZN(ADD_1071_U47) );
  XOR2_X1 U11375 ( .A(n10357), .B(n10356), .Z(ADD_1071_U54) );
  XOR2_X1 U11376 ( .A(n10358), .B(n10359), .Z(ADD_1071_U53) );
  XNOR2_X1 U11377 ( .A(n10361), .B(n10360), .ZN(ADD_1071_U52) );
  INV_X1 U4891 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6283) );
  BUF_X1 U4938 ( .A(n6570), .Z(n4377) );
  CLKBUF_X2 U4882 ( .A(n6736), .Z(n4380) );
  NAND2_X1 U6210 ( .A1(n5350), .A2(n4481), .ZN(n7647) );
  XNOR2_X1 U6306 ( .A(n5886), .B(n5885), .ZN(n8223) );
endmodule

