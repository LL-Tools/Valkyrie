

module b14_C_gen_AntiSAT_k_256_3 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084;

  AND2_X1 U2468 ( .A1(n3448), .A2(n3447), .ZN(n3445) );
  NAND2_X1 U2469 ( .A1(n3237), .A2(n3220), .ZN(n3232) );
  INV_X1 U2470 ( .A(n2501), .ZN(n3863) );
  CLKBUF_X1 U2471 ( .A(n2422), .Z(n2547) );
  AND2_X1 U2472 ( .A1(n2399), .A2(n2400), .ZN(n2422) );
  XNOR2_X1 U2473 ( .A(n2396), .B(IR_REG_29__SCAN_IN), .ZN(n2976) );
  OR2_X1 U2474 ( .A1(n2395), .A2(n2765), .ZN(n2396) );
  OAI21_X1 U2475 ( .B1(n2804), .B2(n3885), .A(n2748), .ZN(n2749) );
  CLKBUF_X2 U2476 ( .A(n2843), .Z(n3727) );
  OR2_X1 U2477 ( .A1(n4208), .A2(n3898), .ZN(n4189) );
  OR2_X1 U2478 ( .A1(n3270), .A2(n3973), .ZN(n2723) );
  NAND2_X1 U2479 ( .A1(n2720), .A2(n3975), .ZN(n3172) );
  INV_X1 U2480 ( .A(n3257), .ZN(n3122) );
  MUX2_X1 U2482 ( .A(REG1_REG_28__SCAN_IN), .B(n2815), .S(n4710), .Z(n2810) );
  MUX2_X1 U2483 ( .A(REG0_REG_28__SCAN_IN), .B(n2815), .S(n4703), .Z(n2816) );
  XNOR2_X1 U2484 ( .A(n2394), .B(IR_REG_30__SCAN_IN), .ZN(n4495) );
  AOI21_X2 U2485 ( .B1(n3758), .B2(n3759), .A(n2367), .ZN(n3765) );
  NAND2_X2 U2486 ( .A1(n2327), .A2(n2242), .ZN(n3758) );
  NAND4_X4 U2487 ( .A1(n2409), .A2(n2408), .A3(n2407), .A4(n2406), .ZN(n2419)
         );
  AND2_X1 U2488 ( .A1(n4164), .A2(n2807), .ZN(n2808) );
  OAI21_X1 U2489 ( .B1(n3795), .B2(n3797), .A(n3796), .ZN(n3775) );
  AND2_X1 U2490 ( .A1(n4513), .A2(n4516), .ZN(n3647) );
  OR2_X1 U2491 ( .A1(n3850), .A2(n4514), .ZN(n3648) );
  AOI21_X1 U2492 ( .B1(n3591), .B2(n2241), .A(n2353), .ZN(n3640) );
  NAND2_X1 U2493 ( .A1(n3109), .A2(n2926), .ZN(n3184) );
  OAI21_X1 U2494 ( .B1(n4260), .B2(n2699), .A(n2644), .ZN(n4402) );
  NAND2_X2 U2495 ( .A1(n4703), .A2(n4357), .ZN(n4492) );
  AND2_X2 U2496 ( .A1(n2894), .A2(n4368), .ZN(n4509) );
  INV_X1 U2497 ( .A(n2433), .ZN(n2432) );
  INV_X2 U2498 ( .A(n2844), .ZN(n2843) );
  INV_X2 U2499 ( .A(n3711), .ZN(n3725) );
  NAND4_X1 U2500 ( .A1(n2427), .A2(n2426), .A3(n2425), .A4(n2424), .ZN(n2433)
         );
  AND2_X2 U2501 ( .A1(n2833), .A2(n2832), .ZN(n3708) );
  NAND2_X2 U2502 ( .A1(n2778), .A2(n2777), .ZN(n2833) );
  AND2_X2 U2503 ( .A1(n2829), .A2(n2832), .ZN(n3711) );
  INV_X1 U2504 ( .A(n2832), .ZN(n3166) );
  NAND2_X1 U2505 ( .A1(n3948), .A2(n4016), .ZN(n2832) );
  INV_X1 U2506 ( .A(n2781), .ZN(n3948) );
  NAND2_X1 U2507 ( .A1(n3738), .A2(IR_REG_31__SCAN_IN), .ZN(n2394) );
  INV_X1 U2508 ( .A(n4496), .ZN(n2796) );
  OR2_X1 U2509 ( .A1(n2768), .A2(n2767), .ZN(n2973) );
  NOR2_X1 U2510 ( .A1(n2703), .A2(IR_REG_21__SCAN_IN), .ZN(n2770) );
  NAND2_X1 U2511 ( .A1(n2700), .A2(IR_REG_31__SCAN_IN), .ZN(n2706) );
  NOR2_X1 U2512 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2263)
         );
  NAND2_X2 U2513 ( .A1(n2556), .A2(n4893), .ZN(n2565) );
  XNOR2_X2 U2514 ( .A(n2773), .B(IR_REG_24__SCAN_IN), .ZN(n2778) );
  NOR2_X2 U2515 ( .A1(n3555), .A2(n3609), .ZN(n3556) );
  NOR3_X2 U2516 ( .A1(n3815), .A2(n3750), .A3(n3749), .ZN(n3748) );
  NOR2_X2 U2517 ( .A1(n3816), .A2(n3817), .ZN(n3815) );
  NOR2_X2 U2518 ( .A1(n3571), .A2(n2259), .ZN(n4356) );
  OR2_X2 U2519 ( .A1(n3474), .A2(n3641), .ZN(n3571) );
  AOI21_X2 U2520 ( .B1(n3714), .B2(n2419), .A(n2848), .ZN(n2858) );
  AOI21_X1 U2521 ( .B1(n3714), .B2(n2838), .A(n2837), .ZN(n2840) );
  AOI21_X1 U2522 ( .B1(n3714), .B2(n2825), .A(n2831), .ZN(n2910) );
  INV_X4 U2523 ( .A(n3724), .ZN(n3714) );
  NOR2_X2 U2524 ( .A1(n4216), .A2(n4197), .ZN(n4196) );
  OR2_X2 U2525 ( .A1(n4229), .A2(n4214), .ZN(n4216) );
  AND2_X4 U2526 ( .A1(n2833), .A2(n3166), .ZN(n2844) );
  NOR2_X4 U2527 ( .A1(n4312), .A2(n4419), .ZN(n4289) );
  NAND2_X1 U2528 ( .A1(n2299), .A2(n2606), .ZN(n2298) );
  INV_X1 U2529 ( .A(n4307), .ZN(n2299) );
  NOR2_X1 U2530 ( .A1(n3931), .A2(n2277), .ZN(n2276) );
  INV_X1 U2531 ( .A(n3786), .ZN(n2332) );
  OR2_X1 U2532 ( .A1(n3797), .A2(n2345), .ZN(n2344) );
  INV_X1 U2533 ( .A(n2421), .ZN(n2695) );
  INV_X1 U2534 ( .A(n2491), .ZN(n2699) );
  XNOR2_X1 U2535 ( .A(n2311), .B(n3004), .ZN(n4063) );
  NAND2_X1 U2536 ( .A1(n4544), .A2(n4545), .ZN(n4543) );
  XNOR2_X1 U2537 ( .A(n4100), .B(n4099), .ZN(n4556) );
  NAND2_X1 U2538 ( .A1(n4565), .A2(n4566), .ZN(n4564) );
  XNOR2_X1 U2539 ( .A(n4078), .B(n4671), .ZN(n4577) );
  AOI21_X1 U2540 ( .B1(n2250), .B2(n4585), .A(n2230), .ZN(n2314) );
  OR2_X1 U2541 ( .A1(n2683), .A2(n2682), .ZN(n4150) );
  INV_X1 U2542 ( .A(n2284), .ZN(n2283) );
  OAI21_X1 U2543 ( .B1(n2286), .B2(n2285), .A(n3943), .ZN(n2284) );
  AOI21_X1 U2544 ( .B1(n4206), .B2(n2664), .A(n2663), .ZN(n4187) );
  NAND2_X1 U2545 ( .A1(n4568), .A2(n4569), .ZN(n4567) );
  NAND2_X1 U2546 ( .A1(n4579), .A2(REG2_REG_12__SCAN_IN), .ZN(n4578) );
  OAI21_X1 U2547 ( .B1(n2356), .B2(n2355), .A(n2354), .ZN(n2353) );
  INV_X1 U2548 ( .A(n3631), .ZN(n2354) );
  INV_X1 U2549 ( .A(n4087), .ZN(n2325) );
  AND2_X1 U2550 ( .A1(n4195), .A2(n4384), .ZN(n3887) );
  OR2_X1 U2551 ( .A1(n4291), .A2(n4279), .ZN(n4250) );
  NOR2_X1 U2552 ( .A1(n2623), .A2(n2622), .ZN(n2624) );
  OR2_X1 U2553 ( .A1(n4353), .A2(n2298), .ZN(n2297) );
  INV_X1 U2554 ( .A(n4308), .ZN(n2622) );
  INV_X1 U2555 ( .A(n4337), .ZN(n2605) );
  OR2_X1 U2556 ( .A1(n4244), .A2(n4243), .ZN(n4328) );
  AND2_X1 U2557 ( .A1(n3641), .A2(n4033), .ZN(n2592) );
  INV_X1 U2558 ( .A(n2577), .ZN(n2266) );
  OAI21_X1 U2559 ( .B1(n2276), .B2(n2274), .A(n2244), .ZN(n2273) );
  INV_X1 U2560 ( .A(n2546), .ZN(n2274) );
  INV_X1 U2561 ( .A(n2488), .ZN(n2291) );
  INV_X1 U2562 ( .A(n2976), .ZN(n2400) );
  NOR2_X1 U2563 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2388)
         );
  NAND2_X1 U2564 ( .A1(n2385), .A2(n2362), .ZN(n2361) );
  INV_X1 U2565 ( .A(n2363), .ZN(n2362) );
  INV_X1 U2566 ( .A(IR_REG_25__SCAN_IN), .ZN(n2390) );
  NAND2_X1 U2567 ( .A1(n3325), .A2(n3324), .ZN(n2350) );
  XNOR2_X1 U2568 ( .A(n2836), .B(n3725), .ZN(n2839) );
  NAND2_X1 U2569 ( .A1(n2838), .A2(n2844), .ZN(n2835) );
  OR2_X1 U2570 ( .A1(n3724), .A2(n2849), .ZN(n2850) );
  NAND2_X1 U2571 ( .A1(n2617), .A2(n2616), .ZN(n2625) );
  AND2_X1 U2572 ( .A1(n3426), .A2(n3425), .ZN(n3529) );
  XNOR2_X1 U2573 ( .A(n2847), .B(n3725), .ZN(n2860) );
  AOI21_X1 U2574 ( .B1(n3646), .B2(n2332), .A(n2246), .ZN(n2331) );
  OR2_X1 U2575 ( .A1(n2331), .A2(n2330), .ZN(n2329) );
  INV_X1 U2576 ( .A(n3829), .ZN(n2330) );
  NAND3_X1 U2577 ( .A1(n3648), .A2(n3647), .A3(n2240), .ZN(n2327) );
  NOR2_X1 U2578 ( .A1(n2471), .A2(n3017), .ZN(n2479) );
  NAND2_X1 U2579 ( .A1(n3776), .A2(n2343), .ZN(n2338) );
  INV_X1 U2580 ( .A(n3700), .ZN(n2335) );
  AND2_X1 U2581 ( .A1(n2342), .A2(n2346), .ZN(n2341) );
  INV_X1 U2582 ( .A(n3777), .ZN(n2346) );
  INV_X1 U2583 ( .A(n4506), .ZN(n3853) );
  NOR2_X1 U2584 ( .A1(n3640), .A2(n3639), .ZN(n3850) );
  OAI21_X1 U2585 ( .B1(n2695), .B2(n2349), .A(n2435), .ZN(n2348) );
  OAI21_X1 U2586 ( .B1(n2990), .B2(n2991), .A(n2306), .ZN(n4050) );
  NAND2_X1 U2587 ( .A1(n2990), .A2(n2991), .ZN(n2306) );
  AOI21_X1 U2588 ( .B1(n4063), .B2(REG2_REG_3__SCAN_IN), .A(n2235), .ZN(n2994)
         );
  OAI22_X1 U2589 ( .A1(n4072), .A2(n4093), .B1(n4071), .B2(n4070), .ZN(n4073)
         );
  OR2_X1 U2590 ( .A1(n4095), .A2(n4094), .ZN(n4096) );
  NOR2_X1 U2591 ( .A1(n4093), .A2(n4092), .ZN(n4094) );
  NAND2_X1 U2592 ( .A1(n4543), .A2(n4075), .ZN(n4076) );
  NAND2_X1 U2593 ( .A1(n4546), .A2(n4098), .ZN(n4100) );
  NAND2_X1 U2594 ( .A1(n4556), .A2(REG2_REG_10__SCAN_IN), .ZN(n4555) );
  NAND2_X1 U2595 ( .A1(n4564), .A2(n2247), .ZN(n4078) );
  NAND2_X1 U2596 ( .A1(n4670), .A2(n2551), .ZN(n2317) );
  NOR2_X1 U2597 ( .A1(n4599), .A2(n2560), .ZN(n4598) );
  NOR2_X1 U2598 ( .A1(n4606), .A2(n2249), .ZN(n4110) );
  NAND2_X1 U2599 ( .A1(n4626), .A2(n2309), .ZN(n4115) );
  NAND2_X1 U2600 ( .A1(n4665), .A2(n2401), .ZN(n2309) );
  NOR2_X1 U2601 ( .A1(n4115), .A2(n4114), .ZN(n4129) );
  OR2_X1 U2602 ( .A1(n2665), .A2(n3842), .ZN(n2683) );
  AOI22_X1 U2603 ( .A1(n4227), .A2(n2654), .B1(n4236), .B2(n4253), .ZN(n4206)
         );
  AOI21_X1 U2604 ( .B1(n4287), .B2(n2631), .A(n2630), .ZN(n4267) );
  AND2_X1 U2605 ( .A1(n3819), .A2(n4298), .ZN(n2630) );
  AND2_X1 U2606 ( .A1(n2594), .A2(REG3_REG_18__SCAN_IN), .ZN(n2617) );
  AOI21_X1 U2607 ( .B1(n3649), .B2(n4511), .A(n2593), .ZN(n4354) );
  NOR2_X1 U2608 ( .A1(n2591), .A2(n2578), .ZN(n2268) );
  NAND2_X1 U2609 ( .A1(n3438), .A2(n2577), .ZN(n2269) );
  NOR2_X1 U2610 ( .A1(n2523), .A2(n3447), .ZN(n2277) );
  NAND2_X1 U2611 ( .A1(n2279), .A2(n2226), .ZN(n2278) );
  INV_X1 U2612 ( .A(n3449), .ZN(n2279) );
  NAND2_X1 U2613 ( .A1(n2278), .A2(n2276), .ZN(n3390) );
  AND2_X1 U2614 ( .A1(n3375), .A2(n3981), .ZN(n3931) );
  AND2_X1 U2615 ( .A1(n2399), .A2(n2976), .ZN(n2421) );
  AND2_X1 U2616 ( .A1(n3227), .A2(n2420), .ZN(n3129) );
  AND2_X1 U2617 ( .A1(n2714), .A2(n3230), .ZN(n3228) );
  AND2_X1 U2618 ( .A1(n2828), .A2(n2781), .ZN(n3221) );
  AND2_X1 U2619 ( .A1(n2873), .A2(n2981), .ZN(n3162) );
  NAND2_X1 U2620 ( .A1(n2833), .A2(n4664), .ZN(n3159) );
  AND2_X1 U2621 ( .A1(n2690), .A2(n2689), .ZN(n4388) );
  NAND2_X1 U2622 ( .A1(n3554), .A2(n4682), .ZN(n4443) );
  AND2_X1 U2623 ( .A1(n3221), .A2(n4498), .ZN(n4430) );
  AND2_X2 U2624 ( .A1(n3221), .A2(n4016), .ZN(n4357) );
  INV_X1 U2625 ( .A(IR_REG_28__SCAN_IN), .ZN(n2754) );
  NAND2_X1 U2626 ( .A1(n2612), .A2(n2611), .ZN(n2700) );
  INV_X1 U2627 ( .A(IR_REG_4__SCAN_IN), .ZN(n2452) );
  NAND2_X1 U2628 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2305)
         );
  NAND2_X1 U2629 ( .A1(n3591), .A2(n2357), .ZN(n2352) );
  INV_X1 U2630 ( .A(n3844), .ZN(n4512) );
  XNOR2_X1 U2631 ( .A(n2990), .B(REG1_REG_1__SCAN_IN), .ZN(n4048) );
  XNOR2_X1 U2632 ( .A(n2994), .B(n2310), .ZN(n3096) );
  NOR2_X1 U2633 ( .A1(n3001), .A2(n3000), .ZN(n4095) );
  NAND2_X1 U2634 ( .A1(n4547), .A2(n4548), .ZN(n4546) );
  NAND2_X1 U2635 ( .A1(n4104), .A2(n4578), .ZN(n4588) );
  XNOR2_X1 U2636 ( .A(n4110), .B(n4085), .ZN(n4617) );
  NAND2_X1 U2637 ( .A1(n4617), .A2(n3476), .ZN(n4616) );
  INV_X1 U2638 ( .A(n3941), .ZN(n2288) );
  NAND2_X1 U2639 ( .A1(n2281), .A2(n2280), .ZN(n2289) );
  AOI21_X1 U2640 ( .B1(n2283), .B2(n2285), .A(n2243), .ZN(n2280) );
  NAND2_X1 U2641 ( .A1(n2282), .A2(n2374), .ZN(n2803) );
  INV_X1 U2642 ( .A(n3902), .ZN(n2623) );
  NAND2_X1 U2643 ( .A1(n2368), .A2(n2364), .ZN(n2363) );
  INV_X1 U2644 ( .A(IR_REG_6__SCAN_IN), .ZN(n2485) );
  INV_X1 U2645 ( .A(IR_REG_10__SCAN_IN), .ZN(n2531) );
  INV_X1 U2646 ( .A(n3590), .ZN(n2358) );
  AND2_X1 U2647 ( .A1(n4388), .A2(n2691), .ZN(n3888) );
  NAND2_X1 U2648 ( .A1(n3073), .A2(n2993), .ZN(n2311) );
  NAND2_X1 U2649 ( .A1(n4504), .A2(REG2_REG_2__SCAN_IN), .ZN(n2993) );
  OR2_X1 U2650 ( .A1(n4585), .A2(n4081), .ZN(n2315) );
  INV_X1 U2651 ( .A(n2317), .ZN(n2316) );
  AND2_X1 U2652 ( .A1(n3936), .A2(n4188), .ZN(n4009) );
  OR2_X1 U2653 ( .A1(n3376), .A2(n3983), .ZN(n2728) );
  NAND2_X1 U2654 ( .A1(n3252), .A2(n2454), .ZN(n3956) );
  NOR2_X1 U2655 ( .A1(n3392), .A2(n3490), .ZN(n2261) );
  NAND2_X1 U2656 ( .A1(n3192), .A2(n3215), .ZN(n3193) );
  AND2_X1 U2657 ( .A1(n3948), .A2(n4497), .ZN(n2988) );
  NOR2_X1 U2658 ( .A1(n2227), .A2(IR_REG_18__SCAN_IN), .ZN(n2351) );
  OR3_X1 U2659 ( .A1(n2510), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2521) );
  INV_X1 U2660 ( .A(IR_REG_19__SCAN_IN), .ZN(n2705) );
  OR2_X1 U2661 ( .A1(n3589), .A2(n2358), .ZN(n2357) );
  NAND2_X1 U2662 ( .A1(n3589), .A2(n2358), .ZN(n2356) );
  NOR2_X1 U2663 ( .A1(n2503), .A2(n2502), .ZN(n2514) );
  AND2_X1 U2664 ( .A1(n2647), .A2(REG3_REG_24__SCAN_IN), .ZN(n2655) );
  NAND2_X1 U2665 ( .A1(n2336), .A2(n2343), .ZN(n3796) );
  INV_X1 U2666 ( .A(n2339), .ZN(n2336) );
  AND2_X1 U2667 ( .A1(n2948), .A2(n2949), .ZN(n3276) );
  OR2_X1 U2668 ( .A1(n2535), .A2(n4865), .ZN(n2549) );
  OR2_X1 U2669 ( .A1(n2549), .A2(n2548), .ZN(n2558) );
  NAND2_X1 U2670 ( .A1(n2524), .A2(REG3_REG_11__SCAN_IN), .ZN(n2535) );
  INV_X1 U2671 ( .A(n2431), .ZN(n3131) );
  NAND2_X1 U2672 ( .A1(n2457), .A2(REG3_REG_5__SCAN_IN), .ZN(n2471) );
  NOR2_X1 U2673 ( .A1(n2558), .A2(n4743), .ZN(n2570) );
  NOR3_X1 U2674 ( .A1(n4050), .A2(n3060), .A3(n2262), .ZN(n4051) );
  NAND2_X1 U2675 ( .A1(n2322), .A2(n2321), .ZN(n2320) );
  NAND2_X1 U2676 ( .A1(n4502), .A2(REG1_REG_5__SCAN_IN), .ZN(n2321) );
  INV_X1 U2677 ( .A(n3024), .ZN(n2322) );
  NAND2_X1 U2678 ( .A1(n3020), .A2(n2319), .ZN(n4069) );
  NAND2_X1 U2679 ( .A1(n2320), .A2(n4501), .ZN(n2319) );
  NAND2_X1 U2680 ( .A1(n4539), .A2(n4074), .ZN(n4544) );
  NAND2_X1 U2681 ( .A1(n4560), .A2(n4077), .ZN(n4565) );
  NAND2_X1 U2682 ( .A1(n4567), .A2(n4102), .ZN(n4103) );
  NAND2_X1 U2683 ( .A1(n4592), .A2(n4080), .ZN(n4082) );
  NAND2_X1 U2684 ( .A1(n4632), .A2(n2251), .ZN(n2323) );
  NAND2_X1 U2685 ( .A1(n2325), .A2(n2251), .ZN(n2324) );
  NAND2_X1 U2686 ( .A1(n2811), .A2(n3886), .ZN(n4378) );
  INV_X1 U2687 ( .A(n2374), .ZN(n2285) );
  NOR2_X1 U2688 ( .A1(n2681), .A2(n2287), .ZN(n2286) );
  INV_X1 U2689 ( .A(n2370), .ZN(n2287) );
  INV_X1 U2690 ( .A(n4173), .ZN(n4170) );
  NAND2_X1 U2691 ( .A1(n4385), .A2(n4197), .ZN(n2672) );
  AND2_X1 U2692 ( .A1(n2679), .A2(n2678), .ZN(n4195) );
  AND2_X1 U2693 ( .A1(n4402), .A2(n2253), .ZN(n2645) );
  AOI21_X1 U2694 ( .B1(n2231), .B2(n2298), .A(n2295), .ZN(n2294) );
  INV_X1 U2695 ( .A(n3903), .ZN(n2295) );
  OR2_X1 U2696 ( .A1(n4328), .A2(n4245), .ZN(n4304) );
  NAND2_X1 U2697 ( .A1(n4352), .A2(n2606), .ZN(n4326) );
  NAND2_X1 U2698 ( .A1(n4354), .A2(n4353), .ZN(n4352) );
  NAND2_X1 U2699 ( .A1(n2732), .A2(n3990), .ZN(n4244) );
  INV_X1 U2700 ( .A(n3863), .ZN(n2986) );
  AOI21_X1 U2701 ( .B1(n2268), .B2(n2266), .A(n2592), .ZN(n2265) );
  INV_X1 U2702 ( .A(n2268), .ZN(n2267) );
  OR2_X1 U2703 ( .A1(n2580), .A2(n5057), .ZN(n2582) );
  NAND2_X1 U2704 ( .A1(n3549), .A2(n3919), .ZN(n3550) );
  INV_X1 U2705 ( .A(n2271), .ZN(n3543) );
  OAI21_X1 U2706 ( .B1(n3449), .B2(n2234), .A(n2272), .ZN(n2271) );
  INV_X1 U2707 ( .A(n2273), .ZN(n2272) );
  INV_X1 U2708 ( .A(n2293), .ZN(n2292) );
  AOI21_X1 U2709 ( .B1(n2293), .B2(n2291), .A(n2232), .ZN(n2290) );
  AOI21_X1 U2710 ( .B1(n3927), .B2(n2488), .A(n2233), .ZN(n2293) );
  INV_X1 U2711 ( .A(REG3_REG_8__SCAN_IN), .ZN(n5056) );
  AND2_X1 U2712 ( .A1(n3961), .A2(n3967), .ZN(n3927) );
  NAND2_X1 U2713 ( .A1(n3150), .A2(n2456), .ZN(n3078) );
  AND2_X1 U2714 ( .A1(n3956), .A2(n3958), .ZN(n3926) );
  NAND2_X1 U2715 ( .A1(n2386), .A2(IR_REG_27__SCAN_IN), .ZN(n2301) );
  NAND2_X1 U2716 ( .A1(n2751), .A2(n2388), .ZN(n2300) );
  NOR2_X1 U2717 ( .A1(n4378), .A2(n4381), .ZN(n4377) );
  NAND2_X1 U2718 ( .A1(n4378), .A2(n2258), .ZN(n4151) );
  OR2_X1 U2719 ( .A1(n2811), .A2(n3886), .ZN(n2258) );
  AND2_X1 U2720 ( .A1(n4175), .A2(n4163), .ZN(n2811) );
  INV_X1 U2721 ( .A(n3704), .ZN(n4214) );
  OR2_X1 U2722 ( .A1(n4259), .A2(n4401), .ZN(n4229) );
  NAND2_X1 U2723 ( .A1(n4289), .A2(n2252), .ZN(n4259) );
  NOR2_X1 U2724 ( .A1(n2254), .A2(n2253), .ZN(n2252) );
  INV_X1 U2725 ( .A(n4279), .ZN(n2254) );
  AND2_X1 U2726 ( .A1(n4289), .A2(n4279), .ZN(n4269) );
  NAND2_X1 U2727 ( .A1(n3790), .A2(n4359), .ZN(n2259) );
  NAND2_X1 U2728 ( .A1(n4356), .A2(n4342), .ZN(n4341) );
  NOR2_X1 U2729 ( .A1(n3571), .A2(n3649), .ZN(n4360) );
  INV_X1 U2730 ( .A(n4508), .ZN(n3641) );
  NAND2_X1 U2731 ( .A1(n3556), .A2(n3856), .ZN(n3474) );
  NAND2_X1 U2732 ( .A1(n2261), .A2(n3510), .ZN(n3555) );
  NAND2_X1 U2733 ( .A1(n3445), .A2(n3430), .ZN(n3392) );
  INV_X1 U2734 ( .A(n2261), .ZN(n3394) );
  MUX2_X1 U2735 ( .A(DATAI_12_), .B(n4575), .S(n2986), .Z(n3490) );
  INV_X1 U2736 ( .A(n4424), .ZN(n4432) );
  NOR2_X1 U2737 ( .A1(n3302), .A2(n3292), .ZN(n3448) );
  OR2_X1 U2738 ( .A1(n3193), .A2(n3308), .ZN(n3302) );
  NOR2_X1 U2739 ( .A1(n3145), .A2(n2255), .ZN(n3192) );
  NAND2_X1 U2740 ( .A1(n3188), .A2(n2256), .ZN(n2255) );
  INV_X1 U2741 ( .A(n3355), .ZN(n3188) );
  OR2_X1 U2742 ( .A1(n3144), .A2(n2454), .ZN(n3145) );
  NOR2_X1 U2743 ( .A1(n3145), .A2(n3246), .ZN(n3176) );
  INV_X1 U2744 ( .A(n4430), .ZN(n4334) );
  INV_X1 U2745 ( .A(n4443), .ZN(n4690) );
  NOR2_X1 U2746 ( .A1(n3232), .A2(n2431), .ZN(n3139) );
  INV_X1 U2747 ( .A(n2875), .ZN(n3163) );
  NAND2_X1 U2748 ( .A1(n2360), .A2(n2392), .ZN(n2359) );
  INV_X1 U2749 ( .A(n2361), .ZN(n2360) );
  XNOR2_X1 U2750 ( .A(n2711), .B(n2769), .ZN(n2828) );
  NAND2_X1 U2751 ( .A1(n2710), .A2(IR_REG_31__SCAN_IN), .ZN(n2711) );
  INV_X1 U2752 ( .A(IR_REG_7__SCAN_IN), .ZN(n2497) );
  NAND2_X1 U2753 ( .A1(n2350), .A2(n2959), .ZN(n2962) );
  INV_X1 U2754 ( .A(n3668), .ZN(n4342) );
  AND2_X1 U2755 ( .A1(n4150), .A2(n2684), .ZN(n4160) );
  AOI21_X1 U2756 ( .B1(n3648), .B2(n3647), .A(n3646), .ZN(n3785) );
  OAI21_X1 U2757 ( .B1(n3280), .B2(n3276), .A(n3277), .ZN(n3325) );
  INV_X1 U2758 ( .A(n3220), .ZN(n3230) );
  AND2_X1 U2759 ( .A1(n3497), .A2(n3526), .ZN(n3498) );
  OR2_X1 U2760 ( .A1(n2897), .A2(n2890), .ZN(n3844) );
  INV_X1 U2761 ( .A(n3054), .ZN(n2866) );
  OR2_X1 U2762 ( .A1(n2897), .A2(n2896), .ZN(n4506) );
  NAND2_X1 U2763 ( .A1(n2328), .A2(n2331), .ZN(n3827) );
  AND2_X1 U2764 ( .A1(n2327), .A2(n2329), .ZN(n3826) );
  NAND2_X1 U2765 ( .A1(n2341), .A2(n2337), .ZN(n2333) );
  NAND2_X1 U2766 ( .A1(n2341), .A2(n2335), .ZN(n2334) );
  AND2_X1 U2767 ( .A1(n2344), .A2(n2338), .ZN(n2337) );
  OR2_X1 U2768 ( .A1(n2897), .A2(n2879), .ZN(n3861) );
  INV_X1 U2769 ( .A(n4522), .ZN(n3859) );
  NAND2_X1 U2770 ( .A1(n2662), .A2(n2661), .ZN(n4231) );
  NAND2_X1 U2771 ( .A1(n2636), .A2(n2635), .ZN(n4291) );
  OAI211_X1 U2772 ( .C1(n4293), .C2(n2699), .A(n2629), .B(n2628), .ZN(n4433)
         );
  OR2_X1 U2773 ( .A1(n2824), .A2(n2833), .ZN(n4031) );
  OAI211_X1 U2774 ( .C1(n2759), .C2(n2621), .A(n2620), .B(n2619), .ZN(n4421)
         );
  OAI211_X1 U2775 ( .C1(n2759), .C2(n4346), .A(n2610), .B(n2609), .ZN(n4032)
         );
  NAND4_X1 U2776 ( .A1(n2600), .A2(n2599), .A3(n2598), .A4(n2597), .ZN(n4337)
         );
  NAND4_X1 U2777 ( .A1(n2496), .A2(n2495), .A3(n2494), .A4(n2493), .ZN(n4041)
         );
  NAND3_X1 U2778 ( .A1(n2347), .A2(n2437), .A3(n2436), .ZN(n2838) );
  NAND2_X1 U2779 ( .A1(n2421), .A2(REG1_REG_1__SCAN_IN), .ZN(n2409) );
  NAND2_X1 U2780 ( .A1(n2422), .A2(REG0_REG_1__SCAN_IN), .ZN(n2408) );
  AND2_X1 U2781 ( .A1(n2415), .A2(n2414), .ZN(n2418) );
  AND2_X1 U2782 ( .A1(n2999), .A2(n2998), .ZN(n4529) );
  NAND2_X1 U2783 ( .A1(n4048), .A2(n4047), .ZN(n4046) );
  INV_X1 U2784 ( .A(IR_REG_2__SCAN_IN), .ZN(n2429) );
  NOR2_X1 U2785 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2428)
         );
  AOI22_X1 U2786 ( .A1(n3096), .A2(REG2_REG_4__SCAN_IN), .B1(n2310), .B2(n2995), .ZN(n3029) );
  NAND2_X1 U2787 ( .A1(n2248), .A2(REG1_REG_6__SCAN_IN), .ZN(n3020) );
  NAND2_X1 U2788 ( .A1(n4534), .A2(n4097), .ZN(n4547) );
  XNOR2_X1 U2789 ( .A(n4076), .B(n4099), .ZN(n4561) );
  NAND2_X1 U2790 ( .A1(n4555), .A2(n4101), .ZN(n4568) );
  XNOR2_X1 U2791 ( .A(n4103), .B(n4671), .ZN(n4579) );
  NAND2_X1 U2792 ( .A1(n4576), .A2(n4079), .ZN(n4593) );
  NAND2_X1 U2793 ( .A1(n4593), .A2(n4594), .ZN(n4592) );
  XNOR2_X1 U2794 ( .A(n4082), .B(n4669), .ZN(n4603) );
  NOR2_X1 U2795 ( .A1(n4598), .A2(n4107), .ZN(n4608) );
  NAND2_X1 U2796 ( .A1(n2318), .A2(n2317), .ZN(n4106) );
  OR2_X1 U2797 ( .A1(n4588), .A2(n4585), .ZN(n2318) );
  NAND2_X1 U2798 ( .A1(n4616), .A2(n4111), .ZN(n4625) );
  NOR2_X1 U2799 ( .A1(n4633), .A2(n4632), .ZN(n4634) );
  XNOR2_X1 U2800 ( .A(n4125), .B(n2326), .ZN(n4088) );
  INV_X1 U2801 ( .A(n4124), .ZN(n2326) );
  AND2_X1 U2802 ( .A1(n4529), .A2(n3009), .ZN(n4631) );
  XNOR2_X1 U2803 ( .A(n2307), .B(n4130), .ZN(n4135) );
  NOR2_X1 U2804 ( .A1(n4129), .A2(n2308), .ZN(n2307) );
  NOR2_X1 U2805 ( .A1(n4123), .A2(n4370), .ZN(n2308) );
  AND2_X1 U2806 ( .A1(n4529), .A2(n4023), .ZN(n4586) );
  INV_X1 U2807 ( .A(n2691), .ZN(n4163) );
  AND2_X1 U2808 ( .A1(n2269), .A2(n2268), .ZN(n3473) );
  INV_X1 U2809 ( .A(n3634), .ZN(n3856) );
  NAND2_X1 U2810 ( .A1(n2278), .A2(n2275), .ZN(n3334) );
  INV_X1 U2811 ( .A(n2277), .ZN(n2275) );
  NAND4_X1 U2812 ( .A1(n2476), .A2(n2475), .A3(n2474), .A4(n2473), .ZN(n4043)
         );
  INV_X1 U2813 ( .A(n4343), .ZN(n4655) );
  INV_X1 U2814 ( .A(n4368), .ZN(n4652) );
  OR2_X1 U2815 ( .A1(n4151), .A2(n4446), .ZN(n2821) );
  NAND2_X1 U2816 ( .A1(n2762), .A2(n2372), .ZN(n2819) );
  NAND2_X1 U2817 ( .A1(n2980), .A2(n3037), .ZN(n4662) );
  XNOR2_X1 U2818 ( .A(n2775), .B(IR_REG_26__SCAN_IN), .ZN(n4496) );
  NAND2_X1 U2819 ( .A1(n2772), .A2(IR_REG_31__SCAN_IN), .ZN(n2773) );
  AND2_X1 U2820 ( .A1(n2987), .A2(STATE_REG_SCAN_IN), .ZN(n4664) );
  INV_X1 U2821 ( .A(IR_REG_3__SCAN_IN), .ZN(n2449) );
  XNOR2_X1 U2822 ( .A(n2450), .B(IR_REG_3__SCAN_IN), .ZN(n4503) );
  NAND2_X1 U2823 ( .A1(n2303), .A2(n2302), .ZN(n2990) );
  NAND2_X1 U2824 ( .A1(n2305), .A2(n2304), .ZN(n2303) );
  INV_X1 U2825 ( .A(IR_REG_1__SCAN_IN), .ZN(n2304) );
  OR2_X1 U2826 ( .A1(n4157), .A2(n4446), .ZN(n2813) );
  OR2_X1 U2827 ( .A1(n4157), .A2(n4492), .ZN(n2817) );
  INV_X1 U2828 ( .A(IR_REG_31__SCAN_IN), .ZN(n2765) );
  OR2_X1 U2829 ( .A1(n4039), .A2(n3451), .ZN(n2226) );
  XNOR2_X1 U2830 ( .A(n2430), .B(n2429), .ZN(n3066) );
  OR2_X1 U2831 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2227)
         );
  AND2_X1 U2832 ( .A1(n2960), .A2(n2959), .ZN(n2228) );
  AND2_X1 U2833 ( .A1(n2455), .A2(n2440), .ZN(n2229) );
  INV_X1 U2834 ( .A(n3479), .ZN(n2591) );
  AND2_X1 U2835 ( .A1(n2316), .A2(n4669), .ZN(n2230) );
  OR2_X2 U2836 ( .A1(n3687), .A2(n4357), .ZN(n3724) );
  INV_X1 U2837 ( .A(n3103), .ZN(n2310) );
  NAND2_X1 U2838 ( .A1(n4495), .A2(n2400), .ZN(n2423) );
  INV_X1 U2839 ( .A(n3246), .ZN(n2256) );
  NAND2_X1 U2840 ( .A1(n2448), .A2(n2447), .ZN(n2825) );
  AOI21_X1 U2841 ( .B1(n4241), .B2(n2646), .A(n2645), .ZN(n4227) );
  AND2_X1 U2842 ( .A1(n2624), .A2(n2297), .ZN(n2231) );
  NOR2_X1 U2843 ( .A1(n2565), .A2(n2361), .ZN(n2763) );
  NAND2_X1 U2844 ( .A1(n2264), .A2(n2262), .ZN(n2438) );
  AND2_X1 U2845 ( .A1(n4041), .A2(n3308), .ZN(n2232) );
  NOR2_X1 U2846 ( .A1(n4041), .A2(n3308), .ZN(n2233) );
  NAND2_X1 U2847 ( .A1(n2546), .A2(n2226), .ZN(n2234) );
  AND2_X1 U2848 ( .A1(n2311), .A2(n4503), .ZN(n2235) );
  XNOR2_X1 U2849 ( .A(n2289), .B(n2288), .ZN(n4145) );
  INV_X1 U2850 ( .A(n2340), .ZN(n3795) );
  INV_X1 U2851 ( .A(IR_REG_18__SCAN_IN), .ZN(n2611) );
  OR2_X1 U2852 ( .A1(n2833), .A2(n2852), .ZN(n2236) );
  NAND2_X1 U2853 ( .A1(n3420), .A2(n3419), .ZN(n3500) );
  OR2_X1 U2854 ( .A1(n2565), .A2(IR_REG_14__SCAN_IN), .ZN(n2237) );
  NOR2_X1 U2855 ( .A1(n4035), .A2(n3609), .ZN(n2238) );
  NAND2_X1 U2856 ( .A1(n2296), .A2(n2294), .ZN(n4287) );
  INV_X1 U2857 ( .A(n2270), .ZN(n3570) );
  NAND2_X1 U2858 ( .A1(n2771), .A2(IR_REG_31__SCAN_IN), .ZN(n2779) );
  NAND2_X1 U2859 ( .A1(n2352), .A2(n2356), .ZN(n3633) );
  AND2_X1 U2860 ( .A1(n2269), .A2(n2579), .ZN(n2239) );
  OAI21_X1 U2861 ( .B1(n3268), .B2(n2513), .A(n2512), .ZN(n3449) );
  INV_X1 U2862 ( .A(n3790), .ZN(n3649) );
  AND2_X1 U2863 ( .A1(n3829), .A2(n2332), .ZN(n2240) );
  NOR2_X1 U2864 ( .A1(n4341), .A2(n4431), .ZN(n2260) );
  AND2_X1 U2865 ( .A1(n2357), .A2(n3632), .ZN(n2241) );
  AND2_X1 U2866 ( .A1(n2329), .A2(n3828), .ZN(n2242) );
  INV_X1 U2867 ( .A(n2578), .ZN(n2579) );
  AND2_X1 U2868 ( .A1(n4030), .A2(n2691), .ZN(n2243) );
  NAND2_X1 U2869 ( .A1(n4037), .A2(n3490), .ZN(n2244) );
  AND2_X1 U2870 ( .A1(n3698), .A2(n3697), .ZN(n2245) );
  INV_X1 U2871 ( .A(n3776), .ZN(n2345) );
  INV_X1 U2872 ( .A(n4710), .ZN(n4711) );
  OR2_X1 U2873 ( .A1(n3201), .A2(n3927), .ZN(n3204) );
  INV_X1 U2874 ( .A(n4257), .ZN(n2253) );
  NAND2_X1 U2875 ( .A1(n3204), .A2(n2488), .ZN(n3305) );
  INV_X1 U2876 ( .A(n3632), .ZN(n2355) );
  AND2_X1 U2877 ( .A1(n3655), .A2(n3654), .ZN(n2246) );
  NAND2_X1 U2878 ( .A1(n2441), .A2(n2440), .ZN(n3151) );
  OR2_X1 U2879 ( .A1(n4672), .A2(n4712), .ZN(n2247) );
  AND2_X1 U2880 ( .A1(n2602), .A2(n2601), .ZN(n2612) );
  AND2_X2 U2881 ( .A1(n2809), .A2(n3163), .ZN(n4703) );
  XNOR2_X1 U2882 ( .A(n2909), .B(n2910), .ZN(n2914) );
  XOR2_X1 U2883 ( .A(n2320), .B(n4501), .Z(n2248) );
  AND2_X1 U2884 ( .A1(n4109), .A2(REG2_REG_15__SCAN_IN), .ZN(n2249) );
  INV_X1 U2885 ( .A(n4085), .ZN(n4666) );
  AND2_X1 U2886 ( .A1(n4081), .A2(n2317), .ZN(n2250) );
  INV_X1 U2887 ( .A(DATAI_0_), .ZN(n2257) );
  INV_X1 U2888 ( .A(IR_REG_14__SCAN_IN), .ZN(n2364) );
  INV_X1 U2889 ( .A(n4112), .ZN(n4665) );
  OR2_X1 U2890 ( .A1(n4112), .A2(REG1_REG_17__SCAN_IN), .ZN(n2251) );
  NOR2_X2 U2891 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2376)
         );
  MUX2_X1 U2892 ( .A(n2257), .B(n2262), .S(n2501), .Z(n3220) );
  NAND2_X2 U2893 ( .A1(n2301), .A2(n2300), .ZN(n2501) );
  AND2_X2 U2894 ( .A1(n4196), .A2(n4182), .ZN(n4175) );
  INV_X1 U2895 ( .A(n2260), .ZN(n4312) );
  NAND3_X1 U2896 ( .A1(n2264), .A2(n2263), .A3(n2262), .ZN(n2466) );
  INV_X2 U2897 ( .A(IR_REG_0__SCAN_IN), .ZN(n2262) );
  NOR2_X2 U2898 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2264)
         );
  OAI21_X1 U2899 ( .B1(n3438), .B2(n2267), .A(n2265), .ZN(n2270) );
  NAND2_X1 U2900 ( .A1(n2673), .A2(n2283), .ZN(n2281) );
  NAND2_X1 U2901 ( .A1(n2673), .A2(n2286), .ZN(n2282) );
  NAND2_X1 U2902 ( .A1(n2673), .A2(n2370), .ZN(n4174) );
  OAI21_X1 U2903 ( .B1(n3201), .B2(n2292), .A(n2290), .ZN(n3268) );
  NAND2_X1 U2904 ( .A1(n4354), .A2(n2231), .ZN(n2296) );
  OR2_X2 U2905 ( .A1(n2766), .A2(IR_REG_26__SCAN_IN), .ZN(n2752) );
  NAND2_X1 U2906 ( .A1(n2763), .A2(n2390), .ZN(n2766) );
  NAND2_X1 U2907 ( .A1(n2441), .A2(n2229), .ZN(n3150) );
  MUX2_X1 U2908 ( .A(DATAI_2_), .B(n4504), .S(n2501), .Z(n2431) );
  NAND3_X1 U2909 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .A3(
        IR_REG_1__SCAN_IN), .ZN(n2302) );
  NAND3_X1 U2910 ( .A1(n2313), .A2(n2314), .A3(n2312), .ZN(n4599) );
  NAND2_X1 U2911 ( .A1(n4588), .A2(n2250), .ZN(n2312) );
  OR2_X1 U2912 ( .A1(n4588), .A2(n2315), .ZN(n2313) );
  OAI21_X1 U2913 ( .B1(n4621), .B2(n2324), .A(n2323), .ZN(n4125) );
  NOR2_X1 U2914 ( .A1(n4621), .A2(n4087), .ZN(n4633) );
  NAND3_X1 U2915 ( .A1(n3648), .A2(n3647), .A3(n2332), .ZN(n2328) );
  OAI21_X1 U2916 ( .B1(n3748), .B2(n2334), .A(n2333), .ZN(n3841) );
  NOR2_X1 U2917 ( .A1(n3748), .A2(n3700), .ZN(n2339) );
  NAND2_X1 U2918 ( .A1(n2339), .A2(n2245), .ZN(n2340) );
  OR2_X1 U2919 ( .A1(n2344), .A2(n2245), .ZN(n2342) );
  INV_X1 U2920 ( .A(n2245), .ZN(n2343) );
  AOI21_X2 U2921 ( .B1(n3841), .B2(n3838), .A(n3837), .ZN(n3742) );
  INV_X1 U2922 ( .A(n2348), .ZN(n2347) );
  INV_X1 U2923 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2349) );
  NAND2_X1 U2924 ( .A1(n2350), .A2(n2228), .ZN(n3420) );
  NAND2_X1 U2925 ( .A1(n2612), .A2(n2351), .ZN(n2703) );
  NOR2_X1 U2926 ( .A1(n2565), .A2(n2363), .ZN(n2602) );
  NOR2_X2 U2927 ( .A1(n2359), .A2(n2565), .ZN(n2395) );
  NAND2_X1 U2928 ( .A1(n2833), .A2(n2832), .ZN(n3687) );
  OR2_X1 U2929 ( .A1(n2423), .A2(n2991), .ZN(n2407) );
  OR2_X1 U2930 ( .A1(n2428), .A2(n2765), .ZN(n2430) );
  NAND2_X1 U2931 ( .A1(n3640), .A2(n3639), .ZN(n4513) );
  OAI21_X2 U2932 ( .B1(n3500), .B2(n3499), .A(n3498), .ZN(n3591) );
  OR2_X1 U2933 ( .A1(STATE_REG_SCAN_IN), .A2(n4116), .ZN(n2365) );
  NAND2_X1 U2934 ( .A1(n3040), .A2(n3041), .ZN(n3039) );
  AND2_X1 U2935 ( .A1(n2491), .A2(n3158), .ZN(n2366) );
  AND2_X1 U2936 ( .A1(n3671), .A2(n3670), .ZN(n2367) );
  AND2_X1 U2937 ( .A1(n4874), .A2(n4987), .ZN(n2368) );
  NOR2_X1 U2938 ( .A1(n2880), .A2(n2914), .ZN(n2369) );
  OR2_X1 U2939 ( .A1(n4385), .A2(n4197), .ZN(n2370) );
  INV_X1 U2940 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2502) );
  INV_X1 U2941 ( .A(n3149), .ZN(n2454) );
  OR2_X1 U2942 ( .A1(n4425), .A2(n4279), .ZN(n2371) );
  AND2_X1 U2943 ( .A1(n4149), .A2(n2761), .ZN(n2372) );
  AND2_X1 U2944 ( .A1(n3682), .A2(n3806), .ZN(n2373) );
  INV_X1 U2945 ( .A(n3843), .ZN(n4197) );
  INV_X1 U2946 ( .A(n4554), .ZN(n4099) );
  OR2_X1 U2947 ( .A1(n4195), .A2(n4182), .ZN(n2374) );
  INV_X1 U2948 ( .A(n4385), .ZN(n4213) );
  NAND2_X1 U2949 ( .A1(n2671), .A2(n2670), .ZN(n4385) );
  INV_X1 U2950 ( .A(n2963), .ZN(n2960) );
  AND2_X1 U2951 ( .A1(n3900), .A2(n4222), .ZN(n4001) );
  INV_X1 U2952 ( .A(IR_REG_13__SCAN_IN), .ZN(n4893) );
  NOR2_X1 U2953 ( .A1(n2828), .A2(n4499), .ZN(n2885) );
  AND4_X1 U2954 ( .A1(n2384), .A2(n2383), .A3(n2382), .A4(n2381), .ZN(n2385)
         );
  NOR2_X1 U2955 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2378)
         );
  NAND2_X1 U2956 ( .A1(n3089), .A2(n2870), .ZN(n2906) );
  OR4_X1 U2957 ( .A1(n3884), .A2(n3888), .A3(n3887), .A4(n3889), .ZN(n3895) );
  INV_X1 U2958 ( .A(n4495), .ZN(n2399) );
  AND2_X1 U2959 ( .A1(n2391), .A2(n2390), .ZN(n2392) );
  INV_X1 U2960 ( .A(n3767), .ZN(n3683) );
  NAND2_X1 U2961 ( .A1(n2655), .A2(REG3_REG_25__SCAN_IN), .ZN(n2665) );
  NOR2_X1 U2962 ( .A1(n2973), .A2(n2796), .ZN(n2777) );
  AND2_X1 U2963 ( .A1(n4231), .A2(n4214), .ZN(n2663) );
  AND2_X1 U2964 ( .A1(n4303), .A2(n2736), .ZN(n4247) );
  NAND2_X1 U2965 ( .A1(n2605), .A2(n4359), .ZN(n2606) );
  INV_X1 U2966 ( .A(n4298), .ZN(n4419) );
  AND2_X1 U2967 ( .A1(n2514), .A2(REG3_REG_10__SCAN_IN), .ZN(n2524) );
  OR2_X1 U2968 ( .A1(n2856), .A2(n3725), .ZN(n2857) );
  INV_X1 U2969 ( .A(n4291), .ZN(n4425) );
  NAND2_X1 U2970 ( .A1(n2842), .A2(n2870), .ZN(n2915) );
  NAND2_X1 U2971 ( .A1(n3684), .A2(n3683), .ZN(n3685) );
  NOR2_X1 U2972 ( .A1(n2582), .A2(n2397), .ZN(n2594) );
  AND2_X1 U2973 ( .A1(n2665), .A2(n2656), .ZN(n4217) );
  INV_X1 U2974 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3017) );
  INV_X1 U2975 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4865) );
  OR2_X1 U2976 ( .A1(n4007), .A2(n3887), .ZN(n4173) );
  OR2_X1 U2977 ( .A1(n2489), .A2(n5056), .ZN(n2503) );
  AND2_X1 U2978 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2457) );
  NAND2_X1 U2979 ( .A1(n3129), .A2(n3128), .ZN(n3127) );
  OR2_X1 U2980 ( .A1(n3159), .A2(n2893), .ZN(n4368) );
  OR2_X1 U2981 ( .A1(n2980), .A2(D_REG_0__SCAN_IN), .ZN(n2798) );
  INV_X1 U2982 ( .A(n4236), .ZN(n4401) );
  NOR2_X1 U2983 ( .A1(n2986), .A2(n5062), .ZN(n4431) );
  INV_X1 U2984 ( .A(n3603), .ZN(n3609) );
  INV_X1 U2985 ( .A(n4366), .ZN(n4339) );
  OR2_X1 U2986 ( .A1(n2980), .A2(n2793), .ZN(n2873) );
  NOR2_X1 U2987 ( .A1(n2639), .A2(n2638), .ZN(n2647) );
  OR2_X1 U2988 ( .A1(n2625), .A2(n5031), .ZN(n2639) );
  INV_X1 U2989 ( .A(n3861), .ZN(n4517) );
  OR2_X1 U2990 ( .A1(n4200), .A2(n2699), .ZN(n2671) );
  OR2_X1 U2991 ( .A1(n2759), .A2(n2516), .ZN(n2517) );
  NAND2_X1 U2992 ( .A1(n4117), .A2(n2365), .ZN(n4118) );
  AOI21_X1 U2993 ( .B1(n4115), .B2(n4114), .A(n4624), .ZN(n4119) );
  INV_X1 U2994 ( .A(n4374), .ZN(n4311) );
  NAND2_X1 U2995 ( .A1(n2750), .A2(n4020), .ZN(n4366) );
  AND2_X1 U2996 ( .A1(n2798), .A2(n2983), .ZN(n2875) );
  INV_X1 U2997 ( .A(n3451), .ZN(n3447) );
  AND2_X1 U2998 ( .A1(n3223), .A2(n2828), .ZN(n4700) );
  AND3_X1 U2999 ( .A1(n2795), .A2(n2794), .A3(n2873), .ZN(n2809) );
  NAND2_X1 U3000 ( .A1(n2776), .A2(n4496), .ZN(n2980) );
  AND2_X1 U3001 ( .A1(n2999), .A2(n2989), .ZN(n4630) );
  AND2_X1 U3002 ( .A1(n2888), .A2(n2887), .ZN(n4522) );
  INV_X1 U3003 ( .A(n4388), .ZN(n4030) );
  OAI21_X1 U3004 ( .B1(n4232), .B2(n2699), .A(n2653), .ZN(n4210) );
  NAND4_X1 U3005 ( .A1(n2587), .A2(n2586), .A3(n2585), .A4(n2584), .ZN(n4033)
         );
  NAND4_X1 U3006 ( .A1(n2520), .A2(n2519), .A3(n2518), .A4(n2517), .ZN(n4039)
         );
  INV_X1 U3007 ( .A(n4586), .ZN(n4624) );
  AOI21_X1 U3008 ( .B1(n4120), .B2(n4119), .A(n4118), .ZN(n4121) );
  NAND2_X1 U3009 ( .A1(n4349), .A2(n3203), .ZN(n4374) );
  AND2_X1 U3010 ( .A1(n2821), .A2(n2820), .ZN(n2822) );
  AND2_X1 U3011 ( .A1(n2800), .A2(n2799), .ZN(n2801) );
  INV_X1 U3012 ( .A(n4703), .ZN(n4701) );
  INV_X1 U3013 ( .A(n4662), .ZN(n4663) );
  XNOR2_X1 U3014 ( .A(n2706), .B(IR_REG_19__SCAN_IN), .ZN(n4499) );
  INV_X1 U3015 ( .A(n4090), .ZN(n4672) );
  INV_X1 U3016 ( .A(DATAI_17_), .ZN(n2387) );
  NOR2_X2 U3017 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2377)
         );
  NOR2_X2 U3018 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2375)
         );
  NAND4_X1 U3019 ( .A1(n2378), .A2(n2377), .A3(n2376), .A4(n2375), .ZN(n2379)
         );
  NOR2_X2 U3020 ( .A1(n2466), .A2(n2379), .ZN(n2556) );
  OR2_X1 U3022 ( .A1(n2602), .A2(n2765), .ZN(n2380) );
  XNOR2_X1 U3023 ( .A(n2380), .B(IR_REG_17__SCAN_IN), .ZN(n4112) );
  NOR2_X1 U3024 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2384)
         );
  NOR2_X1 U3025 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2383)
         );
  NOR2_X1 U3026 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2382)
         );
  NOR2_X1 U3027 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2381)
         );
  NAND2_X2 U3028 ( .A1(n2752), .A2(IR_REG_31__SCAN_IN), .ZN(n2751) );
  NOR2_X1 U3029 ( .A1(n2751), .A2(n2754), .ZN(n2386) );
  MUX2_X1 U3030 ( .A(n2387), .B(n4665), .S(n2986), .Z(n3790) );
  INV_X1 U3031 ( .A(n2388), .ZN(n2389) );
  NOR2_X1 U3032 ( .A1(IR_REG_26__SCAN_IN), .A2(n2389), .ZN(n2391) );
  INV_X1 U3033 ( .A(IR_REG_29__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U3034 ( .A1(n2395), .A2(n2393), .ZN(n3738) );
  AND2_X4 U3035 ( .A1(n4495), .A2(n2976), .ZN(n2491) );
  NAND2_X1 U3036 ( .A1(n2479), .A2(REG3_REG_7__SCAN_IN), .ZN(n2489) );
  INV_X1 U3037 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2548) );
  INV_X1 U3038 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4743) );
  NAND2_X1 U3039 ( .A1(n2570), .A2(REG3_REG_15__SCAN_IN), .ZN(n2580) );
  INV_X1 U3040 ( .A(REG3_REG_16__SCAN_IN), .ZN(n5057) );
  INV_X1 U3041 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2397) );
  AND2_X1 U3042 ( .A1(n2582), .A2(n2397), .ZN(n2398) );
  NOR2_X1 U3043 ( .A1(n2594), .A2(n2398), .ZN(n3792) );
  NAND2_X1 U3044 ( .A1(n2491), .A2(n3792), .ZN(n2405) );
  INV_X2 U3045 ( .A(n2695), .ZN(n3864) );
  NAND2_X1 U3046 ( .A1(n3864), .A2(REG1_REG_17__SCAN_IN), .ZN(n2404) );
  NAND2_X1 U3047 ( .A1(n2547), .A2(REG0_REG_17__SCAN_IN), .ZN(n2403) );
  INV_X1 U3048 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2401) );
  OR2_X1 U3049 ( .A1(n2759), .A2(n2401), .ZN(n2402) );
  NAND4_X1 U3050 ( .A1(n2405), .A2(n2404), .A3(n2403), .A4(n2402), .ZN(n4511)
         );
  INV_X1 U3051 ( .A(n4511), .ZN(n3832) );
  INV_X1 U3052 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2991) );
  NAND2_X1 U3053 ( .A1(n2491), .A2(REG3_REG_1__SCAN_IN), .ZN(n2406) );
  INV_X1 U3054 ( .A(n2419), .ZN(n2413) );
  INV_X1 U3055 ( .A(DATAI_1_), .ZN(n2410) );
  NAND2_X1 U3056 ( .A1(n2501), .A2(n2990), .ZN(n2411) );
  OAI21_X2 U3057 ( .B1(n2501), .B2(DATAI_1_), .A(n2411), .ZN(n3237) );
  NAND2_X1 U3059 ( .A1(n2413), .A2(n3231), .ZN(n2715) );
  NAND2_X1 U3060 ( .A1(n2419), .A2(n3237), .ZN(n3946) );
  NAND2_X1 U3061 ( .A1(n2715), .A2(n3946), .ZN(n2713) );
  NAND2_X1 U3062 ( .A1(n2421), .A2(REG1_REG_0__SCAN_IN), .ZN(n2415) );
  NAND2_X1 U3063 ( .A1(n2491), .A2(REG3_REG_0__SCAN_IN), .ZN(n2414) );
  NAND2_X1 U3064 ( .A1(n2422), .A2(REG0_REG_0__SCAN_IN), .ZN(n2417) );
  INV_X1 U3065 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3060) );
  OR2_X1 U3066 ( .A1(n2423), .A2(n3060), .ZN(n2416) );
  NAND3_X1 U3067 ( .A1(n2418), .A2(n2417), .A3(n2416), .ZN(n2714) );
  NAND2_X1 U3068 ( .A1(n2713), .A2(n3228), .ZN(n3227) );
  INV_X1 U3069 ( .A(n3237), .ZN(n3231) );
  NAND2_X1 U3070 ( .A1(n2419), .A2(n3231), .ZN(n2420) );
  NAND2_X1 U3071 ( .A1(n2421), .A2(REG1_REG_2__SCAN_IN), .ZN(n2427) );
  NAND2_X1 U3072 ( .A1(n2422), .A2(REG0_REG_2__SCAN_IN), .ZN(n2426) );
  NAND2_X1 U3073 ( .A1(n2491), .A2(REG3_REG_2__SCAN_IN), .ZN(n2425) );
  INV_X1 U3074 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2992) );
  OR2_X1 U3075 ( .A1(n2423), .A2(n2992), .ZN(n2424) );
  NAND2_X1 U3076 ( .A1(n2432), .A2(n2431), .ZN(n3950) );
  NAND2_X1 U3077 ( .A1(n2433), .A2(n3131), .ZN(n3953) );
  NAND2_X1 U3078 ( .A1(n3950), .A2(n3953), .ZN(n3128) );
  OR2_X1 U3079 ( .A1(n2433), .A2(n2431), .ZN(n2434) );
  NAND2_X1 U3080 ( .A1(n3127), .A2(n2434), .ZN(n3117) );
  INV_X1 U3081 ( .A(REG2_REG_3__SCAN_IN), .ZN(n4062) );
  OR2_X1 U3082 ( .A1(n2423), .A2(n4062), .ZN(n2437) );
  NAND2_X1 U3083 ( .A1(n2422), .A2(REG0_REG_3__SCAN_IN), .ZN(n2436) );
  INV_X1 U3084 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3091) );
  NAND2_X1 U3085 ( .A1(n2491), .A2(n3091), .ZN(n2435) );
  NAND2_X1 U3086 ( .A1(n2438), .A2(IR_REG_31__SCAN_IN), .ZN(n2450) );
  MUX2_X1 U3087 ( .A(DATAI_3_), .B(n4503), .S(n2501), .Z(n3257) );
  NAND2_X1 U3088 ( .A1(n2838), .A2(n3257), .ZN(n2439) );
  NAND2_X1 U3089 ( .A1(n3117), .A2(n2439), .ZN(n2441) );
  OR2_X1 U3090 ( .A1(n2838), .A2(n3257), .ZN(n2440) );
  NAND2_X1 U3091 ( .A1(n2422), .A2(REG0_REG_4__SCAN_IN), .ZN(n2444) );
  INV_X1 U3092 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2442) );
  OR2_X1 U3093 ( .A1(n2423), .A2(n2442), .ZN(n2443) );
  NAND2_X1 U3094 ( .A1(n2444), .A2(n2443), .ZN(n2446) );
  NOR2_X1 U3095 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2445) );
  NOR2_X1 U3096 ( .A1(n2457), .A2(n2445), .ZN(n3158) );
  NOR2_X1 U3097 ( .A1(n2446), .A2(n2366), .ZN(n2448) );
  NAND2_X1 U3098 ( .A1(n2421), .A2(REG1_REG_4__SCAN_IN), .ZN(n2447) );
  INV_X1 U3099 ( .A(DATAI_4_), .ZN(n2970) );
  NAND2_X1 U3100 ( .A1(n2450), .A2(n2449), .ZN(n2451) );
  NAND2_X1 U3101 ( .A1(n2451), .A2(IR_REG_31__SCAN_IN), .ZN(n2453) );
  XNOR2_X1 U3102 ( .A(n2453), .B(n2452), .ZN(n3103) );
  MUX2_X1 U3103 ( .A(n2970), .B(n3103), .S(n2501), .Z(n3149) );
  NAND2_X1 U3104 ( .A1(n2825), .A2(n3149), .ZN(n3958) );
  INV_X1 U3105 ( .A(n3926), .ZN(n2455) );
  NAND2_X1 U3106 ( .A1(n2825), .A2(n2454), .ZN(n2456) );
  NAND2_X1 U3107 ( .A1(n2547), .A2(REG0_REG_5__SCAN_IN), .ZN(n2465) );
  NAND2_X1 U3108 ( .A1(n3864), .A2(REG1_REG_5__SCAN_IN), .ZN(n2464) );
  INV_X1 U3109 ( .A(n2457), .ZN(n2459) );
  INV_X1 U3110 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2458) );
  NAND2_X1 U3111 ( .A1(n2459), .A2(n2458), .ZN(n2460) );
  AND2_X1 U3112 ( .A1(n2460), .A2(n2471), .ZN(n3247) );
  NAND2_X1 U3113 ( .A1(n2491), .A2(n3247), .ZN(n2463) );
  INV_X1 U3114 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2461) );
  OR2_X1 U3115 ( .A1(n2423), .A2(n2461), .ZN(n2462) );
  NAND4_X1 U3116 ( .A1(n2465), .A2(n2464), .A3(n2463), .A4(n2462), .ZN(n4044)
         );
  NAND2_X1 U3117 ( .A1(n2466), .A2(IR_REG_31__SCAN_IN), .ZN(n2467) );
  XNOR2_X1 U3118 ( .A(n2467), .B(IR_REG_5__SCAN_IN), .ZN(n4502) );
  MUX2_X1 U3119 ( .A(DATAI_5_), .B(n4502), .S(n2501), .Z(n3246) );
  OR2_X1 U3120 ( .A1(n4044), .A2(n3246), .ZN(n2468) );
  NAND2_X1 U3121 ( .A1(n3078), .A2(n2468), .ZN(n2470) );
  NAND2_X1 U3122 ( .A1(n4044), .A2(n3246), .ZN(n2469) );
  NAND2_X1 U3123 ( .A1(n2470), .A2(n2469), .ZN(n3170) );
  NAND2_X1 U3124 ( .A1(n2422), .A2(REG0_REG_6__SCAN_IN), .ZN(n2476) );
  NAND2_X1 U3125 ( .A1(n3864), .A2(REG1_REG_6__SCAN_IN), .ZN(n2475) );
  AND2_X1 U3126 ( .A1(n2471), .A2(n3017), .ZN(n2472) );
  NOR2_X1 U3127 ( .A1(n2479), .A2(n2472), .ZN(n3356) );
  NAND2_X1 U3128 ( .A1(n2491), .A2(n3356), .ZN(n2474) );
  INV_X1 U3129 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3358) );
  OR2_X1 U3130 ( .A1(n2759), .A2(n3358), .ZN(n2473) );
  NOR2_X1 U3131 ( .A1(n2466), .A2(IR_REG_5__SCAN_IN), .ZN(n2486) );
  OR2_X1 U3132 ( .A1(n2486), .A2(n2765), .ZN(n2477) );
  XNOR2_X1 U3133 ( .A(n2477), .B(IR_REG_6__SCAN_IN), .ZN(n4501) );
  MUX2_X1 U3134 ( .A(DATAI_6_), .B(n4501), .S(n2501), .Z(n3355) );
  AND2_X1 U3135 ( .A1(n4043), .A2(n3355), .ZN(n2478) );
  OAI22_X1 U3136 ( .A1(n3170), .A2(n2478), .B1(n3355), .B2(n4043), .ZN(n3201)
         );
  NAND2_X1 U3137 ( .A1(n2422), .A2(REG0_REG_7__SCAN_IN), .ZN(n2484) );
  NAND2_X1 U3138 ( .A1(n3864), .A2(REG1_REG_7__SCAN_IN), .ZN(n2483) );
  OR2_X1 U3139 ( .A1(n2479), .A2(REG3_REG_7__SCAN_IN), .ZN(n2480) );
  AND2_X1 U3140 ( .A1(n2489), .A2(n2480), .ZN(n3217) );
  NAND2_X1 U3141 ( .A1(n2491), .A2(n3217), .ZN(n2482) );
  INV_X1 U3142 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4092) );
  OR2_X1 U3143 ( .A1(n2759), .A2(n4092), .ZN(n2481) );
  NAND4_X1 U3144 ( .A1(n2484), .A2(n2483), .A3(n2482), .A4(n2481), .ZN(n4042)
         );
  INV_X1 U3145 ( .A(DATAI_7_), .ZN(n2487) );
  NAND2_X1 U3146 ( .A1(n2486), .A2(n2485), .ZN(n2510) );
  NAND2_X1 U3147 ( .A1(n2510), .A2(IR_REG_31__SCAN_IN), .ZN(n2498) );
  XNOR2_X1 U31480 ( .A(n2498), .B(n2497), .ZN(n4093) );
  MUX2_X1 U31490 ( .A(n2487), .B(n4093), .S(n2501), .Z(n3215) );
  OR2_X1 U3150 ( .A1(n4042), .A2(n3215), .ZN(n3961) );
  NAND2_X1 U3151 ( .A1(n4042), .A2(n3215), .ZN(n3967) );
  INV_X1 U3152 ( .A(n3215), .ZN(n3195) );
  NAND2_X1 U3153 ( .A1(n4042), .A2(n3195), .ZN(n2488) );
  NAND2_X1 U3154 ( .A1(n2489), .A2(n5056), .ZN(n2490) );
  AND2_X1 U3155 ( .A1(n2503), .A2(n2490), .ZN(n4645) );
  NAND2_X1 U3156 ( .A1(n2491), .A2(n4645), .ZN(n2496) );
  NAND2_X1 U3157 ( .A1(n3864), .A2(REG1_REG_8__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U3158 ( .A1(n2422), .A2(REG0_REG_8__SCAN_IN), .ZN(n2494) );
  INV_X1 U3159 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2492) );
  OR2_X1 U3160 ( .A1(n2759), .A2(n2492), .ZN(n2493) );
  NAND2_X1 U3161 ( .A1(n2498), .A2(n2497), .ZN(n2499) );
  NAND2_X1 U3162 ( .A1(n2499), .A2(IR_REG_31__SCAN_IN), .ZN(n2500) );
  XNOR2_X1 U3163 ( .A(n2500), .B(IR_REG_8__SCAN_IN), .ZN(n4533) );
  MUX2_X1 U3164 ( .A(DATAI_8_), .B(n4533), .S(n2501), .Z(n3308) );
  AND2_X1 U3165 ( .A1(n2503), .A2(n2502), .ZN(n2504) );
  OR2_X1 U3166 ( .A1(n2504), .A2(n2514), .ZN(n3295) );
  INV_X1 U3167 ( .A(n3295), .ZN(n3330) );
  NAND2_X1 U3168 ( .A1(n2491), .A2(n3330), .ZN(n2509) );
  NAND2_X1 U3169 ( .A1(n3864), .A2(REG1_REG_9__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U3170 ( .A1(n2422), .A2(REG0_REG_9__SCAN_IN), .ZN(n2507) );
  INV_X1 U3171 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2505) );
  OR2_X1 U3172 ( .A1(n2759), .A2(n2505), .ZN(n2506) );
  NAND4_X1 U3173 ( .A1(n2509), .A2(n2508), .A3(n2507), .A4(n2506), .ZN(n4040)
         );
  NAND2_X1 U3174 ( .A1(n2521), .A2(IR_REG_31__SCAN_IN), .ZN(n2511) );
  XNOR2_X1 U3175 ( .A(n2511), .B(IR_REG_9__SCAN_IN), .ZN(n4091) );
  MUX2_X1 U3176 ( .A(DATAI_9_), .B(n4091), .S(n2986), .Z(n3292) );
  AND2_X1 U3177 ( .A1(n4040), .A2(n3292), .ZN(n2513) );
  OR2_X1 U3178 ( .A1(n4040), .A2(n3292), .ZN(n2512) );
  NOR2_X1 U3179 ( .A1(n2514), .A2(REG3_REG_10__SCAN_IN), .ZN(n2515) );
  OR2_X1 U3180 ( .A1(n2524), .A2(n2515), .ZN(n2964) );
  INV_X1 U3181 ( .A(n2964), .ZN(n4638) );
  NAND2_X1 U3182 ( .A1(n2491), .A2(n4638), .ZN(n2520) );
  NAND2_X1 U3183 ( .A1(n3864), .A2(REG1_REG_10__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U3184 ( .A1(n2547), .A2(REG0_REG_10__SCAN_IN), .ZN(n2518) );
  INV_X1 U3185 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2516) );
  NOR2_X1 U3186 ( .A1(n2521), .A2(IR_REG_9__SCAN_IN), .ZN(n2532) );
  OR2_X1 U3187 ( .A1(n2532), .A2(n2765), .ZN(n2522) );
  XNOR2_X1 U3188 ( .A(n2522), .B(IR_REG_10__SCAN_IN), .ZN(n4554) );
  MUX2_X1 U3189 ( .A(DATAI_10_), .B(n4554), .S(n2986), .Z(n3451) );
  INV_X1 U3190 ( .A(n4039), .ZN(n2523) );
  NAND2_X1 U3191 ( .A1(n2547), .A2(REG0_REG_11__SCAN_IN), .ZN(n2530) );
  NAND2_X1 U3192 ( .A1(n3864), .A2(REG1_REG_11__SCAN_IN), .ZN(n2529) );
  OR2_X1 U3193 ( .A1(n2524), .A2(REG3_REG_11__SCAN_IN), .ZN(n2525) );
  AND2_X1 U3194 ( .A1(n2535), .A2(n2525), .ZN(n3432) );
  NAND2_X1 U3195 ( .A1(n2491), .A2(n3432), .ZN(n2528) );
  INV_X1 U3196 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2526) );
  OR2_X1 U3197 ( .A1(n2423), .A2(n2526), .ZN(n2527) );
  NAND4_X1 U3198 ( .A1(n2530), .A2(n2529), .A3(n2528), .A4(n2527), .ZN(n4038)
         );
  INV_X1 U3199 ( .A(DATAI_11_), .ZN(n2534) );
  NAND2_X1 U3200 ( .A1(n2532), .A2(n2531), .ZN(n2533) );
  NAND2_X1 U3201 ( .A1(n2533), .A2(IR_REG_31__SCAN_IN), .ZN(n2542) );
  XNOR2_X1 U3202 ( .A(n2542), .B(IR_REG_11__SCAN_IN), .ZN(n4090) );
  MUX2_X1 U3203 ( .A(n2534), .B(n4672), .S(n2986), .Z(n3430) );
  OR2_X1 U3204 ( .A1(n4038), .A2(n3430), .ZN(n3375) );
  NAND2_X1 U3205 ( .A1(n4038), .A2(n3430), .ZN(n3981) );
  INV_X1 U3206 ( .A(n3430), .ZN(n3424) );
  OR2_X1 U3207 ( .A1(n4038), .A2(n3424), .ZN(n3389) );
  NAND2_X1 U3208 ( .A1(n2547), .A2(REG0_REG_12__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U3209 ( .A1(n3864), .A2(REG1_REG_12__SCAN_IN), .ZN(n2539) );
  NAND2_X1 U32100 ( .A1(n2535), .A2(n4865), .ZN(n2536) );
  AND2_X1 U32110 ( .A1(n2549), .A2(n2536), .ZN(n3539) );
  NAND2_X1 U32120 ( .A1(n2491), .A2(n3539), .ZN(n2538) );
  INV_X1 U32130 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3396) );
  OR2_X1 U32140 ( .A1(n2759), .A2(n3396), .ZN(n2537) );
  NAND4_X1 U32150 ( .A1(n2540), .A2(n2539), .A3(n2538), .A4(n2537), .ZN(n4037)
         );
  INV_X1 U32160 ( .A(IR_REG_11__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U32170 ( .A1(n2542), .A2(n2541), .ZN(n2543) );
  NAND2_X1 U32180 ( .A1(n2543), .A2(IR_REG_31__SCAN_IN), .ZN(n2544) );
  XNOR2_X1 U32190 ( .A(n2544), .B(IR_REG_12__SCAN_IN), .ZN(n4575) );
  OR2_X1 U32200 ( .A1(n4037), .A2(n3490), .ZN(n2545) );
  AND2_X1 U32210 ( .A1(n3389), .A2(n2545), .ZN(n2546) );
  NAND2_X1 U32220 ( .A1(n3864), .A2(REG1_REG_13__SCAN_IN), .ZN(n2555) );
  NAND2_X1 U32230 ( .A1(n2547), .A2(REG0_REG_13__SCAN_IN), .ZN(n2554) );
  NAND2_X1 U32240 ( .A1(n2549), .A2(n2548), .ZN(n2550) );
  AND2_X1 U32250 ( .A1(n2558), .A2(n2550), .ZN(n3512) );
  NAND2_X1 U32260 ( .A1(n2491), .A2(n3512), .ZN(n2553) );
  INV_X1 U32270 ( .A(REG2_REG_13__SCAN_IN), .ZN(n2551) );
  OR2_X1 U32280 ( .A1(n2759), .A2(n2551), .ZN(n2552) );
  NAND4_X1 U32290 ( .A1(n2555), .A2(n2554), .A3(n2553), .A4(n2552), .ZN(n4036)
         );
  OR2_X1 U32300 ( .A1(n2556), .A2(n2765), .ZN(n2557) );
  XNOR2_X1 U32310 ( .A(n2557), .B(IR_REG_13__SCAN_IN), .ZN(n4105) );
  MUX2_X1 U32320 ( .A(DATAI_13_), .B(n4105), .S(n2986), .Z(n3504) );
  NOR2_X1 U32330 ( .A1(n4036), .A2(n3504), .ZN(n3542) );
  NAND2_X1 U32340 ( .A1(n2547), .A2(REG0_REG_14__SCAN_IN), .ZN(n2564) );
  NAND2_X1 U32350 ( .A1(n3864), .A2(REG1_REG_14__SCAN_IN), .ZN(n2563) );
  AND2_X1 U32360 ( .A1(n2558), .A2(n4743), .ZN(n2559) );
  NOR2_X1 U32370 ( .A1(n2570), .A2(n2559), .ZN(n3588) );
  NAND2_X1 U32380 ( .A1(n2491), .A2(n3588), .ZN(n2562) );
  INV_X1 U32390 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2560) );
  OR2_X1 U32400 ( .A1(n2759), .A2(n2560), .ZN(n2561) );
  NAND4_X1 U32410 ( .A1(n2564), .A2(n2563), .A3(n2562), .A4(n2561), .ZN(n4035)
         );
  INV_X1 U32420 ( .A(DATAI_14_), .ZN(n4668) );
  NAND2_X1 U32430 ( .A1(n2565), .A2(IR_REG_31__SCAN_IN), .ZN(n2566) );
  XNOR2_X1 U32440 ( .A(n2566), .B(IR_REG_14__SCAN_IN), .ZN(n4081) );
  INV_X1 U32450 ( .A(n4081), .ZN(n4669) );
  MUX2_X1 U32460 ( .A(n4668), .B(n4669), .S(n2986), .Z(n3603) );
  OR2_X1 U32470 ( .A1(n3542), .A2(n2238), .ZN(n2567) );
  NOR2_X1 U32480 ( .A1(n3543), .A2(n2567), .ZN(n2569) );
  OR2_X1 U32490 ( .A1(n4035), .A2(n3603), .ZN(n3868) );
  NAND2_X1 U32500 ( .A1(n4035), .A2(n3603), .ZN(n3869) );
  NAND2_X1 U32510 ( .A1(n3868), .A2(n3869), .ZN(n3552) );
  NAND2_X1 U32520 ( .A1(n4036), .A2(n3504), .ZN(n3544) );
  AND2_X1 U32530 ( .A1(n3552), .A2(n3544), .ZN(n3545) );
  NOR2_X1 U32540 ( .A1(n2238), .A2(n3545), .ZN(n2568) );
  NOR2_X1 U32550 ( .A1(n2569), .A2(n2568), .ZN(n3438) );
  NAND2_X1 U32560 ( .A1(n2547), .A2(REG0_REG_15__SCAN_IN), .ZN(n2576) );
  NAND2_X1 U32570 ( .A1(n3864), .A2(REG1_REG_15__SCAN_IN), .ZN(n2575) );
  OR2_X1 U32580 ( .A1(n2570), .A2(REG3_REG_15__SCAN_IN), .ZN(n2571) );
  AND2_X1 U32590 ( .A1(n2571), .A2(n2580), .ZN(n3858) );
  NAND2_X1 U32600 ( .A1(n2491), .A2(n3858), .ZN(n2574) );
  INV_X1 U32610 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2572) );
  OR2_X1 U32620 ( .A1(n2759), .A2(n2572), .ZN(n2573) );
  NAND4_X1 U32630 ( .A1(n2576), .A2(n2575), .A3(n2574), .A4(n2573), .ZN(n4034)
         );
  NAND2_X1 U32640 ( .A1(n2237), .A2(IR_REG_31__SCAN_IN), .ZN(n2588) );
  XNOR2_X1 U32650 ( .A(n2588), .B(IR_REG_15__SCAN_IN), .ZN(n4109) );
  MUX2_X1 U32660 ( .A(DATAI_15_), .B(n4109), .S(n2986), .Z(n3634) );
  NAND2_X1 U32670 ( .A1(n4034), .A2(n3634), .ZN(n2577) );
  NOR2_X1 U32680 ( .A1(n4034), .A2(n3634), .ZN(n2578) );
  NAND2_X1 U32690 ( .A1(n2580), .A2(n5057), .ZN(n2581) );
  NAND2_X1 U32700 ( .A1(n2582), .A2(n2581), .ZN(n4521) );
  INV_X1 U32710 ( .A(n4521), .ZN(n2583) );
  NAND2_X1 U32720 ( .A1(n2491), .A2(n2583), .ZN(n2587) );
  NAND2_X1 U32730 ( .A1(n3864), .A2(REG1_REG_16__SCAN_IN), .ZN(n2586) );
  NAND2_X1 U32740 ( .A1(n2547), .A2(REG0_REG_16__SCAN_IN), .ZN(n2585) );
  INV_X1 U32750 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3476) );
  OR2_X1 U32760 ( .A1(n2423), .A2(n3476), .ZN(n2584) );
  INV_X1 U32770 ( .A(DATAI_16_), .ZN(n5053) );
  NAND2_X1 U32780 ( .A1(n2588), .A2(n4874), .ZN(n2589) );
  NAND2_X1 U32790 ( .A1(n2589), .A2(IR_REG_31__SCAN_IN), .ZN(n2590) );
  XNOR2_X1 U32800 ( .A(n2590), .B(IR_REG_16__SCAN_IN), .ZN(n4085) );
  MUX2_X1 U32810 ( .A(n5053), .B(n4666), .S(n2986), .Z(n4508) );
  OR2_X1 U32820 ( .A1(n4033), .A2(n4508), .ZN(n3994) );
  NAND2_X1 U32830 ( .A1(n4033), .A2(n4508), .ZN(n3990) );
  NAND2_X1 U32840 ( .A1(n3994), .A2(n3990), .ZN(n3479) );
  AOI21_X1 U32850 ( .B1(n3832), .B2(n3790), .A(n3570), .ZN(n2593) );
  NOR2_X1 U32860 ( .A1(n2594), .A2(REG3_REG_18__SCAN_IN), .ZN(n2595) );
  OR2_X1 U32870 ( .A1(n2617), .A2(n2595), .ZN(n4369) );
  INV_X1 U32880 ( .A(n4369), .ZN(n2596) );
  NAND2_X1 U32890 ( .A1(n2596), .A2(n2491), .ZN(n2600) );
  NAND2_X1 U32900 ( .A1(n2547), .A2(REG0_REG_18__SCAN_IN), .ZN(n2599) );
  NAND2_X1 U32910 ( .A1(n3864), .A2(REG1_REG_18__SCAN_IN), .ZN(n2598) );
  INV_X1 U32920 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4370) );
  OR2_X1 U32930 ( .A1(n2759), .A2(n4370), .ZN(n2597) );
  INV_X1 U32940 ( .A(DATAI_18_), .ZN(n5032) );
  INV_X1 U32950 ( .A(IR_REG_17__SCAN_IN), .ZN(n2601) );
  INV_X1 U32960 ( .A(n2612), .ZN(n2603) );
  NAND2_X1 U32970 ( .A1(n2603), .A2(IR_REG_31__SCAN_IN), .ZN(n2604) );
  XNOR2_X1 U32980 ( .A(n2604), .B(n2611), .ZN(n4123) );
  MUX2_X1 U32990 ( .A(n5032), .B(n4123), .S(n2986), .Z(n4359) );
  OR2_X1 U33000 ( .A1(n4337), .A2(n4359), .ZN(n4329) );
  NAND2_X1 U33010 ( .A1(n4337), .A2(n4359), .ZN(n4330) );
  NAND2_X1 U33020 ( .A1(n4329), .A2(n4330), .ZN(n4353) );
  INV_X1 U33030 ( .A(n4359), .ZN(n4363) );
  INV_X1 U33040 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4346) );
  NAND2_X1 U33050 ( .A1(n3864), .A2(REG1_REG_19__SCAN_IN), .ZN(n2608) );
  NAND2_X1 U33060 ( .A1(n2547), .A2(REG0_REG_19__SCAN_IN), .ZN(n2607) );
  AND2_X1 U33070 ( .A1(n2608), .A2(n2607), .ZN(n2610) );
  INV_X1 U33080 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4824) );
  XNOR2_X1 U33090 ( .A(n2617), .B(n4824), .ZN(n4344) );
  NAND2_X1 U33100 ( .A1(n4344), .A2(n2491), .ZN(n2609) );
  MUX2_X1 U33110 ( .A(DATAI_19_), .B(n4499), .S(n2986), .Z(n3668) );
  NOR2_X1 U33120 ( .A1(n4032), .A2(n3668), .ZN(n4307) );
  INV_X1 U33130 ( .A(REG2_REG_20__SCAN_IN), .ZN(n2621) );
  NAND2_X1 U33140 ( .A1(n2547), .A2(REG0_REG_20__SCAN_IN), .ZN(n2614) );
  NAND2_X1 U33150 ( .A1(n3864), .A2(REG1_REG_20__SCAN_IN), .ZN(n2613) );
  AND2_X1 U33160 ( .A1(n2614), .A2(n2613), .ZN(n2620) );
  NAND2_X1 U33170 ( .A1(n2617), .A2(REG3_REG_19__SCAN_IN), .ZN(n2615) );
  INV_X1 U33180 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3810) );
  NAND2_X1 U33190 ( .A1(n2615), .A2(n3810), .ZN(n2618) );
  AND2_X1 U33200 ( .A1(REG3_REG_19__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2616) );
  NAND2_X1 U33210 ( .A1(n2618), .A2(n2625), .ZN(n4317) );
  OR2_X1 U33220 ( .A1(n4317), .A2(n2699), .ZN(n2619) );
  INV_X1 U33230 ( .A(DATAI_20_), .ZN(n5062) );
  NAND2_X1 U33240 ( .A1(n4421), .A2(n4431), .ZN(n3902) );
  NAND2_X1 U33250 ( .A1(n4032), .A2(n3668), .ZN(n4308) );
  OR2_X1 U33260 ( .A1(n4421), .A2(n4431), .ZN(n3903) );
  INV_X1 U33270 ( .A(REG3_REG_21__SCAN_IN), .ZN(n5031) );
  NAND2_X1 U33280 ( .A1(n2625), .A2(n5031), .ZN(n2626) );
  NAND2_X1 U33290 ( .A1(n2639), .A2(n2626), .ZN(n4293) );
  AOI22_X1 U33300 ( .A1(n2547), .A2(REG0_REG_21__SCAN_IN), .B1(n3864), .B2(
        REG1_REG_21__SCAN_IN), .ZN(n2629) );
  INV_X1 U33310 ( .A(REG2_REG_21__SCAN_IN), .ZN(n2627) );
  OR2_X1 U33320 ( .A1(n2759), .A2(n2627), .ZN(n2628) );
  NAND2_X1 U33330 ( .A1(n3863), .A2(DATAI_21_), .ZN(n4298) );
  NAND2_X1 U33340 ( .A1(n4433), .A2(n4419), .ZN(n2631) );
  INV_X1 U33350 ( .A(n4433), .ZN(n3819) );
  XNOR2_X1 U33360 ( .A(n2639), .B(REG3_REG_22__SCAN_IN), .ZN(n4270) );
  NAND2_X1 U33370 ( .A1(n4270), .A2(n2491), .ZN(n2636) );
  INV_X1 U33380 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4272) );
  NAND2_X1 U33390 ( .A1(n2547), .A2(REG0_REG_22__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U33400 ( .A1(n3864), .A2(REG1_REG_22__SCAN_IN), .ZN(n2632) );
  OAI211_X1 U33410 ( .C1(n4272), .C2(n2423), .A(n2633), .B(n2632), .ZN(n2634)
         );
  INV_X1 U33420 ( .A(n2634), .ZN(n2635) );
  NAND2_X1 U33430 ( .A1(n3863), .A2(DATAI_22_), .ZN(n4279) );
  NAND2_X1 U33440 ( .A1(n4291), .A2(n4279), .ZN(n2741) );
  NAND2_X1 U33450 ( .A1(n4250), .A2(n2741), .ZN(n4275) );
  NAND2_X1 U33460 ( .A1(n4267), .A2(n4275), .ZN(n4266) );
  NAND2_X1 U33470 ( .A1(n4266), .A2(n2371), .ZN(n4241) );
  INV_X1 U33480 ( .A(n2639), .ZN(n2637) );
  AOI21_X1 U33490 ( .B1(n2637), .B2(REG3_REG_22__SCAN_IN), .A(
        REG3_REG_23__SCAN_IN), .ZN(n2640) );
  NAND2_X1 U33500 ( .A1(REG3_REG_23__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2638) );
  OR2_X1 U33510 ( .A1(n2640), .A2(n2647), .ZN(n4260) );
  INV_X1 U33520 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4261) );
  NAND2_X1 U3353 ( .A1(n3864), .A2(REG1_REG_23__SCAN_IN), .ZN(n2642) );
  NAND2_X1 U33540 ( .A1(n2547), .A2(REG0_REG_23__SCAN_IN), .ZN(n2641) );
  OAI211_X1 U3355 ( .C1(n4261), .C2(n2759), .A(n2642), .B(n2641), .ZN(n2643)
         );
  INV_X1 U3356 ( .A(n2643), .ZN(n2644) );
  INV_X1 U3357 ( .A(n4402), .ZN(n3820) );
  NAND2_X1 U3358 ( .A1(n3863), .A2(DATAI_23_), .ZN(n4257) );
  NAND2_X1 U3359 ( .A1(n3820), .A2(n4257), .ZN(n2646) );
  NOR2_X1 U3360 ( .A1(n2647), .A2(REG3_REG_24__SCAN_IN), .ZN(n2648) );
  OR2_X1 U3361 ( .A1(n2655), .A2(n2648), .ZN(n4232) );
  INV_X1 U3362 ( .A(REG2_REG_24__SCAN_IN), .ZN(n2651) );
  NAND2_X1 U3363 ( .A1(n2547), .A2(REG0_REG_24__SCAN_IN), .ZN(n2650) );
  NAND2_X1 U3364 ( .A1(n3864), .A2(REG1_REG_24__SCAN_IN), .ZN(n2649) );
  OAI211_X1 U3365 ( .C1(n2651), .C2(n2759), .A(n2650), .B(n2649), .ZN(n2652)
         );
  INV_X1 U3366 ( .A(n2652), .ZN(n2653) );
  NAND2_X1 U3367 ( .A1(n3863), .A2(DATAI_24_), .ZN(n4236) );
  NAND2_X1 U3368 ( .A1(n4210), .A2(n4401), .ZN(n2654) );
  INV_X1 U3369 ( .A(n4210), .ZN(n4253) );
  OR2_X1 U3370 ( .A1(n2655), .A2(REG3_REG_25__SCAN_IN), .ZN(n2656) );
  NAND2_X1 U3371 ( .A1(n4217), .A2(n2491), .ZN(n2662) );
  INV_X1 U3372 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2659) );
  NAND2_X1 U3373 ( .A1(n3864), .A2(REG1_REG_25__SCAN_IN), .ZN(n2658) );
  NAND2_X1 U3374 ( .A1(n2547), .A2(REG0_REG_25__SCAN_IN), .ZN(n2657) );
  OAI211_X1 U3375 ( .C1(n2659), .C2(n2759), .A(n2658), .B(n2657), .ZN(n2660)
         );
  INV_X1 U3376 ( .A(n2660), .ZN(n2661) );
  INV_X1 U3377 ( .A(n4231), .ZN(n4405) );
  NAND2_X1 U3378 ( .A1(n3863), .A2(DATAI_25_), .ZN(n3704) );
  NAND2_X1 U3379 ( .A1(n4405), .A2(n3704), .ZN(n2664) );
  INV_X1 U3380 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3842) );
  NAND2_X1 U3381 ( .A1(n2665), .A2(n3842), .ZN(n2666) );
  NAND2_X1 U3382 ( .A1(n2683), .A2(n2666), .ZN(n4200) );
  INV_X1 U3383 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4201) );
  NAND2_X1 U3384 ( .A1(n2547), .A2(REG0_REG_26__SCAN_IN), .ZN(n2668) );
  NAND2_X1 U3385 ( .A1(n3864), .A2(REG1_REG_26__SCAN_IN), .ZN(n2667) );
  OAI211_X1 U3386 ( .C1(n4201), .C2(n2759), .A(n2668), .B(n2667), .ZN(n2669)
         );
  INV_X1 U3387 ( .A(n2669), .ZN(n2670) );
  NAND2_X1 U3388 ( .A1(n3863), .A2(DATAI_26_), .ZN(n3843) );
  NAND2_X1 U3389 ( .A1(n4187), .A2(n2672), .ZN(n2673) );
  XNOR2_X1 U3390 ( .A(n2683), .B(REG3_REG_27__SCAN_IN), .ZN(n4179) );
  NAND2_X1 U3391 ( .A1(n4179), .A2(n2491), .ZN(n2679) );
  INV_X1 U3392 ( .A(REG2_REG_27__SCAN_IN), .ZN(n2676) );
  NAND2_X1 U3393 ( .A1(n3864), .A2(REG1_REG_27__SCAN_IN), .ZN(n2675) );
  NAND2_X1 U3394 ( .A1(n2547), .A2(REG0_REG_27__SCAN_IN), .ZN(n2674) );
  OAI211_X1 U3395 ( .C1(n2676), .C2(n2759), .A(n2675), .B(n2674), .ZN(n2677)
         );
  INV_X1 U3396 ( .A(n2677), .ZN(n2678) );
  INV_X1 U3397 ( .A(n4195), .ZN(n4159) );
  INV_X1 U3398 ( .A(DATAI_27_), .ZN(n2680) );
  NOR2_X1 U3399 ( .A1(n2986), .A2(n2680), .ZN(n4384) );
  NOR2_X1 U3400 ( .A1(n4159), .A2(n4384), .ZN(n2681) );
  INV_X1 U3401 ( .A(n4384), .ZN(n4182) );
  NAND2_X1 U3402 ( .A1(REG3_REG_28__SCAN_IN), .A2(REG3_REG_27__SCAN_IN), .ZN(
        n2682) );
  INV_X1 U3403 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3743) );
  INV_X1 U3404 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3733) );
  OAI21_X1 U3405 ( .B1(n2683), .B2(n3743), .A(n3733), .ZN(n2684) );
  NAND2_X1 U3406 ( .A1(n4160), .A2(n2491), .ZN(n2690) );
  INV_X1 U3407 ( .A(REG2_REG_28__SCAN_IN), .ZN(n2687) );
  NAND2_X1 U3408 ( .A1(n2547), .A2(REG0_REG_28__SCAN_IN), .ZN(n2686) );
  NAND2_X1 U3409 ( .A1(n3864), .A2(REG1_REG_28__SCAN_IN), .ZN(n2685) );
  OAI211_X1 U3410 ( .C1(n2687), .C2(n2759), .A(n2686), .B(n2685), .ZN(n2688)
         );
  INV_X1 U3411 ( .A(n2688), .ZN(n2689) );
  INV_X1 U3412 ( .A(DATAI_28_), .ZN(n4847) );
  NOR2_X1 U3413 ( .A1(n2986), .A2(n4847), .ZN(n2691) );
  INV_X1 U3414 ( .A(n3888), .ZN(n2748) );
  NAND2_X1 U3415 ( .A1(n4030), .A2(n4163), .ZN(n2747) );
  NAND2_X1 U3416 ( .A1(n2748), .A2(n2747), .ZN(n3943) );
  INV_X1 U3417 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U3418 ( .A1(n2547), .A2(REG0_REG_29__SCAN_IN), .ZN(n2694) );
  INV_X1 U3419 ( .A(n2759), .ZN(n2692) );
  NAND2_X1 U3420 ( .A1(n2692), .A2(REG2_REG_29__SCAN_IN), .ZN(n2693) );
  OAI211_X1 U3421 ( .C1(n2696), .C2(n2695), .A(n2694), .B(n2693), .ZN(n2697)
         );
  INV_X1 U3422 ( .A(n2697), .ZN(n2698) );
  OAI21_X1 U3423 ( .B1(n4150), .B2(n2699), .A(n2698), .ZN(n4158) );
  NAND2_X1 U3424 ( .A1(n3863), .A2(DATAI_29_), .ZN(n3886) );
  XNOR2_X1 U3425 ( .A(n4158), .B(n3886), .ZN(n3941) );
  NAND2_X1 U3426 ( .A1(n2703), .A2(IR_REG_31__SCAN_IN), .ZN(n2702) );
  INV_X1 U3427 ( .A(IR_REG_21__SCAN_IN), .ZN(n2701) );
  MUX2_X1 U3428 ( .A(n2702), .B(IR_REG_31__SCAN_IN), .S(n2701), .Z(n2704) );
  INV_X1 U3429 ( .A(n2770), .ZN(n2710) );
  NAND2_X1 U3430 ( .A1(n2704), .A2(n2710), .ZN(n2781) );
  NAND2_X1 U3431 ( .A1(n2706), .A2(n2705), .ZN(n2707) );
  NAND2_X1 U3432 ( .A1(n2707), .A2(IR_REG_31__SCAN_IN), .ZN(n2709) );
  INV_X1 U3433 ( .A(IR_REG_20__SCAN_IN), .ZN(n2708) );
  XNOR2_X2 U3434 ( .A(n2709), .B(n2708), .ZN(n4016) );
  INV_X1 U3435 ( .A(IR_REG_22__SCAN_IN), .ZN(n2769) );
  INV_X1 U3436 ( .A(n2828), .ZN(n4497) );
  XNOR2_X1 U3437 ( .A(n2832), .B(n4497), .ZN(n2712) );
  INV_X1 U3438 ( .A(n4499), .ZN(n4133) );
  NAND2_X1 U3439 ( .A1(n2712), .A2(n4133), .ZN(n3554) );
  AND2_X1 U3440 ( .A1(n4016), .A2(n4499), .ZN(n3223) );
  INV_X1 U3441 ( .A(n4700), .ZN(n4682) );
  NAND2_X1 U3442 ( .A1(n4145), .A2(n4443), .ZN(n2762) );
  OR2_X1 U3443 ( .A1(n2714), .A2(n3220), .ZN(n3945) );
  OAI21_X1 U3444 ( .B1(n2713), .B2(n3945), .A(n2715), .ZN(n3130) );
  INV_X1 U3445 ( .A(n3128), .ZN(n3925) );
  NAND2_X1 U3446 ( .A1(n3130), .A2(n3925), .ZN(n2716) );
  NAND2_X1 U3447 ( .A1(n2716), .A2(n3950), .ZN(n3118) );
  OR2_X1 U3448 ( .A1(n2838), .A2(n3122), .ZN(n3955) );
  NAND2_X1 U3449 ( .A1(n2838), .A2(n3122), .ZN(n3952) );
  AND2_X1 U3450 ( .A1(n3955), .A2(n3952), .ZN(n3923) );
  NAND2_X1 U3451 ( .A1(n3118), .A2(n3923), .ZN(n2717) );
  NAND2_X1 U3452 ( .A1(n2717), .A2(n3955), .ZN(n3147) );
  INV_X1 U3453 ( .A(n3956), .ZN(n2718) );
  OR2_X1 U3454 ( .A1(n3147), .A2(n2718), .ZN(n2719) );
  NAND2_X1 U3455 ( .A1(n2719), .A2(n3958), .ZN(n3080) );
  AND2_X1 U3456 ( .A1(n4044), .A2(n2256), .ZN(n3959) );
  OR2_X1 U3457 ( .A1(n3080), .A2(n3959), .ZN(n2720) );
  OR2_X1 U34580 ( .A1(n4044), .A2(n2256), .ZN(n3975) );
  NAND2_X1 U34590 ( .A1(n4043), .A2(n3188), .ZN(n3171) );
  NOR2_X1 U3460 ( .A1(n4043), .A2(n3188), .ZN(n3962) );
  AOI21_X1 U3461 ( .B1(n3172), .B2(n3171), .A(n3962), .ZN(n3196) );
  NAND2_X1 U3462 ( .A1(n3196), .A2(n3961), .ZN(n2721) );
  NAND2_X1 U3463 ( .A1(n2721), .A2(n3967), .ZN(n3306) );
  INV_X1 U3464 ( .A(n3308), .ZN(n3303) );
  OR2_X1 U3465 ( .A1(n4041), .A2(n3303), .ZN(n3968) );
  NAND2_X1 U3466 ( .A1(n3306), .A2(n3968), .ZN(n2722) );
  NAND2_X1 U34670 ( .A1(n4041), .A2(n3303), .ZN(n3966) );
  NAND2_X1 U3468 ( .A1(n2722), .A2(n3966), .ZN(n3270) );
  INV_X1 U34690 ( .A(n3292), .ZN(n3328) );
  AND2_X1 U3470 ( .A1(n4040), .A2(n3328), .ZN(n3973) );
  OR2_X1 U34710 ( .A1(n4040), .A2(n3328), .ZN(n3969) );
  NAND2_X1 U3472 ( .A1(n2723), .A2(n3969), .ZN(n3450) );
  NAND2_X1 U34730 ( .A1(n4039), .A2(n3447), .ZN(n3982) );
  NAND2_X1 U3474 ( .A1(n3450), .A2(n3982), .ZN(n2724) );
  OR2_X1 U34750 ( .A1(n4039), .A2(n3447), .ZN(n3977) );
  NAND2_X1 U3476 ( .A1(n2724), .A2(n3977), .ZN(n3333) );
  NAND2_X1 U34770 ( .A1(n3333), .A2(n3981), .ZN(n3376) );
  INV_X1 U3478 ( .A(n3490), .ZN(n3537) );
  NAND2_X1 U34790 ( .A1(n4037), .A2(n3537), .ZN(n3387) );
  INV_X1 U3480 ( .A(n3504), .ZN(n3510) );
  NAND2_X1 U34810 ( .A1(n4036), .A2(n3510), .ZN(n3373) );
  NAND2_X1 U3482 ( .A1(n3387), .A2(n3373), .ZN(n3983) );
  INV_X1 U34830 ( .A(n3983), .ZN(n2727) );
  OR2_X1 U3484 ( .A1(n4037), .A2(n3537), .ZN(n3388) );
  NAND2_X1 U34850 ( .A1(n3375), .A2(n3388), .ZN(n2726) );
  OR2_X1 U3486 ( .A1(n4036), .A2(n3510), .ZN(n3374) );
  INV_X1 U34870 ( .A(n3374), .ZN(n2725) );
  AOI21_X1 U3488 ( .B1(n2727), .B2(n2726), .A(n2725), .ZN(n3989) );
  NAND2_X1 U34890 ( .A1(n2728), .A2(n3989), .ZN(n3549) );
  INV_X1 U3490 ( .A(n3552), .ZN(n3919) );
  OR2_X1 U34910 ( .A1(n4034), .A2(n3856), .ZN(n3871) );
  NAND2_X1 U3492 ( .A1(n4034), .A2(n3856), .ZN(n3870) );
  NAND2_X1 U34930 ( .A1(n3871), .A2(n3870), .ZN(n3437) );
  INV_X1 U3494 ( .A(n3868), .ZN(n2729) );
  NOR2_X1 U34950 ( .A1(n3437), .A2(n2729), .ZN(n2730) );
  NAND2_X1 U3496 ( .A1(n3550), .A2(n2730), .ZN(n2731) );
  NAND2_X1 U34970 ( .A1(n2731), .A2(n3870), .ZN(n3480) );
  NAND2_X1 U3498 ( .A1(n3480), .A2(n2591), .ZN(n2732) );
  NAND2_X1 U34990 ( .A1(n4032), .A2(n4342), .ZN(n2733) );
  AND2_X1 U3500 ( .A1(n4330), .A2(n2733), .ZN(n2737) );
  OR2_X1 U35010 ( .A1(n4511), .A2(n3790), .ZN(n4327) );
  NAND2_X1 U3502 ( .A1(n4329), .A2(n4327), .ZN(n2735) );
  NOR2_X1 U35030 ( .A1(n4032), .A2(n4342), .ZN(n2734) );
  AOI21_X1 U3504 ( .B1(n2737), .B2(n2735), .A(n2734), .ZN(n4303) );
  INV_X1 U35050 ( .A(n4431), .ZN(n4313) );
  OR2_X1 U35060 ( .A1(n4421), .A2(n4313), .ZN(n2736) );
  NAND2_X1 U35070 ( .A1(n4244), .A2(n4247), .ZN(n2738) );
  INV_X1 U35080 ( .A(n2737), .ZN(n4245) );
  AND2_X1 U35090 ( .A1(n4511), .A2(n3790), .ZN(n4243) );
  OR2_X1 U35100 ( .A1(n4245), .A2(n4243), .ZN(n3993) );
  AND2_X1 U35110 ( .A1(n4421), .A2(n4313), .ZN(n4246) );
  AOI21_X1 U35120 ( .B1(n4247), .B2(n3993), .A(n4246), .ZN(n3875) );
  NAND2_X1 U35130 ( .A1(n2738), .A2(n3875), .ZN(n2740) );
  OR2_X1 U35140 ( .A1(n4433), .A2(n4298), .ZN(n4248) );
  NAND2_X1 U35150 ( .A1(n4250), .A2(n4248), .ZN(n3999) );
  INV_X1 U35160 ( .A(n3999), .ZN(n2739) );
  NAND2_X1 U35170 ( .A1(n2740), .A2(n2739), .ZN(n2744) );
  NAND2_X1 U35180 ( .A1(n4402), .A2(n4257), .ZN(n2742) );
  NAND2_X1 U35190 ( .A1(n2742), .A2(n2741), .ZN(n4002) );
  AND2_X1 U35200 ( .A1(n4433), .A2(n4298), .ZN(n3997) );
  AND2_X1 U35210 ( .A1(n4250), .A2(n3997), .ZN(n2743) );
  NOR2_X1 U35220 ( .A1(n4002), .A2(n2743), .ZN(n3878) );
  NAND2_X1 U35230 ( .A1(n2744), .A2(n3878), .ZN(n4223) );
  OR2_X1 U35240 ( .A1(n4210), .A2(n4236), .ZN(n3900) );
  OR2_X1 U35250 ( .A1(n4402), .A2(n4257), .ZN(n4222) );
  NAND2_X1 U35260 ( .A1(n4223), .A2(n4001), .ZN(n2745) );
  NAND2_X1 U35270 ( .A1(n4210), .A2(n4236), .ZN(n3901) );
  NAND2_X1 U35280 ( .A1(n2745), .A2(n3901), .ZN(n4208) );
  AND2_X1 U35290 ( .A1(n4231), .A2(n3704), .ZN(n3898) );
  NAND2_X1 U35300 ( .A1(n4213), .A2(n4197), .ZN(n3936) );
  OR2_X1 U35310 ( .A1(n4231), .A2(n3704), .ZN(n4188) );
  NAND2_X1 U35320 ( .A1(n4385), .A2(n3843), .ZN(n3935) );
  INV_X1 U35330 ( .A(n3935), .ZN(n2746) );
  AOI21_X2 U35340 ( .B1(n4189), .B2(n4009), .A(n2746), .ZN(n4171) );
  NOR2_X1 U35350 ( .A1(n4195), .A2(n4384), .ZN(n4007) );
  AOI21_X1 U35360 ( .B1(n4171), .B2(n4170), .A(n3887), .ZN(n2804) );
  INV_X1 U35370 ( .A(n2747), .ZN(n3885) );
  XOR2_X1 U35380 ( .A(n3941), .B(n2749), .Z(n2760) );
  NAND2_X1 U35390 ( .A1(n4497), .A2(n4499), .ZN(n2750) );
  INV_X1 U35400 ( .A(n4016), .ZN(n4498) );
  NAND2_X1 U35410 ( .A1(n3948), .A2(n4498), .ZN(n4020) );
  XNOR2_X1 U35420 ( .A(n2751), .B(IR_REG_27__SCAN_IN), .ZN(n4527) );
  OR2_X1 U35430 ( .A1(n2752), .A2(IR_REG_27__SCAN_IN), .ZN(n2753) );
  NAND2_X1 U35440 ( .A1(n2753), .A2(IR_REG_31__SCAN_IN), .ZN(n2755) );
  XNOR2_X1 U35450 ( .A(n2755), .B(n2754), .ZN(n4505) );
  NAND2_X1 U35460 ( .A1(n2988), .A2(n4505), .ZN(n4424) );
  AOI21_X1 U35470 ( .B1(B_REG_SCAN_IN), .B2(n4527), .A(n4424), .ZN(n4139) );
  INV_X1 U35480 ( .A(REG2_REG_30__SCAN_IN), .ZN(n2758) );
  NAND2_X1 U35490 ( .A1(n3864), .A2(REG1_REG_30__SCAN_IN), .ZN(n2757) );
  NAND2_X1 U35500 ( .A1(n2547), .A2(REG0_REG_30__SCAN_IN), .ZN(n2756) );
  OAI211_X1 U35510 ( .C1(n2759), .C2(n2758), .A(n2757), .B(n2756), .ZN(n4029)
         );
  AOI22_X1 U35520 ( .A1(n2760), .A2(n4366), .B1(n4139), .B2(n4029), .ZN(n4149)
         );
  INV_X1 U35530 ( .A(n4505), .ZN(n2895) );
  AND2_X2 U35540 ( .A1(n2988), .A2(n2895), .ZN(n4420) );
  INV_X1 U35550 ( .A(n3886), .ZN(n4148) );
  AOI22_X1 U35560 ( .A1(n4030), .A2(n4420), .B1(n4148), .B2(n4430), .ZN(n2761)
         );
  NOR2_X1 U35570 ( .A1(n2763), .A2(n2765), .ZN(n2764) );
  MUX2_X1 U35580 ( .A(n2765), .B(n2764), .S(IR_REG_25__SCAN_IN), .Z(n2768) );
  INV_X1 U35590 ( .A(n2766), .ZN(n2767) );
  NAND2_X1 U35600 ( .A1(n2973), .A2(B_REG_SCAN_IN), .ZN(n2774) );
  NAND2_X1 U35610 ( .A1(n2770), .A2(n2769), .ZN(n2771) );
  INV_X1 U35620 ( .A(IR_REG_23__SCAN_IN), .ZN(n2780) );
  NAND2_X1 U35630 ( .A1(n2779), .A2(n2780), .ZN(n2772) );
  MUX2_X1 U35640 ( .A(n2774), .B(B_REG_SCAN_IN), .S(n2778), .Z(n2776) );
  NAND2_X1 U35650 ( .A1(n2766), .A2(IR_REG_31__SCAN_IN), .ZN(n2775) );
  OR2_X1 U35660 ( .A1(n2980), .A2(D_REG_1__SCAN_IN), .ZN(n2874) );
  NAND2_X1 U35670 ( .A1(n2796), .A2(n2973), .ZN(n2981) );
  NAND2_X1 U35680 ( .A1(n2874), .A2(n2981), .ZN(n2795) );
  XNOR2_X1 U35690 ( .A(n2779), .B(n2780), .ZN(n2987) );
  NAND2_X1 U35700 ( .A1(n4700), .A2(n2781), .ZN(n2893) );
  NAND2_X1 U35710 ( .A1(n4016), .A2(n4133), .ZN(n2876) );
  NAND2_X1 U35720 ( .A1(n2988), .A2(n2876), .ZN(n3161) );
  NAND2_X1 U35730 ( .A1(n2893), .A2(n3161), .ZN(n2782) );
  NOR2_X1 U35740 ( .A1(n3159), .A2(n2782), .ZN(n2794) );
  NOR2_X1 U35750 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_19__SCAN_IN), .ZN(n2786)
         );
  NOR4_X1 U35760 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2785) );
  NOR4_X1 U35770 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2784) );
  NOR4_X1 U35780 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2783) );
  NAND4_X1 U35790 ( .A1(n2786), .A2(n2785), .A3(n2784), .A4(n2783), .ZN(n2792)
         );
  NOR4_X1 U35800 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2790) );
  NOR4_X1 U35810 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_27__SCAN_IN), .ZN(n2789) );
  NOR4_X1 U3582 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2788) );
  NOR4_X1 U3583 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2787) );
  NAND4_X1 U3584 ( .A1(n2790), .A2(n2789), .A3(n2788), .A4(n2787), .ZN(n2791)
         );
  NOR2_X1 U3585 ( .A1(n2792), .A2(n2791), .ZN(n2793) );
  INV_X1 U3586 ( .A(n2778), .ZN(n2797) );
  NAND2_X1 U3587 ( .A1(n2797), .A2(n2796), .ZN(n2983) );
  NAND2_X1 U3588 ( .A1(n2819), .A2(n4703), .ZN(n2802) );
  NAND2_X1 U3589 ( .A1(n3139), .A2(n3122), .ZN(n3144) );
  OR2_X1 U3590 ( .A1(n4151), .A2(n4492), .ZN(n2800) );
  NAND2_X1 U3591 ( .A1(n4701), .A2(REG0_REG_29__SCAN_IN), .ZN(n2799) );
  NAND2_X1 U3592 ( .A1(n2802), .A2(n2801), .ZN(U3515) );
  XNOR2_X1 U3593 ( .A(n2803), .B(n3943), .ZN(n4169) );
  XNOR2_X1 U3594 ( .A(n2804), .B(n3943), .ZN(n2805) );
  NAND2_X1 U3595 ( .A1(n2805), .A2(n4366), .ZN(n4164) );
  INV_X1 U3596 ( .A(n4158), .ZN(n3732) );
  OAI22_X1 U3597 ( .A1(n3732), .A2(n4424), .B1(n4334), .B2(n4163), .ZN(n2806)
         );
  AOI21_X1 U3598 ( .B1(n4420), .B2(n4159), .A(n2806), .ZN(n2807) );
  OAI21_X1 U3599 ( .B1(n4169), .B2(n4690), .A(n2808), .ZN(n2815) );
  AND2_X2 U3600 ( .A1(n2809), .A2(n2875), .ZN(n4710) );
  INV_X1 U3601 ( .A(n2810), .ZN(n2814) );
  INV_X1 U3602 ( .A(n2811), .ZN(n2812) );
  OAI21_X1 U3603 ( .B1(n4175), .B2(n4163), .A(n2812), .ZN(n4157) );
  NAND2_X2 U3604 ( .A1(n4710), .A2(n4357), .ZN(n4446) );
  NAND2_X1 U3605 ( .A1(n2814), .A2(n2813), .ZN(U3546) );
  INV_X1 U3606 ( .A(n2816), .ZN(n2818) );
  NAND2_X1 U3607 ( .A1(n2818), .A2(n2817), .ZN(U3514) );
  NAND2_X1 U3608 ( .A1(n2819), .A2(n4710), .ZN(n2823) );
  OR2_X1 U3609 ( .A1(n4710), .A2(n2696), .ZN(n2820) );
  NAND2_X1 U3610 ( .A1(n2823), .A2(n2822), .ZN(U3547) );
  INV_X1 U3611 ( .A(n4664), .ZN(n2824) );
  INV_X2 U3612 ( .A(n4031), .ZN(U4043) );
  INV_X2 U3613 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U3614 ( .A1(n2825), .A2(n2844), .ZN(n2827) );
  NAND2_X1 U3615 ( .A1(n3708), .A2(n2454), .ZN(n2826) );
  NAND2_X1 U3616 ( .A1(n2827), .A2(n2826), .ZN(n2830) );
  INV_X1 U3617 ( .A(n2885), .ZN(n2829) );
  XNOR2_X1 U3618 ( .A(n2830), .B(n3711), .ZN(n2909) );
  NOR2_X1 U3619 ( .A1(n2843), .A2(n3149), .ZN(n2831) );
  NAND2_X1 U3620 ( .A1(n3708), .A2(n3257), .ZN(n2834) );
  NAND2_X1 U3621 ( .A1(n2835), .A2(n2834), .ZN(n2836) );
  NOR2_X1 U3622 ( .A1(n2843), .A2(n3122), .ZN(n2837) );
  XNOR2_X1 U3623 ( .A(n2839), .B(n2840), .ZN(n3088) );
  INV_X1 U3624 ( .A(n3088), .ZN(n2842) );
  INV_X1 U3625 ( .A(n2839), .ZN(n2841) );
  NAND2_X1 U3626 ( .A1(n2841), .A2(n2840), .ZN(n2870) );
  NAND2_X1 U3627 ( .A1(n2419), .A2(n2844), .ZN(n2846) );
  NAND2_X1 U3628 ( .A1(n3708), .A2(n3231), .ZN(n2845) );
  NAND2_X1 U3629 ( .A1(n2846), .A2(n2845), .ZN(n2847) );
  NOR2_X1 U3630 ( .A1(n2843), .A2(n3237), .ZN(n2848) );
  XNOR2_X1 U3631 ( .A(n2860), .B(n2858), .ZN(n3048) );
  INV_X1 U3632 ( .A(n2833), .ZN(n2884) );
  AOI22_X1 U3633 ( .A1(n2844), .A2(n3230), .B1(n2884), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2851) );
  INV_X1 U3634 ( .A(n2714), .ZN(n2849) );
  NAND2_X1 U3635 ( .A1(n2851), .A2(n2850), .ZN(n3040) );
  NAND2_X1 U3636 ( .A1(n2714), .A2(n2844), .ZN(n2854) );
  NAND2_X1 U3637 ( .A1(n3708), .A2(n3230), .ZN(n2855) );
  INV_X1 U3638 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2852) );
  AND2_X1 U3639 ( .A1(n2855), .A2(n2236), .ZN(n2853) );
  NAND2_X1 U3640 ( .A1(n2854), .A2(n2853), .ZN(n3041) );
  INV_X1 U3641 ( .A(n2855), .ZN(n2856) );
  NAND2_X1 U3642 ( .A1(n3039), .A2(n2857), .ZN(n3047) );
  NAND2_X1 U3643 ( .A1(n3048), .A2(n3047), .ZN(n3046) );
  INV_X1 U3644 ( .A(n2858), .ZN(n2859) );
  NAND2_X1 U3645 ( .A1(n2860), .A2(n2859), .ZN(n2861) );
  NAND2_X1 U3646 ( .A1(n3046), .A2(n2861), .ZN(n3053) );
  INV_X1 U3647 ( .A(n3053), .ZN(n2867) );
  NAND2_X1 U3648 ( .A1(n2433), .A2(n2844), .ZN(n2863) );
  NAND2_X1 U3649 ( .A1(n3708), .A2(n2431), .ZN(n2862) );
  NAND2_X1 U3650 ( .A1(n2863), .A2(n2862), .ZN(n2864) );
  XNOR2_X1 U3651 ( .A(n2864), .B(n3711), .ZN(n2869) );
  NOR2_X1 U3652 ( .A1(n2843), .A2(n3131), .ZN(n2865) );
  AOI21_X1 U3653 ( .B1(n3714), .B2(n2433), .A(n2865), .ZN(n2868) );
  XNOR2_X1 U3654 ( .A(n2869), .B(n2868), .ZN(n3054) );
  NAND2_X1 U3655 ( .A1(n2867), .A2(n2866), .ZN(n2908) );
  NAND2_X1 U3656 ( .A1(n2869), .A2(n2868), .ZN(n3089) );
  INV_X1 U3657 ( .A(n2906), .ZN(n2871) );
  NAND2_X1 U3658 ( .A1(n2908), .A2(n2871), .ZN(n2872) );
  AND2_X1 U3659 ( .A1(n2915), .A2(n2872), .ZN(n2880) );
  NAND3_X1 U3660 ( .A1(n3162), .A2(n2875), .A3(n2874), .ZN(n2897) );
  INV_X1 U3661 ( .A(n2988), .ZN(n2878) );
  NAND2_X1 U3662 ( .A1(n3221), .A2(n2876), .ZN(n2877) );
  NAND2_X1 U3663 ( .A1(n2878), .A2(n2877), .ZN(n2881) );
  OR2_X1 U3664 ( .A1(n3159), .A2(n2881), .ZN(n2879) );
  AOI211_X1 U3665 ( .C1(n2914), .C2(n2880), .A(n3861), .B(n2369), .ZN(n2901)
         );
  NAND2_X1 U3666 ( .A1(n4334), .A2(n2881), .ZN(n2882) );
  NAND2_X1 U3667 ( .A1(n2897), .A2(n2882), .ZN(n2883) );
  NAND2_X1 U3668 ( .A1(n2883), .A2(n3161), .ZN(n3035) );
  OAI21_X1 U3669 ( .B1(n3035), .B2(n2884), .A(STATE_REG_SCAN_IN), .ZN(n2888)
         );
  NAND2_X1 U3670 ( .A1(n4664), .A2(n2885), .ZN(n2886) );
  NOR2_X1 U3671 ( .A1(n3727), .A2(n2886), .ZN(n4024) );
  NAND2_X1 U3672 ( .A1(n2897), .A2(n4024), .ZN(n3036) );
  OR2_X1 U3673 ( .A1(n2987), .A2(U3149), .ZN(n4027) );
  AND2_X1 U3674 ( .A1(n3036), .A2(n4027), .ZN(n2887) );
  INV_X1 U3675 ( .A(n3158), .ZN(n2889) );
  NOR2_X1 U3676 ( .A1(n4522), .A2(n2889), .ZN(n2900) );
  NAND2_X1 U3677 ( .A1(n4024), .A2(n4505), .ZN(n2890) );
  INV_X1 U3678 ( .A(n4044), .ZN(n2891) );
  NAND2_X1 U3679 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3099) );
  OAI21_X1 U3680 ( .B1(n3844), .B2(n2891), .A(n3099), .ZN(n2899) );
  OR2_X1 U3681 ( .A1(n3159), .A2(n4334), .ZN(n2892) );
  OR2_X1 U3682 ( .A1(n2897), .A2(n2892), .ZN(n2894) );
  INV_X1 U3683 ( .A(n2838), .ZN(n3135) );
  NAND2_X1 U3684 ( .A1(n4024), .A2(n2895), .ZN(n2896) );
  OAI22_X1 U3685 ( .A1(n4509), .A2(n3149), .B1(n3135), .B2(n4506), .ZN(n2898)
         );
  OR4_X1 U3686 ( .A1(n2901), .A2(n2900), .A3(n2899), .A4(n2898), .ZN(U3227) );
  NAND2_X1 U3687 ( .A1(n4039), .A2(n2844), .ZN(n2903) );
  NAND2_X1 U3688 ( .A1(n3708), .A2(n3451), .ZN(n2902) );
  NAND2_X1 U3689 ( .A1(n2903), .A2(n2902), .ZN(n2904) );
  XNOR2_X1 U3690 ( .A(n2904), .B(n3711), .ZN(n3415) );
  NOR2_X1 U3691 ( .A1(n3727), .A2(n3447), .ZN(n2905) );
  AOI21_X1 U3692 ( .B1(n3714), .B2(n4039), .A(n2905), .ZN(n3416) );
  XNOR2_X1 U3693 ( .A(n3415), .B(n3416), .ZN(n2963) );
  NOR2_X1 U3694 ( .A1(n2906), .A2(n2914), .ZN(n2907) );
  NAND2_X1 U3695 ( .A1(n2908), .A2(n2907), .ZN(n2918) );
  INV_X1 U3696 ( .A(n2909), .ZN(n2912) );
  INV_X1 U3697 ( .A(n2910), .ZN(n2911) );
  NAND2_X1 U3698 ( .A1(n2912), .A2(n2911), .ZN(n2913) );
  OAI21_X1 U3699 ( .B1(n2915), .B2(n2914), .A(n2913), .ZN(n2916) );
  INV_X1 U3700 ( .A(n2916), .ZN(n2917) );
  NAND2_X1 U3701 ( .A1(n2918), .A2(n2917), .ZN(n3108) );
  NAND2_X1 U3702 ( .A1(n4044), .A2(n2844), .ZN(n2920) );
  NAND2_X1 U3703 ( .A1(n3708), .A2(n3246), .ZN(n2919) );
  NAND2_X1 U3704 ( .A1(n2920), .A2(n2919), .ZN(n2921) );
  XNOR2_X1 U3705 ( .A(n2921), .B(n3725), .ZN(n2925) );
  NOR2_X1 U3706 ( .A1(n3727), .A2(n2256), .ZN(n2922) );
  AOI21_X1 U3707 ( .B1(n3714), .B2(n4044), .A(n2922), .ZN(n2923) );
  XNOR2_X1 U3708 ( .A(n2925), .B(n2923), .ZN(n3110) );
  NAND2_X1 U3709 ( .A1(n3108), .A2(n3110), .ZN(n3109) );
  INV_X1 U3710 ( .A(n2923), .ZN(n2924) );
  NAND2_X1 U3711 ( .A1(n2925), .A2(n2924), .ZN(n2926) );
  NAND2_X1 U3712 ( .A1(n3714), .A2(n4043), .ZN(n2928) );
  NAND2_X1 U3713 ( .A1(n2844), .A2(n3355), .ZN(n2927) );
  NAND2_X1 U3714 ( .A1(n2928), .A2(n2927), .ZN(n3182) );
  NAND2_X1 U3715 ( .A1(n4043), .A2(n2844), .ZN(n2930) );
  NAND2_X1 U3716 ( .A1(n3708), .A2(n3355), .ZN(n2929) );
  NAND2_X1 U3717 ( .A1(n2930), .A2(n2929), .ZN(n2931) );
  XNOR2_X1 U3718 ( .A(n2931), .B(n3725), .ZN(n3181) );
  OAI21_X1 U3719 ( .B1(n3184), .B2(n3182), .A(n3181), .ZN(n2933) );
  NAND2_X1 U3720 ( .A1(n3184), .A2(n3182), .ZN(n2932) );
  NAND2_X1 U3721 ( .A1(n2933), .A2(n2932), .ZN(n3210) );
  NAND2_X1 U3722 ( .A1(n4042), .A2(n2844), .ZN(n2935) );
  NAND2_X1 U3723 ( .A1(n3708), .A2(n3195), .ZN(n2934) );
  NAND2_X1 U3724 ( .A1(n2935), .A2(n2934), .ZN(n2936) );
  XNOR2_X1 U3725 ( .A(n2936), .B(n3725), .ZN(n2940) );
  NOR2_X1 U3726 ( .A1(n3727), .A2(n3215), .ZN(n2937) );
  AOI21_X1 U3727 ( .B1(n3714), .B2(n4042), .A(n2937), .ZN(n2938) );
  XNOR2_X1 U3728 ( .A(n2940), .B(n2938), .ZN(n3211) );
  NAND2_X1 U3729 ( .A1(n3210), .A2(n3211), .ZN(n2942) );
  INV_X1 U3730 ( .A(n2938), .ZN(n2939) );
  NAND2_X1 U3731 ( .A1(n2940), .A2(n2939), .ZN(n2941) );
  NAND2_X1 U3732 ( .A1(n2942), .A2(n2941), .ZN(n3280) );
  NAND2_X1 U3733 ( .A1(n4041), .A2(n2844), .ZN(n2944) );
  NAND2_X1 U3734 ( .A1(n3708), .A2(n3308), .ZN(n2943) );
  NAND2_X1 U3735 ( .A1(n2944), .A2(n2943), .ZN(n2945) );
  XNOR2_X1 U3736 ( .A(n2945), .B(n3725), .ZN(n2948) );
  NAND2_X1 U3737 ( .A1(n3714), .A2(n4041), .ZN(n2947) );
  NAND2_X1 U3738 ( .A1(n2844), .A2(n3308), .ZN(n2946) );
  NAND2_X1 U3739 ( .A1(n2947), .A2(n2946), .ZN(n2949) );
  INV_X1 U3740 ( .A(n2948), .ZN(n2951) );
  INV_X1 U3741 ( .A(n2949), .ZN(n2950) );
  NAND2_X1 U3742 ( .A1(n2951), .A2(n2950), .ZN(n3277) );
  NAND2_X1 U3743 ( .A1(n4040), .A2(n2844), .ZN(n2953) );
  NAND2_X1 U3744 ( .A1(n3708), .A2(n3292), .ZN(n2952) );
  NAND2_X1 U3745 ( .A1(n2953), .A2(n2952), .ZN(n2954) );
  XNOR2_X1 U3746 ( .A(n2954), .B(n3725), .ZN(n2956) );
  NOR2_X1 U3747 ( .A1(n3727), .A2(n3328), .ZN(n2955) );
  AOI21_X1 U3748 ( .B1(n3714), .B2(n4040), .A(n2955), .ZN(n2957) );
  XNOR2_X1 U3749 ( .A(n2956), .B(n2957), .ZN(n3324) );
  INV_X1 U3750 ( .A(n2956), .ZN(n2958) );
  NAND2_X1 U3751 ( .A1(n2958), .A2(n2957), .ZN(n2959) );
  INV_X1 U3752 ( .A(n3420), .ZN(n2961) );
  AOI211_X1 U3753 ( .C1(n2963), .C2(n2962), .A(n3861), .B(n2961), .ZN(n2968)
         );
  NOR2_X1 U3754 ( .A1(n4522), .A2(n2964), .ZN(n2967) );
  INV_X1 U3755 ( .A(n4040), .ZN(n3311) );
  NAND2_X1 U3756 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4557) );
  OAI21_X1 U3757 ( .B1(n4506), .B2(n3311), .A(n4557), .ZN(n2966) );
  INV_X1 U3758 ( .A(n4038), .ZN(n3453) );
  OAI22_X1 U3759 ( .A1(n4509), .A2(n3447), .B1(n3453), .B2(n3844), .ZN(n2965)
         );
  OR4_X1 U3760 ( .A1(n2968), .A2(n2967), .A3(n2966), .A4(n2965), .ZN(U3214) );
  MUX2_X1 U3761 ( .A(n2990), .B(n2410), .S(U3149), .Z(n2969) );
  INV_X1 U3762 ( .A(n2969), .ZN(U3351) );
  MUX2_X1 U3763 ( .A(n2970), .B(n3103), .S(STATE_REG_SCAN_IN), .Z(n2971) );
  INV_X1 U3764 ( .A(n2971), .ZN(U3348) );
  MUX2_X1 U3765 ( .A(n2487), .B(n4093), .S(STATE_REG_SCAN_IN), .Z(n2972) );
  INV_X1 U3766 ( .A(n2972), .ZN(U3345) );
  INV_X1 U3767 ( .A(DATAI_25_), .ZN(n4819) );
  INV_X1 U3768 ( .A(n2973), .ZN(n2974) );
  NAND2_X1 U3769 ( .A1(n2974), .A2(STATE_REG_SCAN_IN), .ZN(n2975) );
  OAI21_X1 U3770 ( .B1(STATE_REG_SCAN_IN), .B2(n4819), .A(n2975), .ZN(U3327)
         );
  INV_X1 U3771 ( .A(DATAI_29_), .ZN(n4852) );
  NAND2_X1 U3772 ( .A1(n2976), .A2(STATE_REG_SCAN_IN), .ZN(n2977) );
  OAI21_X1 U3773 ( .B1(STATE_REG_SCAN_IN), .B2(n4852), .A(n2977), .ZN(U3323)
         );
  NAND2_X1 U3774 ( .A1(n4527), .A2(STATE_REG_SCAN_IN), .ZN(n2978) );
  OAI21_X1 U3775 ( .B1(STATE_REG_SCAN_IN), .B2(n2680), .A(n2978), .ZN(U3325)
         );
  INV_X1 U3776 ( .A(DATAI_21_), .ZN(n4972) );
  NAND2_X1 U3777 ( .A1(n3948), .A2(STATE_REG_SCAN_IN), .ZN(n2979) );
  OAI21_X1 U3778 ( .B1(STATE_REG_SCAN_IN), .B2(n4972), .A(n2979), .ZN(U3331)
         );
  INV_X1 U3779 ( .A(n3159), .ZN(n3037) );
  INV_X1 U3780 ( .A(D_REG_1__SCAN_IN), .ZN(n5063) );
  INV_X1 U3781 ( .A(n2981), .ZN(n2982) );
  AOI22_X1 U3782 ( .A1(n4662), .A2(n5063), .B1(n2982), .B2(n4664), .ZN(U3459)
         );
  INV_X1 U3783 ( .A(D_REG_0__SCAN_IN), .ZN(n2985) );
  INV_X1 U3784 ( .A(n2983), .ZN(n2984) );
  AOI22_X1 U3785 ( .A1(n4662), .A2(n2985), .B1(n2984), .B2(n4664), .ZN(U3458)
         );
  NAND2_X1 U3786 ( .A1(n3159), .A2(n4027), .ZN(n2999) );
  AOI21_X1 U3787 ( .B1(n2988), .B2(n2987), .A(n2986), .ZN(n2998) );
  INV_X1 U3788 ( .A(n2998), .ZN(n2989) );
  NOR2_X1 U3789 ( .A1(n4630), .A2(U4043), .ZN(U3148) );
  NOR2_X1 U3790 ( .A1(n2990), .A2(n2991), .ZN(n3070) );
  MUX2_X1 U3791 ( .A(n2992), .B(REG2_REG_2__SCAN_IN), .S(n3066), .Z(n3071) );
  OAI21_X1 U3792 ( .B1(n4051), .B2(n3070), .A(n3071), .ZN(n3073) );
  INV_X1 U3793 ( .A(n2994), .ZN(n2995) );
  MUX2_X1 U3794 ( .A(n2461), .B(REG2_REG_5__SCAN_IN), .S(n4502), .Z(n3028) );
  NOR2_X1 U3795 ( .A1(n3029), .A2(n3028), .ZN(n3027) );
  AOI21_X1 U3796 ( .B1(REG2_REG_5__SCAN_IN), .B2(n4502), .A(n3027), .ZN(n2996)
         );
  XNOR2_X1 U3797 ( .A(n2996), .B(n4501), .ZN(n3016) );
  INV_X1 U3798 ( .A(n2996), .ZN(n2997) );
  AOI22_X1 U3799 ( .A1(n3016), .A2(REG2_REG_6__SCAN_IN), .B1(n4501), .B2(n2997), .ZN(n3001) );
  MUX2_X1 U3800 ( .A(REG2_REG_7__SCAN_IN), .B(n4092), .S(n4093), .Z(n3000) );
  INV_X1 U3801 ( .A(n4527), .ZN(n3009) );
  NOR2_X1 U3802 ( .A1(n4505), .A2(n3009), .ZN(n4023) );
  AOI211_X1 U3803 ( .C1(n3001), .C2(n3000), .A(n4624), .B(n4095), .ZN(n3015)
         );
  AND2_X1 U3804 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4047)
         );
  INV_X1 U3805 ( .A(n2990), .ZN(n4045) );
  NAND2_X1 U3806 ( .A1(n4045), .A2(REG1_REG_1__SCAN_IN), .ZN(n3002) );
  NAND2_X1 U3807 ( .A1(n4046), .A2(n3002), .ZN(n3068) );
  XNOR2_X1 U3808 ( .A(n3066), .B(REG1_REG_2__SCAN_IN), .ZN(n3069) );
  NAND2_X1 U3809 ( .A1(n3068), .A2(n3069), .ZN(n3067) );
  INV_X1 U3810 ( .A(n3066), .ZN(n4504) );
  NAND2_X1 U3811 ( .A1(n4504), .A2(REG1_REG_2__SCAN_IN), .ZN(n3003) );
  NAND2_X1 U3812 ( .A1(n3067), .A2(n3003), .ZN(n3005) );
  INV_X1 U3813 ( .A(n4503), .ZN(n3004) );
  XNOR2_X1 U3814 ( .A(n3005), .B(n3004), .ZN(n4061) );
  NAND2_X1 U3815 ( .A1(n4061), .A2(REG1_REG_3__SCAN_IN), .ZN(n4060) );
  NAND2_X1 U3816 ( .A1(n3005), .A2(n4503), .ZN(n3006) );
  NAND2_X1 U3817 ( .A1(n4060), .A2(n3006), .ZN(n3008) );
  XNOR2_X1 U3818 ( .A(n3008), .B(n3103), .ZN(n3098) );
  NAND2_X1 U3819 ( .A1(n3098), .A2(REG1_REG_4__SCAN_IN), .ZN(n3097) );
  INV_X1 U3820 ( .A(n3097), .ZN(n3007) );
  AOI21_X1 U3821 ( .B1(n2310), .B2(n3008), .A(n3007), .ZN(n3026) );
  XNOR2_X1 U3822 ( .A(n4502), .B(REG1_REG_5__SCAN_IN), .ZN(n3025) );
  NOR2_X1 U3823 ( .A1(n3026), .A2(n3025), .ZN(n3024) );
  INV_X1 U3824 ( .A(n4501), .ZN(n3018) );
  INV_X1 U3825 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3368) );
  INV_X1 U3826 ( .A(n4069), .ZN(n4071) );
  XOR2_X1 U3827 ( .A(REG1_REG_7__SCAN_IN), .B(n4093), .Z(n3011) );
  OAI21_X1 U3828 ( .B1(n4071), .B2(n3011), .A(n4631), .ZN(n3010) );
  AOI21_X1 U3829 ( .B1(n4071), .B2(n3011), .A(n3010), .ZN(n3014) );
  NAND2_X1 U3830 ( .A1(n4529), .A2(n4505), .ZN(n4637) );
  INV_X1 U3831 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4985) );
  NOR2_X1 U3832 ( .A1(STATE_REG_SCAN_IN), .A2(n4985), .ZN(n3212) );
  AOI21_X1 U3833 ( .B1(n4630), .B2(ADDR_REG_7__SCAN_IN), .A(n3212), .ZN(n3012)
         );
  OAI21_X1 U3834 ( .B1(n4637), .B2(n4093), .A(n3012), .ZN(n3013) );
  OR3_X1 U3835 ( .A1(n3015), .A2(n3014), .A3(n3013), .ZN(U3247) );
  XNOR2_X1 U3836 ( .A(n3016), .B(REG2_REG_6__SCAN_IN), .ZN(n3023) );
  NOR2_X1 U3837 ( .A1(STATE_REG_SCAN_IN), .A2(n3017), .ZN(n3185) );
  NOR2_X1 U3838 ( .A1(n4637), .A2(n3018), .ZN(n3019) );
  AOI211_X1 U3839 ( .C1(n4630), .C2(ADDR_REG_6__SCAN_IN), .A(n3185), .B(n3019), 
        .ZN(n3022) );
  OAI211_X1 U3840 ( .C1(REG1_REG_6__SCAN_IN), .C2(n2248), .A(n3020), .B(n4631), 
        .ZN(n3021) );
  OAI211_X1 U3841 ( .C1(n3023), .C2(n4624), .A(n3022), .B(n3021), .ZN(U3246)
         );
  INV_X1 U3842 ( .A(n4631), .ZN(n4138) );
  AOI211_X1 U3843 ( .C1(n3026), .C2(n3025), .A(n3024), .B(n4138), .ZN(n3034)
         );
  AOI211_X1 U3844 ( .C1(n3029), .C2(n3028), .A(n3027), .B(n4624), .ZN(n3033)
         );
  INV_X1 U3845 ( .A(n4502), .ZN(n3031) );
  NOR2_X1 U3846 ( .A1(STATE_REG_SCAN_IN), .A2(n2458), .ZN(n3111) );
  AOI21_X1 U3847 ( .B1(n4630), .B2(ADDR_REG_5__SCAN_IN), .A(n3111), .ZN(n3030)
         );
  OAI21_X1 U3848 ( .B1(n4637), .B2(n3031), .A(n3030), .ZN(n3032) );
  OR3_X1 U3849 ( .A1(n3034), .A2(n3033), .A3(n3032), .ZN(U3245) );
  INV_X1 U3850 ( .A(n3035), .ZN(n3038) );
  NAND3_X1 U3851 ( .A1(n3038), .A2(n3037), .A3(n3036), .ZN(n3057) );
  INV_X1 U3852 ( .A(n3057), .ZN(n3051) );
  INV_X1 U3853 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3044) );
  INV_X1 U3854 ( .A(n4509), .ZN(n3799) );
  OAI21_X1 U3855 ( .B1(n3041), .B2(n3040), .A(n3039), .ZN(n3062) );
  OAI22_X1 U3856 ( .A1(n3062), .A2(n3861), .B1(n3844), .B2(n2413), .ZN(n3042)
         );
  AOI21_X1 U3857 ( .B1(n3230), .B2(n3799), .A(n3042), .ZN(n3043) );
  OAI21_X1 U3858 ( .B1(n3051), .B2(n3044), .A(n3043), .ZN(U3229) );
  INV_X1 U3859 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3234) );
  OAI22_X1 U3860 ( .A1(n2849), .A2(n4506), .B1(n3844), .B2(n2432), .ZN(n3045)
         );
  AOI21_X1 U3861 ( .B1(n3231), .B2(n3799), .A(n3045), .ZN(n3050) );
  OAI211_X1 U3862 ( .C1(n3048), .C2(n3047), .A(n3046), .B(n4517), .ZN(n3049)
         );
  OAI211_X1 U3863 ( .C1(n3051), .C2(n3234), .A(n3050), .B(n3049), .ZN(U3219)
         );
  INV_X1 U3864 ( .A(n2908), .ZN(n3052) );
  AOI21_X1 U3865 ( .B1(n3054), .B2(n3053), .A(n3052), .ZN(n3059) );
  AOI22_X1 U3866 ( .A1(n4512), .A2(n2838), .B1(n3853), .B2(n2419), .ZN(n3055)
         );
  OAI21_X1 U3867 ( .B1(n4509), .B2(n3131), .A(n3055), .ZN(n3056) );
  AOI21_X1 U3868 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3057), .A(n3056), .ZN(n3058)
         );
  OAI21_X1 U3869 ( .B1(n3059), .B2(n3861), .A(n3058), .ZN(U3234) );
  AND2_X1 U3870 ( .A1(n4527), .A2(n3060), .ZN(n3061) );
  OR2_X1 U3871 ( .A1(n4505), .A2(n3061), .ZN(n4528) );
  NAND2_X1 U3872 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4049) );
  NOR2_X1 U3873 ( .A1(n3062), .A2(n4527), .ZN(n3063) );
  AOI211_X1 U3874 ( .C1(n4527), .C2(n4049), .A(n4505), .B(n3063), .ZN(n3064)
         );
  AOI211_X1 U3875 ( .C1(n2262), .C2(n4528), .A(n4031), .B(n3064), .ZN(n3104)
         );
  AOI22_X1 U3876 ( .A1(n4630), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3065) );
  OAI21_X1 U3877 ( .B1(n4637), .B2(n3066), .A(n3065), .ZN(n3077) );
  OAI211_X1 U3878 ( .C1(n3069), .C2(n3068), .A(n4631), .B(n3067), .ZN(n3075)
         );
  OR3_X1 U3879 ( .A1(n3071), .A2(n4051), .A3(n3070), .ZN(n3072) );
  NAND3_X1 U3880 ( .A1(n4586), .A2(n3073), .A3(n3072), .ZN(n3074) );
  NAND2_X1 U3881 ( .A1(n3075), .A2(n3074), .ZN(n3076) );
  OR3_X1 U3882 ( .A1(n3104), .A2(n3077), .A3(n3076), .ZN(U3242) );
  XNOR2_X1 U3883 ( .A(n4044), .B(n2256), .ZN(n3915) );
  XNOR2_X1 U3884 ( .A(n3078), .B(n3915), .ZN(n3256) );
  INV_X1 U3885 ( .A(n4043), .ZN(n3079) );
  OAI22_X1 U3886 ( .A1(n3079), .A2(n4424), .B1(n4334), .B2(n2256), .ZN(n3082)
         );
  XOR2_X1 U3887 ( .A(n3915), .B(n3080), .Z(n3081) );
  NOR2_X1 U3888 ( .A1(n3081), .A2(n4339), .ZN(n3254) );
  AOI211_X1 U3889 ( .C1(n4420), .C2(n2825), .A(n3082), .B(n3254), .ZN(n3083)
         );
  OAI21_X1 U3890 ( .B1(n4690), .B2(n3256), .A(n3083), .ZN(n3318) );
  INV_X1 U3891 ( .A(n3318), .ZN(n3087) );
  INV_X1 U3892 ( .A(n4492), .ZN(n3085) );
  AND2_X1 U3893 ( .A1(n3145), .A2(n3246), .ZN(n3084) );
  NOR2_X1 U3894 ( .A1(n3176), .A2(n3084), .ZN(n3319) );
  AOI22_X1 U3895 ( .A1(n3085), .A2(n3319), .B1(REG0_REG_5__SCAN_IN), .B2(n4701), .ZN(n3086) );
  OAI21_X1 U3896 ( .B1(n3087), .B2(n4701), .A(n3086), .ZN(U3477) );
  NAND2_X1 U3897 ( .A1(n2908), .A2(n3089), .ZN(n3090) );
  XOR2_X1 U3898 ( .A(n3088), .B(n3090), .Z(n3095) );
  INV_X1 U3899 ( .A(n2825), .ZN(n3252) );
  OAI22_X1 U3900 ( .A1(n2432), .A2(n4506), .B1(n3844), .B2(n3252), .ZN(n3093)
         );
  MUX2_X1 U3901 ( .A(U3149), .B(n3859), .S(n3091), .Z(n3092) );
  AOI211_X1 U3902 ( .C1(n3257), .C2(n3799), .A(n3093), .B(n3092), .ZN(n3094)
         );
  OAI21_X1 U3903 ( .B1(n3861), .B2(n3095), .A(n3094), .ZN(U3215) );
  XOR2_X1 U3904 ( .A(REG2_REG_4__SCAN_IN), .B(n3096), .Z(n3106) );
  OAI211_X1 U3905 ( .C1(REG1_REG_4__SCAN_IN), .C2(n3098), .A(n4631), .B(n3097), 
        .ZN(n3102) );
  INV_X1 U3906 ( .A(n3099), .ZN(n3100) );
  AOI21_X1 U3907 ( .B1(n4630), .B2(ADDR_REG_4__SCAN_IN), .A(n3100), .ZN(n3101)
         );
  OAI211_X1 U3908 ( .C1(n4637), .C2(n3103), .A(n3102), .B(n3101), .ZN(n3105)
         );
  AOI211_X1 U3909 ( .C1(n4586), .C2(n3106), .A(n3105), .B(n3104), .ZN(n3107)
         );
  INV_X1 U3910 ( .A(n3107), .ZN(U3244) );
  OAI211_X1 U3911 ( .C1(n3108), .C2(n3110), .A(n3109), .B(n4517), .ZN(n3116)
         );
  AOI21_X1 U3912 ( .B1(n3853), .B2(n2825), .A(n3111), .ZN(n3113) );
  NAND2_X1 U3913 ( .A1(n4512), .A2(n4043), .ZN(n3112) );
  OAI211_X1 U3914 ( .C1(n4509), .C2(n2256), .A(n3113), .B(n3112), .ZN(n3114)
         );
  AOI21_X1 U3915 ( .B1(n3859), .B2(n3247), .A(n3114), .ZN(n3115) );
  NAND2_X1 U3916 ( .A1(n3116), .A2(n3115), .ZN(U3224) );
  XNOR2_X1 U3917 ( .A(n3117), .B(n3923), .ZN(n3265) );
  OAI22_X1 U3918 ( .A1(n3252), .A2(n4424), .B1(n4334), .B2(n3122), .ZN(n3120)
         );
  XOR2_X1 U3919 ( .A(n3923), .B(n3118), .Z(n3119) );
  NOR2_X1 U3920 ( .A1(n3119), .A2(n4339), .ZN(n3263) );
  AOI211_X1 U3921 ( .C1(n4420), .C2(n2433), .A(n3120), .B(n3263), .ZN(n3121)
         );
  OAI21_X1 U3922 ( .B1(n4690), .B2(n3265), .A(n3121), .ZN(n3349) );
  OR2_X1 U3923 ( .A1(n3139), .A2(n3122), .ZN(n3123) );
  NAND2_X1 U3924 ( .A1(n3144), .A2(n3123), .ZN(n3347) );
  INV_X1 U3925 ( .A(REG0_REG_3__SCAN_IN), .ZN(n3124) );
  OAI22_X1 U3926 ( .A1(n4492), .A2(n3347), .B1(n4703), .B2(n3124), .ZN(n3125)
         );
  AOI21_X1 U3927 ( .B1(n3349), .B2(n4703), .A(n3125), .ZN(n3126) );
  INV_X1 U3928 ( .A(n3126), .ZN(U3473) );
  OAI21_X1 U3929 ( .B1(n3129), .B2(n3128), .A(n3127), .ZN(n4656) );
  INV_X1 U3930 ( .A(n4656), .ZN(n3138) );
  XNOR2_X1 U3931 ( .A(n3130), .B(n3925), .ZN(n3137) );
  INV_X1 U3932 ( .A(n3554), .ZN(n3339) );
  NAND2_X1 U3933 ( .A1(n4656), .A2(n3339), .ZN(n3134) );
  NOR2_X1 U3934 ( .A1(n4334), .A2(n3131), .ZN(n3132) );
  AOI21_X1 U3935 ( .B1(n2419), .B2(n4420), .A(n3132), .ZN(n3133) );
  OAI211_X1 U3936 ( .C1(n3135), .C2(n4424), .A(n3134), .B(n3133), .ZN(n3136)
         );
  AOI21_X1 U3937 ( .B1(n3137), .B2(n4366), .A(n3136), .ZN(n4660) );
  OAI21_X1 U3938 ( .B1(n3138), .B2(n4682), .A(n4660), .ZN(n3353) );
  AND2_X1 U3939 ( .A1(n3232), .A2(n2431), .ZN(n3140) );
  OR2_X1 U3940 ( .A1(n3140), .A2(n3139), .ZN(n4653) );
  INV_X1 U3941 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3141) );
  OAI22_X1 U3942 ( .A1(n4492), .A2(n4653), .B1(n4703), .B2(n3141), .ZN(n3142)
         );
  AOI21_X1 U3943 ( .B1(n3353), .B2(n4703), .A(n3142), .ZN(n3143) );
  INV_X1 U3944 ( .A(n3143), .ZN(U3471) );
  INV_X1 U3945 ( .A(n3144), .ZN(n3146) );
  OAI211_X1 U3946 ( .C1(n3146), .C2(n3149), .A(n4357), .B(n3145), .ZN(n4686)
         );
  NOR2_X1 U3947 ( .A1(n4686), .A2(n4499), .ZN(n3157) );
  XOR2_X1 U3948 ( .A(n3926), .B(n3147), .Z(n3156) );
  NAND2_X1 U3949 ( .A1(n2838), .A2(n4420), .ZN(n3148) );
  OAI21_X1 U3950 ( .B1(n4334), .B2(n3149), .A(n3148), .ZN(n3154) );
  NAND2_X1 U3951 ( .A1(n3151), .A2(n3926), .ZN(n3152) );
  NAND2_X1 U3952 ( .A1(n3150), .A2(n3152), .ZN(n3165) );
  NOR2_X1 U3953 ( .A1(n3165), .A2(n3554), .ZN(n3153) );
  AOI211_X1 U3954 ( .C1(n4432), .C2(n4044), .A(n3154), .B(n3153), .ZN(n3155)
         );
  OAI21_X1 U3955 ( .B1(n4339), .B2(n3156), .A(n3155), .ZN(n4687) );
  AOI211_X1 U3956 ( .C1(n4652), .C2(n3158), .A(n3157), .B(n4687), .ZN(n3169)
         );
  OAI21_X1 U3957 ( .B1(n5063), .B2(n3159), .A(n4662), .ZN(n3160) );
  NAND4_X1 U3958 ( .A1(n3163), .A2(n3162), .A3(n3161), .A4(n3160), .ZN(n3164)
         );
  NAND2_X2 U3959 ( .A1(n3164), .A2(n4368), .ZN(n4349) );
  INV_X2 U3960 ( .A(n4349), .ZN(n4661) );
  INV_X1 U3961 ( .A(n3165), .ZN(n4689) );
  NAND2_X1 U3962 ( .A1(n3166), .A2(n4499), .ZN(n3202) );
  INV_X1 U3963 ( .A(n3202), .ZN(n3167) );
  NAND2_X1 U3964 ( .A1(n4349), .A2(n3167), .ZN(n3565) );
  INV_X1 U3965 ( .A(n3565), .ZN(n4657) );
  AOI22_X1 U3966 ( .A1(n4689), .A2(n4657), .B1(REG2_REG_4__SCAN_IN), .B2(n4661), .ZN(n3168) );
  OAI21_X1 U3967 ( .B1(n3169), .B2(n4661), .A(n3168), .ZN(U3286) );
  INV_X1 U3968 ( .A(n3171), .ZN(n3972) );
  OR2_X1 U3969 ( .A1(n3972), .A2(n3962), .ZN(n3917) );
  XNOR2_X1 U3970 ( .A(n3170), .B(n3917), .ZN(n3367) );
  INV_X1 U3971 ( .A(n4042), .ZN(n3363) );
  OAI22_X1 U3972 ( .A1(n3363), .A2(n4424), .B1(n4334), .B2(n3188), .ZN(n3174)
         );
  XNOR2_X1 U3973 ( .A(n3172), .B(n3917), .ZN(n3173) );
  NOR2_X1 U3974 ( .A1(n3173), .A2(n4339), .ZN(n3365) );
  AOI211_X1 U3975 ( .C1(n4420), .C2(n4044), .A(n3174), .B(n3365), .ZN(n3175)
         );
  OAI21_X1 U3976 ( .B1(n4690), .B2(n3367), .A(n3175), .ZN(n3371) );
  NOR2_X1 U3977 ( .A1(n3176), .A2(n3188), .ZN(n3177) );
  OR2_X1 U3978 ( .A1(n3192), .A2(n3177), .ZN(n3369) );
  INV_X1 U3979 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3178) );
  OAI22_X1 U3980 ( .A1(n3369), .A2(n4492), .B1(n4703), .B2(n3178), .ZN(n3179)
         );
  AOI21_X1 U3981 ( .B1(n3371), .B2(n4703), .A(n3179), .ZN(n3180) );
  INV_X1 U3982 ( .A(n3180), .ZN(U3479) );
  XOR2_X1 U3983 ( .A(n3182), .B(n3181), .Z(n3183) );
  XNOR2_X1 U3984 ( .A(n3184), .B(n3183), .ZN(n3191) );
  AOI21_X1 U3985 ( .B1(n4512), .B2(n4042), .A(n3185), .ZN(n3187) );
  NAND2_X1 U3986 ( .A1(n3853), .A2(n4044), .ZN(n3186) );
  OAI211_X1 U3987 ( .C1(n4509), .C2(n3188), .A(n3187), .B(n3186), .ZN(n3189)
         );
  AOI21_X1 U3988 ( .B1(n3859), .B2(n3356), .A(n3189), .ZN(n3190) );
  OAI21_X1 U3989 ( .B1(n3191), .B2(n3861), .A(n3190), .ZN(U3236) );
  INV_X1 U3990 ( .A(n3192), .ZN(n3194) );
  INV_X1 U3991 ( .A(n4357), .ZN(n4695) );
  INV_X1 U3992 ( .A(n3193), .ZN(n3304) );
  AOI211_X1 U3993 ( .C1(n3195), .C2(n3194), .A(n4695), .B(n3304), .ZN(n4693)
         );
  XNOR2_X1 U3994 ( .A(n3196), .B(n3927), .ZN(n3200) );
  NOR2_X1 U3995 ( .A1(n4334), .A2(n3215), .ZN(n3197) );
  AOI21_X1 U3996 ( .B1(n4041), .B2(n4432), .A(n3197), .ZN(n3199) );
  NAND2_X1 U3997 ( .A1(n4043), .A2(n4420), .ZN(n3198) );
  OAI211_X1 U3998 ( .C1(n3200), .C2(n4339), .A(n3199), .B(n3198), .ZN(n4692)
         );
  AOI21_X1 U3999 ( .B1(n4693), .B2(n4133), .A(n4692), .ZN(n3209) );
  AND2_X1 U4000 ( .A1(n3201), .A2(n3927), .ZN(n4691) );
  NAND2_X1 U4001 ( .A1(n3554), .A2(n3202), .ZN(n3203) );
  NOR2_X1 U4002 ( .A1(n4691), .A2(n4374), .ZN(n3207) );
  INV_X1 U4003 ( .A(n3217), .ZN(n3205) );
  OAI22_X1 U4004 ( .A1(n4349), .A2(n4092), .B1(n3205), .B2(n4368), .ZN(n3206)
         );
  AOI21_X1 U4005 ( .B1(n3207), .B2(n3204), .A(n3206), .ZN(n3208) );
  OAI21_X1 U4006 ( .B1(n3209), .B2(n4661), .A(n3208), .ZN(U3283) );
  XNOR2_X1 U4007 ( .A(n3210), .B(n3211), .ZN(n3219) );
  AOI21_X1 U4008 ( .B1(n4512), .B2(n4041), .A(n3212), .ZN(n3214) );
  NAND2_X1 U4009 ( .A1(n3853), .A2(n4043), .ZN(n3213) );
  OAI211_X1 U4010 ( .C1(n4509), .C2(n3215), .A(n3214), .B(n3213), .ZN(n3216)
         );
  AOI21_X1 U4011 ( .B1(n3859), .B2(n3217), .A(n3216), .ZN(n3218) );
  OAI21_X1 U4012 ( .B1(n3219), .B2(n3861), .A(n3218), .ZN(U3210) );
  NAND2_X1 U4013 ( .A1(n2714), .A2(n3220), .ZN(n3947) );
  AND2_X1 U4014 ( .A1(n3945), .A2(n3947), .ZN(n4679) );
  NAND2_X1 U4015 ( .A1(n3230), .A2(n3221), .ZN(n4677) );
  AOI21_X1 U4016 ( .B1(n4339), .B2(n3554), .A(n4679), .ZN(n3222) );
  AOI21_X1 U4017 ( .B1(n4432), .B2(n2419), .A(n3222), .ZN(n4678) );
  OAI21_X1 U4018 ( .B1(n3223), .B2(n4677), .A(n4678), .ZN(n3224) );
  AOI22_X1 U4019 ( .A1(n3224), .A2(n4349), .B1(REG3_REG_0__SCAN_IN), .B2(n4652), .ZN(n3226) );
  NAND2_X1 U4020 ( .A1(n4661), .A2(REG2_REG_0__SCAN_IN), .ZN(n3225) );
  OAI211_X1 U4021 ( .C1(n4679), .C2(n3565), .A(n3226), .B(n3225), .ZN(U3290)
         );
  OAI21_X1 U4022 ( .B1(n2713), .B2(n3228), .A(n3227), .ZN(n4683) );
  INV_X1 U4023 ( .A(n4683), .ZN(n3244) );
  AND2_X1 U4024 ( .A1(n4357), .A2(n4133), .ZN(n3229) );
  NAND2_X1 U4025 ( .A1(n4349), .A2(n3229), .ZN(n4343) );
  NAND2_X1 U4026 ( .A1(n3231), .A2(n3230), .ZN(n3233) );
  NAND2_X1 U4027 ( .A1(n3233), .A2(n3232), .ZN(n4681) );
  OAI22_X1 U4028 ( .A1(n4343), .A2(n4681), .B1(n3234), .B2(n4368), .ZN(n3243)
         );
  NAND2_X1 U4029 ( .A1(n2714), .A2(n4420), .ZN(n3236) );
  NAND2_X1 U4030 ( .A1(n2433), .A2(n4432), .ZN(n3235) );
  OAI211_X1 U4031 ( .C1(n4334), .C2(n3237), .A(n3236), .B(n3235), .ZN(n3238)
         );
  INV_X1 U4032 ( .A(n3238), .ZN(n3241) );
  XNOR2_X1 U4033 ( .A(n2713), .B(n3945), .ZN(n3239) );
  NAND2_X1 U4034 ( .A1(n3239), .A2(n4366), .ZN(n3240) );
  OAI211_X1 U4035 ( .C1(n4683), .C2(n3554), .A(n3241), .B(n3240), .ZN(n4685)
         );
  MUX2_X1 U4036 ( .A(n4685), .B(REG2_REG_1__SCAN_IN), .S(n4661), .Z(n3242) );
  AOI211_X1 U4037 ( .C1(n3244), .C2(n4657), .A(n3243), .B(n3242), .ZN(n3245)
         );
  INV_X1 U4038 ( .A(n3245), .ZN(U3289) );
  NAND2_X1 U4039 ( .A1(n4349), .A2(n4420), .ZN(n4321) );
  AND2_X1 U4040 ( .A1(n4349), .A2(n4430), .ZN(n4316) );
  AND2_X1 U4041 ( .A1(n4349), .A2(n4432), .ZN(n4315) );
  AOI22_X1 U4042 ( .A1(n4316), .A2(n3246), .B1(n4315), .B2(n4043), .ZN(n3251)
         );
  INV_X1 U40430 ( .A(n3247), .ZN(n3248) );
  OAI22_X1 U4044 ( .A1(n4349), .A2(n2461), .B1(n3248), .B2(n4368), .ZN(n3249)
         );
  AOI21_X1 U4045 ( .B1(n4655), .B2(n3319), .A(n3249), .ZN(n3250) );
  OAI211_X1 U4046 ( .C1(n3252), .C2(n4321), .A(n3251), .B(n3250), .ZN(n3253)
         );
  AOI21_X1 U4047 ( .B1(n3254), .B2(n4349), .A(n3253), .ZN(n3255) );
  OAI21_X1 U4048 ( .B1(n4374), .B2(n3256), .A(n3255), .ZN(U3285) );
  AOI22_X1 U4049 ( .A1(n4316), .A2(n3257), .B1(n4315), .B2(n2825), .ZN(n3261)
         );
  INV_X1 U4050 ( .A(n3347), .ZN(n3259) );
  OAI22_X1 U4051 ( .A1(n4349), .A2(n4062), .B1(REG3_REG_3__SCAN_IN), .B2(n4368), .ZN(n3258) );
  AOI21_X1 U4052 ( .B1(n4655), .B2(n3259), .A(n3258), .ZN(n3260) );
  OAI211_X1 U4053 ( .C1(n2432), .C2(n4321), .A(n3261), .B(n3260), .ZN(n3262)
         );
  AOI21_X1 U4054 ( .B1(n3263), .B2(n4349), .A(n3262), .ZN(n3264) );
  OAI21_X1 U4055 ( .B1(n3265), .B2(n4374), .A(n3264), .ZN(U3287) );
  INV_X1 U4056 ( .A(n3302), .ZN(n3267) );
  INV_X1 U4057 ( .A(n3448), .ZN(n3266) );
  OAI21_X1 U4058 ( .B1(n3267), .B2(n3328), .A(n3266), .ZN(n3291) );
  INV_X1 U4059 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3274) );
  INV_X1 U4060 ( .A(n3973), .ZN(n3269) );
  NAND2_X1 U4061 ( .A1(n3269), .A2(n3969), .ZN(n3918) );
  XOR2_X1 U4062 ( .A(n3268), .B(n3918), .Z(n3290) );
  INV_X1 U4063 ( .A(n4041), .ZN(n3294) );
  INV_X1 U4064 ( .A(n4420), .ZN(n4436) );
  XNOR2_X1 U4065 ( .A(n3270), .B(n3918), .ZN(n3271) );
  NAND2_X1 U4066 ( .A1(n3271), .A2(n4366), .ZN(n3301) );
  AOI22_X1 U4067 ( .A1(n4039), .A2(n4432), .B1(n4430), .B2(n3292), .ZN(n3272)
         );
  OAI211_X1 U4068 ( .C1(n3294), .C2(n4436), .A(n3301), .B(n3272), .ZN(n3273)
         );
  AOI21_X1 U4069 ( .B1(n3290), .B2(n4443), .A(n3273), .ZN(n3287) );
  MUX2_X1 U4070 ( .A(n3274), .B(n3287), .S(n4703), .Z(n3275) );
  OAI21_X1 U4071 ( .B1(n3291), .B2(n4492), .A(n3275), .ZN(U3485) );
  INV_X1 U4072 ( .A(n4645), .ZN(n3286) );
  INV_X1 U4073 ( .A(n3276), .ZN(n3278) );
  NAND2_X1 U4074 ( .A1(n3278), .A2(n3277), .ZN(n3279) );
  XNOR2_X1 U4075 ( .A(n3280), .B(n3279), .ZN(n3281) );
  NAND2_X1 U4076 ( .A1(n3281), .A2(n4517), .ZN(n3285) );
  OAI22_X1 U4077 ( .A1(n4509), .A2(n3303), .B1(n3363), .B2(n4506), .ZN(n3283)
         );
  NAND2_X1 U4078 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4536) );
  OAI21_X1 U4079 ( .B1(n3844), .B2(n3311), .A(n4536), .ZN(n3282) );
  NOR2_X1 U4080 ( .A1(n3283), .A2(n3282), .ZN(n3284) );
  OAI211_X1 U4081 ( .C1(n4522), .C2(n3286), .A(n3285), .B(n3284), .ZN(U3218)
         );
  INV_X1 U4082 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3288) );
  MUX2_X1 U4083 ( .A(n3288), .B(n3287), .S(n4710), .Z(n3289) );
  OAI21_X1 U4084 ( .B1(n4446), .B2(n3291), .A(n3289), .ZN(U3527) );
  NAND2_X1 U4085 ( .A1(n3290), .A2(n4311), .ZN(n3300) );
  INV_X1 U4086 ( .A(n3291), .ZN(n3298) );
  AOI22_X1 U4087 ( .A1(n4316), .A2(n3292), .B1(n4315), .B2(n4039), .ZN(n3293)
         );
  OAI21_X1 U4088 ( .B1(n3294), .B2(n4321), .A(n3293), .ZN(n3297) );
  OAI22_X1 U4089 ( .A1(n3295), .A2(n4368), .B1(n2505), .B2(n4349), .ZN(n3296)
         );
  AOI211_X1 U4090 ( .C1(n3298), .C2(n4655), .A(n3297), .B(n3296), .ZN(n3299)
         );
  OAI211_X1 U4091 ( .C1(n4661), .C2(n3301), .A(n3300), .B(n3299), .ZN(U3281)
         );
  OAI21_X1 U4092 ( .B1(n3304), .B2(n3303), .A(n3302), .ZN(n4646) );
  INV_X1 U4093 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3314) );
  NAND2_X1 U4094 ( .A1(n3968), .A2(n3966), .ZN(n3928) );
  XOR2_X1 U4095 ( .A(n3928), .B(n3305), .Z(n4648) );
  XNOR2_X1 U4096 ( .A(n3306), .B(n3928), .ZN(n3307) );
  NAND2_X1 U4097 ( .A1(n3307), .A2(n4366), .ZN(n3310) );
  AOI22_X1 U4098 ( .A1(n4042), .A2(n4420), .B1(n4430), .B2(n3308), .ZN(n3309)
         );
  OAI211_X1 U4099 ( .C1(n3311), .C2(n4424), .A(n3310), .B(n3309), .ZN(n3312)
         );
  AOI21_X1 U4100 ( .B1(n4648), .B2(n3339), .A(n3312), .ZN(n4651) );
  INV_X1 U4101 ( .A(n4651), .ZN(n3313) );
  AOI21_X1 U4102 ( .B1(n4700), .B2(n4648), .A(n3313), .ZN(n3316) );
  MUX2_X1 U4103 ( .A(n3314), .B(n3316), .S(n4710), .Z(n3315) );
  OAI21_X1 U4104 ( .B1(n4646), .B2(n4446), .A(n3315), .ZN(U3526) );
  INV_X1 U4105 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4996) );
  MUX2_X1 U4106 ( .A(n4996), .B(n3316), .S(n4703), .Z(n3317) );
  OAI21_X1 U4107 ( .B1(n4646), .B2(n4492), .A(n3317), .ZN(U3483) );
  INV_X1 U4108 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3323) );
  NAND2_X1 U4109 ( .A1(n3318), .A2(n4710), .ZN(n3322) );
  INV_X1 U4110 ( .A(n4446), .ZN(n3320) );
  NAND2_X1 U4111 ( .A1(n3320), .A2(n3319), .ZN(n3321) );
  OAI211_X1 U4112 ( .C1(n4710), .C2(n3323), .A(n3322), .B(n3321), .ZN(U3523)
         );
  XOR2_X1 U4113 ( .A(n3325), .B(n3324), .Z(n3332) );
  NOR2_X1 U4114 ( .A1(STATE_REG_SCAN_IN), .A2(n2502), .ZN(n4552) );
  AOI21_X1 U4115 ( .B1(n4512), .B2(n4039), .A(n4552), .ZN(n3327) );
  NAND2_X1 U4116 ( .A1(n3853), .A2(n4041), .ZN(n3326) );
  OAI211_X1 U4117 ( .C1(n4509), .C2(n3328), .A(n3327), .B(n3326), .ZN(n3329)
         );
  AOI21_X1 U4118 ( .B1(n3859), .B2(n3330), .A(n3329), .ZN(n3331) );
  OAI21_X1 U4119 ( .B1(n3332), .B2(n3861), .A(n3331), .ZN(U3228) );
  XOR2_X1 U4120 ( .A(n3931), .B(n3333), .Z(n3341) );
  NAND2_X1 U4121 ( .A1(n3334), .A2(n3931), .ZN(n3335) );
  NAND2_X1 U4122 ( .A1(n3390), .A2(n3335), .ZN(n4699) );
  NAND2_X1 U4123 ( .A1(n4039), .A2(n4420), .ZN(n3337) );
  NAND2_X1 U4124 ( .A1(n4037), .A2(n4432), .ZN(n3336) );
  OAI211_X1 U4125 ( .C1(n4334), .C2(n3430), .A(n3337), .B(n3336), .ZN(n3338)
         );
  AOI21_X1 U4126 ( .B1(n4699), .B2(n3339), .A(n3338), .ZN(n3340) );
  OAI21_X1 U4127 ( .B1(n4339), .B2(n3341), .A(n3340), .ZN(n4697) );
  INV_X1 U4128 ( .A(n4697), .ZN(n3346) );
  OAI21_X1 U4129 ( .B1(n3445), .B2(n3430), .A(n3392), .ZN(n4696) );
  NOR2_X1 U4130 ( .A1(n4696), .A2(n4343), .ZN(n3344) );
  INV_X1 U4131 ( .A(n3432), .ZN(n3342) );
  OAI22_X1 U4132 ( .A1(n4349), .A2(n2526), .B1(n3342), .B2(n4368), .ZN(n3343)
         );
  AOI211_X1 U4133 ( .C1(n4699), .C2(n4657), .A(n3344), .B(n3343), .ZN(n3345)
         );
  OAI21_X1 U4134 ( .B1(n3346), .B2(n4661), .A(n3345), .ZN(U3279) );
  OAI22_X1 U4135 ( .A1(n4446), .A2(n3347), .B1(n4710), .B2(n2349), .ZN(n3348)
         );
  AOI21_X1 U4136 ( .B1(n3349), .B2(n4710), .A(n3348), .ZN(n3350) );
  INV_X1 U4137 ( .A(n3350), .ZN(U3521) );
  INV_X1 U4138 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3351) );
  OAI22_X1 U4139 ( .A1(n4446), .A2(n4653), .B1(n4710), .B2(n3351), .ZN(n3352)
         );
  AOI21_X1 U4140 ( .B1(n3353), .B2(n4710), .A(n3352), .ZN(n3354) );
  INV_X1 U4141 ( .A(n3354), .ZN(U3520) );
  INV_X1 U4142 ( .A(n4315), .ZN(n4177) );
  INV_X1 U4143 ( .A(n4321), .ZN(n4292) );
  AOI22_X1 U4144 ( .A1(n4292), .A2(n4044), .B1(n4316), .B2(n3355), .ZN(n3362)
         );
  INV_X1 U4145 ( .A(n3369), .ZN(n3360) );
  INV_X1 U4146 ( .A(n3356), .ZN(n3357) );
  OAI22_X1 U4147 ( .A1(n4349), .A2(n3358), .B1(n3357), .B2(n4368), .ZN(n3359)
         );
  AOI21_X1 U4148 ( .B1(n3360), .B2(n4655), .A(n3359), .ZN(n3361) );
  OAI211_X1 U4149 ( .C1(n3363), .C2(n4177), .A(n3362), .B(n3361), .ZN(n3364)
         );
  AOI21_X1 U4150 ( .B1(n3365), .B2(n4349), .A(n3364), .ZN(n3366) );
  OAI21_X1 U4151 ( .B1(n4374), .B2(n3367), .A(n3366), .ZN(U3284) );
  OAI22_X1 U4152 ( .A1(n3369), .A2(n4446), .B1(n4710), .B2(n3368), .ZN(n3370)
         );
  AOI21_X1 U4153 ( .B1(n3371), .B2(n4710), .A(n3370), .ZN(n3372) );
  INV_X1 U4154 ( .A(n3372), .ZN(U3524) );
  AND2_X1 U4155 ( .A1(n3374), .A2(n3373), .ZN(n3910) );
  XOR2_X1 U4156 ( .A(n3910), .B(n3543), .Z(n3465) );
  INV_X1 U4157 ( .A(n3465), .ZN(n3386) );
  NAND2_X1 U4158 ( .A1(n3376), .A2(n3375), .ZN(n3400) );
  INV_X1 U4159 ( .A(n3388), .ZN(n3377) );
  OAI21_X1 U4160 ( .B1(n3400), .B2(n3377), .A(n3387), .ZN(n3378) );
  XNOR2_X1 U4161 ( .A(n3378), .B(n3910), .ZN(n3381) );
  INV_X1 U4162 ( .A(n4035), .ZN(n3517) );
  OAI22_X1 U4163 ( .A1(n3517), .A2(n4424), .B1(n4334), .B2(n3510), .ZN(n3379)
         );
  AOI21_X1 U4164 ( .B1(n4420), .B2(n4037), .A(n3379), .ZN(n3380) );
  OAI21_X1 U4165 ( .B1(n3381), .B2(n4339), .A(n3380), .ZN(n3464) );
  NAND2_X1 U4166 ( .A1(n3394), .A2(n3504), .ZN(n3382) );
  NAND2_X1 U4167 ( .A1(n3555), .A2(n3382), .ZN(n3471) );
  AOI22_X1 U4168 ( .A1(n4661), .A2(REG2_REG_13__SCAN_IN), .B1(n3512), .B2(
        n4652), .ZN(n3383) );
  OAI21_X1 U4169 ( .B1(n3471), .B2(n4343), .A(n3383), .ZN(n3384) );
  AOI21_X1 U4170 ( .B1(n3464), .B2(n4349), .A(n3384), .ZN(n3385) );
  OAI21_X1 U4171 ( .B1(n3386), .B2(n4374), .A(n3385), .ZN(U3277) );
  AND2_X1 U4172 ( .A1(n3388), .A2(n3387), .ZN(n3911) );
  NAND2_X1 U4173 ( .A1(n3390), .A2(n3389), .ZN(n3391) );
  XOR2_X1 U4174 ( .A(n3911), .B(n3391), .Z(n3408) );
  NAND2_X1 U4175 ( .A1(n3392), .A2(n3490), .ZN(n3393) );
  NAND2_X1 U4176 ( .A1(n3394), .A2(n3393), .ZN(n3414) );
  INV_X1 U4177 ( .A(n3539), .ZN(n3395) );
  OAI22_X1 U4178 ( .A1(n4349), .A2(n3396), .B1(n3395), .B2(n4368), .ZN(n3397)
         );
  AOI21_X1 U4179 ( .B1(n3490), .B2(n4316), .A(n3397), .ZN(n3399) );
  AOI22_X1 U4180 ( .A1(n4292), .A2(n4038), .B1(n4315), .B2(n4036), .ZN(n3398)
         );
  OAI211_X1 U4181 ( .C1(n3414), .C2(n4343), .A(n3399), .B(n3398), .ZN(n3403)
         );
  XNOR2_X1 U4182 ( .A(n3400), .B(n3911), .ZN(n3401) );
  NAND2_X1 U4183 ( .A1(n3401), .A2(n4366), .ZN(n3406) );
  NOR2_X1 U4184 ( .A1(n3406), .A2(n4661), .ZN(n3402) );
  AOI211_X1 U4185 ( .C1(n3408), .C2(n4311), .A(n3403), .B(n3402), .ZN(n3404)
         );
  INV_X1 U4186 ( .A(n3404), .ZN(U3278) );
  INV_X1 U4187 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4188 ( .A1(n4036), .A2(n4432), .B1(n4430), .B2(n3490), .ZN(n3405)
         );
  OAI211_X1 U4189 ( .C1(n3453), .C2(n4436), .A(n3406), .B(n3405), .ZN(n3407)
         );
  AOI21_X1 U4190 ( .B1(n3408), .B2(n4443), .A(n3407), .ZN(n3411) );
  MUX2_X1 U4191 ( .A(n3409), .B(n3411), .S(n4710), .Z(n3410) );
  OAI21_X1 U4192 ( .B1(n4446), .B2(n3414), .A(n3410), .ZN(U3530) );
  INV_X1 U4193 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3412) );
  MUX2_X1 U4194 ( .A(n3412), .B(n3411), .S(n4703), .Z(n3413) );
  OAI21_X1 U4195 ( .B1(n3414), .B2(n4492), .A(n3413), .ZN(U3491) );
  INV_X1 U4196 ( .A(n3415), .ZN(n3418) );
  INV_X1 U4197 ( .A(n3416), .ZN(n3417) );
  NAND2_X1 U4198 ( .A1(n3418), .A2(n3417), .ZN(n3419) );
  NAND2_X1 U4199 ( .A1(n4038), .A2(n2844), .ZN(n3422) );
  NAND2_X1 U4200 ( .A1(n3708), .A2(n3424), .ZN(n3421) );
  NAND2_X1 U4201 ( .A1(n3422), .A2(n3421), .ZN(n3423) );
  XNOR2_X1 U4202 ( .A(n3423), .B(n3711), .ZN(n3531) );
  NAND2_X1 U4203 ( .A1(n3714), .A2(n4038), .ZN(n3426) );
  NAND2_X1 U4204 ( .A1(n2844), .A2(n3424), .ZN(n3425) );
  INV_X1 U4205 ( .A(n3529), .ZN(n3528) );
  XNOR2_X1 U4206 ( .A(n3531), .B(n3528), .ZN(n3427) );
  XNOR2_X1 U4207 ( .A(n3500), .B(n3427), .ZN(n3434) );
  AND2_X1 U4208 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4573) );
  AOI21_X1 U4209 ( .B1(n3853), .B2(n4039), .A(n4573), .ZN(n3429) );
  NAND2_X1 U4210 ( .A1(n4512), .A2(n4037), .ZN(n3428) );
  OAI211_X1 U4211 ( .C1(n4509), .C2(n3430), .A(n3429), .B(n3428), .ZN(n3431)
         );
  AOI21_X1 U4212 ( .B1(n3859), .B2(n3432), .A(n3431), .ZN(n3433) );
  OAI21_X1 U4213 ( .B1(n3434), .B2(n3861), .A(n3433), .ZN(U3233) );
  NAND2_X1 U4214 ( .A1(n3550), .A2(n3868), .ZN(n3435) );
  INV_X1 U4215 ( .A(n3437), .ZN(n3920) );
  XNOR2_X1 U4216 ( .A(n3435), .B(n3920), .ZN(n3436) );
  NAND2_X1 U4217 ( .A1(n3436), .A2(n4366), .ZN(n3516) );
  XNOR2_X1 U4218 ( .A(n3438), .B(n3437), .ZN(n3519) );
  NAND2_X1 U4219 ( .A1(n3519), .A2(n4311), .ZN(n3444) );
  OAI21_X1 U4220 ( .B1(n3556), .B2(n3856), .A(n3474), .ZN(n3525) );
  INV_X1 U4221 ( .A(n3525), .ZN(n3442) );
  INV_X1 U4222 ( .A(n4316), .ZN(n4297) );
  AOI22_X1 U4223 ( .A1(n4292), .A2(n4035), .B1(n4315), .B2(n4033), .ZN(n3440)
         );
  AOI22_X1 U4224 ( .A1(n4661), .A2(REG2_REG_15__SCAN_IN), .B1(n3858), .B2(
        n4652), .ZN(n3439) );
  OAI211_X1 U4225 ( .C1(n3856), .C2(n4297), .A(n3440), .B(n3439), .ZN(n3441)
         );
  AOI21_X1 U4226 ( .B1(n3442), .B2(n4655), .A(n3441), .ZN(n3443) );
  OAI211_X1 U4227 ( .C1(n4661), .C2(n3516), .A(n3444), .B(n3443), .ZN(U3275)
         );
  INV_X1 U4228 ( .A(n3445), .ZN(n3446) );
  OAI21_X1 U4229 ( .B1(n3448), .B2(n3447), .A(n3446), .ZN(n4639) );
  INV_X1 U4230 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3459) );
  NAND2_X1 U4231 ( .A1(n3977), .A2(n3982), .ZN(n3929) );
  XOR2_X1 U4232 ( .A(n3929), .B(n3449), .Z(n3454) );
  INV_X1 U4233 ( .A(n3454), .ZN(n4641) );
  XOR2_X1 U4234 ( .A(n3929), .B(n3450), .Z(n3457) );
  AOI22_X1 U4235 ( .A1(n4040), .A2(n4420), .B1(n3451), .B2(n4430), .ZN(n3452)
         );
  OAI21_X1 U4236 ( .B1(n3453), .B2(n4424), .A(n3452), .ZN(n3456) );
  NOR2_X1 U4237 ( .A1(n3454), .A2(n3554), .ZN(n3455) );
  AOI211_X1 U4238 ( .C1(n3457), .C2(n4366), .A(n3456), .B(n3455), .ZN(n4644)
         );
  INV_X1 U4239 ( .A(n4644), .ZN(n3458) );
  AOI21_X1 U4240 ( .B1(n4700), .B2(n4641), .A(n3458), .ZN(n3461) );
  MUX2_X1 U4241 ( .A(n3459), .B(n3461), .S(n4703), .Z(n3460) );
  OAI21_X1 U4242 ( .B1(n4639), .B2(n4492), .A(n3460), .ZN(U3487) );
  INV_X1 U4243 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3462) );
  MUX2_X1 U4244 ( .A(n3462), .B(n3461), .S(n4710), .Z(n3463) );
  OAI21_X1 U4245 ( .B1(n4639), .B2(n4446), .A(n3463), .ZN(U3528) );
  INV_X1 U4246 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3466) );
  AOI21_X1 U4247 ( .B1(n3465), .B2(n4443), .A(n3464), .ZN(n3468) );
  MUX2_X1 U4248 ( .A(n3466), .B(n3468), .S(n4703), .Z(n3467) );
  OAI21_X1 U4249 ( .B1(n3471), .B2(n4492), .A(n3467), .ZN(U3493) );
  INV_X1 U4250 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3469) );
  MUX2_X1 U4251 ( .A(n3469), .B(n3468), .S(n4710), .Z(n3470) );
  OAI21_X1 U4252 ( .B1(n4446), .B2(n3471), .A(n3470), .ZN(U3531) );
  NOR2_X1 U4253 ( .A1(n2239), .A2(n3479), .ZN(n3472) );
  OR2_X1 U4254 ( .A1(n3473), .A2(n3472), .ZN(n3581) );
  NAND2_X1 U4255 ( .A1(n3474), .A2(n3641), .ZN(n3475) );
  NAND2_X1 U4256 ( .A1(n3571), .A2(n3475), .ZN(n3587) );
  INV_X1 U4257 ( .A(n3587), .ZN(n3478) );
  OAI22_X1 U4258 ( .A1(n4349), .A2(n3476), .B1(n4521), .B2(n4368), .ZN(n3477)
         );
  AOI21_X1 U4259 ( .B1(n3478), .B2(n4655), .A(n3477), .ZN(n3486) );
  XNOR2_X1 U4260 ( .A(n3480), .B(n3479), .ZN(n3484) );
  NAND2_X1 U4261 ( .A1(n4034), .A2(n4420), .ZN(n3482) );
  NAND2_X1 U4262 ( .A1(n4511), .A2(n4432), .ZN(n3481) );
  OAI211_X1 U4263 ( .C1(n4334), .C2(n4508), .A(n3482), .B(n3481), .ZN(n3483)
         );
  AOI21_X1 U4264 ( .B1(n3484), .B2(n4366), .A(n3483), .ZN(n3580) );
  OR2_X1 U4265 ( .A1(n3580), .A2(n4661), .ZN(n3485) );
  OAI211_X1 U4266 ( .C1(n3581), .C2(n4374), .A(n3486), .B(n3485), .ZN(U3274)
         );
  NAND2_X1 U4267 ( .A1(n4037), .A2(n2844), .ZN(n3488) );
  NAND2_X1 U4268 ( .A1(n3708), .A2(n3490), .ZN(n3487) );
  NAND2_X1 U4269 ( .A1(n3488), .A2(n3487), .ZN(n3489) );
  XNOR2_X1 U4270 ( .A(n3489), .B(n3725), .ZN(n3493) );
  NAND2_X1 U4271 ( .A1(n3714), .A2(n4037), .ZN(n3492) );
  NAND2_X1 U4272 ( .A1(n2844), .A2(n3490), .ZN(n3491) );
  NAND2_X1 U4273 ( .A1(n3492), .A2(n3491), .ZN(n3494) );
  NAND2_X1 U4274 ( .A1(n3493), .A2(n3494), .ZN(n3527) );
  OAI21_X1 U4275 ( .B1(n3531), .B2(n3529), .A(n3527), .ZN(n3499) );
  NAND3_X1 U4276 ( .A1(n3527), .A2(n3529), .A3(n3531), .ZN(n3497) );
  INV_X1 U4277 ( .A(n3493), .ZN(n3496) );
  INV_X1 U4278 ( .A(n3494), .ZN(n3495) );
  NAND2_X1 U4279 ( .A1(n3496), .A2(n3495), .ZN(n3526) );
  NAND2_X1 U4280 ( .A1(n4036), .A2(n2844), .ZN(n3502) );
  NAND2_X1 U4281 ( .A1(n3708), .A2(n3504), .ZN(n3501) );
  NAND2_X1 U4282 ( .A1(n3502), .A2(n3501), .ZN(n3503) );
  XNOR2_X1 U4283 ( .A(n3503), .B(n3711), .ZN(n3589) );
  INV_X1 U4284 ( .A(n3589), .ZN(n3592) );
  NAND2_X1 U4285 ( .A1(n3714), .A2(n4036), .ZN(n3506) );
  NAND2_X1 U4286 ( .A1(n2844), .A2(n3504), .ZN(n3505) );
  NAND2_X1 U4287 ( .A1(n3506), .A2(n3505), .ZN(n3590) );
  XNOR2_X1 U4288 ( .A(n3592), .B(n3590), .ZN(n3507) );
  XNOR2_X1 U4289 ( .A(n3591), .B(n3507), .ZN(n3514) );
  NOR2_X1 U4290 ( .A1(STATE_REG_SCAN_IN), .A2(n2548), .ZN(n4590) );
  AOI21_X1 U4291 ( .B1(n3853), .B2(n4037), .A(n4590), .ZN(n3509) );
  NAND2_X1 U4292 ( .A1(n4512), .A2(n4035), .ZN(n3508) );
  OAI211_X1 U4293 ( .C1(n4509), .C2(n3510), .A(n3509), .B(n3508), .ZN(n3511)
         );
  AOI21_X1 U4294 ( .B1(n3859), .B2(n3512), .A(n3511), .ZN(n3513) );
  OAI21_X1 U4295 ( .B1(n3514), .B2(n3861), .A(n3513), .ZN(U3231) );
  AOI22_X1 U4296 ( .A1(n4033), .A2(n4432), .B1(n4430), .B2(n3634), .ZN(n3515)
         );
  OAI211_X1 U4297 ( .C1(n3517), .C2(n4436), .A(n3516), .B(n3515), .ZN(n3518)
         );
  AOI21_X1 U4298 ( .B1(n3519), .B2(n4443), .A(n3518), .ZN(n3523) );
  INV_X1 U4299 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3520) );
  MUX2_X1 U4300 ( .A(n3523), .B(n3520), .S(n4701), .Z(n3521) );
  OAI21_X1 U4301 ( .B1(n3525), .B2(n4492), .A(n3521), .ZN(U3497) );
  INV_X1 U4302 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3522) );
  MUX2_X1 U4303 ( .A(n3523), .B(n3522), .S(n4711), .Z(n3524) );
  OAI21_X1 U4304 ( .B1(n4446), .B2(n3525), .A(n3524), .ZN(U3533) );
  NAND2_X1 U4305 ( .A1(n3527), .A2(n3526), .ZN(n3534) );
  NOR2_X1 U4306 ( .A1(n3500), .A2(n3528), .ZN(n3532) );
  INV_X1 U4307 ( .A(n3500), .ZN(n3530) );
  OAI22_X1 U4308 ( .A1(n3532), .A2(n3531), .B1(n3530), .B2(n3529), .ZN(n3533)
         );
  XOR2_X1 U4309 ( .A(n3534), .B(n3533), .Z(n3541) );
  NOR2_X1 U4310 ( .A1(STATE_REG_SCAN_IN), .A2(n4865), .ZN(n4583) );
  AOI21_X1 U4311 ( .B1(n3853), .B2(n4038), .A(n4583), .ZN(n3536) );
  NAND2_X1 U4312 ( .A1(n4512), .A2(n4036), .ZN(n3535) );
  OAI211_X1 U4313 ( .C1(n4509), .C2(n3537), .A(n3536), .B(n3535), .ZN(n3538)
         );
  AOI21_X1 U4314 ( .B1(n3859), .B2(n3539), .A(n3538), .ZN(n3540) );
  OAI21_X1 U4315 ( .B1(n3541), .B2(n3861), .A(n3540), .ZN(U3221) );
  OR2_X1 U4316 ( .A1(n3543), .A2(n3542), .ZN(n3546) );
  AND2_X1 U4317 ( .A1(n3546), .A2(n3544), .ZN(n3548) );
  NAND2_X1 U4318 ( .A1(n3546), .A2(n3545), .ZN(n3547) );
  OAI21_X1 U4319 ( .B1(n3548), .B2(n3552), .A(n3547), .ZN(n3614) );
  INV_X1 U4320 ( .A(n3614), .ZN(n3566) );
  INV_X1 U4321 ( .A(n3549), .ZN(n3872) );
  INV_X1 U4322 ( .A(n3550), .ZN(n3551) );
  AOI21_X1 U4323 ( .B1(n3872), .B2(n3552), .A(n3551), .ZN(n3553) );
  OAI22_X1 U4324 ( .A1(n3566), .A2(n3554), .B1(n4339), .B2(n3553), .ZN(n3612)
         );
  NAND2_X1 U4325 ( .A1(n3612), .A2(n4349), .ZN(n3564) );
  INV_X1 U4326 ( .A(n3555), .ZN(n3558) );
  INV_X1 U4327 ( .A(n3556), .ZN(n3557) );
  OAI21_X1 U4328 ( .B1(n3558), .B2(n3603), .A(n3557), .ZN(n3620) );
  INV_X1 U4329 ( .A(n3620), .ZN(n3562) );
  AOI22_X1 U4330 ( .A1(n4292), .A2(n4036), .B1(n4315), .B2(n4034), .ZN(n3560)
         );
  AOI22_X1 U4331 ( .A1(n4661), .A2(REG2_REG_14__SCAN_IN), .B1(n3588), .B2(
        n4652), .ZN(n3559) );
  OAI211_X1 U4332 ( .C1(n3603), .C2(n4297), .A(n3560), .B(n3559), .ZN(n3561)
         );
  AOI21_X1 U4333 ( .B1(n3562), .B2(n4655), .A(n3561), .ZN(n3563) );
  OAI211_X1 U4334 ( .C1(n3566), .C2(n3565), .A(n3564), .B(n3563), .ZN(U3276)
         );
  INV_X1 U4335 ( .A(n4243), .ZN(n3567) );
  AND2_X1 U4336 ( .A1(n3567), .A2(n4327), .ZN(n3912) );
  INV_X1 U4337 ( .A(n3912), .ZN(n3568) );
  XNOR2_X1 U4338 ( .A(n4244), .B(n3568), .ZN(n3569) );
  NAND2_X1 U4339 ( .A1(n3569), .A2(n4366), .ZN(n3622) );
  XOR2_X1 U4340 ( .A(n3912), .B(n3570), .Z(n3624) );
  NAND2_X1 U4341 ( .A1(n3624), .A2(n4311), .ZN(n3579) );
  INV_X1 U4342 ( .A(n3571), .ZN(n3573) );
  INV_X1 U4343 ( .A(n4360), .ZN(n3572) );
  OAI21_X1 U4344 ( .B1(n3573), .B2(n3790), .A(n3572), .ZN(n3630) );
  INV_X1 U4345 ( .A(n3630), .ZN(n3577) );
  AOI22_X1 U4346 ( .A1(n4292), .A2(n4033), .B1(n4315), .B2(n4337), .ZN(n3575)
         );
  AOI22_X1 U4347 ( .A1(n4661), .A2(REG2_REG_17__SCAN_IN), .B1(n3792), .B2(
        n4652), .ZN(n3574) );
  OAI211_X1 U4348 ( .C1(n3790), .C2(n4297), .A(n3575), .B(n3574), .ZN(n3576)
         );
  AOI21_X1 U4349 ( .B1(n3577), .B2(n4655), .A(n3576), .ZN(n3578) );
  OAI211_X1 U4350 ( .C1(n4661), .C2(n3622), .A(n3579), .B(n3578), .ZN(U3273)
         );
  OAI21_X1 U4351 ( .B1(n3581), .B2(n4690), .A(n3580), .ZN(n3584) );
  MUX2_X1 U4352 ( .A(REG1_REG_16__SCAN_IN), .B(n3584), .S(n4710), .Z(n3582) );
  INV_X1 U4353 ( .A(n3582), .ZN(n3583) );
  OAI21_X1 U4354 ( .B1(n4446), .B2(n3587), .A(n3583), .ZN(U3534) );
  MUX2_X1 U4355 ( .A(REG0_REG_16__SCAN_IN), .B(n3584), .S(n4703), .Z(n3585) );
  INV_X1 U4356 ( .A(n3585), .ZN(n3586) );
  OAI21_X1 U4357 ( .B1(n3587), .B2(n4492), .A(n3586), .ZN(U3499) );
  INV_X1 U4358 ( .A(n3588), .ZN(n3608) );
  NAND2_X1 U4359 ( .A1(n4035), .A2(n2844), .ZN(n3594) );
  NAND2_X1 U4360 ( .A1(n3708), .A2(n3609), .ZN(n3593) );
  NAND2_X1 U4361 ( .A1(n3594), .A2(n3593), .ZN(n3595) );
  XNOR2_X1 U4362 ( .A(n3595), .B(n3711), .ZN(n3600) );
  INV_X1 U4363 ( .A(n3600), .ZN(n3598) );
  NOR2_X1 U4364 ( .A1(n3727), .A2(n3603), .ZN(n3596) );
  AOI21_X1 U4365 ( .B1(n3714), .B2(n4035), .A(n3596), .ZN(n3599) );
  INV_X1 U4366 ( .A(n3599), .ZN(n3597) );
  NAND2_X1 U4367 ( .A1(n3598), .A2(n3597), .ZN(n3632) );
  AND2_X1 U4368 ( .A1(n3600), .A2(n3599), .ZN(n3631) );
  NOR2_X1 U4369 ( .A1(n2355), .A2(n3631), .ZN(n3601) );
  XNOR2_X1 U4370 ( .A(n3633), .B(n3601), .ZN(n3602) );
  NAND2_X1 U4371 ( .A1(n3602), .A2(n4517), .ZN(n3607) );
  INV_X1 U4372 ( .A(n4036), .ZN(n3611) );
  OAI22_X1 U4373 ( .A1(n4509), .A2(n3603), .B1(n3611), .B2(n4506), .ZN(n3605)
         );
  INV_X1 U4374 ( .A(n4034), .ZN(n4507) );
  NAND2_X1 U4375 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4597) );
  OAI21_X1 U4376 ( .B1(n3844), .B2(n4507), .A(n4597), .ZN(n3604) );
  NOR2_X1 U4377 ( .A1(n3605), .A2(n3604), .ZN(n3606) );
  OAI211_X1 U4378 ( .C1(n4522), .C2(n3608), .A(n3607), .B(n3606), .ZN(U3212)
         );
  INV_X1 U4379 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4380 ( .A1(n4034), .A2(n4432), .B1(n3609), .B2(n4430), .ZN(n3610)
         );
  OAI21_X1 U4381 ( .B1(n3611), .B2(n4436), .A(n3610), .ZN(n3613) );
  AOI211_X1 U4382 ( .C1(n4700), .C2(n3614), .A(n3613), .B(n3612), .ZN(n3617)
         );
  MUX2_X1 U4383 ( .A(n3615), .B(n3617), .S(n4703), .Z(n3616) );
  OAI21_X1 U4384 ( .B1(n3620), .B2(n4492), .A(n3616), .ZN(U3495) );
  INV_X1 U4385 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3618) );
  MUX2_X1 U4386 ( .A(n3618), .B(n3617), .S(n4710), .Z(n3619) );
  OAI21_X1 U4387 ( .B1(n4446), .B2(n3620), .A(n3619), .ZN(U3532) );
  INV_X1 U4388 ( .A(REG0_REG_17__SCAN_IN), .ZN(n3625) );
  INV_X1 U4389 ( .A(n4033), .ZN(n3643) );
  AOI22_X1 U4390 ( .A1(n4337), .A2(n4432), .B1(n4430), .B2(n3649), .ZN(n3621)
         );
  OAI211_X1 U4391 ( .C1(n3643), .C2(n4436), .A(n3622), .B(n3621), .ZN(n3623)
         );
  AOI21_X1 U4392 ( .B1(n3624), .B2(n4443), .A(n3623), .ZN(n3627) );
  MUX2_X1 U4393 ( .A(n3625), .B(n3627), .S(n4703), .Z(n3626) );
  OAI21_X1 U4394 ( .B1(n3630), .B2(n4492), .A(n3626), .ZN(U3501) );
  INV_X1 U4395 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3628) );
  MUX2_X1 U4396 ( .A(n3628), .B(n3627), .S(n4710), .Z(n3629) );
  OAI21_X1 U4397 ( .B1(n4446), .B2(n3630), .A(n3629), .ZN(U3535) );
  NAND2_X1 U4398 ( .A1(n4034), .A2(n2844), .ZN(n3636) );
  NAND2_X1 U4399 ( .A1(n3708), .A2(n3634), .ZN(n3635) );
  NAND2_X1 U4400 ( .A1(n3636), .A2(n3635), .ZN(n3637) );
  XNOR2_X1 U4401 ( .A(n3637), .B(n3725), .ZN(n3639) );
  NOR2_X1 U4402 ( .A1(n3727), .A2(n3856), .ZN(n3638) );
  AOI21_X1 U4403 ( .B1(n3714), .B2(n4034), .A(n3638), .ZN(n4514) );
  AOI22_X1 U4404 ( .A1(n4033), .A2(n2844), .B1(n3641), .B2(n3708), .ZN(n3642)
         );
  XOR2_X1 U4405 ( .A(n3725), .B(n3642), .Z(n3645) );
  OAI22_X1 U4406 ( .A1(n3643), .A2(n3724), .B1(n4508), .B2(n3727), .ZN(n3644)
         );
  NOR2_X1 U4407 ( .A1(n3645), .A2(n3644), .ZN(n3646) );
  AOI21_X1 U4408 ( .B1(n3645), .B2(n3644), .A(n3646), .ZN(n4516) );
  NAND2_X1 U4409 ( .A1(n4511), .A2(n2844), .ZN(n3651) );
  NAND2_X1 U4410 ( .A1(n3708), .A2(n3649), .ZN(n3650) );
  NAND2_X1 U4411 ( .A1(n3651), .A2(n3650), .ZN(n3652) );
  XNOR2_X1 U4412 ( .A(n3652), .B(n3711), .ZN(n3655) );
  NOR2_X1 U4413 ( .A1(n3727), .A2(n3790), .ZN(n3653) );
  AOI21_X1 U4414 ( .B1(n3714), .B2(n4511), .A(n3653), .ZN(n3654) );
  NOR2_X1 U4415 ( .A1(n3655), .A2(n3654), .ZN(n3786) );
  NAND2_X1 U4416 ( .A1(n4337), .A2(n2844), .ZN(n3657) );
  NAND2_X1 U4417 ( .A1(n3708), .A2(n4363), .ZN(n3656) );
  NAND2_X1 U4418 ( .A1(n3657), .A2(n3656), .ZN(n3658) );
  XNOR2_X1 U4419 ( .A(n3658), .B(n3725), .ZN(n3661) );
  NAND2_X1 U4420 ( .A1(n4337), .A2(n3714), .ZN(n3660) );
  NAND2_X1 U4421 ( .A1(n2844), .A2(n4363), .ZN(n3659) );
  NAND2_X1 U4422 ( .A1(n3660), .A2(n3659), .ZN(n3662) );
  NAND2_X1 U4423 ( .A1(n3661), .A2(n3662), .ZN(n3829) );
  INV_X1 U4424 ( .A(n3661), .ZN(n3664) );
  INV_X1 U4425 ( .A(n3662), .ZN(n3663) );
  NAND2_X1 U4426 ( .A1(n3664), .A2(n3663), .ZN(n3828) );
  NAND2_X1 U4427 ( .A1(n4032), .A2(n2844), .ZN(n3666) );
  NAND2_X1 U4428 ( .A1(n3708), .A2(n3668), .ZN(n3665) );
  NAND2_X1 U4429 ( .A1(n3666), .A2(n3665), .ZN(n3667) );
  XNOR2_X1 U4430 ( .A(n3667), .B(n3725), .ZN(n3669) );
  AOI22_X1 U4431 ( .A1(n4032), .A2(n3714), .B1(n2844), .B2(n3668), .ZN(n3670)
         );
  XNOR2_X1 U4432 ( .A(n3669), .B(n3670), .ZN(n3759) );
  INV_X1 U4433 ( .A(n3669), .ZN(n3671) );
  NAND2_X1 U4434 ( .A1(n4421), .A2(n2844), .ZN(n3673) );
  NAND2_X1 U4435 ( .A1(n3708), .A2(n4431), .ZN(n3672) );
  NAND2_X1 U4436 ( .A1(n3673), .A2(n3672), .ZN(n3674) );
  XNOR2_X1 U4437 ( .A(n3674), .B(n3711), .ZN(n3681) );
  NOR2_X1 U4438 ( .A1(n3727), .A2(n4313), .ZN(n3675) );
  AOI21_X1 U4439 ( .B1(n4421), .B2(n3714), .A(n3675), .ZN(n3680) );
  NOR2_X1 U4440 ( .A1(n3681), .A2(n3680), .ZN(n3805) );
  NAND2_X1 U4441 ( .A1(n4433), .A2(n2844), .ZN(n3677) );
  NAND2_X1 U4442 ( .A1(n3708), .A2(n4419), .ZN(n3676) );
  NAND2_X1 U4443 ( .A1(n3677), .A2(n3676), .ZN(n3678) );
  XNOR2_X1 U4444 ( .A(n3678), .B(n3711), .ZN(n3766) );
  NOR2_X1 U4445 ( .A1(n3727), .A2(n4298), .ZN(n3679) );
  AOI21_X1 U4446 ( .B1(n4433), .B2(n3714), .A(n3679), .ZN(n3767) );
  NAND2_X1 U4447 ( .A1(n3766), .A2(n3767), .ZN(n3682) );
  NAND2_X1 U4448 ( .A1(n3681), .A2(n3680), .ZN(n3806) );
  OAI21_X1 U4449 ( .B1(n3765), .B2(n3805), .A(n2373), .ZN(n3686) );
  INV_X1 U4450 ( .A(n3766), .ZN(n3684) );
  NAND2_X1 U4451 ( .A1(n3686), .A2(n3685), .ZN(n3816) );
  OAI22_X1 U4452 ( .A1(n4425), .A2(n3727), .B1(n4279), .B2(n3687), .ZN(n3688)
         );
  XNOR2_X1 U4453 ( .A(n3688), .B(n3725), .ZN(n3690) );
  OAI22_X1 U4454 ( .A1(n4425), .A2(n3724), .B1(n4279), .B2(n3727), .ZN(n3689)
         );
  XNOR2_X1 U4455 ( .A(n3690), .B(n3689), .ZN(n3817) );
  NOR2_X1 U4456 ( .A1(n3690), .A2(n3689), .ZN(n3750) );
  NAND2_X1 U4457 ( .A1(n4402), .A2(n2844), .ZN(n3692) );
  NAND2_X1 U4458 ( .A1(n3708), .A2(n2253), .ZN(n3691) );
  NAND2_X1 U4459 ( .A1(n3692), .A2(n3691), .ZN(n3693) );
  XNOR2_X1 U4460 ( .A(n3693), .B(n3711), .ZN(n3696) );
  NOR2_X1 U4461 ( .A1(n3727), .A2(n4257), .ZN(n3694) );
  AOI21_X1 U4462 ( .B1(n4402), .B2(n3714), .A(n3694), .ZN(n3695) );
  XNOR2_X1 U4463 ( .A(n3696), .B(n3695), .ZN(n3749) );
  NOR2_X1 U4464 ( .A1(n3696), .A2(n3695), .ZN(n3700) );
  NAND2_X1 U4465 ( .A1(n4210), .A2(n3714), .ZN(n3698) );
  NAND2_X1 U4466 ( .A1(n2844), .A2(n4401), .ZN(n3697) );
  OAI22_X1 U4467 ( .A1(n4253), .A2(n3727), .B1(n4236), .B2(n3687), .ZN(n3699)
         );
  XOR2_X1 U4468 ( .A(n3725), .B(n3699), .Z(n3797) );
  NAND2_X1 U4469 ( .A1(n4231), .A2(n2844), .ZN(n3702) );
  NAND2_X1 U4470 ( .A1(n3708), .A2(n4214), .ZN(n3701) );
  NAND2_X1 U4471 ( .A1(n3702), .A2(n3701), .ZN(n3703) );
  XNOR2_X1 U4472 ( .A(n3703), .B(n3711), .ZN(n3707) );
  NOR2_X1 U4473 ( .A1(n3727), .A2(n3704), .ZN(n3705) );
  AOI21_X1 U4474 ( .B1(n4231), .B2(n3714), .A(n3705), .ZN(n3706) );
  NAND2_X1 U4475 ( .A1(n3707), .A2(n3706), .ZN(n3776) );
  NOR2_X1 U4476 ( .A1(n3707), .A2(n3706), .ZN(n3777) );
  NAND2_X1 U4477 ( .A1(n4385), .A2(n2844), .ZN(n3710) );
  NAND2_X1 U4478 ( .A1(n3708), .A2(n4197), .ZN(n3709) );
  NAND2_X1 U4479 ( .A1(n3710), .A2(n3709), .ZN(n3712) );
  XNOR2_X1 U4480 ( .A(n3712), .B(n3711), .ZN(n3718) );
  INV_X1 U4481 ( .A(n3718), .ZN(n3716) );
  NOR2_X1 U4482 ( .A1(n3727), .A2(n3843), .ZN(n3713) );
  AOI21_X1 U4483 ( .B1(n4385), .B2(n3714), .A(n3713), .ZN(n3717) );
  INV_X1 U4484 ( .A(n3717), .ZN(n3715) );
  NAND2_X1 U4485 ( .A1(n3716), .A2(n3715), .ZN(n3838) );
  AND2_X1 U4486 ( .A1(n3718), .A2(n3717), .ZN(n3837) );
  OR2_X1 U4487 ( .A1(n4195), .A2(n3724), .ZN(n3720) );
  NAND2_X1 U4488 ( .A1(n2844), .A2(n4384), .ZN(n3719) );
  NAND2_X1 U4489 ( .A1(n3720), .A2(n3719), .ZN(n3723) );
  OAI22_X1 U4490 ( .A1(n4195), .A2(n3727), .B1(n3687), .B2(n4182), .ZN(n3721)
         );
  XNOR2_X1 U4491 ( .A(n3721), .B(n3725), .ZN(n3722) );
  XOR2_X1 U4492 ( .A(n3723), .B(n3722), .Z(n3741) );
  AOI22_X1 U4493 ( .A1(n3742), .A2(n3741), .B1(n3723), .B2(n3722), .ZN(n3731)
         );
  OAI22_X1 U4494 ( .A1(n4388), .A2(n3724), .B1(n4163), .B2(n3727), .ZN(n3726)
         );
  XNOR2_X1 U4495 ( .A(n3726), .B(n3725), .ZN(n3729) );
  OAI22_X1 U4496 ( .A1(n4388), .A2(n2843), .B1(n4163), .B2(n3687), .ZN(n3728)
         );
  XNOR2_X1 U4497 ( .A(n3729), .B(n3728), .ZN(n3730) );
  XNOR2_X1 U4498 ( .A(n3731), .B(n3730), .ZN(n3737) );
  OAI22_X1 U4499 ( .A1(n3732), .A2(n3844), .B1(n4509), .B2(n4163), .ZN(n3735)
         );
  OAI22_X1 U4500 ( .A1(n4195), .A2(n4506), .B1(STATE_REG_SCAN_IN), .B2(n3733), 
        .ZN(n3734) );
  AOI211_X1 U4501 ( .C1(n4160), .C2(n3859), .A(n3735), .B(n3734), .ZN(n3736)
         );
  OAI21_X1 U4502 ( .B1(n3737), .B2(n3861), .A(n3736), .ZN(U3217) );
  INV_X1 U4503 ( .A(IR_REG_30__SCAN_IN), .ZN(n3739) );
  NAND3_X1 U4504 ( .A1(n3739), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3740) );
  INV_X1 U4505 ( .A(DATAI_31_), .ZN(n4973) );
  OAI22_X1 U4506 ( .A1(n3738), .A2(n3740), .B1(STATE_REG_SCAN_IN), .B2(n4973), 
        .ZN(U3321) );
  XNOR2_X1 U4507 ( .A(n3742), .B(n3741), .ZN(n3747) );
  OAI22_X1 U4508 ( .A1(n4213), .A2(n4506), .B1(n4509), .B2(n4182), .ZN(n3745)
         );
  OAI22_X1 U4509 ( .A1(n4388), .A2(n3844), .B1(STATE_REG_SCAN_IN), .B2(n3743), 
        .ZN(n3744) );
  AOI211_X1 U4510 ( .C1(n4179), .C2(n3859), .A(n3745), .B(n3744), .ZN(n3746)
         );
  OAI21_X1 U4511 ( .B1(n3747), .B2(n3861), .A(n3746), .ZN(U3211) );
  INV_X1 U4512 ( .A(n3748), .ZN(n3752) );
  OAI21_X1 U4513 ( .B1(n3815), .B2(n3750), .A(n3749), .ZN(n3751) );
  NAND3_X1 U4514 ( .A1(n3752), .A2(n4517), .A3(n3751), .ZN(n3757) );
  NAND2_X1 U4515 ( .A1(n4512), .A2(n4210), .ZN(n3753) );
  OAI21_X1 U4516 ( .B1(n4509), .B2(n4257), .A(n3753), .ZN(n3755) );
  INV_X1 U4517 ( .A(REG3_REG_23__SCAN_IN), .ZN(n5054) );
  OAI22_X1 U4518 ( .A1(n4506), .A2(n4425), .B1(STATE_REG_SCAN_IN), .B2(n5054), 
        .ZN(n3754) );
  NOR2_X1 U4519 ( .A1(n3755), .A2(n3754), .ZN(n3756) );
  OAI211_X1 U4520 ( .C1(n4522), .C2(n4260), .A(n3757), .B(n3756), .ZN(U3213)
         );
  XOR2_X1 U4521 ( .A(n3759), .B(n3758), .Z(n3764) );
  AND2_X1 U4522 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4131) );
  AOI21_X1 U4523 ( .B1(n3853), .B2(n4337), .A(n4131), .ZN(n3761) );
  NAND2_X1 U4524 ( .A1(n4512), .A2(n4421), .ZN(n3760) );
  OAI211_X1 U4525 ( .C1(n4509), .C2(n4342), .A(n3761), .B(n3760), .ZN(n3762)
         );
  AOI21_X1 U4526 ( .B1(n3859), .B2(n4344), .A(n3762), .ZN(n3763) );
  OAI21_X1 U4527 ( .B1(n3764), .B2(n3861), .A(n3763), .ZN(U3216) );
  AOI21_X1 U4528 ( .B1(n3765), .B2(n3806), .A(n3805), .ZN(n3769) );
  XOR2_X1 U4529 ( .A(n3767), .B(n3766), .Z(n3768) );
  XNOR2_X1 U4530 ( .A(n3769), .B(n3768), .ZN(n3770) );
  NAND2_X1 U4531 ( .A1(n3770), .A2(n4517), .ZN(n3774) );
  OAI22_X1 U4532 ( .A1(n4509), .A2(n4298), .B1(n4425), .B2(n3844), .ZN(n3772)
         );
  INV_X1 U4533 ( .A(n4421), .ZN(n4335) );
  OAI22_X1 U4534 ( .A1(n4506), .A2(n4335), .B1(STATE_REG_SCAN_IN), .B2(n5031), 
        .ZN(n3771) );
  NOR2_X1 U4535 ( .A1(n3772), .A2(n3771), .ZN(n3773) );
  OAI211_X1 U4536 ( .C1(n4522), .C2(n4293), .A(n3774), .B(n3773), .ZN(U3220)
         );
  NOR2_X1 U4537 ( .A1(n3777), .A2(n2345), .ZN(n3778) );
  XNOR2_X1 U4538 ( .A(n3775), .B(n3778), .ZN(n3784) );
  INV_X1 U4539 ( .A(n4217), .ZN(n3781) );
  AOI22_X1 U4540 ( .A1(n3853), .A2(n4210), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3780) );
  AOI22_X1 U4541 ( .A1(n4214), .A2(n3799), .B1(n4385), .B2(n4512), .ZN(n3779)
         );
  OAI211_X1 U4542 ( .C1(n4522), .C2(n3781), .A(n3780), .B(n3779), .ZN(n3782)
         );
  INV_X1 U4543 ( .A(n3782), .ZN(n3783) );
  OAI21_X1 U4544 ( .B1(n3784), .B2(n3861), .A(n3783), .ZN(U3222) );
  NOR2_X1 U4545 ( .A1(n3786), .A2(n2246), .ZN(n3787) );
  XNOR2_X1 U4546 ( .A(n3785), .B(n3787), .ZN(n3794) );
  NOR2_X1 U4547 ( .A1(STATE_REG_SCAN_IN), .A2(n2397), .ZN(n4629) );
  AOI21_X1 U4548 ( .B1(n3853), .B2(n4033), .A(n4629), .ZN(n3789) );
  NAND2_X1 U4549 ( .A1(n4512), .A2(n4337), .ZN(n3788) );
  OAI211_X1 U4550 ( .C1(n4509), .C2(n3790), .A(n3789), .B(n3788), .ZN(n3791)
         );
  AOI21_X1 U4551 ( .B1(n3859), .B2(n3792), .A(n3791), .ZN(n3793) );
  OAI21_X1 U4552 ( .B1(n3794), .B2(n3861), .A(n3793), .ZN(U3225) );
  NAND2_X1 U4553 ( .A1(n2340), .A2(n3796), .ZN(n3798) );
  XNOR2_X1 U4554 ( .A(n3798), .B(n3797), .ZN(n3804) );
  AOI22_X1 U4555 ( .A1(n3853), .A2(n4402), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3801) );
  AOI22_X1 U4556 ( .A1(n3799), .A2(n4401), .B1(n4512), .B2(n4231), .ZN(n3800)
         );
  OAI211_X1 U4557 ( .C1(n4522), .C2(n4232), .A(n3801), .B(n3800), .ZN(n3802)
         );
  INV_X1 U4558 ( .A(n3802), .ZN(n3803) );
  OAI21_X1 U4559 ( .B1(n3804), .B2(n3861), .A(n3803), .ZN(U3226) );
  INV_X1 U4560 ( .A(n3805), .ZN(n3807) );
  NAND2_X1 U4561 ( .A1(n3807), .A2(n3806), .ZN(n3808) );
  XNOR2_X1 U4562 ( .A(n3765), .B(n3808), .ZN(n3809) );
  NAND2_X1 U4563 ( .A1(n3809), .A2(n4517), .ZN(n3814) );
  OAI22_X1 U4564 ( .A1(n4509), .A2(n4313), .B1(n3819), .B2(n3844), .ZN(n3812)
         );
  INV_X1 U4565 ( .A(n4032), .ZN(n4437) );
  OAI22_X1 U4566 ( .A1(n4506), .A2(n4437), .B1(STATE_REG_SCAN_IN), .B2(n3810), 
        .ZN(n3811) );
  NOR2_X1 U4567 ( .A1(n3812), .A2(n3811), .ZN(n3813) );
  OAI211_X1 U4568 ( .C1(n4522), .C2(n4317), .A(n3814), .B(n3813), .ZN(U3230)
         );
  AOI21_X1 U4569 ( .B1(n3817), .B2(n3816), .A(n3815), .ZN(n3824) );
  INV_X1 U4570 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3818) );
  OAI22_X1 U4571 ( .A1(n4506), .A2(n3819), .B1(STATE_REG_SCAN_IN), .B2(n3818), 
        .ZN(n3822) );
  OAI22_X1 U4572 ( .A1(n4509), .A2(n4279), .B1(n3820), .B2(n3844), .ZN(n3821)
         );
  AOI211_X1 U4573 ( .C1(n3859), .C2(n4270), .A(n3822), .B(n3821), .ZN(n3823)
         );
  OAI21_X1 U4574 ( .B1(n3824), .B2(n3861), .A(n3823), .ZN(U3232) );
  INV_X1 U4575 ( .A(n3828), .ZN(n3825) );
  NOR2_X1 U4576 ( .A1(n3826), .A2(n3825), .ZN(n3831) );
  AOI21_X1 U4577 ( .B1(n3829), .B2(n3828), .A(n3827), .ZN(n3830) );
  OAI21_X1 U4578 ( .B1(n3831), .B2(n3830), .A(n4517), .ZN(n3836) );
  OAI22_X1 U4579 ( .A1(n4509), .A2(n4359), .B1(n4437), .B2(n3844), .ZN(n3834)
         );
  INV_X1 U4580 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4116) );
  OAI22_X1 U4581 ( .A1(n4506), .A2(n3832), .B1(STATE_REG_SCAN_IN), .B2(n4116), 
        .ZN(n3833) );
  NOR2_X1 U4582 ( .A1(n3834), .A2(n3833), .ZN(n3835) );
  OAI211_X1 U4583 ( .C1(n4522), .C2(n4369), .A(n3836), .B(n3835), .ZN(U3235)
         );
  INV_X1 U4584 ( .A(n3837), .ZN(n3839) );
  NAND2_X1 U4585 ( .A1(n3839), .A2(n3838), .ZN(n3840) );
  XNOR2_X1 U4586 ( .A(n3841), .B(n3840), .ZN(n3849) );
  INV_X1 U4587 ( .A(n4200), .ZN(n3847) );
  OAI22_X1 U4588 ( .A1(n4405), .A2(n4506), .B1(STATE_REG_SCAN_IN), .B2(n3842), 
        .ZN(n3846) );
  OAI22_X1 U4589 ( .A1(n4195), .A2(n3844), .B1(n4509), .B2(n3843), .ZN(n3845)
         );
  AOI211_X1 U4590 ( .C1(n3847), .C2(n3859), .A(n3846), .B(n3845), .ZN(n3848)
         );
  OAI21_X1 U4591 ( .B1(n3849), .B2(n3861), .A(n3848), .ZN(U3237) );
  INV_X1 U4592 ( .A(n3850), .ZN(n3851) );
  NAND2_X1 U4593 ( .A1(n3851), .A2(n4513), .ZN(n3852) );
  XNOR2_X1 U4594 ( .A(n3852), .B(n4514), .ZN(n3862) );
  AND2_X1 U4595 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4610) );
  AOI21_X1 U4596 ( .B1(n4512), .B2(n4033), .A(n4610), .ZN(n3855) );
  NAND2_X1 U4597 ( .A1(n3853), .A2(n4035), .ZN(n3854) );
  OAI211_X1 U4598 ( .C1(n4509), .C2(n3856), .A(n3855), .B(n3854), .ZN(n3857)
         );
  AOI21_X1 U4599 ( .B1(n3859), .B2(n3858), .A(n3857), .ZN(n3860) );
  OAI21_X1 U4600 ( .B1(n3862), .B2(n3861), .A(n3860), .ZN(U3238) );
  NAND2_X1 U4601 ( .A1(n3863), .A2(DATAI_31_), .ZN(n4141) );
  INV_X1 U4602 ( .A(n4141), .ZN(n3897) );
  NAND2_X1 U4603 ( .A1(n3863), .A2(DATAI_30_), .ZN(n3892) );
  AND2_X1 U4604 ( .A1(n4029), .A2(n3892), .ZN(n3905) );
  INV_X1 U4605 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4142) );
  NAND2_X1 U4606 ( .A1(n3864), .A2(REG1_REG_31__SCAN_IN), .ZN(n3866) );
  NAND2_X1 U4607 ( .A1(n2547), .A2(REG0_REG_31__SCAN_IN), .ZN(n3865) );
  OAI211_X1 U4608 ( .C1(n2423), .C2(n4142), .A(n3866), .B(n3865), .ZN(n4140)
         );
  NOR2_X1 U4609 ( .A1(n4140), .A2(n4141), .ZN(n3904) );
  INV_X1 U4610 ( .A(n3901), .ZN(n3867) );
  NOR2_X1 U4611 ( .A1(n3898), .A2(n3867), .ZN(n4005) );
  INV_X1 U4612 ( .A(n4005), .ZN(n3881) );
  AND2_X1 U4613 ( .A1(n3868), .A2(n3871), .ZN(n3988) );
  NAND2_X1 U4614 ( .A1(n3870), .A2(n3869), .ZN(n3971) );
  AND2_X1 U4615 ( .A1(n3971), .A2(n3871), .ZN(n3987) );
  AOI21_X1 U4616 ( .B1(n3872), .B2(n3988), .A(n3987), .ZN(n3874) );
  INV_X1 U4617 ( .A(n3994), .ZN(n3873) );
  OAI21_X1 U4618 ( .B1(n3874), .B2(n3873), .A(n3990), .ZN(n3877) );
  INV_X1 U4619 ( .A(n3875), .ZN(n3876) );
  AOI21_X1 U4620 ( .B1(n3877), .B2(n4247), .A(n3876), .ZN(n3879) );
  OAI21_X1 U4621 ( .B1(n3879), .B2(n3999), .A(n3878), .ZN(n3880) );
  OAI221_X1 U4622 ( .B1(n3881), .B2(n4001), .C1(n3881), .C2(n3880), .A(n4009), 
        .ZN(n3884) );
  OR2_X1 U4623 ( .A1(n4158), .A2(n3886), .ZN(n3883) );
  NAND2_X1 U4624 ( .A1(n4140), .A2(n4141), .ZN(n4013) );
  OR2_X1 U4625 ( .A1(n4029), .A2(n3892), .ZN(n3882) );
  AND2_X1 U4626 ( .A1(n4013), .A2(n3882), .ZN(n3908) );
  NAND2_X1 U4627 ( .A1(n3883), .A2(n3908), .ZN(n3889) );
  AOI21_X1 U4628 ( .B1(n4158), .B2(n3886), .A(n3885), .ZN(n3890) );
  NAND2_X1 U4629 ( .A1(n3890), .A2(n3935), .ZN(n4006) );
  OR2_X1 U4630 ( .A1(n3888), .A2(n3887), .ZN(n3891) );
  AOI21_X1 U4631 ( .B1(n3891), .B2(n3890), .A(n3889), .ZN(n4010) );
  OAI21_X1 U4632 ( .B1(n4006), .B2(n4173), .A(n4010), .ZN(n3894) );
  INV_X1 U4633 ( .A(n4140), .ZN(n3893) );
  INV_X1 U4634 ( .A(n3892), .ZN(n4381) );
  AOI22_X1 U4635 ( .A1(n3895), .A2(n3894), .B1(n3893), .B2(n4381), .ZN(n3896)
         );
  AOI211_X1 U4636 ( .C1(n3897), .C2(n3905), .A(n3904), .B(n3896), .ZN(n4021)
         );
  INV_X1 U4637 ( .A(n3898), .ZN(n3899) );
  NAND2_X1 U4638 ( .A1(n3899), .A2(n4188), .ZN(n4207) );
  XNOR2_X1 U4639 ( .A(n4032), .B(n4342), .ZN(n4333) );
  NOR3_X1 U4640 ( .A1(n4207), .A2(n4275), .A3(n4333), .ZN(n3940) );
  NAND2_X1 U4641 ( .A1(n3901), .A2(n3900), .ZN(n4228) );
  NAND2_X1 U4642 ( .A1(n3903), .A2(n3902), .ZN(n4309) );
  INV_X1 U4643 ( .A(n3904), .ZN(n3907) );
  INV_X1 U4644 ( .A(n3905), .ZN(n3906) );
  NAND2_X1 U4645 ( .A1(n3907), .A2(n3906), .ZN(n4014) );
  INV_X1 U4646 ( .A(n4014), .ZN(n3909) );
  NAND4_X1 U4647 ( .A1(n3910), .A2(n4309), .A3(n3909), .A4(n3908), .ZN(n3914)
         );
  NAND2_X1 U4648 ( .A1(n3912), .A2(n3911), .ZN(n3913) );
  NOR4_X1 U4649 ( .A1(n4228), .A2(n3915), .A3(n3914), .A4(n3913), .ZN(n3939)
         );
  INV_X1 U4650 ( .A(n3997), .ZN(n3916) );
  AND2_X1 U4651 ( .A1(n3916), .A2(n4248), .ZN(n4288) );
  NOR2_X1 U4652 ( .A1(n3918), .A2(n3917), .ZN(n3922) );
  AND4_X1 U4653 ( .A1(n2591), .A2(n4679), .A3(n3920), .A4(n3919), .ZN(n3921)
         );
  NAND4_X1 U4654 ( .A1(n4288), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(n3934)
         );
  INV_X1 U4655 ( .A(n2713), .ZN(n3924) );
  AND4_X1 U4656 ( .A1(n3927), .A2(n3926), .A3(n3925), .A4(n3924), .ZN(n3932)
         );
  INV_X1 U4657 ( .A(n4353), .ZN(n4361) );
  NOR2_X1 U4658 ( .A1(n3929), .A2(n3928), .ZN(n3930) );
  NAND4_X1 U4659 ( .A1(n3932), .A2(n4361), .A3(n3931), .A4(n3930), .ZN(n3933)
         );
  NOR2_X1 U4660 ( .A1(n3934), .A2(n3933), .ZN(n3938) );
  NAND2_X1 U4661 ( .A1(n3936), .A2(n3935), .ZN(n4191) );
  XNOR2_X1 U4662 ( .A(n4402), .B(n2253), .ZN(n4242) );
  INV_X1 U4663 ( .A(n4242), .ZN(n4251) );
  NOR2_X1 U4664 ( .A1(n4191), .A2(n4251), .ZN(n3937) );
  NAND4_X1 U4665 ( .A1(n3940), .A2(n3939), .A3(n3938), .A4(n3937), .ZN(n3942)
         );
  NOR4_X1 U4666 ( .A1(n3943), .A2(n3942), .A3(n4173), .A4(n3941), .ZN(n3944)
         );
  OR2_X1 U4667 ( .A1(n3944), .A2(n3948), .ZN(n4018) );
  INV_X1 U4668 ( .A(n3945), .ZN(n3949) );
  OAI211_X1 U4669 ( .C1(n3949), .C2(n3948), .A(n3947), .B(n3946), .ZN(n3951)
         );
  NAND3_X1 U4670 ( .A1(n3951), .A2(n3950), .A3(n2715), .ZN(n3954) );
  NAND3_X1 U4671 ( .A1(n3954), .A2(n3953), .A3(n3952), .ZN(n3957) );
  NAND3_X1 U4672 ( .A1(n3957), .A2(n3956), .A3(n3955), .ZN(n3965) );
  INV_X1 U4673 ( .A(n3958), .ZN(n3960) );
  NOR3_X1 U4674 ( .A1(n3972), .A2(n3960), .A3(n3959), .ZN(n3964) );
  INV_X1 U4675 ( .A(n3961), .ZN(n3963) );
  AOI211_X1 U4676 ( .C1(n3965), .C2(n3964), .A(n3963), .B(n3962), .ZN(n3970)
         );
  NAND2_X1 U4677 ( .A1(n3967), .A2(n3966), .ZN(n3974) );
  OAI211_X1 U4678 ( .C1(n3970), .C2(n3974), .A(n3969), .B(n3968), .ZN(n3980)
         );
  NOR2_X1 U4679 ( .A1(n3971), .A2(n3973), .ZN(n3979) );
  OR4_X1 U4680 ( .A1(n3975), .A2(n3974), .A3(n3973), .A4(n3972), .ZN(n3976) );
  AOI21_X1 U4681 ( .B1(n3977), .B2(n3976), .A(n3987), .ZN(n3978) );
  AOI21_X1 U4682 ( .B1(n3980), .B2(n3979), .A(n3978), .ZN(n3986) );
  INV_X1 U4683 ( .A(n3981), .ZN(n3985) );
  INV_X1 U4684 ( .A(n3982), .ZN(n3984) );
  NOR4_X1 U4685 ( .A1(n3986), .A2(n3985), .A3(n3984), .A4(n3983), .ZN(n3992)
         );
  AOI21_X1 U4686 ( .B1(n3989), .B2(n3988), .A(n3987), .ZN(n3991) );
  OAI21_X1 U4687 ( .B1(n3992), .B2(n3991), .A(n3990), .ZN(n3995) );
  AOI21_X1 U4688 ( .B1(n3995), .B2(n3994), .A(n3993), .ZN(n3996) );
  INV_X1 U4689 ( .A(n3996), .ZN(n3998) );
  AOI211_X1 U4690 ( .C1(n3998), .C2(n4247), .A(n3997), .B(n4246), .ZN(n4000)
         );
  NOR2_X1 U4691 ( .A1(n4000), .A2(n3999), .ZN(n4003) );
  OAI21_X1 U4692 ( .B1(n4003), .B2(n4002), .A(n4001), .ZN(n4004) );
  NAND2_X1 U4693 ( .A1(n4005), .A2(n4004), .ZN(n4008) );
  AOI211_X1 U4694 ( .C1(n4009), .C2(n4008), .A(n4007), .B(n4006), .ZN(n4012)
         );
  INV_X1 U4695 ( .A(n4010), .ZN(n4011) );
  NOR2_X1 U4696 ( .A1(n4012), .A2(n4011), .ZN(n4015) );
  OAI21_X1 U4697 ( .B1(n4015), .B2(n4014), .A(n4013), .ZN(n4017) );
  MUX2_X1 U4698 ( .A(n4018), .B(n4017), .S(n4016), .Z(n4019) );
  OAI21_X1 U4699 ( .B1(n4021), .B2(n4020), .A(n4019), .ZN(n4022) );
  XNOR2_X1 U4700 ( .A(n4022), .B(n4133), .ZN(n4028) );
  NAND2_X1 U4701 ( .A1(n4024), .A2(n4023), .ZN(n4025) );
  OAI211_X1 U4702 ( .C1(n4497), .C2(n4027), .A(n4025), .B(B_REG_SCAN_IN), .ZN(
        n4026) );
  OAI21_X1 U4703 ( .B1(n4028), .B2(n4027), .A(n4026), .ZN(U3239) );
  MUX2_X1 U4704 ( .A(DATAO_REG_31__SCAN_IN), .B(n4140), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4705 ( .A(DATAO_REG_30__SCAN_IN), .B(n4029), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4706 ( .A(DATAO_REG_29__SCAN_IN), .B(n4158), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4707 ( .A(DATAO_REG_28__SCAN_IN), .B(n4030), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4708 ( .A(DATAO_REG_27__SCAN_IN), .B(n4159), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4709 ( .A(n4385), .B(DATAO_REG_26__SCAN_IN), .S(n4031), .Z(U3576)
         );
  MUX2_X1 U4710 ( .A(DATAO_REG_25__SCAN_IN), .B(n4231), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4711 ( .A(n4210), .B(DATAO_REG_24__SCAN_IN), .S(n4031), .Z(U3574)
         );
  MUX2_X1 U4712 ( .A(n4402), .B(DATAO_REG_23__SCAN_IN), .S(n4031), .Z(U3573)
         );
  MUX2_X1 U4713 ( .A(n4291), .B(DATAO_REG_22__SCAN_IN), .S(n4031), .Z(U3572)
         );
  MUX2_X1 U4714 ( .A(n4433), .B(DATAO_REG_21__SCAN_IN), .S(n4031), .Z(U3571)
         );
  MUX2_X1 U4715 ( .A(DATAO_REG_20__SCAN_IN), .B(n4421), .S(U4043), .Z(U3570)
         );
  MUX2_X1 U4716 ( .A(DATAO_REG_19__SCAN_IN), .B(n4032), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4717 ( .A(DATAO_REG_18__SCAN_IN), .B(n4337), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4718 ( .A(DATAO_REG_17__SCAN_IN), .B(n4511), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4719 ( .A(DATAO_REG_16__SCAN_IN), .B(n4033), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4720 ( .A(DATAO_REG_15__SCAN_IN), .B(n4034), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4721 ( .A(DATAO_REG_14__SCAN_IN), .B(n4035), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4722 ( .A(DATAO_REG_13__SCAN_IN), .B(n4036), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4723 ( .A(DATAO_REG_12__SCAN_IN), .B(n4037), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4724 ( .A(DATAO_REG_11__SCAN_IN), .B(n4038), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4725 ( .A(DATAO_REG_10__SCAN_IN), .B(n4039), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4726 ( .A(DATAO_REG_9__SCAN_IN), .B(n4040), .S(U4043), .Z(U3559) );
  MUX2_X1 U4727 ( .A(DATAO_REG_8__SCAN_IN), .B(n4041), .S(U4043), .Z(U3558) );
  MUX2_X1 U4728 ( .A(DATAO_REG_7__SCAN_IN), .B(n4042), .S(U4043), .Z(U3557) );
  MUX2_X1 U4729 ( .A(DATAO_REG_6__SCAN_IN), .B(n4043), .S(U4043), .Z(U3556) );
  MUX2_X1 U4730 ( .A(DATAO_REG_5__SCAN_IN), .B(n4044), .S(U4043), .Z(U3555) );
  MUX2_X1 U4731 ( .A(DATAO_REG_4__SCAN_IN), .B(n2825), .S(U4043), .Z(U3554) );
  MUX2_X1 U4732 ( .A(DATAO_REG_3__SCAN_IN), .B(n2838), .S(U4043), .Z(U3553) );
  MUX2_X1 U4733 ( .A(DATAO_REG_2__SCAN_IN), .B(n2433), .S(U4043), .Z(U3552) );
  MUX2_X1 U4734 ( .A(DATAO_REG_1__SCAN_IN), .B(n2419), .S(U4043), .Z(U3551) );
  MUX2_X1 U4735 ( .A(DATAO_REG_0__SCAN_IN), .B(n2714), .S(U4043), .Z(U3550) );
  INV_X1 U4736 ( .A(n4637), .ZN(n4059) );
  NAND2_X1 U4737 ( .A1(n4059), .A2(n4045), .ZN(n4058) );
  OAI211_X1 U4738 ( .C1(n4048), .C2(n4047), .A(n4631), .B(n4046), .ZN(n4057)
         );
  INV_X1 U4739 ( .A(n4049), .ZN(n4054) );
  INV_X1 U4740 ( .A(n4050), .ZN(n4053) );
  INV_X1 U4741 ( .A(n4051), .ZN(n4052) );
  OAI211_X1 U4742 ( .C1(n4054), .C2(n4053), .A(n4586), .B(n4052), .ZN(n4056)
         );
  AOI22_X1 U4743 ( .A1(n4630), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4055) );
  NAND4_X1 U4744 ( .A1(n4058), .A2(n4057), .A3(n4056), .A4(n4055), .ZN(U3241)
         );
  NAND2_X1 U4745 ( .A1(n4059), .A2(n4503), .ZN(n4068) );
  OAI211_X1 U4746 ( .C1(REG1_REG_3__SCAN_IN), .C2(n4061), .A(n4631), .B(n4060), 
        .ZN(n4067) );
  AOI22_X1 U4747 ( .A1(n4630), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n4066) );
  XNOR2_X1 U4748 ( .A(n4063), .B(n4062), .ZN(n4064) );
  NAND2_X1 U4749 ( .A1(n4586), .A2(n4064), .ZN(n4065) );
  NAND4_X1 U4750 ( .A1(n4068), .A2(n4067), .A3(n4066), .A4(n4065), .ZN(U3243)
         );
  XNOR2_X1 U4751 ( .A(n4123), .B(REG1_REG_18__SCAN_IN), .ZN(n4124) );
  NAND2_X1 U4752 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4109), .ZN(n4084) );
  INV_X1 U4753 ( .A(n4109), .ZN(n4667) );
  AOI22_X1 U4754 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4109), .B1(n4667), .B2(
        n3522), .ZN(n4613) );
  NAND2_X1 U4755 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4105), .ZN(n4080) );
  INV_X1 U4756 ( .A(n4105), .ZN(n4670) );
  AOI22_X1 U4757 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4105), .B1(n4670), .B2(
        n3469), .ZN(n4594) );
  INV_X1 U4758 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4712) );
  AOI22_X1 U4759 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4090), .B1(n4672), .B2(
        n4712), .ZN(n4566) );
  NAND2_X1 U4760 ( .A1(n4091), .A2(REG1_REG_9__SCAN_IN), .ZN(n4075) );
  INV_X1 U4761 ( .A(n4091), .ZN(n4674) );
  AOI22_X1 U4762 ( .A1(n4091), .A2(REG1_REG_9__SCAN_IN), .B1(n3288), .B2(n4674), .ZN(n4545) );
  NOR2_X1 U4763 ( .A1(n4069), .A2(REG1_REG_7__SCAN_IN), .ZN(n4072) );
  INV_X1 U4764 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4070) );
  NAND2_X1 U4765 ( .A1(n4533), .A2(n4073), .ZN(n4074) );
  XOR2_X1 U4766 ( .A(n4533), .B(n4073), .Z(n4540) );
  NAND2_X1 U4767 ( .A1(REG1_REG_8__SCAN_IN), .A2(n4540), .ZN(n4539) );
  NAND2_X1 U4768 ( .A1(n4554), .A2(n4076), .ZN(n4077) );
  NAND2_X1 U4769 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4561), .ZN(n4560) );
  NAND2_X1 U4770 ( .A1(n4575), .A2(n4078), .ZN(n4079) );
  NAND2_X1 U4771 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4577), .ZN(n4576) );
  NAND2_X1 U4772 ( .A1(n4081), .A2(n4082), .ZN(n4083) );
  NAND2_X1 U4773 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4603), .ZN(n4602) );
  NAND2_X1 U4774 ( .A1(n4083), .A2(n4602), .ZN(n4612) );
  NAND2_X1 U4775 ( .A1(n4613), .A2(n4612), .ZN(n4611) );
  NAND2_X1 U4776 ( .A1(n4084), .A2(n4611), .ZN(n4086) );
  NOR2_X1 U4777 ( .A1(n4085), .A2(n4086), .ZN(n4087) );
  XNOR2_X1 U4778 ( .A(n4086), .B(n4085), .ZN(n4620) );
  NOR2_X1 U4779 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4620), .ZN(n4621) );
  AOI22_X1 U4780 ( .A1(n4112), .A2(n3628), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4665), .ZN(n4632) );
  NAND2_X1 U4781 ( .A1(n4088), .A2(n4631), .ZN(n4122) );
  NOR2_X1 U4782 ( .A1(n4112), .A2(REG2_REG_17__SCAN_IN), .ZN(n4089) );
  AOI21_X1 U4783 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4112), .A(n4089), .ZN(n4627) );
  NOR2_X1 U4784 ( .A1(n2551), .A2(n4670), .ZN(n4585) );
  NAND2_X1 U4785 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4090), .ZN(n4102) );
  AOI22_X1 U4786 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4090), .B1(n4672), .B2(
        n2526), .ZN(n4569) );
  NAND2_X1 U4787 ( .A1(n4091), .A2(REG2_REG_9__SCAN_IN), .ZN(n4098) );
  AOI22_X1 U4788 ( .A1(n4091), .A2(REG2_REG_9__SCAN_IN), .B1(n2505), .B2(n4674), .ZN(n4548) );
  NAND2_X1 U4789 ( .A1(n4533), .A2(n4096), .ZN(n4097) );
  XOR2_X1 U4790 ( .A(n4096), .B(n4533), .Z(n4535) );
  NAND2_X1 U4791 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4535), .ZN(n4534) );
  NAND2_X1 U4792 ( .A1(n4554), .A2(n4100), .ZN(n4101) );
  NAND2_X1 U4793 ( .A1(n4575), .A2(n4103), .ZN(n4104) );
  NOR2_X1 U4794 ( .A1(n4669), .A2(n4106), .ZN(n4107) );
  NAND2_X1 U4795 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4109), .ZN(n4108) );
  OAI21_X1 U4796 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4109), .A(n4108), .ZN(n4607) );
  NOR2_X1 U4797 ( .A1(n4608), .A2(n4607), .ZN(n4606) );
  NAND2_X1 U4798 ( .A1(n4110), .A2(n4666), .ZN(n4111) );
  NAND2_X1 U4799 ( .A1(n4627), .A2(n4625), .ZN(n4626) );
  INV_X1 U4800 ( .A(n4123), .ZN(n4500) );
  NOR2_X1 U4801 ( .A1(n4500), .A2(n4370), .ZN(n4113) );
  AOI21_X1 U4802 ( .B1(n4500), .B2(n4370), .A(n4113), .ZN(n4114) );
  INV_X1 U4803 ( .A(n4129), .ZN(n4120) );
  NAND2_X1 U4804 ( .A1(n4630), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4117) );
  OAI211_X1 U4805 ( .C1(n4637), .C2(n4123), .A(n4122), .B(n4121), .ZN(U3258)
         );
  AOI22_X1 U4806 ( .A1(n4125), .A2(n4124), .B1(n4500), .B2(
        REG1_REG_18__SCAN_IN), .ZN(n4128) );
  INV_X1 U4807 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4126) );
  MUX2_X1 U4808 ( .A(n4126), .B(REG1_REG_19__SCAN_IN), .S(n4499), .Z(n4127) );
  XNOR2_X1 U4809 ( .A(n4128), .B(n4127), .ZN(n4137) );
  MUX2_X1 U4810 ( .A(REG2_REG_19__SCAN_IN), .B(n4346), .S(n4499), .Z(n4130) );
  AOI21_X1 U4811 ( .B1(n4630), .B2(ADDR_REG_19__SCAN_IN), .A(n4131), .ZN(n4132) );
  OAI21_X1 U4812 ( .B1(n4637), .B2(n4133), .A(n4132), .ZN(n4134) );
  AOI21_X1 U4813 ( .B1(n4135), .B2(n4586), .A(n4134), .ZN(n4136) );
  OAI21_X1 U4814 ( .B1(n4138), .B2(n4137), .A(n4136), .ZN(U3259) );
  XNOR2_X1 U4815 ( .A(n4377), .B(n4141), .ZN(n4453) );
  NAND2_X1 U4816 ( .A1(n4140), .A2(n4139), .ZN(n4379) );
  OAI21_X1 U4817 ( .B1(n4141), .B2(n4334), .A(n4379), .ZN(n4450) );
  NOR2_X1 U4818 ( .A1(n4349), .A2(n4142), .ZN(n4143) );
  AOI21_X1 U4819 ( .B1(n4349), .B2(n4450), .A(n4143), .ZN(n4144) );
  OAI21_X1 U4820 ( .B1(n4453), .B2(n4343), .A(n4144), .ZN(U3260) );
  INV_X1 U4821 ( .A(n4145), .ZN(n4156) );
  INV_X1 U4822 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4146) );
  OAI22_X1 U4823 ( .A1(n4388), .A2(n4321), .B1(n4146), .B2(n4349), .ZN(n4147)
         );
  AOI21_X1 U4824 ( .B1(n4148), .B2(n4316), .A(n4147), .ZN(n4155) );
  INV_X1 U4825 ( .A(n4149), .ZN(n4153) );
  OAI22_X1 U4826 ( .A1(n4151), .A2(n4343), .B1(n4150), .B2(n4368), .ZN(n4152)
         );
  OAI21_X1 U4827 ( .B1(n4153), .B2(n4152), .A(n4349), .ZN(n4154) );
  OAI211_X1 U4828 ( .C1(n4156), .C2(n4374), .A(n4155), .B(n4154), .ZN(U3354)
         );
  INV_X1 U4829 ( .A(n4157), .ZN(n4167) );
  AOI22_X1 U4830 ( .A1(n4159), .A2(n4292), .B1(n4315), .B2(n4158), .ZN(n4162)
         );
  AOI22_X1 U4831 ( .A1(n4160), .A2(n4652), .B1(n4661), .B2(
        REG2_REG_28__SCAN_IN), .ZN(n4161) );
  OAI211_X1 U4832 ( .C1(n4163), .C2(n4297), .A(n4162), .B(n4161), .ZN(n4166)
         );
  NOR2_X1 U4833 ( .A1(n4164), .A2(n4661), .ZN(n4165) );
  AOI211_X1 U4834 ( .C1(n4655), .C2(n4167), .A(n4166), .B(n4165), .ZN(n4168)
         );
  OAI21_X1 U4835 ( .B1(n4169), .B2(n4374), .A(n4168), .ZN(U3262) );
  XNOR2_X1 U4836 ( .A(n4171), .B(n4170), .ZN(n4172) );
  NAND2_X1 U4837 ( .A1(n4172), .A2(n4366), .ZN(n4387) );
  XNOR2_X1 U4838 ( .A(n4174), .B(n4173), .ZN(n4390) );
  NAND2_X1 U4839 ( .A1(n4390), .A2(n4311), .ZN(n4186) );
  INV_X1 U4840 ( .A(n4175), .ZN(n4176) );
  OAI21_X1 U4841 ( .B1(n4196), .B2(n4182), .A(n4176), .ZN(n4460) );
  INV_X1 U4842 ( .A(n4460), .ZN(n4184) );
  OAI22_X1 U4843 ( .A1(n4388), .A2(n4177), .B1(n4213), .B2(n4321), .ZN(n4178)
         );
  INV_X1 U4844 ( .A(n4178), .ZN(n4181) );
  AOI22_X1 U4845 ( .A1(n4179), .A2(n4652), .B1(n4661), .B2(
        REG2_REG_27__SCAN_IN), .ZN(n4180) );
  OAI211_X1 U4846 ( .C1(n4182), .C2(n4297), .A(n4181), .B(n4180), .ZN(n4183)
         );
  AOI21_X1 U4847 ( .B1(n4184), .B2(n4655), .A(n4183), .ZN(n4185) );
  OAI211_X1 U4848 ( .C1(n4661), .C2(n4387), .A(n4186), .B(n4185), .ZN(U3263)
         );
  XNOR2_X1 U4849 ( .A(n4187), .B(n4191), .ZN(n4394) );
  INV_X1 U4850 ( .A(n4394), .ZN(n4205) );
  NAND2_X1 U4851 ( .A1(n4189), .A2(n4188), .ZN(n4190) );
  XOR2_X1 U4852 ( .A(n4191), .B(n4190), .Z(n4192) );
  NAND2_X1 U4853 ( .A1(n4192), .A2(n4366), .ZN(n4194) );
  AOI22_X1 U4854 ( .A1(n4231), .A2(n4420), .B1(n4197), .B2(n4430), .ZN(n4193)
         );
  OAI211_X1 U4855 ( .C1(n4195), .C2(n4424), .A(n4194), .B(n4193), .ZN(n4393)
         );
  INV_X1 U4856 ( .A(n4196), .ZN(n4199) );
  NAND2_X1 U4857 ( .A1(n4216), .A2(n4197), .ZN(n4198) );
  NAND2_X1 U4858 ( .A1(n4199), .A2(n4198), .ZN(n4464) );
  NOR2_X1 U4859 ( .A1(n4464), .A2(n4343), .ZN(n4203) );
  OAI22_X1 U4860 ( .A1(n4201), .A2(n4349), .B1(n4200), .B2(n4368), .ZN(n4202)
         );
  AOI211_X1 U4861 ( .C1(n4393), .C2(n4349), .A(n4203), .B(n4202), .ZN(n4204)
         );
  OAI21_X1 U4862 ( .B1(n4205), .B2(n4374), .A(n4204), .ZN(U3264) );
  XOR2_X1 U4863 ( .A(n4207), .B(n4206), .Z(n4398) );
  INV_X1 U4864 ( .A(n4398), .ZN(n4221) );
  XNOR2_X1 U4865 ( .A(n4208), .B(n4207), .ZN(n4209) );
  NAND2_X1 U4866 ( .A1(n4209), .A2(n4366), .ZN(n4212) );
  AOI22_X1 U4867 ( .A1(n4210), .A2(n4420), .B1(n4214), .B2(n4430), .ZN(n4211)
         );
  OAI211_X1 U4868 ( .C1(n4213), .C2(n4424), .A(n4212), .B(n4211), .ZN(n4397)
         );
  NAND2_X1 U4869 ( .A1(n4229), .A2(n4214), .ZN(n4215) );
  NAND2_X1 U4870 ( .A1(n4216), .A2(n4215), .ZN(n4468) );
  AOI22_X1 U4871 ( .A1(n4661), .A2(REG2_REG_25__SCAN_IN), .B1(n4217), .B2(
        n4652), .ZN(n4218) );
  OAI21_X1 U4872 ( .B1(n4468), .B2(n4343), .A(n4218), .ZN(n4219) );
  AOI21_X1 U4873 ( .B1(n4397), .B2(n4349), .A(n4219), .ZN(n4220) );
  OAI21_X1 U4874 ( .B1(n4221), .B2(n4374), .A(n4220), .ZN(U3265) );
  NAND2_X1 U4875 ( .A1(n4223), .A2(n4222), .ZN(n4225) );
  INV_X1 U4876 ( .A(n4228), .ZN(n4224) );
  XNOR2_X1 U4877 ( .A(n4225), .B(n4224), .ZN(n4226) );
  NAND2_X1 U4878 ( .A1(n4226), .A2(n4366), .ZN(n4404) );
  XNOR2_X1 U4879 ( .A(n4227), .B(n4228), .ZN(n4407) );
  NAND2_X1 U4880 ( .A1(n4407), .A2(n4311), .ZN(n4240) );
  INV_X1 U4881 ( .A(n4259), .ZN(n4230) );
  OAI21_X1 U4882 ( .B1(n4230), .B2(n4236), .A(n4229), .ZN(n4472) );
  INV_X1 U4883 ( .A(n4472), .ZN(n4238) );
  AOI22_X1 U4884 ( .A1(n4292), .A2(n4402), .B1(n4315), .B2(n4231), .ZN(n4235)
         );
  INV_X1 U4885 ( .A(n4232), .ZN(n4233) );
  AOI22_X1 U4886 ( .A1(n4661), .A2(REG2_REG_24__SCAN_IN), .B1(n4233), .B2(
        n4652), .ZN(n4234) );
  OAI211_X1 U4887 ( .C1(n4236), .C2(n4297), .A(n4235), .B(n4234), .ZN(n4237)
         );
  AOI21_X1 U4888 ( .B1(n4238), .B2(n4655), .A(n4237), .ZN(n4239) );
  OAI211_X1 U4889 ( .C1(n4661), .C2(n4404), .A(n4240), .B(n4239), .ZN(U3266)
         );
  XNOR2_X1 U4890 ( .A(n4241), .B(n4242), .ZN(n4411) );
  INV_X1 U4891 ( .A(n4411), .ZN(n4265) );
  AOI21_X1 U4892 ( .B1(n4304), .B2(n4247), .A(n4246), .ZN(n4285) );
  INV_X1 U4893 ( .A(n4248), .ZN(n4249) );
  AOI21_X1 U4894 ( .B1(n4285), .B2(n4288), .A(n4249), .ZN(n4276) );
  OAI21_X1 U4895 ( .B1(n4276), .B2(n4275), .A(n4250), .ZN(n4252) );
  XNOR2_X1 U4896 ( .A(n4252), .B(n4251), .ZN(n4256) );
  OAI22_X1 U4897 ( .A1(n4253), .A2(n4424), .B1(n4334), .B2(n4257), .ZN(n4254)
         );
  AOI21_X1 U4898 ( .B1(n4420), .B2(n4291), .A(n4254), .ZN(n4255) );
  OAI21_X1 U4899 ( .B1(n4256), .B2(n4339), .A(n4255), .ZN(n4410) );
  OR2_X1 U4900 ( .A1(n4269), .A2(n4257), .ZN(n4258) );
  NAND2_X1 U4901 ( .A1(n4259), .A2(n4258), .ZN(n4476) );
  NOR2_X1 U4902 ( .A1(n4476), .A2(n4343), .ZN(n4263) );
  OAI22_X1 U4903 ( .A1(n4349), .A2(n4261), .B1(n4260), .B2(n4368), .ZN(n4262)
         );
  AOI211_X1 U4904 ( .C1(n4410), .C2(n4349), .A(n4263), .B(n4262), .ZN(n4264)
         );
  OAI21_X1 U4905 ( .B1(n4265), .B2(n4374), .A(n4264), .ZN(U3267) );
  OAI21_X1 U4906 ( .B1(n4267), .B2(n4275), .A(n4266), .ZN(n4414) );
  NOR2_X1 U4907 ( .A1(n4289), .A2(n4279), .ZN(n4268) );
  OR2_X1 U4908 ( .A1(n4269), .A2(n4268), .ZN(n4480) );
  INV_X1 U4909 ( .A(n4480), .ZN(n4274) );
  INV_X1 U4910 ( .A(n4270), .ZN(n4271) );
  OAI22_X1 U4911 ( .A1(n4349), .A2(n4272), .B1(n4271), .B2(n4368), .ZN(n4273)
         );
  AOI21_X1 U4912 ( .B1(n4274), .B2(n4655), .A(n4273), .ZN(n4284) );
  XNOR2_X1 U4913 ( .A(n4276), .B(n4275), .ZN(n4277) );
  NAND2_X1 U4914 ( .A1(n4277), .A2(n4366), .ZN(n4282) );
  NAND2_X1 U4915 ( .A1(n4433), .A2(n4420), .ZN(n4278) );
  OAI21_X1 U4916 ( .B1(n4334), .B2(n4279), .A(n4278), .ZN(n4280) );
  AOI21_X1 U4917 ( .B1(n4402), .B2(n4432), .A(n4280), .ZN(n4281) );
  NAND2_X1 U4918 ( .A1(n4282), .A2(n4281), .ZN(n4415) );
  NAND2_X1 U4919 ( .A1(n4415), .A2(n4349), .ZN(n4283) );
  OAI211_X1 U4920 ( .C1(n4414), .C2(n4374), .A(n4284), .B(n4283), .ZN(U3268)
         );
  XNOR2_X1 U4921 ( .A(n4285), .B(n4288), .ZN(n4286) );
  NAND2_X1 U4922 ( .A1(n4286), .A2(n4366), .ZN(n4423) );
  XOR2_X1 U4923 ( .A(n4288), .B(n4287), .Z(n4427) );
  NAND2_X1 U4924 ( .A1(n4427), .A2(n4311), .ZN(n4302) );
  INV_X1 U4925 ( .A(n4289), .ZN(n4290) );
  OAI21_X1 U4926 ( .B1(n2260), .B2(n4298), .A(n4290), .ZN(n4484) );
  INV_X1 U4927 ( .A(n4484), .ZN(n4300) );
  AOI22_X1 U4928 ( .A1(n4292), .A2(n4421), .B1(n4315), .B2(n4291), .ZN(n4296)
         );
  INV_X1 U4929 ( .A(n4293), .ZN(n4294) );
  AOI22_X1 U4930 ( .A1(n4661), .A2(REG2_REG_21__SCAN_IN), .B1(n4294), .B2(
        n4652), .ZN(n4295) );
  OAI211_X1 U4931 ( .C1(n4298), .C2(n4297), .A(n4296), .B(n4295), .ZN(n4299)
         );
  AOI21_X1 U4932 ( .B1(n4300), .B2(n4655), .A(n4299), .ZN(n4301) );
  OAI211_X1 U4933 ( .C1(n4661), .C2(n4423), .A(n4302), .B(n4301), .ZN(U3269)
         );
  NAND2_X1 U4934 ( .A1(n4304), .A2(n4303), .ZN(n4305) );
  XNOR2_X1 U4935 ( .A(n4305), .B(n4309), .ZN(n4306) );
  NAND2_X1 U4936 ( .A1(n4306), .A2(n4366), .ZN(n4435) );
  AOI21_X1 U4937 ( .B1(n4326), .B2(n4308), .A(n4307), .ZN(n4310) );
  XNOR2_X1 U4938 ( .A(n4310), .B(n4309), .ZN(n4439) );
  NAND2_X1 U4939 ( .A1(n4439), .A2(n4311), .ZN(n4325) );
  INV_X1 U4940 ( .A(n4341), .ZN(n4314) );
  OAI21_X1 U4941 ( .B1(n4314), .B2(n4313), .A(n4312), .ZN(n4488) );
  INV_X1 U4942 ( .A(n4488), .ZN(n4323) );
  AOI22_X1 U4943 ( .A1(n4431), .A2(n4316), .B1(n4315), .B2(n4433), .ZN(n4320)
         );
  INV_X1 U4944 ( .A(n4317), .ZN(n4318) );
  AOI22_X1 U4945 ( .A1(n4661), .A2(REG2_REG_20__SCAN_IN), .B1(n4318), .B2(
        n4652), .ZN(n4319) );
  OAI211_X1 U4946 ( .C1(n4437), .C2(n4321), .A(n4320), .B(n4319), .ZN(n4322)
         );
  AOI21_X1 U4947 ( .B1(n4323), .B2(n4655), .A(n4322), .ZN(n4324) );
  OAI211_X1 U4948 ( .C1(n4661), .C2(n4435), .A(n4325), .B(n4324), .ZN(U3270)
         );
  XNOR2_X1 U4949 ( .A(n4326), .B(n4333), .ZN(n4444) );
  INV_X1 U4950 ( .A(n4444), .ZN(n4351) );
  NAND2_X1 U4951 ( .A1(n4328), .A2(n4327), .ZN(n4362) );
  INV_X1 U4952 ( .A(n4329), .ZN(n4331) );
  OAI21_X1 U4953 ( .B1(n4362), .B2(n4331), .A(n4330), .ZN(n4332) );
  XOR2_X1 U4954 ( .A(n4333), .B(n4332), .Z(n4340) );
  OAI22_X1 U4955 ( .A1(n4335), .A2(n4424), .B1(n4334), .B2(n4342), .ZN(n4336)
         );
  AOI21_X1 U4956 ( .B1(n4420), .B2(n4337), .A(n4336), .ZN(n4338) );
  OAI21_X1 U4957 ( .B1(n4340), .B2(n4339), .A(n4338), .ZN(n4442) );
  OAI21_X1 U4958 ( .B1(n4356), .B2(n4342), .A(n4341), .ZN(n4493) );
  NOR2_X1 U4959 ( .A1(n4493), .A2(n4343), .ZN(n4348) );
  INV_X1 U4960 ( .A(n4344), .ZN(n4345) );
  OAI22_X1 U4961 ( .A1(n4349), .A2(n4346), .B1(n4345), .B2(n4368), .ZN(n4347)
         );
  AOI211_X1 U4962 ( .C1(n4442), .C2(n4349), .A(n4348), .B(n4347), .ZN(n4350)
         );
  OAI21_X1 U4963 ( .B1(n4351), .B2(n4374), .A(n4350), .ZN(U3271) );
  OAI21_X1 U4964 ( .B1(n4354), .B2(n4353), .A(n4352), .ZN(n4355) );
  INV_X1 U4965 ( .A(n4355), .ZN(n4449) );
  INV_X1 U4966 ( .A(n4356), .ZN(n4358) );
  OAI211_X1 U4967 ( .C1(n4360), .C2(n4359), .A(n4358), .B(n4357), .ZN(n4447)
         );
  XNOR2_X1 U4968 ( .A(n4362), .B(n4361), .ZN(n4367) );
  AOI22_X1 U4969 ( .A1(n4511), .A2(n4420), .B1(n4363), .B2(n4430), .ZN(n4364)
         );
  OAI21_X1 U4970 ( .B1(n4437), .B2(n4424), .A(n4364), .ZN(n4365) );
  AOI21_X1 U4971 ( .B1(n4367), .B2(n4366), .A(n4365), .ZN(n4448) );
  OAI21_X1 U4972 ( .B1(n4499), .B2(n4447), .A(n4448), .ZN(n4372) );
  OAI22_X1 U4973 ( .A1(n4349), .A2(n4370), .B1(n4369), .B2(n4368), .ZN(n4371)
         );
  AOI21_X1 U4974 ( .B1(n4372), .B2(n4349), .A(n4371), .ZN(n4373) );
  OAI21_X1 U4975 ( .B1(n4449), .B2(n4374), .A(n4373), .ZN(U3272) );
  NAND2_X1 U4976 ( .A1(n4710), .A2(n4450), .ZN(n4376) );
  NAND2_X1 U4977 ( .A1(n4711), .A2(REG1_REG_31__SCAN_IN), .ZN(n4375) );
  OAI211_X1 U4978 ( .C1(n4453), .C2(n4446), .A(n4376), .B(n4375), .ZN(U3549)
         );
  AOI21_X1 U4979 ( .B1(n4381), .B2(n4378), .A(n4377), .ZN(n4523) );
  INV_X1 U4980 ( .A(n4523), .ZN(n4456) );
  INV_X1 U4981 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4382) );
  INV_X1 U4982 ( .A(n4379), .ZN(n4380) );
  AOI21_X1 U4983 ( .B1(n4381), .B2(n4430), .A(n4380), .ZN(n4525) );
  MUX2_X1 U4984 ( .A(n4382), .B(n4525), .S(n4710), .Z(n4383) );
  OAI21_X1 U4985 ( .B1(n4456), .B2(n4446), .A(n4383), .ZN(U3548) );
  INV_X1 U4986 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4391) );
  AOI22_X1 U4987 ( .A1(n4385), .A2(n4420), .B1(n4384), .B2(n4430), .ZN(n4386)
         );
  OAI211_X1 U4988 ( .C1(n4388), .C2(n4424), .A(n4387), .B(n4386), .ZN(n4389)
         );
  AOI21_X1 U4989 ( .B1(n4390), .B2(n4443), .A(n4389), .ZN(n4457) );
  MUX2_X1 U4990 ( .A(n4391), .B(n4457), .S(n4710), .Z(n4392) );
  OAI21_X1 U4991 ( .B1(n4446), .B2(n4460), .A(n4392), .ZN(U3545) );
  INV_X1 U4992 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4395) );
  AOI21_X1 U4993 ( .B1(n4394), .B2(n4443), .A(n4393), .ZN(n4461) );
  MUX2_X1 U4994 ( .A(n4395), .B(n4461), .S(n4710), .Z(n4396) );
  OAI21_X1 U4995 ( .B1(n4446), .B2(n4464), .A(n4396), .ZN(U3544) );
  INV_X1 U4996 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4399) );
  AOI21_X1 U4997 ( .B1(n4398), .B2(n4443), .A(n4397), .ZN(n4465) );
  MUX2_X1 U4998 ( .A(n4399), .B(n4465), .S(n4710), .Z(n4400) );
  OAI21_X1 U4999 ( .B1(n4446), .B2(n4468), .A(n4400), .ZN(U3543) );
  INV_X1 U5000 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4408) );
  AOI22_X1 U5001 ( .A1(n4402), .A2(n4420), .B1(n4401), .B2(n4430), .ZN(n4403)
         );
  OAI211_X1 U5002 ( .C1(n4405), .C2(n4424), .A(n4404), .B(n4403), .ZN(n4406)
         );
  AOI21_X1 U5003 ( .B1(n4407), .B2(n4443), .A(n4406), .ZN(n4469) );
  MUX2_X1 U5004 ( .A(n4408), .B(n4469), .S(n4710), .Z(n4409) );
  OAI21_X1 U5005 ( .B1(n4446), .B2(n4472), .A(n4409), .ZN(U3542) );
  INV_X1 U5006 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4412) );
  AOI21_X1 U5007 ( .B1(n4411), .B2(n4443), .A(n4410), .ZN(n4473) );
  MUX2_X1 U5008 ( .A(n4412), .B(n4473), .S(n4710), .Z(n4413) );
  OAI21_X1 U5009 ( .B1(n4446), .B2(n4476), .A(n4413), .ZN(U3541) );
  INV_X1 U5010 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4417) );
  INV_X1 U5011 ( .A(n4414), .ZN(n4416) );
  AOI21_X1 U5012 ( .B1(n4416), .B2(n4443), .A(n4415), .ZN(n4477) );
  MUX2_X1 U5013 ( .A(n4417), .B(n4477), .S(n4710), .Z(n4418) );
  OAI21_X1 U5014 ( .B1(n4446), .B2(n4480), .A(n4418), .ZN(U3540) );
  INV_X1 U5015 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4428) );
  AOI22_X1 U5016 ( .A1(n4421), .A2(n4420), .B1(n4430), .B2(n4419), .ZN(n4422)
         );
  OAI211_X1 U5017 ( .C1(n4425), .C2(n4424), .A(n4423), .B(n4422), .ZN(n4426)
         );
  AOI21_X1 U5018 ( .B1(n4427), .B2(n4443), .A(n4426), .ZN(n4481) );
  MUX2_X1 U5019 ( .A(n4428), .B(n4481), .S(n4710), .Z(n4429) );
  OAI21_X1 U5020 ( .B1(n4446), .B2(n4484), .A(n4429), .ZN(U3539) );
  INV_X1 U5021 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4440) );
  AOI22_X1 U5022 ( .A1(n4433), .A2(n4432), .B1(n4431), .B2(n4430), .ZN(n4434)
         );
  OAI211_X1 U5023 ( .C1(n4437), .C2(n4436), .A(n4435), .B(n4434), .ZN(n4438)
         );
  AOI21_X1 U5024 ( .B1(n4439), .B2(n4443), .A(n4438), .ZN(n4485) );
  MUX2_X1 U5025 ( .A(n4440), .B(n4485), .S(n4710), .Z(n4441) );
  OAI21_X1 U5026 ( .B1(n4446), .B2(n4488), .A(n4441), .ZN(U3538) );
  AOI21_X1 U5027 ( .B1(n4444), .B2(n4443), .A(n4442), .ZN(n4489) );
  MUX2_X1 U5028 ( .A(n4126), .B(n4489), .S(n4710), .Z(n4445) );
  OAI21_X1 U5029 ( .B1(n4446), .B2(n4493), .A(n4445), .ZN(U3537) );
  OAI211_X1 U5030 ( .C1(n4449), .C2(n4690), .A(n4448), .B(n4447), .ZN(n4494)
         );
  MUX2_X1 U5031 ( .A(REG1_REG_18__SCAN_IN), .B(n4494), .S(n4710), .Z(U3536) );
  NAND2_X1 U5032 ( .A1(n4703), .A2(n4450), .ZN(n4452) );
  NAND2_X1 U5033 ( .A1(n4701), .A2(REG0_REG_31__SCAN_IN), .ZN(n4451) );
  OAI211_X1 U5034 ( .C1(n4453), .C2(n4492), .A(n4452), .B(n4451), .ZN(U3517)
         );
  INV_X1 U5035 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4454) );
  MUX2_X1 U5036 ( .A(n4454), .B(n4525), .S(n4703), .Z(n4455) );
  OAI21_X1 U5037 ( .B1(n4456), .B2(n4492), .A(n4455), .ZN(U3516) );
  INV_X1 U5038 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4458) );
  MUX2_X1 U5039 ( .A(n4458), .B(n4457), .S(n4703), .Z(n4459) );
  OAI21_X1 U5040 ( .B1(n4460), .B2(n4492), .A(n4459), .ZN(U3513) );
  INV_X1 U5041 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4462) );
  MUX2_X1 U5042 ( .A(n4462), .B(n4461), .S(n4703), .Z(n4463) );
  OAI21_X1 U5043 ( .B1(n4464), .B2(n4492), .A(n4463), .ZN(U3512) );
  INV_X1 U5044 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4466) );
  MUX2_X1 U5045 ( .A(n4466), .B(n4465), .S(n4703), .Z(n4467) );
  OAI21_X1 U5046 ( .B1(n4468), .B2(n4492), .A(n4467), .ZN(U3511) );
  INV_X1 U5047 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4470) );
  MUX2_X1 U5048 ( .A(n4470), .B(n4469), .S(n4703), .Z(n4471) );
  OAI21_X1 U5049 ( .B1(n4472), .B2(n4492), .A(n4471), .ZN(U3510) );
  INV_X1 U5050 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4474) );
  MUX2_X1 U5051 ( .A(n4474), .B(n4473), .S(n4703), .Z(n4475) );
  OAI21_X1 U5052 ( .B1(n4476), .B2(n4492), .A(n4475), .ZN(U3509) );
  INV_X1 U5053 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4478) );
  MUX2_X1 U5054 ( .A(n4478), .B(n4477), .S(n4703), .Z(n4479) );
  OAI21_X1 U5055 ( .B1(n4480), .B2(n4492), .A(n4479), .ZN(U3508) );
  INV_X1 U5056 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4482) );
  MUX2_X1 U5057 ( .A(n4482), .B(n4481), .S(n4703), .Z(n4483) );
  OAI21_X1 U5058 ( .B1(n4484), .B2(n4492), .A(n4483), .ZN(U3507) );
  INV_X1 U5059 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4486) );
  MUX2_X1 U5060 ( .A(n4486), .B(n4485), .S(n4703), .Z(n4487) );
  OAI21_X1 U5061 ( .B1(n4488), .B2(n4492), .A(n4487), .ZN(U3506) );
  INV_X1 U5062 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4490) );
  MUX2_X1 U5063 ( .A(n4490), .B(n4489), .S(n4703), .Z(n4491) );
  OAI21_X1 U5064 ( .B1(n4493), .B2(n4492), .A(n4491), .ZN(U3505) );
  MUX2_X1 U5065 ( .A(REG0_REG_18__SCAN_IN), .B(n4494), .S(n4703), .Z(U3503) );
  MUX2_X1 U5066 ( .A(n4495), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5067 ( .A(DATAI_26_), .B(n4496), .S(STATE_REG_SCAN_IN), .Z(U3326)
         );
  MUX2_X1 U5068 ( .A(DATAI_24_), .B(n2778), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U5069 ( .A(DATAI_22_), .B(n4497), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5070 ( .A(DATAI_20_), .B(n4498), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5071 ( .A(DATAI_19_), .B(n4499), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5072 ( .A(DATAI_18_), .B(n4500), .S(STATE_REG_SCAN_IN), .Z(U3334)
         );
  MUX2_X1 U5073 ( .A(n4501), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5074 ( .A(n4502), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5075 ( .A(DATAI_3_), .B(n4503), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5076 ( .A(n4504), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  AOI22_X1 U5077 ( .A1(STATE_REG_SCAN_IN), .A2(n4505), .B1(n4847), .B2(U3149), 
        .ZN(U3324) );
  NOR2_X1 U5078 ( .A1(STATE_REG_SCAN_IN), .A2(n5057), .ZN(n4619) );
  OAI22_X1 U5079 ( .A1(n4509), .A2(n4508), .B1(n4507), .B2(n4506), .ZN(n4510)
         );
  AOI211_X1 U5080 ( .C1(n4512), .C2(n4511), .A(n4619), .B(n4510), .ZN(n4520)
         );
  AOI21_X1 U5081 ( .B1(n4514), .B2(n4513), .A(n3850), .ZN(n4515) );
  XOR2_X1 U5082 ( .A(n4516), .B(n4515), .Z(n4518) );
  NAND2_X1 U5083 ( .A1(n4518), .A2(n4517), .ZN(n4519) );
  OAI211_X1 U5084 ( .C1(n4522), .C2(n4521), .A(n4520), .B(n4519), .ZN(U3223)
         );
  AOI22_X1 U5085 ( .A1(n4523), .A2(n4655), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4661), .ZN(n4524) );
  OAI21_X1 U5086 ( .B1(n4661), .B2(n4525), .A(n4524), .ZN(U3261) );
  INV_X1 U5087 ( .A(n4528), .ZN(n4526) );
  OAI211_X1 U5088 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4527), .A(n4529), .B(n4526), 
        .ZN(n4532) );
  AOI22_X1 U5089 ( .A1(n4529), .A2(n4528), .B1(n4631), .B2(n2852), .ZN(n4531)
         );
  AOI22_X1 U5090 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4630), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4530) );
  OAI221_X1 U5091 ( .B1(IR_REG_0__SCAN_IN), .B2(n4532), .C1(n2262), .C2(n4531), 
        .A(n4530), .ZN(U3240) );
  INV_X1 U5092 ( .A(n4533), .ZN(n4676) );
  OAI211_X1 U5093 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4535), .A(n4586), .B(n4534), 
        .ZN(n4537) );
  NAND2_X1 U5094 ( .A1(n4537), .A2(n4536), .ZN(n4538) );
  AOI21_X1 U5095 ( .B1(n4630), .B2(ADDR_REG_8__SCAN_IN), .A(n4538), .ZN(n4542)
         );
  OAI211_X1 U5096 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4540), .A(n4631), .B(n4539), 
        .ZN(n4541) );
  OAI211_X1 U5097 ( .C1(n4637), .C2(n4676), .A(n4542), .B(n4541), .ZN(U3248)
         );
  OAI211_X1 U5098 ( .C1(n4545), .C2(n4544), .A(n4631), .B(n4543), .ZN(n4550)
         );
  OAI211_X1 U5099 ( .C1(n4548), .C2(n4547), .A(n4586), .B(n4546), .ZN(n4549)
         );
  OAI211_X1 U5100 ( .C1(n4637), .C2(n4674), .A(n4550), .B(n4549), .ZN(n4551)
         );
  AOI211_X1 U5101 ( .C1(n4630), .C2(ADDR_REG_9__SCAN_IN), .A(n4552), .B(n4551), 
        .ZN(n4553) );
  INV_X1 U5102 ( .A(n4553), .ZN(U3249) );
  OAI211_X1 U5103 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4556), .A(n4586), .B(n4555), .ZN(n4558) );
  NAND2_X1 U5104 ( .A1(n4558), .A2(n4557), .ZN(n4559) );
  AOI21_X1 U5105 ( .B1(n4630), .B2(ADDR_REG_10__SCAN_IN), .A(n4559), .ZN(n4563) );
  OAI211_X1 U5106 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4561), .A(n4631), .B(n4560), .ZN(n4562) );
  OAI211_X1 U5107 ( .C1(n4637), .C2(n4099), .A(n4563), .B(n4562), .ZN(U3250)
         );
  OAI211_X1 U5108 ( .C1(n4566), .C2(n4565), .A(n4631), .B(n4564), .ZN(n4571)
         );
  OAI211_X1 U5109 ( .C1(n4569), .C2(n4568), .A(n4586), .B(n4567), .ZN(n4570)
         );
  OAI211_X1 U5110 ( .C1(n4637), .C2(n4672), .A(n4571), .B(n4570), .ZN(n4572)
         );
  AOI211_X1 U5111 ( .C1(n4630), .C2(ADDR_REG_11__SCAN_IN), .A(n4573), .B(n4572), .ZN(n4574) );
  INV_X1 U5112 ( .A(n4574), .ZN(U3251) );
  INV_X1 U5113 ( .A(n4575), .ZN(n4671) );
  OAI211_X1 U5114 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4577), .A(n4631), .B(n4576), .ZN(n4581) );
  OAI211_X1 U5115 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4579), .A(n4586), .B(n4578), .ZN(n4580) );
  OAI211_X1 U5116 ( .C1(n4637), .C2(n4671), .A(n4581), .B(n4580), .ZN(n4582)
         );
  AOI211_X1 U5117 ( .C1(n4630), .C2(ADDR_REG_12__SCAN_IN), .A(n4583), .B(n4582), .ZN(n4584) );
  INV_X1 U5118 ( .A(n4584), .ZN(U3252) );
  AOI21_X1 U5119 ( .B1(n2551), .B2(n4670), .A(n4585), .ZN(n4589) );
  OAI21_X1 U5120 ( .B1(n4589), .B2(n4588), .A(n4586), .ZN(n4587) );
  AOI21_X1 U5121 ( .B1(n4589), .B2(n4588), .A(n4587), .ZN(n4591) );
  AOI211_X1 U5122 ( .C1(n4630), .C2(ADDR_REG_13__SCAN_IN), .A(n4591), .B(n4590), .ZN(n4596) );
  OAI211_X1 U5123 ( .C1(n4594), .C2(n4593), .A(n4631), .B(n4592), .ZN(n4595)
         );
  OAI211_X1 U5124 ( .C1(n4637), .C2(n4670), .A(n4596), .B(n4595), .ZN(U3253)
         );
  INV_X1 U5125 ( .A(n4597), .ZN(n4601) );
  AOI211_X1 U5126 ( .C1(n2560), .C2(n4599), .A(n4598), .B(n4624), .ZN(n4600)
         );
  AOI211_X1 U5127 ( .C1(n4630), .C2(ADDR_REG_14__SCAN_IN), .A(n4601), .B(n4600), .ZN(n4605) );
  OAI211_X1 U5128 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4603), .A(n4631), .B(n4602), .ZN(n4604) );
  OAI211_X1 U5129 ( .C1(n4637), .C2(n4669), .A(n4605), .B(n4604), .ZN(U3254)
         );
  AOI211_X1 U5130 ( .C1(n4608), .C2(n4607), .A(n4606), .B(n4624), .ZN(n4609)
         );
  AOI211_X1 U5131 ( .C1(n4630), .C2(ADDR_REG_15__SCAN_IN), .A(n4610), .B(n4609), .ZN(n4615) );
  OAI211_X1 U5132 ( .C1(n4613), .C2(n4612), .A(n4631), .B(n4611), .ZN(n4614)
         );
  OAI211_X1 U5133 ( .C1(n4637), .C2(n4667), .A(n4615), .B(n4614), .ZN(U3255)
         );
  AOI221_X1 U5134 ( .B1(n4617), .B2(n4616), .C1(n3476), .C2(n4616), .A(n4624), 
        .ZN(n4618) );
  AOI211_X1 U5135 ( .C1(n4630), .C2(ADDR_REG_16__SCAN_IN), .A(n4619), .B(n4618), .ZN(n4623) );
  OAI221_X1 U5136 ( .B1(n4621), .B2(REG1_REG_16__SCAN_IN), .C1(n4621), .C2(
        n4620), .A(n4631), .ZN(n4622) );
  OAI211_X1 U5137 ( .C1(n4637), .C2(n4666), .A(n4623), .B(n4622), .ZN(U3256)
         );
  AOI221_X1 U5138 ( .B1(n4627), .B2(n4626), .C1(n4626), .C2(n4625), .A(n4624), 
        .ZN(n4628) );
  AOI211_X1 U5139 ( .C1(n4630), .C2(ADDR_REG_17__SCAN_IN), .A(n4629), .B(n4628), .ZN(n4636) );
  OAI221_X1 U5140 ( .B1(n4634), .B2(n4633), .C1(n4634), .C2(n4632), .A(n4631), 
        .ZN(n4635) );
  OAI211_X1 U5141 ( .C1(n4637), .C2(n4665), .A(n4636), .B(n4635), .ZN(U3257)
         );
  AOI22_X1 U5142 ( .A1(n4638), .A2(n4652), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4661), .ZN(n4643) );
  INV_X1 U5143 ( .A(n4639), .ZN(n4640) );
  AOI22_X1 U5144 ( .A1(n4641), .A2(n4657), .B1(n4655), .B2(n4640), .ZN(n4642)
         );
  OAI211_X1 U5145 ( .C1(n4661), .C2(n4644), .A(n4643), .B(n4642), .ZN(U3280)
         );
  AOI22_X1 U5146 ( .A1(n4645), .A2(n4652), .B1(REG2_REG_8__SCAN_IN), .B2(n4661), .ZN(n4650) );
  INV_X1 U5147 ( .A(n4646), .ZN(n4647) );
  AOI22_X1 U5148 ( .A1(n4648), .A2(n4657), .B1(n4655), .B2(n4647), .ZN(n4649)
         );
  OAI211_X1 U5149 ( .C1(n4661), .C2(n4651), .A(n4650), .B(n4649), .ZN(U3282)
         );
  AOI22_X1 U5150 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4661), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4652), .ZN(n4659) );
  INV_X1 U5151 ( .A(n4653), .ZN(n4654) );
  AOI22_X1 U5152 ( .A1(n4657), .A2(n4656), .B1(n4655), .B2(n4654), .ZN(n4658)
         );
  OAI211_X1 U5153 ( .C1(n4661), .C2(n4660), .A(n4659), .B(n4658), .ZN(U3288)
         );
  AND2_X1 U5154 ( .A1(n4662), .A2(D_REG_31__SCAN_IN), .ZN(U3291) );
  INV_X1 U5155 ( .A(D_REG_30__SCAN_IN), .ZN(n5002) );
  NOR2_X1 U5156 ( .A1(n4663), .A2(n5002), .ZN(U3292) );
  INV_X1 U5157 ( .A(D_REG_29__SCAN_IN), .ZN(n5014) );
  NOR2_X1 U5158 ( .A1(n4663), .A2(n5014), .ZN(U3293) );
  INV_X1 U5159 ( .A(D_REG_28__SCAN_IN), .ZN(n5022) );
  NOR2_X1 U5160 ( .A1(n4663), .A2(n5022), .ZN(U3294) );
  INV_X1 U5161 ( .A(D_REG_27__SCAN_IN), .ZN(n4845) );
  NOR2_X1 U5162 ( .A1(n4663), .A2(n4845), .ZN(U3295) );
  INV_X1 U5163 ( .A(D_REG_26__SCAN_IN), .ZN(n4796) );
  NOR2_X1 U5164 ( .A1(n4663), .A2(n4796), .ZN(U3296) );
  INV_X1 U5165 ( .A(D_REG_25__SCAN_IN), .ZN(n4808) );
  NOR2_X1 U5166 ( .A1(n4663), .A2(n4808), .ZN(U3297) );
  INV_X1 U5167 ( .A(D_REG_24__SCAN_IN), .ZN(n4826) );
  NOR2_X1 U5168 ( .A1(n4663), .A2(n4826), .ZN(U3298) );
  INV_X1 U5169 ( .A(D_REG_23__SCAN_IN), .ZN(n5020) );
  NOR2_X1 U5170 ( .A1(n4663), .A2(n5020), .ZN(U3299) );
  INV_X1 U5171 ( .A(D_REG_22__SCAN_IN), .ZN(n4823) );
  NOR2_X1 U5172 ( .A1(n4663), .A2(n4823), .ZN(U3300) );
  INV_X1 U5173 ( .A(D_REG_21__SCAN_IN), .ZN(n5019) );
  NOR2_X1 U5174 ( .A1(n4663), .A2(n5019), .ZN(U3301) );
  INV_X1 U5175 ( .A(D_REG_20__SCAN_IN), .ZN(n5017) );
  NOR2_X1 U5176 ( .A1(n4663), .A2(n5017), .ZN(U3302) );
  AND2_X1 U5177 ( .A1(n4662), .A2(D_REG_19__SCAN_IN), .ZN(U3303) );
  INV_X1 U5178 ( .A(D_REG_18__SCAN_IN), .ZN(n5077) );
  NOR2_X1 U5179 ( .A1(n4663), .A2(n5077), .ZN(U3304) );
  AND2_X1 U5180 ( .A1(n4662), .A2(D_REG_17__SCAN_IN), .ZN(U3305) );
  INV_X1 U5181 ( .A(D_REG_16__SCAN_IN), .ZN(n5016) );
  NOR2_X1 U5182 ( .A1(n4663), .A2(n5016), .ZN(U3306) );
  AND2_X1 U5183 ( .A1(n4662), .A2(D_REG_15__SCAN_IN), .ZN(U3307) );
  AND2_X1 U5184 ( .A1(n4662), .A2(D_REG_14__SCAN_IN), .ZN(U3308) );
  INV_X1 U5185 ( .A(D_REG_13__SCAN_IN), .ZN(n5000) );
  NOR2_X1 U5186 ( .A1(n4663), .A2(n5000), .ZN(U3309) );
  AND2_X1 U5187 ( .A1(n4662), .A2(D_REG_12__SCAN_IN), .ZN(U3310) );
  INV_X1 U5188 ( .A(D_REG_11__SCAN_IN), .ZN(n5003) );
  NOR2_X1 U5189 ( .A1(n4663), .A2(n5003), .ZN(U3311) );
  INV_X1 U5190 ( .A(D_REG_10__SCAN_IN), .ZN(n4839) );
  NOR2_X1 U5191 ( .A1(n4663), .A2(n4839), .ZN(U3312) );
  AND2_X1 U5192 ( .A1(n4662), .A2(D_REG_9__SCAN_IN), .ZN(U3313) );
  AND2_X1 U5193 ( .A1(n4662), .A2(D_REG_8__SCAN_IN), .ZN(U3314) );
  AND2_X1 U5194 ( .A1(n4662), .A2(D_REG_7__SCAN_IN), .ZN(U3315) );
  INV_X1 U5195 ( .A(D_REG_6__SCAN_IN), .ZN(n5023) );
  NOR2_X1 U5196 ( .A1(n4663), .A2(n5023), .ZN(U3316) );
  INV_X1 U5197 ( .A(D_REG_5__SCAN_IN), .ZN(n5013) );
  NOR2_X1 U5198 ( .A1(n4663), .A2(n5013), .ZN(U3317) );
  INV_X1 U5199 ( .A(D_REG_4__SCAN_IN), .ZN(n4999) );
  NOR2_X1 U5200 ( .A1(n4663), .A2(n4999), .ZN(U3318) );
  AND2_X1 U5201 ( .A1(n4662), .A2(D_REG_3__SCAN_IN), .ZN(U3319) );
  INV_X1 U5202 ( .A(D_REG_2__SCAN_IN), .ZN(n4849) );
  NOR2_X1 U5203 ( .A1(n4663), .A2(n4849), .ZN(U3320) );
  INV_X1 U5204 ( .A(DATAI_23_), .ZN(n5036) );
  AOI21_X1 U5205 ( .B1(U3149), .B2(n5036), .A(n4664), .ZN(U3329) );
  AOI22_X1 U5206 ( .A1(STATE_REG_SCAN_IN), .A2(n4665), .B1(n2387), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5207 ( .A1(STATE_REG_SCAN_IN), .A2(n4666), .B1(n5053), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5208 ( .A(DATAI_15_), .ZN(n5044) );
  AOI22_X1 U5209 ( .A1(STATE_REG_SCAN_IN), .A2(n4667), .B1(n5044), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U5210 ( .A1(STATE_REG_SCAN_IN), .A2(n4669), .B1(n4668), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5211 ( .A(DATAI_13_), .ZN(n4811) );
  AOI22_X1 U5212 ( .A1(STATE_REG_SCAN_IN), .A2(n4670), .B1(n4811), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5213 ( .A(DATAI_12_), .ZN(n5034) );
  AOI22_X1 U5214 ( .A1(STATE_REG_SCAN_IN), .A2(n4671), .B1(n5034), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5215 ( .A1(STATE_REG_SCAN_IN), .A2(n4672), .B1(n2534), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5216 ( .A(DATAI_10_), .ZN(n4871) );
  AOI22_X1 U5217 ( .A1(STATE_REG_SCAN_IN), .A2(n4099), .B1(n4871), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5218 ( .A(DATAI_9_), .ZN(n4673) );
  AOI22_X1 U5219 ( .A1(STATE_REG_SCAN_IN), .A2(n4674), .B1(n4673), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5220 ( .A(DATAI_8_), .ZN(n4675) );
  AOI22_X1 U5221 ( .A1(STATE_REG_SCAN_IN), .A2(n4676), .B1(n4675), .B2(U3149), 
        .ZN(U3344) );
  OAI211_X1 U5222 ( .C1(n4679), .C2(n4682), .A(n4678), .B(n4677), .ZN(n4680)
         );
  INV_X1 U5223 ( .A(n4680), .ZN(n4704) );
  INV_X1 U5224 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4983) );
  AOI22_X1 U5225 ( .A1(n4703), .A2(n4704), .B1(n4983), .B2(n4701), .ZN(U3467)
         );
  OAI22_X1 U5226 ( .A1(n4683), .A2(n4682), .B1(n4695), .B2(n4681), .ZN(n4684)
         );
  NOR2_X1 U5227 ( .A1(n4685), .A2(n4684), .ZN(n4706) );
  INV_X1 U5228 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4982) );
  AOI22_X1 U5229 ( .A1(n4703), .A2(n4706), .B1(n4982), .B2(n4701), .ZN(U3469)
         );
  INV_X1 U5230 ( .A(n4686), .ZN(n4688) );
  AOI211_X1 U5231 ( .C1(n4689), .C2(n4700), .A(n4688), .B(n4687), .ZN(n4708)
         );
  INV_X1 U5232 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4988) );
  AOI22_X1 U5233 ( .A1(n4703), .A2(n4708), .B1(n4988), .B2(n4701), .ZN(U3475)
         );
  NOR2_X1 U5234 ( .A1(n4691), .A2(n4690), .ZN(n4694) );
  AOI211_X1 U5235 ( .C1(n4694), .C2(n3204), .A(n4693), .B(n4692), .ZN(n4709)
         );
  INV_X1 U5236 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4742) );
  AOI22_X1 U5237 ( .A1(n4703), .A2(n4709), .B1(n4742), .B2(n4701), .ZN(U3481)
         );
  NOR2_X1 U5238 ( .A1(n4696), .A2(n4695), .ZN(n4698) );
  AOI211_X1 U5239 ( .C1(n4700), .C2(n4699), .A(n4698), .B(n4697), .ZN(n4713)
         );
  INV_X1 U5240 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4702) );
  AOI22_X1 U5241 ( .A1(n4703), .A2(n4713), .B1(n4702), .B2(n4701), .ZN(U3489)
         );
  AOI22_X1 U5242 ( .A1(n4710), .A2(n4704), .B1(n2852), .B2(n4711), .ZN(U3518)
         );
  INV_X1 U5243 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4705) );
  AOI22_X1 U5244 ( .A1(n4710), .A2(n4706), .B1(n4705), .B2(n4711), .ZN(U3519)
         );
  INV_X1 U5245 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4707) );
  AOI22_X1 U5246 ( .A1(n4710), .A2(n4708), .B1(n4707), .B2(n4711), .ZN(U3522)
         );
  AOI22_X1 U5247 ( .A1(n4710), .A2(n4709), .B1(n4070), .B2(n4711), .ZN(U3525)
         );
  AOI22_X1 U5248 ( .A1(n4710), .A2(n4713), .B1(n4712), .B2(n4711), .ZN(U3529)
         );
  OAI22_X1 U5249 ( .A1(DATAI_1_), .A2(keyinput_g30), .B1(DATAI_30_), .B2(
        keyinput_g1), .ZN(n4714) );
  AOI221_X1 U5250 ( .B1(DATAI_1_), .B2(keyinput_g30), .C1(keyinput_g1), .C2(
        DATAI_30_), .A(n4714), .ZN(n4721) );
  OAI22_X1 U5251 ( .A1(D_REG_19__SCAN_IN), .A2(keyinput_g106), .B1(
        keyinput_g14), .B2(DATAI_17_), .ZN(n4715) );
  AOI221_X1 U5252 ( .B1(D_REG_19__SCAN_IN), .B2(keyinput_g106), .C1(DATAI_17_), 
        .C2(keyinput_g14), .A(n4715), .ZN(n4720) );
  OAI22_X1 U5253 ( .A1(D_REG_12__SCAN_IN), .A2(keyinput_g99), .B1(
        D_REG_0__SCAN_IN), .B2(keyinput_g87), .ZN(n4716) );
  AOI221_X1 U5254 ( .B1(D_REG_12__SCAN_IN), .B2(keyinput_g99), .C1(
        keyinput_g87), .C2(D_REG_0__SCAN_IN), .A(n4716), .ZN(n4719) );
  OAI22_X1 U5255 ( .A1(D_REG_1__SCAN_IN), .A2(keyinput_g88), .B1(keyinput_g12), 
        .B2(DATAI_19_), .ZN(n4717) );
  AOI221_X1 U5256 ( .B1(D_REG_1__SCAN_IN), .B2(keyinput_g88), .C1(DATAI_19_), 
        .C2(keyinput_g12), .A(n4717), .ZN(n4718) );
  NAND4_X1 U5257 ( .A1(n4721), .A2(n4720), .A3(n4719), .A4(n4718), .ZN(n4751)
         );
  OAI22_X1 U5258 ( .A1(IR_REG_0__SCAN_IN), .A2(keyinput_g55), .B1(
        D_REG_15__SCAN_IN), .B2(keyinput_g102), .ZN(n4722) );
  AOI221_X1 U5259 ( .B1(IR_REG_0__SCAN_IN), .B2(keyinput_g55), .C1(
        keyinput_g102), .C2(D_REG_15__SCAN_IN), .A(n4722), .ZN(n4729) );
  OAI22_X1 U5260 ( .A1(IR_REG_18__SCAN_IN), .A2(keyinput_g73), .B1(
        keyinput_g96), .B2(D_REG_9__SCAN_IN), .ZN(n4723) );
  AOI221_X1 U5261 ( .B1(IR_REG_18__SCAN_IN), .B2(keyinput_g73), .C1(
        D_REG_9__SCAN_IN), .C2(keyinput_g96), .A(n4723), .ZN(n4728) );
  OAI22_X1 U5262 ( .A1(IR_REG_12__SCAN_IN), .A2(keyinput_g67), .B1(
        keyinput_g22), .B2(DATAI_9_), .ZN(n4724) );
  AOI221_X1 U5263 ( .B1(IR_REG_12__SCAN_IN), .B2(keyinput_g67), .C1(DATAI_9_), 
        .C2(keyinput_g22), .A(n4724), .ZN(n4727) );
  OAI22_X1 U5264 ( .A1(IR_REG_21__SCAN_IN), .A2(keyinput_g76), .B1(
        keyinput_g107), .B2(D_REG_20__SCAN_IN), .ZN(n4725) );
  AOI221_X1 U5265 ( .B1(IR_REG_21__SCAN_IN), .B2(keyinput_g76), .C1(
        D_REG_20__SCAN_IN), .C2(keyinput_g107), .A(n4725), .ZN(n4726) );
  NAND4_X1 U5266 ( .A1(n4729), .A2(n4728), .A3(n4727), .A4(n4726), .ZN(n4750)
         );
  OAI22_X1 U5267 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput_g34), .B1(DATAI_21_), .B2(keyinput_g10), .ZN(n4730) );
  AOI221_X1 U5268 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_g34), .C1(
        keyinput_g10), .C2(DATAI_21_), .A(n4730), .ZN(n4737) );
  OAI22_X1 U5269 ( .A1(D_REG_31__SCAN_IN), .A2(keyinput_g118), .B1(
        keyinput_g82), .B2(IR_REG_27__SCAN_IN), .ZN(n4731) );
  AOI221_X1 U5270 ( .B1(D_REG_31__SCAN_IN), .B2(keyinput_g118), .C1(
        IR_REG_27__SCAN_IN), .C2(keyinput_g82), .A(n4731), .ZN(n4736) );
  OAI22_X1 U5271 ( .A1(IR_REG_3__SCAN_IN), .A2(keyinput_g58), .B1(keyinput_g95), .B2(D_REG_8__SCAN_IN), .ZN(n4732) );
  AOI221_X1 U5272 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput_g58), .C1(
        D_REG_8__SCAN_IN), .C2(keyinput_g95), .A(n4732), .ZN(n4735) );
  OAI22_X1 U5273 ( .A1(D_REG_5__SCAN_IN), .A2(keyinput_g92), .B1(
        REG3_REG_17__SCAN_IN), .B2(keyinput_g48), .ZN(n4733) );
  AOI221_X1 U5274 ( .B1(D_REG_5__SCAN_IN), .B2(keyinput_g92), .C1(keyinput_g48), .C2(REG3_REG_17__SCAN_IN), .A(n4733), .ZN(n4734) );
  NAND4_X1 U5275 ( .A1(n4737), .A2(n4736), .A3(n4735), .A4(n4734), .ZN(n4749)
         );
  OAI22_X1 U5276 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_g42), .B1(
        keyinput_g0), .B2(DATAI_31_), .ZN(n4738) );
  AOI221_X1 U5277 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_g42), .C1(DATAI_31_), .C2(keyinput_g0), .A(n4738), .ZN(n4747) );
  OAI22_X1 U5278 ( .A1(D_REG_17__SCAN_IN), .A2(keyinput_g104), .B1(
        D_REG_3__SCAN_IN), .B2(keyinput_g90), .ZN(n4739) );
  AOI221_X1 U5279 ( .B1(D_REG_17__SCAN_IN), .B2(keyinput_g104), .C1(
        keyinput_g90), .C2(D_REG_3__SCAN_IN), .A(n4739), .ZN(n4746) );
  OAI22_X1 U5280 ( .A1(IR_REG_29__SCAN_IN), .A2(keyinput_g84), .B1(DATAI_8_), 
        .B2(keyinput_g23), .ZN(n4740) );
  AOI221_X1 U5281 ( .B1(IR_REG_29__SCAN_IN), .B2(keyinput_g84), .C1(
        keyinput_g23), .C2(DATAI_8_), .A(n4740), .ZN(n4745) );
  OAI22_X1 U5282 ( .A1(n4743), .A2(keyinput_g35), .B1(n4742), .B2(
        keyinput_g126), .ZN(n4741) );
  AOI221_X1 U5283 ( .B1(n4743), .B2(keyinput_g35), .C1(keyinput_g126), .C2(
        n4742), .A(n4741), .ZN(n4744) );
  NAND4_X1 U5284 ( .A1(n4747), .A2(n4746), .A3(n4745), .A4(n4744), .ZN(n4748)
         );
  NOR4_X1 U5285 ( .A1(n4751), .A2(n4750), .A3(n4749), .A4(n4748), .ZN(n5082)
         );
  OAI22_X1 U5286 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput_g37), .B1(
        REG3_REG_8__SCAN_IN), .B2(keyinput_g41), .ZN(n4752) );
  AOI221_X1 U5287 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput_g37), .C1(
        keyinput_g41), .C2(REG3_REG_8__SCAN_IN), .A(n4752), .ZN(n4759) );
  OAI22_X1 U5288 ( .A1(D_REG_14__SCAN_IN), .A2(keyinput_g101), .B1(
        keyinput_g53), .B2(REG3_REG_20__SCAN_IN), .ZN(n4753) );
  AOI221_X1 U5289 ( .B1(D_REG_14__SCAN_IN), .B2(keyinput_g101), .C1(
        REG3_REG_20__SCAN_IN), .C2(keyinput_g53), .A(n4753), .ZN(n4758) );
  OAI22_X1 U5290 ( .A1(IR_REG_31__SCAN_IN), .A2(keyinput_g86), .B1(DATAI_14_), 
        .B2(keyinput_g17), .ZN(n4754) );
  AOI221_X1 U5291 ( .B1(IR_REG_31__SCAN_IN), .B2(keyinput_g86), .C1(
        keyinput_g17), .C2(DATAI_14_), .A(n4754), .ZN(n4757) );
  OAI22_X1 U5292 ( .A1(REG3_REG_13__SCAN_IN), .A2(keyinput_g54), .B1(
        keyinput_g125), .B2(REG0_REG_6__SCAN_IN), .ZN(n4755) );
  AOI221_X1 U5293 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_g54), .C1(
        REG0_REG_6__SCAN_IN), .C2(keyinput_g125), .A(n4755), .ZN(n4756) );
  NAND4_X1 U5294 ( .A1(n4759), .A2(n4758), .A3(n4757), .A4(n4756), .ZN(n4889)
         );
  OAI22_X1 U5295 ( .A1(D_REG_7__SCAN_IN), .A2(keyinput_g94), .B1(
        REG0_REG_1__SCAN_IN), .B2(keyinput_g120), .ZN(n4760) );
  AOI221_X1 U5296 ( .B1(D_REG_7__SCAN_IN), .B2(keyinput_g94), .C1(
        keyinput_g120), .C2(REG0_REG_1__SCAN_IN), .A(n4760), .ZN(n4785) );
  OAI22_X1 U5297 ( .A1(IR_REG_22__SCAN_IN), .A2(keyinput_g77), .B1(
        REG3_REG_16__SCAN_IN), .B2(keyinput_g46), .ZN(n4761) );
  AOI221_X1 U5298 ( .B1(IR_REG_22__SCAN_IN), .B2(keyinput_g77), .C1(
        keyinput_g46), .C2(REG3_REG_16__SCAN_IN), .A(n4761), .ZN(n4764) );
  OAI22_X1 U5299 ( .A1(IR_REG_20__SCAN_IN), .A2(keyinput_g75), .B1(
        keyinput_g56), .B2(IR_REG_1__SCAN_IN), .ZN(n4762) );
  AOI221_X1 U5300 ( .B1(IR_REG_20__SCAN_IN), .B2(keyinput_g75), .C1(
        IR_REG_1__SCAN_IN), .C2(keyinput_g56), .A(n4762), .ZN(n4763) );
  OAI211_X1 U5301 ( .C1(n2601), .C2(keyinput_g72), .A(n4764), .B(n4763), .ZN(
        n4765) );
  AOI21_X1 U5302 ( .B1(n2601), .B2(keyinput_g72), .A(n4765), .ZN(n4784) );
  AOI22_X1 U5303 ( .A1(REG0_REG_2__SCAN_IN), .A2(keyinput_g121), .B1(
        IR_REG_2__SCAN_IN), .B2(keyinput_g57), .ZN(n4766) );
  OAI221_X1 U5304 ( .B1(REG0_REG_2__SCAN_IN), .B2(keyinput_g121), .C1(
        IR_REG_2__SCAN_IN), .C2(keyinput_g57), .A(n4766), .ZN(n4773) );
  AOI22_X1 U5305 ( .A1(REG0_REG_8__SCAN_IN), .A2(keyinput_g127), .B1(
        IR_REG_8__SCAN_IN), .B2(keyinput_g63), .ZN(n4767) );
  OAI221_X1 U5306 ( .B1(REG0_REG_8__SCAN_IN), .B2(keyinput_g127), .C1(
        IR_REG_8__SCAN_IN), .C2(keyinput_g63), .A(n4767), .ZN(n4772) );
  AOI22_X1 U5307 ( .A1(D_REG_6__SCAN_IN), .A2(keyinput_g93), .B1(
        D_REG_30__SCAN_IN), .B2(keyinput_g117), .ZN(n4768) );
  OAI221_X1 U5308 ( .B1(D_REG_6__SCAN_IN), .B2(keyinput_g93), .C1(
        D_REG_30__SCAN_IN), .C2(keyinput_g117), .A(n4768), .ZN(n4771) );
  AOI22_X1 U5309 ( .A1(DATAI_23_), .A2(keyinput_g8), .B1(D_REG_28__SCAN_IN), 
        .B2(keyinput_g115), .ZN(n4769) );
  OAI221_X1 U5310 ( .B1(DATAI_23_), .B2(keyinput_g8), .C1(D_REG_28__SCAN_IN), 
        .C2(keyinput_g115), .A(n4769), .ZN(n4770) );
  NOR4_X1 U5311 ( .A1(n4773), .A2(n4772), .A3(n4771), .A4(n4770), .ZN(n4783)
         );
  AOI22_X1 U5312 ( .A1(DATAI_15_), .A2(keyinput_g16), .B1(DATAI_22_), .B2(
        keyinput_g9), .ZN(n4774) );
  OAI221_X1 U5313 ( .B1(DATAI_15_), .B2(keyinput_g16), .C1(DATAI_22_), .C2(
        keyinput_g9), .A(n4774), .ZN(n4781) );
  AOI22_X1 U5314 ( .A1(DATAI_2_), .A2(keyinput_g29), .B1(REG3_REG_23__SCAN_IN), 
        .B2(keyinput_g36), .ZN(n4775) );
  OAI221_X1 U5315 ( .B1(DATAI_2_), .B2(keyinput_g29), .C1(REG3_REG_23__SCAN_IN), .C2(keyinput_g36), .A(n4775), .ZN(n4780) );
  AOI22_X1 U5316 ( .A1(DATAI_3_), .A2(keyinput_g28), .B1(DATAI_16_), .B2(
        keyinput_g15), .ZN(n4776) );
  OAI221_X1 U5317 ( .B1(DATAI_3_), .B2(keyinput_g28), .C1(DATAI_16_), .C2(
        keyinput_g15), .A(n4776), .ZN(n4779) );
  AOI22_X1 U5318 ( .A1(DATAI_20_), .A2(keyinput_g11), .B1(IR_REG_5__SCAN_IN), 
        .B2(keyinput_g60), .ZN(n4777) );
  OAI221_X1 U5319 ( .B1(DATAI_20_), .B2(keyinput_g11), .C1(IR_REG_5__SCAN_IN), 
        .C2(keyinput_g60), .A(n4777), .ZN(n4778) );
  NOR4_X1 U5320 ( .A1(n4781), .A2(n4780), .A3(n4779), .A4(n4778), .ZN(n4782)
         );
  NAND4_X1 U5321 ( .A1(n4785), .A2(n4784), .A3(n4783), .A4(n4782), .ZN(n4888)
         );
  AOI22_X1 U5322 ( .A1(n2485), .A2(keyinput_g61), .B1(keyinput_g108), .B2(
        n5019), .ZN(n4786) );
  OAI221_X1 U5323 ( .B1(n2485), .B2(keyinput_g61), .C1(n5019), .C2(
        keyinput_g108), .A(n4786), .ZN(n4794) );
  AOI22_X1 U5324 ( .A1(n2680), .A2(keyinput_g4), .B1(n3739), .B2(keyinput_g85), 
        .ZN(n4787) );
  OAI221_X1 U5325 ( .B1(n2680), .B2(keyinput_g4), .C1(n3739), .C2(keyinput_g85), .A(n4787), .ZN(n4793) );
  XOR2_X1 U5326 ( .A(n2364), .B(keyinput_g69), .Z(n4791) );
  XOR2_X1 U5327 ( .A(n4985), .B(keyinput_g33), .Z(n4790) );
  XNOR2_X1 U5328 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_g80), .ZN(n4789) );
  XNOR2_X1 U5329 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_g78), .ZN(n4788) );
  NAND4_X1 U5330 ( .A1(n4791), .A2(n4790), .A3(n4789), .A4(n4788), .ZN(n4792)
         );
  NOR3_X1 U5331 ( .A1(n4794), .A2(n4793), .A3(n4792), .ZN(n4834) );
  INV_X1 U5332 ( .A(DATAI_26_), .ZN(n4797) );
  AOI22_X1 U5333 ( .A1(n4797), .A2(keyinput_g5), .B1(n4796), .B2(keyinput_g113), .ZN(n4795) );
  OAI221_X1 U5334 ( .B1(n4797), .B2(keyinput_g5), .C1(n4796), .C2(
        keyinput_g113), .A(n4795), .ZN(n4806) );
  INV_X1 U5335 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4799) );
  AOI22_X1 U5336 ( .A1(n2531), .A2(keyinput_g65), .B1(keyinput_g49), .B2(n4799), .ZN(n4798) );
  OAI221_X1 U5337 ( .B1(n2531), .B2(keyinput_g65), .C1(n4799), .C2(
        keyinput_g49), .A(n4798), .ZN(n4805) );
  XNOR2_X1 U5338 ( .A(n5020), .B(keyinput_g110), .ZN(n4804) );
  XOR2_X1 U5339 ( .A(n2502), .B(keyinput_g51), .Z(n4802) );
  XNOR2_X1 U5340 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_g50), .ZN(n4801) );
  XNOR2_X1 U5341 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_g38), .ZN(n4800) );
  NAND3_X1 U5342 ( .A1(n4802), .A2(n4801), .A3(n4800), .ZN(n4803) );
  NOR4_X1 U5343 ( .A1(n4806), .A2(n4805), .A3(n4804), .A4(n4803), .ZN(n4833)
         );
  AOI22_X1 U5344 ( .A1(n4808), .A2(keyinput_g112), .B1(keyinput_g24), .B2(
        n2487), .ZN(n4807) );
  OAI221_X1 U5345 ( .B1(n4808), .B2(keyinput_g112), .C1(n2487), .C2(
        keyinput_g24), .A(n4807), .ZN(n4817) );
  AOI22_X1 U5346 ( .A1(n5016), .A2(keyinput_g103), .B1(keyinput_g47), .B2(
        n2458), .ZN(n4809) );
  OAI221_X1 U5347 ( .B1(n5016), .B2(keyinput_g103), .C1(n2458), .C2(
        keyinput_g47), .A(n4809), .ZN(n4816) );
  AOI22_X1 U5348 ( .A1(n2257), .A2(keyinput_g31), .B1(n4811), .B2(keyinput_g18), .ZN(n4810) );
  OAI221_X1 U5349 ( .B1(n2257), .B2(keyinput_g31), .C1(n4811), .C2(
        keyinput_g18), .A(n4810), .ZN(n4815) );
  XNOR2_X1 U5350 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_g83), .ZN(n4813) );
  XNOR2_X1 U5351 ( .A(STATE_REG_SCAN_IN), .B(keyinput_g32), .ZN(n4812) );
  NAND2_X1 U5352 ( .A1(n4813), .A2(n4812), .ZN(n4814) );
  NOR4_X1 U5353 ( .A1(n4817), .A2(n4816), .A3(n4815), .A4(n4814), .ZN(n4832)
         );
  AOI22_X1 U5354 ( .A1(n4819), .A2(keyinput_g6), .B1(n2497), .B2(keyinput_g62), 
        .ZN(n4818) );
  OAI221_X1 U5355 ( .B1(n4819), .B2(keyinput_g6), .C1(n2497), .C2(keyinput_g62), .A(n4818), .ZN(n4830) );
  INV_X1 U5356 ( .A(DATAI_6_), .ZN(n4821) );
  AOI22_X1 U5357 ( .A1(n4821), .A2(keyinput_g25), .B1(keyinput_g123), .B2(
        n4988), .ZN(n4820) );
  OAI221_X1 U5358 ( .B1(n4821), .B2(keyinput_g25), .C1(n4988), .C2(
        keyinput_g123), .A(n4820), .ZN(n4829) );
  AOI22_X1 U5359 ( .A1(n4824), .A2(keyinput_g39), .B1(n4823), .B2(
        keyinput_g109), .ZN(n4822) );
  OAI221_X1 U5360 ( .B1(n4824), .B2(keyinput_g39), .C1(n4823), .C2(
        keyinput_g109), .A(n4822), .ZN(n4828) );
  AOI22_X1 U5361 ( .A1(n4826), .A2(keyinput_g111), .B1(n4987), .B2(
        keyinput_g71), .ZN(n4825) );
  OAI221_X1 U5362 ( .B1(n4826), .B2(keyinput_g111), .C1(n4987), .C2(
        keyinput_g71), .A(n4825), .ZN(n4827) );
  NOR4_X1 U5363 ( .A1(n4830), .A2(n4829), .A3(n4828), .A4(n4827), .ZN(n4831)
         );
  NAND4_X1 U5364 ( .A1(n4834), .A2(n4833), .A3(n4832), .A4(n4831), .ZN(n4887)
         );
  AOI22_X1 U5365 ( .A1(n5003), .A2(keyinput_g98), .B1(n2705), .B2(keyinput_g74), .ZN(n4835) );
  OAI221_X1 U5366 ( .B1(n5003), .B2(keyinput_g98), .C1(n2705), .C2(
        keyinput_g74), .A(n4835), .ZN(n4843) );
  AOI22_X1 U5367 ( .A1(n5034), .A2(keyinput_g19), .B1(keyinput_g122), .B2(
        n3124), .ZN(n4836) );
  OAI221_X1 U5368 ( .B1(n5034), .B2(keyinput_g19), .C1(n3124), .C2(
        keyinput_g122), .A(n4836), .ZN(n4842) );
  AOI22_X1 U5369 ( .A1(n4999), .A2(keyinput_g91), .B1(keyinput_g119), .B2(
        n4983), .ZN(n4837) );
  OAI221_X1 U5370 ( .B1(n4999), .B2(keyinput_g91), .C1(n4983), .C2(
        keyinput_g119), .A(n4837), .ZN(n4841) );
  AOI22_X1 U5371 ( .A1(n4839), .A2(keyinput_g97), .B1(n2541), .B2(keyinput_g66), .ZN(n4838) );
  OAI221_X1 U5372 ( .B1(n4839), .B2(keyinput_g97), .C1(n2541), .C2(
        keyinput_g66), .A(n4838), .ZN(n4840) );
  NOR4_X1 U5373 ( .A1(n4843), .A2(n4842), .A3(n4841), .A4(n4840), .ZN(n4885)
         );
  AOI22_X1 U5374 ( .A1(n4845), .A2(keyinput_g114), .B1(keyinput_g100), .B2(
        n5000), .ZN(n4844) );
  OAI221_X1 U5375 ( .B1(n4845), .B2(keyinput_g114), .C1(n5000), .C2(
        keyinput_g100), .A(n4844), .ZN(n4856) );
  AOI22_X1 U5376 ( .A1(n4847), .A2(keyinput_g3), .B1(n3733), .B2(keyinput_g40), 
        .ZN(n4846) );
  OAI221_X1 U5377 ( .B1(n4847), .B2(keyinput_g3), .C1(n3733), .C2(keyinput_g40), .A(n4846), .ZN(n4855) );
  INV_X1 U5378 ( .A(DATAI_5_), .ZN(n4850) );
  AOI22_X1 U5379 ( .A1(n4850), .A2(keyinput_g26), .B1(n4849), .B2(keyinput_g89), .ZN(n4848) );
  OAI221_X1 U5380 ( .B1(n4850), .B2(keyinput_g26), .C1(n4849), .C2(
        keyinput_g89), .A(n4848), .ZN(n4854) );
  AOI22_X1 U5381 ( .A1(n2452), .A2(keyinput_g59), .B1(keyinput_g2), .B2(n4852), 
        .ZN(n4851) );
  OAI221_X1 U5382 ( .B1(n2452), .B2(keyinput_g59), .C1(n4852), .C2(keyinput_g2), .A(n4851), .ZN(n4853) );
  NOR4_X1 U5383 ( .A1(n4856), .A2(n4855), .A3(n4854), .A4(n4853), .ZN(n4884)
         );
  XOR2_X1 U5384 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_g52), .Z(n4859) );
  XOR2_X1 U5385 ( .A(DATAI_24_), .B(keyinput_g7), .Z(n4858) );
  XNOR2_X1 U5386 ( .A(n5031), .B(keyinput_g43), .ZN(n4857) );
  NOR3_X1 U5387 ( .A1(n4859), .A2(n4858), .A3(n4857), .ZN(n4862) );
  XNOR2_X1 U5388 ( .A(DATAI_4_), .B(keyinput_g27), .ZN(n4861) );
  XNOR2_X1 U5389 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_g79), .ZN(n4860) );
  NAND3_X1 U5390 ( .A1(n4862), .A2(n4861), .A3(n4860), .ZN(n4868) );
  INV_X1 U5391 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4864) );
  AOI22_X1 U5392 ( .A1(n4865), .A2(keyinput_g44), .B1(keyinput_g124), .B2(
        n4864), .ZN(n4863) );
  OAI221_X1 U5393 ( .B1(n4865), .B2(keyinput_g44), .C1(n4864), .C2(
        keyinput_g124), .A(n4863), .ZN(n4867) );
  XNOR2_X1 U5394 ( .A(n5014), .B(keyinput_g116), .ZN(n4866) );
  NOR3_X1 U5395 ( .A1(n4868), .A2(n4867), .A3(n4866), .ZN(n4883) );
  INV_X1 U5396 ( .A(IR_REG_26__SCAN_IN), .ZN(n4870) );
  AOI22_X1 U5397 ( .A1(n4871), .A2(keyinput_g21), .B1(n4870), .B2(keyinput_g81), .ZN(n4869) );
  OAI221_X1 U5398 ( .B1(n4871), .B2(keyinput_g21), .C1(n4870), .C2(
        keyinput_g81), .A(n4869), .ZN(n4881) );
  INV_X1 U5399 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4873) );
  AOI22_X1 U5400 ( .A1(n5032), .A2(keyinput_g13), .B1(n4873), .B2(keyinput_g45), .ZN(n4872) );
  OAI221_X1 U5401 ( .B1(n5032), .B2(keyinput_g13), .C1(n4873), .C2(
        keyinput_g45), .A(n4872), .ZN(n4880) );
  INV_X1 U5402 ( .A(IR_REG_15__SCAN_IN), .ZN(n4874) );
  XOR2_X1 U5403 ( .A(n4874), .B(keyinput_g70), .Z(n4878) );
  XOR2_X1 U5404 ( .A(n2534), .B(keyinput_g20), .Z(n4877) );
  XNOR2_X1 U5405 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_g64), .ZN(n4876) );
  XNOR2_X1 U5406 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_g68), .ZN(n4875) );
  NAND4_X1 U5407 ( .A1(n4878), .A2(n4877), .A3(n4876), .A4(n4875), .ZN(n4879)
         );
  NOR3_X1 U5408 ( .A1(n4881), .A2(n4880), .A3(n4879), .ZN(n4882) );
  NAND4_X1 U5409 ( .A1(n4885), .A2(n4884), .A3(n4883), .A4(n4882), .ZN(n4886)
         );
  NOR4_X1 U5410 ( .A1(n4889), .A2(n4888), .A3(n4887), .A4(n4886), .ZN(n5081)
         );
  XOR2_X1 U5411 ( .A(keyinput_g105), .B(keyinput_f105), .Z(n5079) );
  AOI22_X1 U5412 ( .A1(REG3_REG_24__SCAN_IN), .A2(keyinput_f49), .B1(
        REG3_REG_27__SCAN_IN), .B2(keyinput_f34), .ZN(n4890) );
  OAI221_X1 U5413 ( .B1(REG3_REG_24__SCAN_IN), .B2(keyinput_f49), .C1(
        REG3_REG_27__SCAN_IN), .C2(keyinput_f34), .A(n4890), .ZN(n4897) );
  AOI22_X1 U5414 ( .A1(DATAI_1_), .A2(keyinput_f30), .B1(STATE_REG_SCAN_IN), 
        .B2(keyinput_f32), .ZN(n4891) );
  OAI221_X1 U5415 ( .B1(DATAI_1_), .B2(keyinput_f30), .C1(STATE_REG_SCAN_IN), 
        .C2(keyinput_f32), .A(n4891), .ZN(n4896) );
  AOI22_X1 U5416 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(REG3_REG_0__SCAN_IN), 
        .B2(keyinput_f52), .ZN(n4892) );
  OAI221_X1 U5417 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(REG3_REG_0__SCAN_IN), 
        .C2(keyinput_f52), .A(n4892), .ZN(n4895) );
  XNOR2_X1 U5418 ( .A(n4893), .B(keyinput_f68), .ZN(n4894) );
  NOR4_X1 U5419 ( .A1(n4897), .A2(n4896), .A3(n4895), .A4(n4894), .ZN(n4925)
         );
  AOI22_X1 U5420 ( .A1(DATAI_29_), .A2(keyinput_f2), .B1(REG3_REG_20__SCAN_IN), 
        .B2(keyinput_f53), .ZN(n4898) );
  OAI221_X1 U5421 ( .B1(DATAI_29_), .B2(keyinput_f2), .C1(REG3_REG_20__SCAN_IN), .C2(keyinput_f53), .A(n4898), .ZN(n4905) );
  AOI22_X1 U5422 ( .A1(DATAI_17_), .A2(keyinput_f14), .B1(REG3_REG_3__SCAN_IN), 
        .B2(keyinput_f38), .ZN(n4899) );
  OAI221_X1 U5423 ( .B1(DATAI_17_), .B2(keyinput_f14), .C1(REG3_REG_3__SCAN_IN), .C2(keyinput_f38), .A(n4899), .ZN(n4904) );
  AOI22_X1 U5424 ( .A1(REG3_REG_14__SCAN_IN), .A2(keyinput_f35), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput_f55), .ZN(n4900) );
  OAI221_X1 U5425 ( .B1(REG3_REG_14__SCAN_IN), .B2(keyinput_f35), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput_f55), .A(n4900), .ZN(n4903) );
  AOI22_X1 U5426 ( .A1(D_REG_19__SCAN_IN), .A2(keyinput_f106), .B1(
        D_REG_31__SCAN_IN), .B2(keyinput_f118), .ZN(n4901) );
  OAI221_X1 U5427 ( .B1(D_REG_19__SCAN_IN), .B2(keyinput_f106), .C1(
        D_REG_31__SCAN_IN), .C2(keyinput_f118), .A(n4901), .ZN(n4902) );
  NOR4_X1 U5428 ( .A1(n4905), .A2(n4904), .A3(n4903), .A4(n4902), .ZN(n4924)
         );
  AOI22_X1 U5429 ( .A1(D_REG_15__SCAN_IN), .A2(keyinput_f102), .B1(
        D_REG_17__SCAN_IN), .B2(keyinput_f104), .ZN(n4906) );
  OAI221_X1 U5430 ( .B1(D_REG_15__SCAN_IN), .B2(keyinput_f102), .C1(
        D_REG_17__SCAN_IN), .C2(keyinput_f104), .A(n4906), .ZN(n4913) );
  AOI22_X1 U5431 ( .A1(D_REG_12__SCAN_IN), .A2(keyinput_f99), .B1(
        D_REG_14__SCAN_IN), .B2(keyinput_f101), .ZN(n4907) );
  OAI221_X1 U5432 ( .B1(D_REG_12__SCAN_IN), .B2(keyinput_f99), .C1(
        D_REG_14__SCAN_IN), .C2(keyinput_f101), .A(n4907), .ZN(n4912) );
  AOI22_X1 U5433 ( .A1(D_REG_8__SCAN_IN), .A2(keyinput_f95), .B1(
        D_REG_9__SCAN_IN), .B2(keyinput_f96), .ZN(n4908) );
  OAI221_X1 U5434 ( .B1(D_REG_8__SCAN_IN), .B2(keyinput_f95), .C1(
        D_REG_9__SCAN_IN), .C2(keyinput_f96), .A(n4908), .ZN(n4911) );
  AOI22_X1 U5435 ( .A1(D_REG_3__SCAN_IN), .A2(keyinput_f90), .B1(
        D_REG_7__SCAN_IN), .B2(keyinput_f94), .ZN(n4909) );
  OAI221_X1 U5436 ( .B1(D_REG_3__SCAN_IN), .B2(keyinput_f90), .C1(
        D_REG_7__SCAN_IN), .C2(keyinput_f94), .A(n4909), .ZN(n4910) );
  NOR4_X1 U5437 ( .A1(n4913), .A2(n4912), .A3(n4911), .A4(n4910), .ZN(n4923)
         );
  AOI22_X1 U5438 ( .A1(IR_REG_30__SCAN_IN), .A2(keyinput_f85), .B1(
        IR_REG_31__SCAN_IN), .B2(keyinput_f86), .ZN(n4914) );
  OAI221_X1 U5439 ( .B1(IR_REG_30__SCAN_IN), .B2(keyinput_f85), .C1(
        IR_REG_31__SCAN_IN), .C2(keyinput_f86), .A(n4914), .ZN(n4921) );
  AOI22_X1 U5440 ( .A1(IR_REG_15__SCAN_IN), .A2(keyinput_f70), .B1(
        IR_REG_18__SCAN_IN), .B2(keyinput_f73), .ZN(n4915) );
  OAI221_X1 U5441 ( .B1(IR_REG_15__SCAN_IN), .B2(keyinput_f70), .C1(
        IR_REG_18__SCAN_IN), .C2(keyinput_f73), .A(n4915), .ZN(n4920) );
  AOI22_X1 U5442 ( .A1(DATAI_9_), .A2(keyinput_f22), .B1(DATAI_14_), .B2(
        keyinput_f17), .ZN(n4916) );
  OAI221_X1 U5443 ( .B1(DATAI_9_), .B2(keyinput_f22), .C1(DATAI_14_), .C2(
        keyinput_f17), .A(n4916), .ZN(n4919) );
  AOI22_X1 U5444 ( .A1(REG0_REG_6__SCAN_IN), .A2(keyinput_f125), .B1(
        IR_REG_12__SCAN_IN), .B2(keyinput_f67), .ZN(n4917) );
  OAI221_X1 U5445 ( .B1(REG0_REG_6__SCAN_IN), .B2(keyinput_f125), .C1(
        IR_REG_12__SCAN_IN), .C2(keyinput_f67), .A(n4917), .ZN(n4918) );
  NOR4_X1 U5446 ( .A1(n4921), .A2(n4920), .A3(n4919), .A4(n4918), .ZN(n4922)
         );
  NAND4_X1 U5447 ( .A1(n4925), .A2(n4924), .A3(n4923), .A4(n4922), .ZN(n5075)
         );
  AOI22_X1 U5448 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(IR_REG_11__SCAN_IN), 
        .B2(keyinput_f66), .ZN(n4926) );
  OAI221_X1 U5449 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(IR_REG_11__SCAN_IN), 
        .C2(keyinput_f66), .A(n4926), .ZN(n4933) );
  AOI22_X1 U5450 ( .A1(REG0_REG_5__SCAN_IN), .A2(keyinput_f124), .B1(
        REG0_REG_7__SCAN_IN), .B2(keyinput_f126), .ZN(n4927) );
  OAI221_X1 U5451 ( .B1(REG0_REG_5__SCAN_IN), .B2(keyinput_f124), .C1(
        REG0_REG_7__SCAN_IN), .C2(keyinput_f126), .A(n4927), .ZN(n4932) );
  AOI22_X1 U5452 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput_f47), .B1(
        IR_REG_3__SCAN_IN), .B2(keyinput_f58), .ZN(n4928) );
  OAI221_X1 U5453 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput_f47), .C1(
        IR_REG_3__SCAN_IN), .C2(keyinput_f58), .A(n4928), .ZN(n4931) );
  AOI22_X1 U5454 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput_f50), .B1(
        IR_REG_1__SCAN_IN), .B2(keyinput_f56), .ZN(n4929) );
  OAI221_X1 U5455 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput_f50), .C1(
        IR_REG_1__SCAN_IN), .C2(keyinput_f56), .A(n4929), .ZN(n4930) );
  NOR4_X1 U5456 ( .A1(n4933), .A2(n4932), .A3(n4931), .A4(n4930), .ZN(n4961)
         );
  AOI22_X1 U5457 ( .A1(REG0_REG_2__SCAN_IN), .A2(keyinput_f121), .B1(
        IR_REG_2__SCAN_IN), .B2(keyinput_f57), .ZN(n4934) );
  OAI221_X1 U5458 ( .B1(REG0_REG_2__SCAN_IN), .B2(keyinput_f121), .C1(
        IR_REG_2__SCAN_IN), .C2(keyinput_f57), .A(n4934), .ZN(n4941) );
  AOI22_X1 U5459 ( .A1(IR_REG_8__SCAN_IN), .A2(keyinput_f63), .B1(
        IR_REG_20__SCAN_IN), .B2(keyinput_f75), .ZN(n4935) );
  OAI221_X1 U5460 ( .B1(IR_REG_8__SCAN_IN), .B2(keyinput_f63), .C1(
        IR_REG_20__SCAN_IN), .C2(keyinput_f75), .A(n4935), .ZN(n4940) );
  AOI22_X1 U5461 ( .A1(D_REG_22__SCAN_IN), .A2(keyinput_f109), .B1(
        IR_REG_22__SCAN_IN), .B2(keyinput_f77), .ZN(n4936) );
  OAI221_X1 U5462 ( .B1(D_REG_22__SCAN_IN), .B2(keyinput_f109), .C1(
        IR_REG_22__SCAN_IN), .C2(keyinput_f77), .A(n4936), .ZN(n4939) );
  AOI22_X1 U5463 ( .A1(D_REG_26__SCAN_IN), .A2(keyinput_f113), .B1(
        D_REG_24__SCAN_IN), .B2(keyinput_f111), .ZN(n4937) );
  OAI221_X1 U5464 ( .B1(D_REG_26__SCAN_IN), .B2(keyinput_f113), .C1(
        D_REG_24__SCAN_IN), .C2(keyinput_f111), .A(n4937), .ZN(n4938) );
  NOR4_X1 U5465 ( .A1(n4941), .A2(n4940), .A3(n4939), .A4(n4938), .ZN(n4960)
         );
  AOI22_X1 U5466 ( .A1(D_REG_10__SCAN_IN), .A2(keyinput_f97), .B1(
        D_REG_25__SCAN_IN), .B2(keyinput_f112), .ZN(n4942) );
  OAI221_X1 U5467 ( .B1(D_REG_10__SCAN_IN), .B2(keyinput_f97), .C1(
        D_REG_25__SCAN_IN), .C2(keyinput_f112), .A(n4942), .ZN(n4949) );
  AOI22_X1 U5468 ( .A1(D_REG_2__SCAN_IN), .A2(keyinput_f89), .B1(
        D_REG_27__SCAN_IN), .B2(keyinput_f114), .ZN(n4943) );
  OAI221_X1 U5469 ( .B1(D_REG_2__SCAN_IN), .B2(keyinput_f89), .C1(
        D_REG_27__SCAN_IN), .C2(keyinput_f114), .A(n4943), .ZN(n4948) );
  AOI22_X1 U5470 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput_f45), .B1(
        D_REG_0__SCAN_IN), .B2(keyinput_f87), .ZN(n4944) );
  OAI221_X1 U5471 ( .B1(REG3_REG_25__SCAN_IN), .B2(keyinput_f45), .C1(
        D_REG_0__SCAN_IN), .C2(keyinput_f87), .A(n4944), .ZN(n4947) );
  AOI22_X1 U5472 ( .A1(DATAI_5_), .A2(keyinput_f26), .B1(IR_REG_29__SCAN_IN), 
        .B2(keyinput_f84), .ZN(n4945) );
  OAI221_X1 U5473 ( .B1(DATAI_5_), .B2(keyinput_f26), .C1(IR_REG_29__SCAN_IN), 
        .C2(keyinput_f84), .A(n4945), .ZN(n4946) );
  NOR4_X1 U5474 ( .A1(n4949), .A2(n4948), .A3(n4947), .A4(n4946), .ZN(n4959)
         );
  AOI22_X1 U5475 ( .A1(DATAI_28_), .A2(keyinput_f3), .B1(IR_REG_21__SCAN_IN), 
        .B2(keyinput_f76), .ZN(n4950) );
  OAI221_X1 U5476 ( .B1(DATAI_28_), .B2(keyinput_f3), .C1(IR_REG_21__SCAN_IN), 
        .C2(keyinput_f76), .A(n4950), .ZN(n4957) );
  AOI22_X1 U5477 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(IR_REG_24__SCAN_IN), 
        .B2(keyinput_f79), .ZN(n4951) );
  OAI221_X1 U5478 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(IR_REG_24__SCAN_IN), 
        .C2(keyinput_f79), .A(n4951), .ZN(n4956) );
  AOI22_X1 U5479 ( .A1(DATAI_10_), .A2(keyinput_f21), .B1(REG3_REG_12__SCAN_IN), .B2(keyinput_f44), .ZN(n4952) );
  OAI221_X1 U5480 ( .B1(DATAI_10_), .B2(keyinput_f21), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput_f44), .A(n4952), .ZN(n4955) );
  AOI22_X1 U5481 ( .A1(IR_REG_9__SCAN_IN), .A2(keyinput_f64), .B1(
        IR_REG_26__SCAN_IN), .B2(keyinput_f81), .ZN(n4953) );
  OAI221_X1 U5482 ( .B1(IR_REG_9__SCAN_IN), .B2(keyinput_f64), .C1(
        IR_REG_26__SCAN_IN), .C2(keyinput_f81), .A(n4953), .ZN(n4954) );
  NOR4_X1 U5483 ( .A1(n4957), .A2(n4956), .A3(n4955), .A4(n4954), .ZN(n4958)
         );
  NAND4_X1 U5484 ( .A1(n4961), .A2(n4960), .A3(n4959), .A4(n4958), .ZN(n5074)
         );
  AOI22_X1 U5485 ( .A1(DATAI_11_), .A2(keyinput_f20), .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_f39), .ZN(n4962) );
  OAI221_X1 U5486 ( .B1(DATAI_11_), .B2(keyinput_f20), .C1(
        REG3_REG_19__SCAN_IN), .C2(keyinput_f39), .A(n4962), .ZN(n4969) );
  AOI22_X1 U5487 ( .A1(DATAI_6_), .A2(keyinput_f25), .B1(DATAI_25_), .B2(
        keyinput_f6), .ZN(n4963) );
  OAI221_X1 U5488 ( .B1(DATAI_6_), .B2(keyinput_f25), .C1(DATAI_25_), .C2(
        keyinput_f6), .A(n4963), .ZN(n4968) );
  AOI22_X1 U5489 ( .A1(IR_REG_10__SCAN_IN), .A2(keyinput_f65), .B1(
        IR_REG_25__SCAN_IN), .B2(keyinput_f80), .ZN(n4964) );
  OAI221_X1 U5490 ( .B1(IR_REG_10__SCAN_IN), .B2(keyinput_f65), .C1(
        IR_REG_25__SCAN_IN), .C2(keyinput_f80), .A(n4964), .ZN(n4967) );
  AOI22_X1 U5491 ( .A1(DATAI_27_), .A2(keyinput_f4), .B1(IR_REG_6__SCAN_IN), 
        .B2(keyinput_f61), .ZN(n4965) );
  OAI221_X1 U5492 ( .B1(DATAI_27_), .B2(keyinput_f4), .C1(IR_REG_6__SCAN_IN), 
        .C2(keyinput_f61), .A(n4965), .ZN(n4966) );
  NOR4_X1 U5493 ( .A1(n4969), .A2(n4968), .A3(n4967), .A4(n4966), .ZN(n5011)
         );
  AOI22_X1 U5494 ( .A1(IR_REG_23__SCAN_IN), .A2(keyinput_f78), .B1(n3733), 
        .B2(keyinput_f40), .ZN(n4970) );
  OAI221_X1 U5495 ( .B1(IR_REG_23__SCAN_IN), .B2(keyinput_f78), .C1(n3733), 
        .C2(keyinput_f40), .A(n4970), .ZN(n4980) );
  AOI22_X1 U5496 ( .A1(n4973), .A2(keyinput_f0), .B1(n4972), .B2(keyinput_f10), 
        .ZN(n4971) );
  OAI221_X1 U5497 ( .B1(n4973), .B2(keyinput_f0), .C1(n4972), .C2(keyinput_f10), .A(n4971), .ZN(n4979) );
  AOI22_X1 U5498 ( .A1(DATAI_26_), .A2(keyinput_f5), .B1(IR_REG_17__SCAN_IN), 
        .B2(keyinput_f72), .ZN(n4974) );
  OAI221_X1 U5499 ( .B1(DATAI_26_), .B2(keyinput_f5), .C1(IR_REG_17__SCAN_IN), 
        .C2(keyinput_f72), .A(n4974), .ZN(n4978) );
  XNOR2_X1 U5500 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_f82), .ZN(n4976) );
  XNOR2_X1 U5501 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_f42), .ZN(n4975) );
  NAND2_X1 U5502 ( .A1(n4976), .A2(n4975), .ZN(n4977) );
  NOR4_X1 U5503 ( .A1(n4980), .A2(n4979), .A3(n4978), .A4(n4977), .ZN(n5010)
         );
  AOI22_X1 U5504 ( .A1(n4983), .A2(keyinput_f119), .B1(n4982), .B2(
        keyinput_f120), .ZN(n4981) );
  OAI221_X1 U5505 ( .B1(n4983), .B2(keyinput_f119), .C1(n4982), .C2(
        keyinput_f120), .A(n4981), .ZN(n4994) );
  AOI22_X1 U5506 ( .A1(n2548), .A2(keyinput_f54), .B1(keyinput_f33), .B2(n4985), .ZN(n4984) );
  OAI221_X1 U5507 ( .B1(n2548), .B2(keyinput_f54), .C1(n4985), .C2(
        keyinput_f33), .A(n4984), .ZN(n4993) );
  AOI22_X1 U5508 ( .A1(n2364), .A2(keyinput_f69), .B1(keyinput_f71), .B2(n4987), .ZN(n4986) );
  OAI221_X1 U5509 ( .B1(n2364), .B2(keyinput_f69), .C1(n4987), .C2(
        keyinput_f71), .A(n4986), .ZN(n4992) );
  XOR2_X1 U5510 ( .A(n4988), .B(keyinput_f123), .Z(n4990) );
  XNOR2_X1 U5511 ( .A(DATAI_4_), .B(keyinput_f27), .ZN(n4989) );
  NAND2_X1 U5512 ( .A1(n4990), .A2(n4989), .ZN(n4991) );
  NOR4_X1 U5513 ( .A1(n4994), .A2(n4993), .A3(n4992), .A4(n4991), .ZN(n5009)
         );
  AOI22_X1 U5514 ( .A1(n3124), .A2(keyinput_f122), .B1(n4996), .B2(
        keyinput_f127), .ZN(n4995) );
  OAI221_X1 U5515 ( .B1(n3124), .B2(keyinput_f122), .C1(n4996), .C2(
        keyinput_f127), .A(n4995), .ZN(n5007) );
  AOI22_X1 U5516 ( .A1(n2497), .A2(keyinput_f62), .B1(keyinput_f51), .B2(n2502), .ZN(n4997) );
  OAI221_X1 U5517 ( .B1(n2497), .B2(keyinput_f62), .C1(n2502), .C2(
        keyinput_f51), .A(n4997), .ZN(n5006) );
  AOI22_X1 U5518 ( .A1(n5000), .A2(keyinput_f100), .B1(keyinput_f91), .B2(
        n4999), .ZN(n4998) );
  OAI221_X1 U5519 ( .B1(n5000), .B2(keyinput_f100), .C1(n4999), .C2(
        keyinput_f91), .A(n4998), .ZN(n5005) );
  AOI22_X1 U5520 ( .A1(n5003), .A2(keyinput_f98), .B1(keyinput_f117), .B2(
        n5002), .ZN(n5001) );
  OAI221_X1 U5521 ( .B1(n5003), .B2(keyinput_f98), .C1(n5002), .C2(
        keyinput_f117), .A(n5001), .ZN(n5004) );
  NOR4_X1 U5522 ( .A1(n5007), .A2(n5006), .A3(n5005), .A4(n5004), .ZN(n5008)
         );
  NAND4_X1 U5523 ( .A1(n5011), .A2(n5010), .A3(n5009), .A4(n5008), .ZN(n5073)
         );
  AOI22_X1 U5524 ( .A1(n5014), .A2(keyinput_f116), .B1(keyinput_f92), .B2(
        n5013), .ZN(n5012) );
  OAI221_X1 U5525 ( .B1(n5014), .B2(keyinput_f116), .C1(n5013), .C2(
        keyinput_f92), .A(n5012), .ZN(n5027) );
  AOI22_X1 U5526 ( .A1(n5017), .A2(keyinput_f107), .B1(keyinput_f103), .B2(
        n5016), .ZN(n5015) );
  OAI221_X1 U5527 ( .B1(n5017), .B2(keyinput_f107), .C1(n5016), .C2(
        keyinput_f103), .A(n5015), .ZN(n5026) );
  AOI22_X1 U5528 ( .A1(n5020), .A2(keyinput_f110), .B1(keyinput_f108), .B2(
        n5019), .ZN(n5018) );
  OAI221_X1 U5529 ( .B1(n5020), .B2(keyinput_f110), .C1(n5019), .C2(
        keyinput_f108), .A(n5018), .ZN(n5025) );
  AOI22_X1 U5530 ( .A1(n5023), .A2(keyinput_f93), .B1(n5022), .B2(
        keyinput_f115), .ZN(n5021) );
  OAI221_X1 U5531 ( .B1(n5023), .B2(keyinput_f93), .C1(n5022), .C2(
        keyinput_f115), .A(n5021), .ZN(n5024) );
  NOR4_X1 U5532 ( .A1(n5027), .A2(n5026), .A3(n5025), .A4(n5024), .ZN(n5071)
         );
  INV_X1 U5533 ( .A(DATAI_19_), .ZN(n5029) );
  AOI22_X1 U5534 ( .A1(n2397), .A2(keyinput_f48), .B1(keyinput_f12), .B2(n5029), .ZN(n5028) );
  OAI221_X1 U5535 ( .B1(n2397), .B2(keyinput_f48), .C1(n5029), .C2(
        keyinput_f12), .A(n5028), .ZN(n5040) );
  AOI22_X1 U5536 ( .A1(n5032), .A2(keyinput_f13), .B1(n5031), .B2(keyinput_f43), .ZN(n5030) );
  OAI221_X1 U5537 ( .B1(n5032), .B2(keyinput_f13), .C1(n5031), .C2(
        keyinput_f43), .A(n5030), .ZN(n5039) );
  AOI22_X1 U5538 ( .A1(n2452), .A2(keyinput_f59), .B1(keyinput_f19), .B2(n5034), .ZN(n5033) );
  OAI221_X1 U5539 ( .B1(n2452), .B2(keyinput_f59), .C1(n5034), .C2(
        keyinput_f19), .A(n5033), .ZN(n5038) );
  AOI22_X1 U5540 ( .A1(n2705), .A2(keyinput_f74), .B1(keyinput_f8), .B2(n5036), 
        .ZN(n5035) );
  OAI221_X1 U5541 ( .B1(n2705), .B2(keyinput_f74), .C1(n5036), .C2(keyinput_f8), .A(n5035), .ZN(n5037) );
  NOR4_X1 U5542 ( .A1(n5040), .A2(n5039), .A3(n5038), .A4(n5037), .ZN(n5070)
         );
  AOI22_X1 U5543 ( .A1(n2487), .A2(keyinput_f24), .B1(keyinput_f31), .B2(n2257), .ZN(n5041) );
  OAI221_X1 U5544 ( .B1(n2487), .B2(keyinput_f24), .C1(n2257), .C2(
        keyinput_f31), .A(n5041), .ZN(n5051) );
  INV_X1 U5545 ( .A(DATAI_22_), .ZN(n5043) );
  AOI22_X1 U5546 ( .A1(n5044), .A2(keyinput_f16), .B1(n5043), .B2(keyinput_f9), 
        .ZN(n5042) );
  OAI221_X1 U5547 ( .B1(n5044), .B2(keyinput_f16), .C1(n5043), .C2(keyinput_f9), .A(n5042), .ZN(n5050) );
  XNOR2_X1 U5548 ( .A(DATAI_8_), .B(keyinput_f23), .ZN(n5048) );
  XNOR2_X1 U5549 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_f83), .ZN(n5047) );
  XNOR2_X1 U5550 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_f60), .ZN(n5046) );
  XNOR2_X1 U5551 ( .A(DATAI_2_), .B(keyinput_f29), .ZN(n5045) );
  NAND4_X1 U5552 ( .A1(n5048), .A2(n5047), .A3(n5046), .A4(n5045), .ZN(n5049)
         );
  NOR3_X1 U5553 ( .A1(n5051), .A2(n5050), .A3(n5049), .ZN(n5069) );
  AOI22_X1 U5554 ( .A1(n5054), .A2(keyinput_f36), .B1(keyinput_f15), .B2(n5053), .ZN(n5052) );
  OAI221_X1 U5555 ( .B1(n5054), .B2(keyinput_f36), .C1(n5053), .C2(
        keyinput_f15), .A(n5052), .ZN(n5067) );
  AOI22_X1 U5556 ( .A1(n5057), .A2(keyinput_f46), .B1(keyinput_f41), .B2(n5056), .ZN(n5055) );
  OAI221_X1 U5557 ( .B1(n5057), .B2(keyinput_f46), .C1(n5056), .C2(
        keyinput_f41), .A(n5055), .ZN(n5066) );
  INV_X1 U5558 ( .A(REG3_REG_10__SCAN_IN), .ZN(n5060) );
  INV_X1 U5559 ( .A(DATAI_3_), .ZN(n5059) );
  AOI22_X1 U5560 ( .A1(n5060), .A2(keyinput_f37), .B1(keyinput_f28), .B2(n5059), .ZN(n5058) );
  OAI221_X1 U5561 ( .B1(n5060), .B2(keyinput_f37), .C1(n5059), .C2(
        keyinput_f28), .A(n5058), .ZN(n5065) );
  AOI22_X1 U5562 ( .A1(n5063), .A2(keyinput_f88), .B1(keyinput_f11), .B2(n5062), .ZN(n5061) );
  OAI221_X1 U5563 ( .B1(n5063), .B2(keyinput_f88), .C1(n5062), .C2(
        keyinput_f11), .A(n5061), .ZN(n5064) );
  NOR4_X1 U5564 ( .A1(n5067), .A2(n5066), .A3(n5065), .A4(n5064), .ZN(n5068)
         );
  NAND4_X1 U5565 ( .A1(n5071), .A2(n5070), .A3(n5069), .A4(n5068), .ZN(n5072)
         );
  NOR4_X1 U5566 ( .A1(n5075), .A2(n5074), .A3(n5073), .A4(n5072), .ZN(n5078)
         );
  NAND2_X1 U5567 ( .A1(keyinput_g105), .A2(n5077), .ZN(n5076) );
  OAI221_X1 U5568 ( .B1(n5079), .B2(n5078), .C1(keyinput_g105), .C2(n5077), 
        .A(n5076), .ZN(n5080) );
  AOI21_X1 U5569 ( .B1(n5082), .B2(n5081), .A(n5080), .ZN(n5084) );
  AOI22_X1 U5570 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n5083) );
  XNOR2_X1 U5571 ( .A(n5084), .B(n5083), .ZN(U3352) );
  INV_X1 U2481 ( .A(IR_REG_16__SCAN_IN), .ZN(n4987) );
  CLKBUF_X1 U3021 ( .A(n2423), .Z(n2759) );
endmodule

